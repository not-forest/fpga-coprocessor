// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
xZMOwtVumKb+SCLkrOB+ut0IT5kAeqshseNF3FIHKvS98U290bh/wwZjooLTFBln
dPFtcRuXRjEn5/FrC0wE1XIlKJP7J+QFcykW4u2ws3LeEUveYZxFRxmcS1ygpbyA
IXOXT0yvhlyRuxd/FRFQCTvIMV7TL+G4aoXTs6TDZyk=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 52352 )
`pragma protect data_block
DqB4p2Bq9RY2A4KcpsJnCCIsvTKoJJYQnp9tZWpdo2XBk19qbShY0gpLgWR7BRLd
yLGl4iMKK7mb7gxvAbaCkrwB9Ffg1UxdIzko6tU1NhrMAFMq5WJQQzbYqkXT6/OF
sfgTVSsVdU2fn/glBSvZtJBOMVtAFQnYbXctbRPRck5y3DCogRhs6cR0Dj3hjPDW
RbHBsTkHwY0rb1ELJrccMbhgs85zcNA1Naz5AQT8+jjeIIbEiRUmC+Wj8tztYVCT
3yo9KcM0AUty5JErjjNUWlfZdVRwBQSbjSuKIF/aREpem7pDlJokIh1I5bmWVm/s
TIJpn5FllbGm8urTvY4vz/sbgis3ll0z/1OkUva0ITwDsg16MkzydoLpGX6s4LG/
guIMWbW6Inmlm3qwLJhSm35mPcfypvS5DlkY0WHjprc08sl+ZaH2k1Ssh6kjU97Y
/koBEwhWpomzICobOm3BBzF1p40EG7b1n9lwVhJiDmxqE49RclroTIxsWOAAoZQl
R6v/cchdZesvPqrKMDYJJi/8zMbu1+BGnbe+F93X3Exn5hj6TKBAPWM3tZ7mDez3
fWEtulHuzc4dUvhASTguDEojZXv7TFYtLe1cDYkUhEGrV54405CPwxVtrl54XGL7
mSfgpaoEeW/ne+H4QBwQOovxv/kL4oZ/J+hl5Vi5pyMlvExx55H+UY6w3CtHjcQY
XU2G2atvmCenSiik6PchzmVinamz0KfpzbFyaGq9vxjiY6BJQ5FxW4+e5toFYWLf
5CJ7UnIhklYbkuZoFoJ0AXqfScJ0u1haZ4cJ4h19klKSqbqQlvNTBYJ2n9uJjEXq
4yC/2wzMXQ6WiwIEs6+XzJMHaE05I/YK7qJ/ofiTTpP7O8euSL62uh6r6QXoGx5o
4n9MM4P2GCtJ1BjA64VPUbkrTqiLCz0stT9XCoVB3LOVt5BIruP2OVLKx60o2Bch
uf/Wx09e8eaxzEoqHirDhpYrnfIIcqjN63pmK3ky+sdiWx+w8srLTwNjisCN6zs9
QlMMZDsa9ugAxM8ROiyYORHZQDnrg8AKfzovnkmJ5eclvv2Y34pdnY/E07MiRsjr
3gTg/5It8fEiMpKa0FBa584V9Ka5L/6kVnlYlgGjcWAqAHjtZkAXZlbe0qQ0ETxQ
5A+EH/h9IP+elg9Kg5yRgW7RT45Fcpa0iLFPa/P58AFbkV9iZuNcUHBgAIjZt4eb
tEmEtDz0UhrPuH8xyy1lyASYu0pUMLSlNrnPgiKC9NfeNF6zZk/6ihR/hA61peYl
7T0y9dCOSEFCdvh42lhUCNaysPSGMLMDbTTk4Fki+kJs6lbtuaGlOopW67GQJpei
NbRqJmh/TEmbFOVSsu+LTzNTdk31TSM1emELhqtJcMIUlq8b3uB5wG6G97HDTtVB
TFiCaAAqai0hskblNKBiyoNqQKPRh+D3amTWvfYVGJC88jtzqlBYg/kL8U+KzIV2
RxjFBFZW7iHmaXJYK5nUNCKUWrxL344dwODTVJweI6wFrGIxw5b7WOJf/Guxc1dI
ZXi7ydoZgCP7WHRXaEhVmEj1fKPJ+to85V5qAQeVKlHHCsyS/oeWje0MPNs8AxWB
Jv3l1bbRkib5sWHJortqkBxr7XaI36bkNBODnHuXnsedjVyo7XyKVwZDfSLL+Pzo
NddoF8+m5+g4sB7wfx6CTtn3jKyZ6SsTiYKO97iacHBeJiHASE3Dw82qDaXT7aM+
JF1lKiUJcu0wgLWoybcY1fJGCQ5psloWSYh57KFlvoZa2g3zFieuYXt4qHhXK/Wo
VG1cBB/DYGdXzPWoVoC+f5Zq56e1LXmkneuZVjV8L+2FyVmJBF+BNGjnWG9gsJ1G
TapipWUYuONRlD9sOD5BhkLbQ0uhEPqYAEe7ahG/iSndZPfQ1QbVVlPtDsgQO6TF
85vC8RlIn5boRjammyN6CIHfljARlwFLNrw2wIBPT3zDvhvOt05KJhR+Km9F3r1U
kPVjtEzLcAWtmtZGz9afqs9RAO1VLbNCBa7GJGk+iGdUsLrKVxplPBaVy/5dorrm
+156b/lc1522nkkqQMVV9xkyTndfftEv+MFUYfYX6TOCls+YgABkz3te9lPiey3o
8QUk/o8y/hj5R/HRpXOZqTswNR9ZE6POyFks3tBt3Q9amC3kl2k1ewEf2UpLSz+b
EzJv4L7aMeEPKYoeaeVYO1vx4HQBlAC7rAKWNRidqMIZG5rwkpn6ju2/DZQ6rtJT
hAoZ8SDxYp89TAq/4EMQcJYvgwpmYbHGGeVEiEtZ0EHDuy4hT1+E/jNe/JFPKgwS
RVSgoPCc79GeZW0C3p1GX/k1YuHg4B9Icxwdkq6V+5V0wLg8msdlLt32QrCxTzeq
fURe7KPLoaS0KOEG1rT72N9yKyiIle5S3SSPmedyX1hKNi8kgY0nd45PoHoBpu1+
HI/ZbNDVGm+1givvP/cAD9dl1VBflbwpAKFIfVGOB2Zd5s007HCx3qfkb6H6munS
XqKEsWd4F4ahR9iYF1ebu1FthHTyVm6f3mWmSNNwd7cBWYF/rglENwHBrF7sNlF9
MsWa2cRNTWQnEpFxROmnNAQ7cBwLGIEdNvljmDno/l1ECdHRiQiaI9+Uy4sjSFi6
qS2OCsbREqc1UTKh9NCOUqtldw7A++cCnE+D9XtD841Ob2KGgjlnQ5Ukb8wvYIvG
fsbaruYqpqu0tmQoLYKrY9G9Rg0Zq1Q76+rB5tc9Iynn8wDjMXtJbchE+rSs60PA
4oRLOpbXgJSoUnTo9+lL2DV/Nbz3VaUKARRFEsGailIonjgE64HVkLSXhqj6IYey
uGTWOjsgVTLrOYnBfxPM+VD6OcDFwFCn0klT3OgqXjaadNNsWIHLhAEtP5LVPhL7
INnoZNpNBcMn0/uwyt6pz5oT9pEKG923w0waXFsjK5X2TU6jnvgFLiGF5Se7k4NS
HFPJUKDbs8eh3Uz3A50NNIIwC9bdyaqOpWGzyJ5t+UY6HK5Wim6xA56UNWi8de5u
YGu50LlRDwGLbvnc4vg7LJYSa+vii0ZyhTq+xh6jI88EP0H59lqD6glpA34eqn0x
YcjTF5MZZbDsBk4p06z0BvXgpdqlwLLT71xWVW0GRQvRJlKifB+7vMBJQGxOnNN5
PudPYaALqEDTExWcI9/ZbaXvSiv+bwnx6mfyrMW3MY/NBSHj7bbyo4K5skvabMxJ
YRWyB7PnV7/erfqDWHf9hSJto5ofZl99Ijsq++xZdgFEW66hyiuBVKmPpb/0nAPc
/VZRmxeWpbSrJcvaOBZ1YeIZEIIa5HmeoCEq66keBeVi11YfFlG6GK9g7agv+acc
je/Wo+Elij8pyGMrVpsJ3Ly7jm6KAUvplb3SvZ1RbUdamjMZpgilEevyFLjTP2Vt
+CT3AxdjhKZI3Gc9mjqmCgaldHKpj1cqPx3oQT0IDj4utJ5HKIQffVMmwrKpI6wN
ykiaj0awsLzmlaCZON2+xcVCDazG5MRek7UkYvLiIanwMD62AtN7wzGtXpqB376j
8dgzdsO2luAWz7g7um9VW2RrBedKsCnd7I3KYnTPxllsDFT1wHfsFTdzDx/5lzS3
EKIrWnGAJQdcI5DV0m35fKUwbNQ6S6FLX1ZtO5sql0qM/yUzlnCcxCw/dAPfYRUg
ICbIzXlTNQp09K6hJs5LkFRMwGs6bTL2pBG/LW86aW7DY6bJIPAocX8jdna9ikZ8
+mVKPqDohX+X/5ffRmr/VErUosJAi5x8t8W1YL4V42CAP8DMCTX5JI6XVAsMUB8t
7szA9+7642Ld2b6gWiE5rWyeeYtUeWKSabPJ1dT0IFe7rcjR+qOq+8lS7agREhFI
Dg+hG7ouj001LivEochV4SRbltRjYAvOryZl3LIlhXq4MUCpXSnta+LPA0Ek5lZW
212xO8xugQ1W+hzPFmI+UQ5vq0pRrnL2fA6IcpKYGGL8nc9Qybw6w2KSUMN57G9T
s6baoiAVyGC58evp/+LJPTiqxvM3sBr7kC6AUSpP1NOV42uE/zcMi1b+ja0nSMZ3
nJF2AHHGfuKcHboOKlHz5gtwG6p+kSSG5Mkyv/PXY/tOJPCmPWMqAnMqEUNFjHGL
lXRBTO/e2wuB5bKCB7VoiOqMzXasSRDqHnX8jo0+Pq3GGMvfrpocnRACVJd27aYm
UoWtmMQx7WIHUOKSMiJrKzHhcBIW5Ykt4GYBLopBKjOukgL/cOarLjEG+f9nKh7i
6EVtB2I2RqhEDcIWqtt8wlJSlxQYudWgqN2xLRDIsnJc0ZJLo8pvFr82gJSld4Jy
l+YFQeJrfzPOi5pOXNqauVNoC8ut7rfqC0FpU5VPyhFWZ1UYwAR8FOllWekIt3Hg
mNnuI1At7Di/t3+oyviZ5cIOxtkRe27VbTdKRtVyynCWyfWDox9kjGjyFKYxGCF5
Z2zvEmHfH9AYQWPMehVqnXO13KdyNkRohfryxP1qvkXrBwXzrwBmBid4j3x+upJH
4WEvE5WAj24Syn88C6mt21KF/WF4x16w2gd/+fBluh9Q/joU5yWlB8kUMeDndLkk
UGkWietfYDnPqAUSZLKUCGwpbWPoJISdiwF3bG/N/YFKAEXLfQ5wJAfWYPy4WMu1
3bSk2UuZfHo+KXzTA+MLqwFFSBf88K1IZsrWACk9vlEPX4sPZ4oxZXwpsWfSIurA
Ond+AHYD7N4UUtHdZEkc+9nNrBx+aBC2tZ3231uBFfVS7sgS7UMjL8lX37V+wQnB
AdUriEIrbiJL/XLDNGfjJCbT7vBwFZEDWgnqTZ3MsxNBBR/qq+BMDKaGpad7D6A/
cFqDG2O6hoDVI5p9f/yyfzIy6ygDXXrMa/+Z8S/L26Uy83rNHsYpuV3CEJpb/j1o
PyMuZo1twQrUAVCogf8aTGaqedk5YQeq52TQXlC65dH9MfSrd7VvSW0tp63VnTuR
RJMenC2aZExI2ZUrbTXMbZsiVr4IFdxpNz0WXuhjZREPvfUpvUiKOuBYjid82cII
cOUpRNwBzzjtnuT5XLsqKSN0/Z27j8q2j+48sdv8wNmj5q6NILGVBJLkK5dZPQsz
MzIQror2fg/mZuUXkZIqW3EwgZtptJB0P5SUHXysMstKImRHoSgY4VqIykpxhPcG
9zuUIYdK4snP0XBA+mhdJIIZcid55P2mrheon3Sl2uiIEUAPLfHjBb66xiwY2sxU
RaEjsFD+cuXfudMV9X2MDPfTBoqO6y64yLy4Xz+KlpAPjgyPSBACVVcFAzxBEqE6
p8O/Nl30ENZo1yl2IXYy3QH53hhf04S16RO+mynBZhoyqaRDmwUPNGZ/0rrI9B5/
oYCFSjSxNANhNF6dj/bgZFKyxZVm5Ftvoe0tAtR75WuofxyqgYRNgvC4v/fbceTH
hTGTvm13ekAHbx4aDa1EqKqCkdUjDNxwRli6aonNx6OTT2mpXClMnoEthqgxXA4L
oVUQCNNLGR5z58TTrJc8zxi1IdFjOPnChAajClwjkWoN/YGro4VzJup84C8w3EW2
/PzyqifdUDAB0RpWF4B8yLXowjRdU7cVFQgiWPSYwR/4M8//EAHxhpJut+LQq0VO
7wk8d2l4d6qy4cTyxaxeIv55ZheyuXVEZCre1vYTl7rLUjlErng+7JMeT5HGO15K
JWAVOwj97GQD+Gyihy6tsmmEzup6T5i30sYTuW1MOwqEzLl5qzBW1oDck5Rh3S8F
CcUlpHC/nMATEkrhDEG2BzZva8aK8TMVGtjiEpdKwGcwVaE90bnWorbmR1AmuFmv
898UAUSus4lQ7tdGR7bE1etkkyTpNUb07YlawFUTcCkSBGCEArAMJSvVMYE8Srdy
tiSrMlsCvzeGlrIorQsZmYO9HGeVI6z2/izP3eCQ9tEv+3CI5x5ouj2oQh95sq0m
tD80oxbTaYJGsQKBmP3HtLTcXrvrlYP+nX+y2kOW10M4SyTUtY7XsUQWinHKfL45
cDbgLG8ytyPs+4CReFLME6500PpQ63ccl0jcouZ95OID0WZ0MaPBb1BQSqYHa2Hi
fw81zplpXhxCx6lU0+BJ3eGIN1LU1lRUgzSGE4IggZrnCkAR/4xuQq+NeFDso6jh
fh9lvjOkfYq9x0dlKD0Y9a3a0mbLBRxr/1hGEsGaEOsGHpTc0BBdauqGOHsQmBJ4
TTPa3EQ8sPMw8wfWYHsNtk1JBMfnMug3H2WLXIvVOnoGwY69WmQ00vaB1kF7o2qs
f/4MGyp8qwd6I7TGabFt+uBPMdSI0cRghL4iybLQizsBYnL9P/EQS5r/5mEgPxMU
0/+xCob2aoGPjD4j2aWljnXZ8tSx8Dn4i9W5YE3C/YfBIFeGJQNgXryNa+PePYWG
rgbnpmT9Y7sFmWJPU7XlXgcwfAOlYGwX0p4jj0v4Y746IWab00/ya9PgP4Na/+V3
7/0AZh01lEEOgCsomp7adJlktgqcqrRCvvCUDOU6sWFkE/cq3O2ROrDOdqUy5NXT
W5ZUgAS+AncYTmt95EK3WHysmm34NiMKQ+DXKvKCKrHsA8h2dwcdEyzUJLFiN3pb
cZ8TBQMi7dyzt5iEzNWlRBkhFNSZaXOVCMhyQSA4C0VJE7mi4BN0SrpM3NUIippR
DbcQBUQ5fahMBAYEusXou0UJOS+IITs5KJRNRfvFSc614SEMYoqJ9Sw+hkXGV0Lz
Is33givF6Y0eW01QyJiKp71gbEGWpHVdtcX1bvpLqiAkj2LevaXWTmfJBiDFicWL
3n0YuBGHJRd8y9MvAkD/tKz6r5NBfi4p7r8hiKqyK+4Eer5JMzDjP188GHSt9oNL
pgljxxxgTDNQTVCveDwK6/t6Koo9IhxpQOhwpLyvfcKFFijg+xPnS2hWNReSlzvD
WJfFJbKQU9nuoEXLpndMkJ0Nqw29zIt8njx9CZCrG9yE/7Dwa3Dne37paWI5fbFr
r4690M9ysMNGY0xO3hMyhmUTGuPWwQeLr1qbJhT/VwYGKS1XxZVEeB47EMbzOTAu
efx2NLrxmsCJEEOCafVPDNtUa5aON3VE1b3cQnWpJIgP58KSg+uBhEicAFIGEvlh
vnzC+J57auQe9i2PODy8bwT9PXGuKW0oxpcLap7RTz3W/qesjk47DGU8wcECU1TJ
cb5nC1pjnlF++5ToR0gYCisqtuedDxQG4ooy1uovWvjWSifyRaQlzWmHdZxaq3eW
Gk8GQZIUG9O5y6EuzbxCW5xLGOLJk1Iim05KSyzgAiTlAZQXLQIVzE7ovdIrFbLu
4dnmCo3ysBPjl8nuZymtDAOs3DxS3khXVVHXuaxdtI1KgioC4CZbXOS8GJnOUs0Y
vUPsiFTBwtBj/XY8rmVdq2KwCp3V872QC4NAc8qfGvoXGGXHoRIEMB1LfO947ziF
/QaFJyA0I4Nko9Dk1kr6sdk1Tv8wN5KoDH+IqJkEQAla98JNrM+wHSIUO7zwYl5I
l+Q2glQY4OzthFXVy9ZQ4PJ6GLI6UvEOGOsg537RqfimtaCWFk2f6qLmxSPwf+GE
Cm4eshrBtQJB1Vy+AWkOP+5gN37hkqbk7AT1Ucnd5kLkzwXLcosWz9Zu0xn6LrC3
CA1T2VEk1JfbE2+8aNRE5h8kUIovfqaNkwqG91UiP+PBKYkY+1TKBr95YEKsX3MK
6eewbmz3edZ4WLtv7uYLw3O/1g5vLKuCZrU+XHiWPC+xMXC9UYDndMk/CpUVyYb3
CsPNEXO69zlVmXLMAYTKxyJt/FtOzn7WBL0evzzIIe8yRqnhF+qlAe5I9mxvdGPl
j/pT+WKPM36whTkX3rKENNc9xftBUle4E71aqMcImIwoKHT3ck0iZR4JcsDHPQHA
h9CwUTxA79TfDwOZm3K7N0R2NcXUvkC/ji4RDvO/NfUOijbyvYqkLGf1ob4OGjai
oEnMORnwsX+misBkHYeK1TArhSX1LOZAfAqid8f7D5f+L7hct2g+oqScM8pBl2r/
NR7M1bb/jgGHWm6RHFeACIeDoo1GIEknEjig19F7FUgWW46J+BOqvd5iNkE4kctZ
rbjtR7CV3nVjAFcn29CUzKzxXt/dWMHmSJxSoTTxK/Cxgsyc652znBqjHOvF2h+i
SYcMoiadOe8yLRUx22p3roOHk5nwKyH97bXJua8/2QpwBQ7be5i4qSVaFkrMpbOl
BrvEWz3G5U6j1FJ9z3GCnP8oGwimlfn6iDx54Y0URFBFRWa1WC+umG+pKY1cQ0SR
2fRkDiysJKqQj9xLu6Vc84gd1aQJEBtslFJ7pXXmAQnlBoXl0seK/G9/nidaUIOL
XphbM1e13PIi/I1ySJo9BDNZvv52Xrnmh278J0RhfeutePLZxKJ4yl5TKjL0P/P6
3QzrffL1Wxeyy8HaJGbqBDau5FkmZjAUnG4TYdvZTuVFGUefVn9I1UYxSTGbxWd5
08UVuKu4Lpu9nzFvvNTVm6g+B7luOxGXnszs2jYzceP/g/+QE02+XtmpaMyi358Z
PquGHYLBqfJHDTuu/Bt6sTOMwskzkj62PjXXKpDPWolNeBP+ZMu65yrZoYorzuxB
sLfHJERc4x3L6+bbCfxxzf91MY2SEZpJgwkRBLEVEIB5SHbCRMxVWyUUsTkiabi3
13CHJEir7vgp5Vy6Lz1IyMVsB2Ij4uzUuo5sIdD6baUZZoRviaAtuxYuHVBLdufl
4xnkzSUzK+MrNjsWcutYQ+tHWWnMO3cuPLVYz8T7/flxAEuAeA76rqunZKNgnjtG
bMTF47XUScCQCswVuxXvwkIxV7DOLpPUv4Wh3Job0YpXdvpWk0u6WK0+AIYILBlg
xUyHGjdJfcimrsyH65izKiu6RmyzkmiOPQKv5OT3L0Xu6hwU6ZGvO8to7tkLCaQS
l1ySVaD0bmcYVomuOlC6RynE5Ginrf9CCuhb5GiM7uP1qinbEGXZtNx72uo51vxO
zte2ZkGotcCoLFHqLkIggDc4srpN3CD9ixdKXS450AID67lO3NAoEdwJuaM4Svk5
EbeeWAx5O5c/IFcKLoeS78StzLRtn3BS+tuN115uvSCHRs8ahX8Sk67DQFlIyWUU
0KI+0QUVpPuAyIvc5WMA90HFAaeGFOv0TyhUoe7M14/uwbwbA6YjDbcvmY13sOJI
XJss1IBaXheLfdv74dLg0yZCUtB7RAbPAklke1bB+1fIBx8mnBXBs8qfMUB5UEiL
aRFtgpuA129RX7v6rvZgWc4ULN7s6aeiMpEjrXwlQi4yt8DJQzhERdaf3nQcihId
yPTL0GNh6ysazaUkKCmyLs7syFsgIzdUqHHbxd5g+13KK9dFZ7nx3of9ga3m9Co+
BME9lHb/i+O7Ms4H6kQxoTmnoEwdD8d9VkDusA8I8vVgLJAUjgHnrpM71ljw9CgN
2uSXRO2KvmS0qtjkVv5tqhl8/6GIDUcvd+aGdUQ8JUJOQDCPUsPy7wi3MrpzCqUf
eZFUo78jTl8mVqVYL2RNhbo34FOd6yo0lyxx5y4pBraQ0dCK0iavhy6C65rHnW9P
H+B/9ekNkL3me8i71tFYHdJLzfwHXAffzYVyR9hdD01e787MlzsIOlyxYWMb1/6/
3xhsK0sdfJ0H7ClvfyxLM5cvYBthWc23jNDA0sImRRSUGbGCDhyhl2MFqO2aXXTj
tl9Ktilcyym86yXi6pK952CPqf4MsfjcUmcvYo5Gg4AyukqI2cuzDs7GlSGVRXV5
1FLtxScix8aCWkflwdyxzNTfUl0MGqCjLZ4b1WA/TO8EFcOWOe6ovDyO4rB4+xY7
Qp1eaTBRpZ7i7LobdNYeqaW4c2aJWEvRmoby+la2gbggoryZ0DLhGHyxwlcNiXNY
FYq6vVUTcCHKo7AseAE8OdAFPrMEP/VG8B7FyX2NkWPTvoj2+/nofSaK3ZXPYjL2
AZvL59BPeihFes+zwOYrmK1Vpc5203q7dI0Y5YrZoYpD9b1FO1P49tuTFD3guKhv
s1Oz3h7iXrXeql3Qch03ESO8CTeyjgWWcgzptpQDeFglejwLJNs8Zt5FX+1RlphR
vKSi3BXpjzCMylsOYczIOhmHxuvv9VS+hKonSFNBuwTyZgM0BsMmhqSyzapihdoQ
SLTqCnVCYWW8pQlLVOFMgrfuBOSG62xxI5zfudamIDHKmH7TmfS4Nqb1pscOCFar
RrZu9jolQp3GtqXcV3InTXQQha6mMXx1NJIlEc0p617E0Ro4sdfNmgR6sw1+5LFM
d3c57iHR0RnaL805fD8+g0tfFeKJai0Vwf+AIVjdfe99gHfM72TvFCU11gb1QaNA
m5iJierlMT2y9WjLSY0Kb+5YIn5yB6zfVxDVMF8qvgc99dDkg5JIjs7FVCg/pxyG
K1erZuGlZQWvK/OnHa/ZtwVnFH6ezdGr2+thqJP2MuyyjQDtCzkz7U6nverlJ0nF
o3gqM7evW2s6I/zu1YXR7mmEs4XO8MvsirD2M5k5JQ04xpy4fdRuj8+Zw5mbEuL0
vTjEWPwWA/fAwHsS4DHpyeIOko3Y27UDTeFS2ifNN8d2py8tPNkQzX90KdA+DnQ9
KowQXVn5SrscwcD5+b1Ux2LjdI0cuaBE3nYy/paNGPHNl/J6PlP/qAni11jWohp8
l8dGrdVKFyre80PeB4duSOqukW3kIe19rnDWYpsxPnNERFY5VZbj8x4U9kdiVwx5
l9nOrC+Sd0h3HGhkQk0vNdsK11Ct2OlJACMF5QMIKNxIw9vwbZ62TWkM5E24EpnP
qEgZlKGnphkjPxuazW3kQh++Gjr4wuKfi3z04PfitAEeE6vY+SWoOw4WPCrPPBae
/zcTE06q/oQcEJshqQODH8pCz85Eu00xdFQ3MewnfbeHc7ovHR6m7XIsF96a5lEA
U2vYb7jZxS8qfFxwWHEeoM22LWGO93AqkofHeQxCOQdLwBeeAPlLvib0e/nPSAX+
r/+Lve4fyRASSuiW0LX566+ICFs6R1AL5M3W8bsLWZot5H83SFWOupYPEPtQ0JmH
9sCfSFd7DddK7wvxUTi+jg34In9GIokcwNOR9EteVO2NJhALATxwIyzMKl3gYq7V
+L5AvbS25pkeBWLrUAppisIjK5UWKMGZ11JgCRNkWmOu7wh2lZBpe1q8ZGAlGIhI
Y2aTrT6CxHDS0Jxe7HDo+i5CyzbkhuX/IJOTcjfcOeOrnri9IzO8aDWJGOdqoI4/
1ezXEqwcBbZuMybp1/cgDsOdXWGZEdnej8WXbH5f3nGaX6F/1duROQpA7YoNqScC
YahHksfQ8bCxCpwgNuBBU1QlHaS6UAxsv4D6b4WM+NlgHmDH4H36D4V4tc8F+sSW
ZhhBfAjWkhfvmCZCxow479uBd6ARamjMqvhZhVOqbC1QE5U8/J4j3POz/OvlP2up
64nAwQZOhxr0/MUxG6/JgV3NCJKq8PDHH7YMIg3Ed8leZhFf+gAAJF83T83J97Gg
SiXZLgrxbb/wmYiST3ivV3DAQF0qvRi5x0N2LyYxZlBbJU4z0xiTZUOI5/+q/5Z3
ZA/KbHqDIRlqfpbiBYwbicrR0iWRo3BMY0zIaNL9oAj9tfJPObO8v+HJys1TNahV
zi/0BEq/gkmTlYo+PnXzha3skzBtfMVcbDShQR9b4WFaZM6oOUiuBYn6nKa55GFg
sf9cA5HoxSfb6mXxSBXR7SBh2xNQNp4nl1sbIkavEp2lqcBgg28uQ7QqSZubCU3I
psEUz8xHCV7AJmnmFVGOb/sGTEBx2z9xxImOYXMk89vxM11tW5UWhJALewU446Zp
a2VawhqkrgBSD8F6ooOIKu7XPYmC6e3l7xYAkdZwxvWOkFYhoNKOBw9ZSDob+FY9
Lj2sADwcSKuUqUr4V/prTJPNE40kb7ZCDWjnkHA5IuGNa0XsJ/Tryr292I5UzeH8
vKDyFnNu2UCH5yi6NIHTs8UzwN3f/g1tLbvYCkxxI1izHNgXrTTLRF8m7CLvvWeM
TprSa+5CSlQFgUOB+2QDdVX4wQ6V6e9tla7+J2Tq8qtNOorfWWTU6bK7UEqiooLG
k/U1JwFF0meaaQ1g6E+OqvAoRTW/XOvRcUwYHIOBIQMipZTDFVMVMp8doMZyIDs8
Splso0TamUrJJqZfAMMQESttKty+8abydN6Hv+JaEn2slwFD1WhPtDdC8YmXkkjN
4MHgSF5y3yKrzBz4jUQwj74/Q9GLfo797aYZ1eR11fDlkzH5PUuEr8bAshFqV13y
VtHWiM20t3ilGWzJPgywLG9m1AayR4moTpjwjMDSa8IEd2yG1K1ri3036LjgpNH7
zs0Yjc0pYLyE85Thrn2Y5k8gQffsGdxklFDUk/n/zGk2hf5uYbIUW4i4nmM58ICs
qcBmZkCtlqEyAqRph/bS5fPdWF4CFCozaRu7XMva7LTLRm29H38WZRETqPV9fQZB
aQJO7ji2ebZr43KZ+5nal12Ein8QUwk3F9hoRf0nTksZBmj9gihfVMl1UmH37XhK
zMsQQyaMoXgQ0I1bGvcppKfAZKBFNSylrikmq1nCQwlG2QCbraD2uPnysUJ8b2d3
sRwfByXthKfcBs+ZZWPCRgWuHyI+VmuraEsK2vE+32xXoDq6vlRFzkLtAqf7G0rO
cCVKZIUf6UTHas2U8ThP7FayEsgFCeuUQ4EEVafur4xoE+XOY+deMcIRuovSBR8B
CeNcpuj4WxsrcIQriVxrt8tOub1s4m1V6xIpwD512GfkDKktWpmWOhFKgaA4EqVJ
o70gQH8U2ppNTUJy5mbxY3b4c3BTgMZkl1+293e1N3S3w6iDeOLE8FCYp8ZodnoW
ooJwK+Br7BiKqSREmxd879WNsWRBhKDEWon/+2FKzHAJCo42LjAxtfQ7D+H3S+pv
SqjAPjKMTTWdjY3rsuyCOVPt5FNG+6m7xPP4rHnZVNFz4p0iX/OrEInMn2KlUOdk
OEh9dW00uVaBzQmJiJBIj+Aq+rUgJEgqGU9ZNNSIzwoNy8qOleUdwMfjlAQmWBkQ
sTdCsEeIt3+PPj0oQIEWfGn7IfWnkar4FfypOrE+31jqpE8oeby4ONhnSqmhUizQ
QEeSYQ9xLKCrUkdpeXTny58CGwp3MyEDSaYP8CdVt24DM4ymQAAd4bKu9EGbUEBq
ORWMkCVexHxwtheyjMGhhAxEUjoqxkqXW5g9kxuNXa6Qy/ZlkdwbeexwZquJLJZ0
QaR9Kj+tq0OuFdkMk/dtL6QcZ+U84G6KCJ564lsMOo3pJY28kE4MJhy2MV2ijRZ6
jfWUrqbs2O5UFReLv8jFjNGP0XvZLrnooj7NZDo5JSJI5V5WymYqahOBQ9QCRY2h
b2Q5d18WYJaLAsrv2zcAxD8JlLWo8VhTiEr9ZwBtW3rlsMGQxT/+WFu5eoJ5+j8w
JM3aDrw9rypLyeiFwpCA+3wsxRVY6KLS+W/fpU0FxKOvjIHGUzPgqm4S0i7axiSt
CUSPknFN0cNoDzJ0xitTjFJ1BgOSpwWOoVT9+VpZc7L+6fNEZqDDTkOAWA81F8Xx
JPTMIEEKPPeAsM7kURtB/N/5+KiIMzIipt+rrblUPoKGh7gp0B3BF9LthpSeUjNF
0r1lpynkf6gGIuAJPPPYxvq6LKpqMDyV085Bv6EhS274LBUq9/pRCn6JpxPTDX38
rr4X7ngsxQJYizkZMe+x7UXTq/d2ZDR6P4STJHz+uHNxuj02/451/rJWM8ogxSs2
YrvVlt7ef1rNQmujNMHz8c2fUyj6pcZfK0PRrqxAocXZphBwuTacWW2Dwl/WAFMo
zkJPOKSj/O98uocXgoRZIIJ2v+NE9jDxbyaYzMXbxb7qknc+0U3znkuDeUqcQcxR
LUCiwYUz0BATffh0IejJmgSOphZ8YCe1Z3e2oRx/FnJkJcIlKP4a6plIJ3/2la6Y
7yP6nwNElHLbA/TpmMngfd3BM84dAD0BVMXo6kVzVeqk8RsUU7JA4u3AZRcCh3gT
uBUVLcp+Y3TPTac1CtEFz7Spw74ppo0ldhZlFCdltxBa8wL9OG1LFIYwDz0mhHVu
9sg/iC23XL8Aa5ztElclbk0n8k9mRql/7p1t6iThJo4SJzF6LHHzYI+UUmiVzhQw
6I5NboIwti+aXel6sJESlUgj/C9OV0ZxqC+wkvj/UvDeZKcQRAiYmb94M/In9p5e
Es+kfVo1K/X82WKT3KTAkKpVUjp+N3Quv+aBqACkD3gq9hEqVb2TWmsTSioXzu1J
3Z/zWRsoJyVVNWwGVt2s+DGVVlaPqZIIqcfeSbwhQlwSCxBJqGYZ86n59sdCxgWJ
3V5uP/L1DKhuJNETeEdT5J9ILbMeDcPi88jBUTjVYx9eHn2jLW7GwpkF8bu34Agx
kbfnMm/b7MUi4q1WAl1qrnEscnvpr8HOxcK0ahjYlci3Jtwk8pgT9t+41731Zhgr
Iy25wRo1vT8yHnOTthtXv2OLAHdcunMzrFduuFoBeDeEyVRT7mglQwSqk+8OogJl
yTIH0geq8R211utybe+zSrxZXk2kNqg44B8D8ADfrpEYtpilmaamxW9zRMLFQGFz
74AODdF0WQx14l0zYRv+RJMsdafBuEmrAuMSeeT+bMaUtMZw5sdQxqauRBONaToz
fi2ugUYCk+gS3rLZRiTsXwrpe9ft9q0uDNr9YypB/ku8HYw5Ez4IajkAmSpr1iu7
UW3TI445P+mwXeEH4JqkdPiLwb1qwZvQuK+gJX+WW1gZycHfMjcj0UlOMymMMFpR
w8/d0mIgokrsDk4+dM7dVq0HJ2WEqP8uW1AQtaoB5kHRuXYvGE7kQ8DOs2ClmKKj
17vmSHHcxZDCYlSPgz4lRWgOaUYzL9SydvMxMJ3j3xWR0Dtz/rWMeK9Kbdy4/tZz
V4dw70qPOfTOrHb+/D2wDPB7V0NqnYxpX5SazCiQ58/KZOq80IZ8hGy6bG1nkj0E
/MMvXfVPlAzlSE4xj+qzTB6Xu+QbZSCeqRu6ZIE0Vr0QXv+YekyLVU8npexG6ErJ
UhBys9mDSwidvDfpcOsIDNhXUpfcqQ+o2aawF0bGsX4V0K5C6gDIAiXINjF/dEWq
zpdutl5mO3hFueKGmp3zNtHsya/PQzXUYYMWl4BFtn5GsFchDRnymnb07IejnaMa
JBlBsSA/sFt3rCaWCOEbrkc3/TqAXj8TRX75gmTC8+36rVKLadqTc5EZzuph9z03
M/SNIJ1kvnOX5kUjdQgt1tYoz125VC0iGe5s+OVBmTeK3vjhmTp0nP9+soDZdma1
UVjzqGUG0Ros30qmUk8L0UPFMLK8V3roX1DekBAUUB0Nq1M9NcWUh0rAu0RjTcOF
7YONI4AEqGbEX1/JyUxyUOvXeUt8hORx2LnVVcDr4K4s4vp3e97ugcjQgsIQYKBU
or81JEetxNLDLVqDIy04AdeuwDWnVZlndMEw7kLSt9MqCnZVT4mSHfNXOpuZ3+ec
N9IADIuZ3O7D2Se5IlkULIGb10rAQ2ElN38/IzeHjD0d8aoJt3GyCxN1+0JFvHGP
IYQW2pd0wtMK0UvtOVP8j7jfL+SYt6HFPtXWHlgasipnGCSQovAelXunkYomNz9r
ZCSOJ3/st+S7LQCkQw9TFkY+PvCaWr6luHVRNpS5MKsmlGAzUkR1lb4oFCDwpPlb
SERHFyLpu9kh/p/c9EUCi4uYV+qRkyorYG3eNTuYb9uvuxxmtBQXpq8Vopu3Ricd
1YEpjfFJ99Ndey0dGe5+dFWuT/0pgxtg9huQHDeoVJ4FQ362UVbDNHUSQZcFsOYT
jAPE8JZmlpsuNUvHgWW0atv9etL8PkmMsm+rQArcchgQo9ysk8mLz1d5QuzsVj9H
R3edU2OakRsfQIc+6T3nUGQ4bWMyizGg1ERRt5JxTuSVGW7PxU0ZtAq0N8CUgkLJ
hf7yVGAWEwBGE9DPenFv00w7/4Nsc3Rxt4vSHkr90fCdoCbQ/xrE068+NF6qzbq6
Klqz7gSAwooZT1FklD8a2Gr9jxw1KP6Tp43C6LsdpNkkR6e7TiodENhqnJGHAsLE
9SCacvwITL3eTFgsB6JyH5dTqG58YqX9MF8pbxeyebbzuINLmIa170YRRMcfqC/V
BBqOAUrJnutwyAwCApfFH7vdJkGYQzj7btcHGKjpqEGIXVR6AJpRTj1JJ9CDclx8
w2M8h0MRMA+oUIymOUGQFMpGiVGTu1/C1qC5Sq5UAGfqOGBeuAfp5gLBME/rpoEk
SXgdjpfQWiTyu0h/f+9073MSWLnW0QBYxR/DFJK0+L25sMLNHclqzs6eIk31JIem
3ExCqnMbzsVYDYEnU6TlCCw1UqU35LLjGiuz7Mqc/Hj2JlwRhP71VozMLRfdZnSX
+UTRRZTQwiBMPP4F4n5I7qc4fNhvaPYjZy7QiK60A7wDil4B9+D9aVhEWR3eVx7a
yxlDTVj63GfgpBYPNahcEMULD3Ej4e8t3edU/v7FkAER2heMM5rNIRm8Nw8dq5nA
Qdrr/JQ/IPd2UM0H+qnFt7VJj5HBzYL7vwG1vDBkZn5YUdQYvMtmPERn3uL2PhcP
NAhOnW2QvuiUFkCyDoNThkVOcBifSIUlItb2/8i56lwjDHc9m02oIJIw+Bx6CbFZ
NJrMsCluhbsV1CPYEXtQCn5ws+pv4XiBIg8cSOtsyL3e4RPuBtLHwz7hLe66ab3+
RRklinkx3wQxz59YrBjWGM+9nCj7WcVVpUNfP7LvJZKe766DKNarezJvVjky/zyw
PDarCIfy3Y9kS2CPCG2ar4UH7zrT2A6KveFCkLinq061rAs0Fs4MHKZXH5v8ii+9
4O67rMhjgQuoMtV5K0GlM7APUlJrjIS48OIQSiShrShI17twcPxOz+V1pdt96Ebc
VpY8KzhtBD7D6+mf+voaZahG2QDxORMsVpsOOiO6wl1zQXGRMnQ6qRELuoCbq+pp
WQ/8kxxDmiqb2rHyqbQPPVYjzVZOKyrXrVEk2OO+blPOW4ydh2+6xBhN/xPP1DYO
9xv9vkctqyaxH2TQJt2ALCgfQdznuBwedB4hSNIOY7X5z9Mb2vJuqLyGSuXxMfEF
UqdPn3IqbmDG1/0+HuhYPR2DFBmxPIm00o6Kk9ilJrATLYm1WGnWSUq+akzseE+J
Xwb9PIGv4Ya0QKnxco7X7AmRleM/N0g1n/bCJQh/+EDk388XZxELf5O2HBj2XWjp
BKMy02RHFPLV5yuVsw3Wrx+M0iuUDex+5D76rIlxdLQqw5/ge+/4Ni/qIJq6fy4t
kUGw3GQRMO8GYw9FNpaTa11gv1UxMTOpJIeqoecI6Ff9kfT+FrH1gfyiAr1W3Fsv
cE1r9Dyyz1V33SMtji/CcUBeGBLtw1vzdKQf3G5jOufuIuBWK9ZbGk8BBCVONDb8
XheAujTWAyOI6iuAwaijw4bvZZRZKT+harLDWLOAFofuB7mFYuL9WSc5xdWHPJM0
7SDg7bN5VEGQYNIcVdyecfKJUP5xSQFW3TZbrl2POlgixGcNRwBjv0i7X677HLGd
N5ofD8UoIMLhS+GpGQSWvsbAW5hSpA3Y7tylUbpRAFALSa6Ndi9cZoxPZZYt/62U
KkjeHmIXJwIk+TwEfOzIbykdI/u6+YD9RWoB/h3a9qPstCpY0InyfnQqbPe3rrDS
fWJNHShRQjXbiIJXt3AulWz4aixiTG8AA/0AhmGjJXjzeh0MiGOMPVIh6BRzecDb
RzcHxtV6IfTDwG9MGlGDrK2+Kf8b69XTKlYmbktkizWl1pFlPw9DAeW+XjkIxdtE
SlkpXF4vVITDsX8KNI1BRZa3/EAbjvkHGK1ilWWfkSiMYGxBSTWeYfDv1HwVPm/0
CepBtkT+DNXpFIFrePm9ib3zGkIeKdA3NnhMN4XTRAlI1gXCzzKyAqacFWbqTpgV
skPgHmO40NLkfvsl3gwrfLBFtLhKoEsyrYLcdH9XwOtnF0vw3yy/Y+Fc07RZlfEB
3NvYX6V10b8D9Dp5DAlOlWppb8tuEwGkpno7PiulfjucDMWi4FphFqOm/vSfc0F/
/kgqWWJC3IOVVrflN/ZyDoURoo3TrhEPsFGvFlPWpbBwlKF1dtp28C7I2wZvpAaK
BZNY+HZ6h4FkaKe5OaeYPz/SdupL2CSq2+m9PN8fe7xHSupKiiMoJSXaLmUFBVXz
7kQqwgbsOKWTsqOQcjFFN2o5BzvQRsdZkzbAcgTtaCt97ASZZbPNM/A6DFecWx7N
H1WgGKB4jyLEo2uzi/EYQ+6GTlw0AQ1MOEjFX4N6MolGTtvzR2W04BGk3bnnogik
Jt61gsBF4q4T0ZeSoF440GBpWXbT1bN9BGXzYQKwhXiuOhWek02ewC7RSWUu+4m3
rpO/t3IwAgQoNXfhCrOHBIrNiBAQI7BeHiwS4yiuvj56+YxVj84isVWuVhDipgge
hlRTMJgvARsaHrmsnfFk0OUjahtGKBZsje7JtTqBrbwQNA60jd5Rf46UWt8jEK9C
OGi/Cc8qMvG/j+K1LQ8ZSwg3mAmfTNiLUmd2atVyp+aGXppnf0dFAoHEuq8O8SF8
99zKzZhN00aytEI5IRItML7dBOzNdYPEC07v0N022EJl1lNHw74NHWHe8h4/WUkp
4LmViNJepyhgt/nZPO3evKbds7zw/AxRi6MIYmvo/V8Iof/1VZQqvVTZrQ0zzylm
SOmpVrebTbAX3gG15NjSIPz8b7SwLDvHLoLRsLYyKXAcEPwIWxW/fsRiHVkH9G0R
INFqJLgrApn+AtW9q662INx/Oy9oOGLvbmb8k5XF5QgY0xO9z/4toH4Ya/cVtBi3
z1+/Dk6XWkryfEcw6OOCDa9loZcP6NxvIWeVwwrwbsjURbr3zgMhcFyLD0JA++fj
Fqlutghs637HKhbaSiKtgIsG8EFw5ykp1HiNwbsjwiUhQIsfDD4sz8eosM/5tFBC
qgGK6UJ0oze0vAa+u18tnT6hUM3hv5SoZy+c4bRZEJgQurSMHmDS2f5gMkYHzN/8
6gj2bKoi1UyO9Na2/Ij7OkTWVe7FjBiMM3gaWX64b78Zq/5oJpIi2v0+bRU08d4o
+VRTxuCsAVKLoYlfLIh9EseKcO5TJD1WfHh/HilqOlU5X/bA95YVPqs/geW0E08c
62SGoCR9WxcJ4l0FA/ogVDH6t2e3aTbuW+UhKxWU7D85T2enF4QBgMhjFpyPrpPM
T9TgocEM8uvskNobIBNY3nQ5XBFrOcGi7JoEEbbRMqEVRDGG9yQ+cEfUYUHznbvm
lAz3oFmiLKvB4c3lp9rFwmpldIgsy69h3U5J+ZF/B0crHbQdpsDhsmtN5Q7DE4xZ
CzZ5pECXeRbicKiM+GKHS4DOoSjdkDdbAvSoezuzspAkvRjKSwZy1oYvbvi5GIXE
pFumsHuveobAL1/MZ3k9JJd5FPKYe3PEjtPtqq1id3E2dD3NjHo5r52tEBf2bfyG
PaqM3IGRFbLkIy7g4PTupgh6HC20Qahy4w8Jx7v0YlSvgKNGwmfe4I8kZMoyiit2
ANpMHZNlm6Jxi3KISQf88gCRSh+ZL8uqBUGks7NNkPa1NO/o4Va9mE82OGUwTjnC
urcgzrJkNBi5y7zSyX7ruvsJLOFwbVAb5RsjZgCZz34HUC+Qn0CDf5Sv2Lov/Sn3
CBh0WDpdDJ1G4y90fvAJEN6deDTfTwGlGhdnEtvjqBfYoJ9b4ZFDbygMAzwTeGiw
fvKh58Jf59NPGvtIWopHNs8gH1gAQU50V1NfAneVxYXBnQLeBQ07OuDvD+ZUksLt
KlsubUOS4jILPayVE17JMyV2FHRGrlkeZ6OkETpLGvDzaUl+2Ygu46PMxWRBU5Te
2yMDJH0ozR/qmNtMV8HGPcvgyLsZJlwgNsRIOOiQZSnPbd0Cfr3AzOaSSl2kzFg2
OFSJI1bWEyo12OV4QgholSO8aIcdWJ2unGYNYTmvmSUUgzKTtt269erIiQ7jptFw
HPcFmjmZn22iHWsr3HFc19fm0dLacnGTWRiBawItSg5lXfF3fmBmLlR9/3Mv41KY
+WflzK4Hpm0Fv2ckQqUjGNNXv+X5gpGHWWriFRLpYVoUXzIARQm6ljFc9ZeFg5tf
XGikfLOtE6DPoFsNRSjzkY3rrgylDM73FXSQPkdpj/qhYjs4QhcLxx7Pl7qRVv0d
R0g7SA3ZjIikMH5JeT0fnZ8dw44HHTNPaR4x6ShKTNFeTgDDbox5u21grIua10dD
UD0V0ajOxgbRIae7+Nv3d+wy8XCJ8nqoU/gzvlWpG4QHSKN12oxLwNDClknfq2dF
p42AE6ktZe+kvCmLA+oykiqsC4IK+0QMJMBSsLAbyk4SahWd2NPvR3N4YchlRNUh
v1SCm7wmrRFSA+hN509STopa/B4iN6etBspv749Cgn5LX3G4jjijsqHci1cxtT6o
OcahXVsyrgvqZJCcRdl9LbG7tdVUFWGzSfv443l3PWUpvqCFAD3FJHGcuUPrEpkh
APD00eMUClylwn7l/bscLhdtjWnMXDF9/7PDjacsKk0HjdB4+Bfiq86tXxC4HEm1
+lPu49oy3CyrHCOK0sKNExmNhmwkUGWv6hbwvWox5rkfNYgrVAO4+Kkt1kTvIA7p
3kalGRvFW9o/u0hxhT3YpkwLxYNA7l7LCUg3sKXZJ9/nYT/5LMQgp+BHz2OrQ7sb
Zw/BLvDIVjWztHnnkeXZrJEKOMWnV70IT7uU0Z4DcJIMPE58AMoNaKZ7rR4mnHCd
1Joj+wWgFOBEo/+icEAd9Fn/roR/gA+/lyIPi3K6vdAzv8c8Zt5Zir54W5/ThPTH
HyY3cFmj/bNy0RL1gxZzv0wwLKZE4WmvhDCiVqlHZRpK43brhNOneNUFCqwcEnfO
dHNmRPXwCkYglUoGawF/aSnH66UdgNVQR7sqmwKtluhZjkjvxuKmsDoE9mDf1Ara
UDszz96+xp7kJKych62jUQweS50hm2nLmTazrNOT5666i6q9nagKuYlLRdG3WDQD
pzgs4JQi6yibAQHQuJO51uB2rVoFEzmX6bAdI8BCLGB5oZ1IKoV0a3JKLk7wdRJs
evfpPPS3e0HRtIVMvWl+w0nFha2GymGCbwvB/kzRtjHeW2HMBLlMFZ9/z4/rMcoc
NmUMRLOG6cFyJwabcrV0d5A2eBmJJECZm9ubNIrJpyk49QlXLd67w88kVtRJZj6R
uHbNLxmQY/hvnWTSI5gsZ4DrQ+nBVEmX5xfPouzINtFEB5Q/lvJLQ0OGxUXtxYdQ
FKSTJexektrXgmXQ6XiM+k8KqGOtZmZZXg3sqR5EXqP4c8quplDm4l72+610nG7Z
bVLzNQkcQNMZsYyopd3ImWpcsIhHDlGY5hx575CxwJ08zEUVuqv++ZdrtIxRnQKN
50Va5VVgR4G1M1/ts4e3V5pkoIdej/HobYHdMf4QxlsjLvBOJsbzZyytNa5Gwt6p
bQAGh0SCGpCdSADQL4kDPW7iQOQDrZLLjFa616Lg3sXZxsxImTp3hXZMVBSKVQGx
v+9g/tF4VcfH3S6xbiRkBl5hAHP4s9oClSE8xwOls/81ibeodo9AfPd2PA326XBe
TTpL5S2Wid/kk8ZfT5vQo0c7XTaDHjmpZjVDQ3Rt/cSUFC5T1eMJ8uUGS8yv0Z7P
H1IFGaKVcyFYGe+2v94gdXmzSHpX3VJ3tGoL21/o6WHEHkiFZpfAJs739i723fx3
elLvySdmVvlxM+kMOhgIsYIszGnqJFsBGx1t/FMqzHZ2hU3P+L0M06nfVlg9HXyj
Vy89DG6fC+cwtsBGHmHfhEYmHophVHXNKzquWIrPaxkhTAUHILhZtG1bu5/qyxit
1MRkWMaV/xwOSkNCUBL177I8S8pILD8DVuZpuIS87lAjP390h1gLdTxxM5TbAIxi
Tw/AouNCAPQ0QOMRwfyBEunKifAJf9W68X1278Z+gChv3d2QerXhJuDxqTROILD1
zqRgdSaJJpEasUUxcOavp3t+nppUjNpGXh4CySfrBMuNvdPDksAJyshDQkyswFQr
3wXbxDXenrZVFuoWBjKaNxoQUQI+mwtn4ku2Cm/qGv1avN0TyEEhZMRN8HMmriaN
EMi40AJ2VZKNYDpTgSdxcn29YDqP+2RprrOp92iBxe66T4tUzJWNs1YBW76K7kQt
itTBNFkdWZh4sGdlcOMUyZ+47MFX/vrF52vLU4Lj+AB4cHiFpmdb3lHSKWaXleo6
ZWj9zO9u/Op+myvYZmH2jNQdRm0jRbvNrtwTu8+bAzGI0RKK5tCVlnbvpOTKWawt
zxsb0tNzfsdazV7j4lTSpP5XnBX6deIGQ5vEwtk3INECbvZU5e+uFKZgFu8hbwjP
ylcy45LnpsTcLmd3ths0x54Sh7Wa3Kp5Q0tolHWqhfKzp2dlhhWyf1Na2kH7GTqc
5K1umbiMp/cGz/Jnx2ZjUVeWACbA57DN6C+W/0iU6Q060MdSXgBTx3lgzTQM3Ysh
57m95hqjiY9z293gtmuHH8NY1d4qksuFF1Lkwjogn/Z1J2Rn5tzd5orgTIVNytyQ
PCriaK/I6mUBhHCaUQvcL6Xgzp/x7TyxSaw9lzim9j7MaSzG+oxUQH+0DasXA/+G
x+tnh9yb57UUKfi//jwiMvmuVitLtSm4KEy2s3cgsiCtXZ5Pf9MxkcLIVTSKUD9t
KMyyqbTTKjV2lCBZ8Klw70BgDLYiwDnOkDOVpRndjnOK0WZ2+nb4Qzt6ZTS8VIBJ
mpx8jFToeKtC4svkXJ6VrtnUQME3FJe8yjDGUt1b83mNGSbzLDDODx29bGlgSKJ8
0QUCSMKiu5Oj04hZIKhhnU+GXpr16m64n/t16Pe5y+DmEno1ctlHAtARAQkpGsjF
9cK2qk5gvaTeHa5h7IBtvdNVpMLoC6ZTQnPXiGYj3LjH48cVFodf7AlpvZGifZWX
3kYrQLTyzT68VtJfBHQDqqf8Hm+GnZkFRv5Diz6tdYtJR5jLPe8tSB7/xdd0DuCV
w+hPN6E4erfYMYrcziaOtj8+ReglF/wDphfodPieCfY5CxdbGyhHQGX8e9+uIxNB
TUOG9Fq6v6CGgM+V2fl1SzVFWuDDVwxmMhjCZpRQfYNwL/Yzyjcssq1i6liHfQIZ
DgoWN7GLlHXkqWjJR9atdqo1AfCEFghrD7ssafc0jF/Ais8W8MoH0KXqC/GDLkK2
hFR21Suq0YuXqo2MdQuMU/mqgtB75l584dtJD7oJa1MINNTtIFQvvAXuRlnzzBE/
WIsjyM3psd309yL09f4ib+9CixD2QWprpE4rkkf9ohH0+kwErpURhYZELQWFHa7o
ugQg5YACnW92hL3p+TFVlh9zMMeL/IduslsHPaMB1+Mmfs2xHknAxRImJemDxJS8
tUNoNugNg0p5kZtKpWo6h18gX6vU0phqI1/kGg2xS4WlzfbyLz0Rs2Ojqe+atvIO
JGvdFGWoOqoRXSxvYFxD/hetq3oTAvj/THLpq7sBzkEdG8mhNEVlYFAriuCT0gb2
P0ik4dC8Hszxu2/9aUVKMwUWA4ooZ/9UOpEse9/Bm7ScvczRjqch2qINTdQibpce
GoDOIeJ2ydSVRK8tbupB170qG0xb405c2cep3iH6lQICNt/xhpkqhRkDB6ZVzJKQ
1OaaVZYOEB6LXSt18jkGYLu3gnZHPmKKO70upqdihYRj8Mf1Ajnnf/mI27QYUm9v
rN3MA7VP7dzpYbLZPamJ6aqvJsDtMope2rN0rlJ4GEUT1wJPlUIg4gOdZfibFuV2
B/YyCHvT7uE5fEslxsJqgVQXCSptLBG03i6+1SBnSyFUPrQp8EzUkIfTcwTNuHp+
8nqtyHY2/JiRChTj+R6iRAeMu+zXhPuFqco2BfKknVq/2YlzSDpgIC6yyFLYUh3z
naXUsqy2h2XPpB2Tav6U7PM/6uqIuDUT7f5dJDU7KAXYCuyqwV2o3ZUXjz7OlWn7
tRq8T+t5iZX2agJWpAWJAtUmdk3hv8uoSynyC1iCbZUCDAzCiutF6LM2oUXRlT7n
bSmYJJXL3rFPj9ZGQnNMpeQYKfx8Xiw+WCKm16NHadzKje333dJp5jHwZbaVR/hZ
ps29FxD5Emqp+44I7y3+Ot0/j20ExziEtB5HCKRsR9QR47UtueU79dt8PxO/ZWk4
0/euKwm8X3rMZDgPPiXUqmMQ2xE6N5NeSwNYY529GWQ+B2TtAiGBpZlPZnF01Ifw
DOld5lXumdbVuoWvaCVItOuLwIkCXFp4gzxQ0GTWkumQKJWwVrQDndAIf4gL23yk
76IHjm7GaK/Ik6sVXlnSyp7ZMZCP/l2zxUcvGMRtqoNNtr25ioFqzYa6DVElNiPF
kG4Hrv34/qQ87JiNlKN68X5dJGg72+CdY+GHU+q/5Vs2QCMZjaQwCHq+2LJyhrNc
aptU+MCr1gmHBnVrxvKLx1jnz2KOy+4glCVxJ1iWW37GKJt0MS2R69s6pPFS02Xv
7qTKWjGVT/YzTx5wu4NpkI0YOTz+ivPRt/ATMLPWzAdIDqnEsQMmDQYxbMZi98gn
hMbGF6OXaas291Dlvlcx1+11BggByD6JQTFQQ7VpUTCl1NuH7Hu+NwO6W0umqfZW
GR90NXOsK0bP9aCIlSNEalAIVCXiMqkDBokWIm8tMhGLXtzgWejIaRWIeVL928sF
G/uWrD31GoKdn5A0sfl+w/cgmyt95nHZ9irzj08CN5iU9Kctf+RgxbYMjxAs6lkA
O0cybQClZn95/XeP9vBHaDxvNLS8U1sWcxdsubQ2tAijilC/Jdjmkm82ehqSqdZu
f5blEJtiHIphlKvGi1wlajDl+gnMewmpuuo/QXDAQd7GHOhJR5nW5cTlwkgzoK7w
QkWwE1/5D+KffdU71EJ+dxwQWCoX8a2hI8AcjtgzaL3RzTkGz/2zknHTm4lfUXMr
Ht/szj6NLLNdWn6UEmbkv02K+9RuT2SWds/V4SCA4xF+wgedfFEl6YWkp3r0+rBm
GSScS8uF6BY+fzMrgdDZHX7935oxA3H5fhkYkkaEoEMF2DgEdAMjRXjV/sN9Aeof
W+mJkL64pwKBiLw3e1yygLcszKNhU3UKHU6DI9rbsFSXlW+4pRyEicKwM9NN4QWd
BpQF9+BINWpD2ekpMXn1Oc+BamDHwCKa4oLF1UexWSgBE8WuTUqUnJfuO4prMQ6b
sLWCkWezHrEHTyCeYHAvR5Q7eMA4i/T14rJgU9nfAmZa7H0rJoc0OTc+kKsEIbPk
RStL95WcQBo2B0OE4HO460cUJMItQVc6c/yKzZrjlaXqBunXWzooB/l/+bwo1gmZ
dO6Zo+ZZ/TXt6pfpGGDN+bo4KA2ZL9GiIIJNkk+vl0hEBfycYVHfn8tSdJzsDoR1
oZSzzxN1xctuc24aSKQuOFCn4pC6MfQAPx/UZC2tpBHs7cHTKkI/QCoa9iwy2ioZ
e1RRoJMPDw6adSA07wlWbEVaOMuArKILu/C8CYRDJKfGwTfBIbBJDi2GiCWRYKqV
ByCA6cTaGZd3JYs634ggR+2yi2vBB0BCXo01PvEf1rCs6zKg7BlRnKktxguzDrFE
f6TQVptldsVobGhLA9QUTyXD7yuqgow3F+VePcwJDQ7mw9khpm5oOF0MnaT/6cEA
HVAv7mjNDNBVxY+Svo1tHqgRyyX2eO6m7dP5JM2nuRdqF7yD5aTe7UK13BX5QyQ1
oTF/AUNsBLc+mAw3a0rKk7a7XTMJiDP8ROF9DkorTTniLJ2UP28Mtvub4QgsRUOM
sJf+NnEYTPurmMCOHwqpmu9cG5vJrSKywOVGCQELxa3bdxRURBsLwgriXer0JlqK
HOurnbKNbnLwnBiHCOoFHKW/fb5dHkaxjdTfIcs2YnSboR+/AkXhjPv0fsGrKkKC
ZwQ18W8buH/7CKSQ9xVI/xJl5/tTKOttiZ5/ZUYGIlt5orI+N7gswz3alLvcPjJ4
a2M+VF19QGRxv/nFplt8WTPbHOvW4XI5nCLtMc+W5gIQrQ99sA6+vyN3AGpdbYWv
fpWWpB/AHTFUppXhmaqhj/I6FP55/bOKzufk1dVLKSY7h3vDHnfw1mVqOQ+LevhU
1GEqOXBcItO9mo/PLwbVX0c+qmuAiRpYkE7SgfcksmaqOyikl7B/ClvFeniMdUSS
H0epljdDF//DMm4qte/sNldmvMamAf5zI4COr78086CJYtfDO8wdyYn0lpx+PQGe
dNdV0dH3hjhgWL6xl4tNrVmsAMlKtUhgdlGYQ+UPar4fpyH/QGy6fW/m+ANiTszo
7pFBVk0W5uqB351ENaY3qESFqI5MWDXIn1p7KDM/QQk4LE1nd/H3vVDioJwIrKUM
ThISwPQW/fCy4eo4M5FzAG7t6zyP7l4A0GGPBKbsaHQHxpqQp/PMC5M9W6pzEh1o
EfEN+WMqN5BZ6H4U9Bd+jzLUau4lO4aSgMtF846+JMEdFRcltcwQa5eHYQ5NrJ/x
8uLduMjP4VF/mCaEOyCmb1dJjea5krhb/GSaAqYOya+jQVk4VwOIeGc5t7OYdvpU
sLxLY9/CtvveFaqVR5IzJNbszXeXAQ9Am9V7si0ivbbOCj0PN/SVm+FbbZ7ngUec
mesYESlTsHKx3GPHpYdmpN3XGmIxDFv4U5iE33QcSvkp8K9l2SA7RFPx4//8XKKm
0AqH7knbK0kMtr9R94QSJ0s9uGz1u9rAayQGTK43YeHYwOsUPv7rscPP1YrwB3WD
eF1KER8+VNzskCmdffXkLii4BiJRr9W0A9W7I6dnEfXp3U3CUU0aoUOCZRiNcFXW
F/XmKkJrv6GXStWIcZgMYQZ/Mf36Pz7dowpdzGfFVwcgq8szFXvBtjVMc47JWJWF
zMrraAbtxl/lok/mM0McbpUw5VZImXZ0eRyEB/f7d/JHmNRlujUt7GdrwWJbJgjc
IIZFF9KS6+YMgEA8L5ORCef4bUIGlivB5z3p61npBb2flyvastR+SUH3rBwDGu5B
xK4T1nIVRJrY1glmALloxMIWHmuvVDy2J9qaCXf73PXKCSGeNy3gZHUKE/bgEZhI
O10vIZhmmdB8YQy4qTgKSynS4EvEgyPzfc+i2eva/JJNMwIzKdJqcwvGxw1AaLmG
LuPeX5JshQKg5vguozWoblcUWgCHOi3EjSSsAEWIaHnPHOIoD3CSi8TNYotmJ34z
SFdpWYl7jpa5AvCwtm/lOF3fhlaU8n90UZ23l4Fyqi2xLizJWTQJYMGyD4lhl7Dk
LAHVd6bPuNsWn6pYNR7jdnexsFV9We3NuTkH+Ym2CLlf3VJrpxV8xg+dqocXK1s4
YaASNFwRjRpvXMSFQpUJ4kQel0ZBQwr/JHdPCWCgsJ62syU+cPmnJyWJ3wDsUzo1
sJZ2zZYLReo3lMF4CdNtFtYd5NQyqj/NeWrtvV70W0+zjg48pkHUgpgxhN6qxRD9
4tqYUmevFIGei2/BYSJONUdALZk2+T3dYIXJMbgoqZB2llWrIsQD/ebjQm4HcGEY
wpogL8xdljDrDWxvuVbmsMfnPqwc0qaHVpm2mNkdUmKPOd6YCLcDWbqT6Brqey4i
LWyEYJWOtbjclnRHvJwvIz3fntNZZAF9Vwad/otcMFA5OZU2tmtmCuGMdeKKFi0w
FjF6vzaA/C61V3cy4F5vRTupxbmBjOJVCkFMR8WH4IjtKqQJb5r2mpFpaVKwnxBt
VyUw2QeGmPm1anAzwWRgZjbPM9O6brdWxNLNG9iN0aNq4pBxGtnI1D9ALvkcnt8s
aBCewTXUT5AiP1e7+nm3jnqs+5oMsx/YnXa+/sLhttjG2xzBi+y8tEP79/hB3R7J
Vunuqg91psUQaN7WisdU16LT/xPM1WcN71v5UV08ajQhkXUrgBQyEMWmSdJhxFVK
3YeFgdK0Ke+lPN5L9wpNwz3ni+vsb4OJXtakBDZrdeIPRjTuMAkq1rRV5ok/KpBx
2dnF/YNl7ypI4z5bsCDyoRD5wtWcNABDJhrpoKF1thwkIJCkndOSSzvUISs+gHXT
ZJ+JWWkcUAyuuOvKuG7HUR/cgiWxjSis1fphycFOiXfsOEi4GK+r7vSbn8gHHunp
a7+YtSLMmKfsEgtBVDIismxQk+JaFcfIgklNgilvBffF1Gfu7zCqGK9G92sdoyqp
KRgOYgDD4DMyj7vjn7KXSRl3XOMhPMvOuo/PPbw0Og4KZocjYwCeVbO+fsnyRu/7
75zQ7KJhXNAzz+o0jUKOgsLk4ATcDq0njY1c+8oJOwLL9/x3fpMZpUVO59EGO+2i
jQEm2AOYzkhCh1SUsoSctTitdYycrjm1yOA9VOTXK+Dt7Mly9oLD0bf6j3nTn1IT
kNkZdN1YWGx52CmnlZ0V2dVRF9F+meGUpdZZELTDra/clmcofv8RcZF5FBsBSgzG
OudNm/yndbO11YamhbdAgFq7xEbvNJqdcQrMu6F1XLtEjYr2MWrb8AAexSWku4Hs
UtUVIRf0Cu3BM6JNjaH4zmfDA81ASulWRB0U/vNbBZEmtzx6szUrrgan7ShPZlTO
LlXfvOK+VjfW6G0IHCRfOsVkv4zPLdh0dB4UeUHbAbUbWJTmHpDEg/T6hUmdADkG
eBn1sA9IVgtM+4imgMF+KZ+4Zq0C4uQkClHEY70rqB5pUUyRFTEkDjm2XfmyC+dE
Db0j18K8/gg5qH96UnKzgdTFHS9GOmF0G61IS3XRDiPp+AZ0NPTyEi+u5Af7GRVE
Hh2KeKNrtTqibOST0rLmu1Yc9wXtAKRT7Awjz2JH6tq+QTGmkSLQM3uEp+DrCbAr
AqtSVbXPKhbWTZa4rIG9SLZK2Cq1zE1xzwRg0vOvfRbcf/dfoXK1vlEHg7S/Mo/Z
RfGpH9D0Y4/lE/QQaazYjFVJ5WfODdomiWT2ZHG5f+FvxmBcn1h2njtRPcBGGbdn
Q22b4Y/O8SxM7QzZdADg5hPgav884Ch5EFrbMPscG+axB9GE5HADg0EMVykyK5JU
7v1/+NbdWTlVgikRFJWTAfeXicvcC+DNklpZLj8IEGQeJXcX+ZX9RRzOsAe+m78t
hVxDK24UNkS70fmxQ127cNXj/04Yi5y80XmDBE1JctyL8E7AJjm+4VQehLfU1Jm6
KScvTh1MQCZJuMNJGhdji8bNEqVyBQ1IJK4c3o2/jdsA7I7FC4ok7cCpW1VUh5/y
e3NClfbYQDxuTxveMjM3na4rmiOvfextdl3uNOrXRUwl6+G8VNC6+QXVkcKwf7y6
gY5ggSc9lKrUpAlfWhfc6WiBl2UU+eiTT1D2/CQUNXlVh2SjqJt1wfyoe9HDU007
6ArTqgbODSm/5Cn/NgQI0RR2Y1P4wqp/N3z1VxgJzpKttc9ZKgwx8WyEAdhQPuQI
ibDh9+I9d4QuBYdk01TUzP3PqZPU36rLVwmoQ4izbAFHcxR2ZYZorLW/sg84Zdio
+fk5Z2SO50A+aCdQO1QcKvEWpvFbOzf8BNTu+TQNcpFREHVSb0Mxr2lICsti6YB6
Jo1v5YbIEO0/rvmCGshN4IT4+46WOLO8lPSyPhSBEF5r3UtHXeUamdYE8cCcfgaR
G0Grp9ujzhIlXWIvTIe7+ZdeTvfFZOYRuNj4/kikx3Ks6nPBj4Ron9Apt0sn7CtT
tNJya95O1CXbtxuhrjeNpSCZDtDt5CquqE1niZSSZMAgAIpgYumYBic4/me+bUJb
f020pvRQoUDyEHL0YPidOTyfRtKMzJeoNCrHLIGNakR+Ii2ez6NR5QzK3OOlD/rI
TJMyEbQ7MiIo21WMkWWAzsfu3cTKT9Y0IB0bCXIyFKd0XpC2LCeY7Kt/1d2pm5rr
3M9AsLpJYmdhqYhD1AxzSl8X6TDIY6s1LlIDyVEY/a28qeU49Q5twzKXzT2ijtIq
IvDI6V60cmQm/O0AK+rwjpHtC7Ibc6tyDgWuTH0XKKcZkWCfHaQALh7V1mo3rdoO
fwTFGOvzBMZngeqTlYpTDv/5fGMqPQBhY4QIQZNVWzE1zGytCTlW/nArz4ue6GYs
fJvERdvv/refGKXdqGUzYC7is6zy4QsAxdKdSUvNprCxQcx4OgPBfPMvPAKN6+3+
cttURNrxeDzYI6kW9Z9204hoD654tnpFsrnr/zxDMQ9xSufPW/MiqrgtUPQUVNX8
ejUJMPU/utBNBg1qZnShCf44dwqXEBRrocLEh9RzLoFqvb6M2510zzqhUNI5NH17
RyI7yZnwJp7PN8R4VxK0L8kBmLl2SjTYc+9uGgfliPUkS4pOUaqYuI99tTgEw/n1
/tn/7T44/me/AhzlmQ6ggswE1KX84sIOY475U+oeArAofTybFyishfEN9NSWWTMq
9i9kKhcuU7CwpZR72P9k0+UlsQnRKZnF7/RDF1m0BeQkpcJPMWta8xvClgW2u8jy
1ZbXDIU5Ci0Br3kK2A/kB2ii2oksoFaYadOTGoykthEWpKL6ZxDetZaDIvM6i9uz
fGYlRii/S6S0mIQFbfQQBSMFzBHby2qozCV/rTH7NFLOU+Rv8fc6toHpDPsst9Cm
OJ+PsZBMjAWgPN+87pH+omehlynKzbPg0HfiSsmIneLUf06tS1PTCRoidTc3ErsW
FDG45m5v5yp2sfIOkN/RPCCUrLDM/PDb/4r80r455JNaNEIyqz3O3YM719d9lqy4
lt0+jv5j3XpIALeDO4Hy1cEcfiLqISMKNAxkjVTwcP9kAnNDqPbSd33xdjsR7moo
nKyS1m8HneiA8M3aQCdIdaiGJh7EupzAxmEyx/1U+mpb4DO14DfKWzfeNPti5WhH
P1UyOtRLSTAtDWZwS8mSRapWX/HKaLa4z6Ufw53O+pGETSYQgbNU66AxhtJ+lb4a
g2k4Auc62ahxKA9mTu2szh1w1UV04dHuSgGzTMWclA3JGKk+qqn59A58ryjVSwJ3
NZu0fXhVlI073j23gyL/J2s8eakBEzCRlfoefwzIER3gt5n23svCWHznra+EHmpT
Uq1yjAYG8gJoVU8UsKH9ClE/MfySk73COvhoGJKpk6YBuKBvepePJeTsIZkYHcoJ
uSTtgToglnV289KnKzk4JVJ1Yl6g0/JKaNGma5077IVmabcEkuZt1HLzuvAuGouN
XKT1c8F2dSf4eYXtRv0oRhMr4B0VlAo2BeVNR0gk5IGg5+Pq1BPM4nZqUWC/Otau
eRC8pbooYAIxNKnpio1VGqkkiLcecPoVj/P0jSwp3wCzc/DVnFJHu6n8jz1aL4HR
Cw1eGk/YnC9YOE8julah7CHuLvQAGLpqE9o6/iWxlPgds7sMr3MowlP//5XlUED/
dgZ9BFcCfqBNUv4DBzMgDYuQwjH1S3U/23laDRVhcO1JgQ0WTaH7V7dnF7yl8aMg
i4laYwWmDqrkDWA3EOZ+zXRTbQnEFLM1M8KmMkaOLxVo8SSbO1tAY9Ndif0Jge+4
QqDgdkOW2SYAQr+qveKSnocbrPWMJhGUiNfRtQzsaf3ykl0xsy6vwSc/GP1yTabt
6k7mWXhbk+KHppL33/NL6mgdiQaOhLc5CD/8l8wRlCvykqdDdKxFVvIYEjN+PLaG
+EEcVpBkCyLwwQy3ilTUzo++JI7giLQ0x0kAMmD/MfrkgZavRxWGXzoOMR975jn6
snghgZyYttMiqOV2ZTCExVLiYIkH6AaXR9L9DQk0C/YB45PyexF+FoJBNDlpkfpt
BHwkXW1SU9zzLYA0qR3W0l8NnAHYfOfzAPm6v2aDhozp2R1eua4bBKf5bGgBvH0s
WmcvHMhVo28EK3C+97agaZabJNXWwatCzcuJN7NGJMRnVIfb4ONCeVTgf6NUAR23
hcs1NSvqkS5PQYVRO+UnpWqdoSB5P5ocE9syve9jHLH89+mtGA5/bUAO28qUabI/
bszhB5PVzTDQlX5JgVas5aMOMCqMWyXgDRzdThishE6Yo3zJJEa2syQkwTqCK3ko
AiA+IzMV7jTV18Ft3wf+zI7nlmjmbplnCgdRNm3JGFfO/5MF03XUHuKWWX5lLw7I
xe9xRsYpI4Sqz/pd2rKlhyoLRkoCqmBhtlqq4hcDgbgGvf48QrhGPt8gmNyhnUaL
IPvNstzyrTQ+3pJW1rxftmGbWu0at/QV46XrSXYxLecd/9/zkyPAoShElycEGo0F
93zT0TfmI4A0Hb4Nzd2i/DMg5otHoLXSK9l6FVmA2/kYA7t2nPwxMCvZ78JKHBou
DWZqTPhc050hNmqV+K6pW416BsY/RyVw6BPWBosUiFs3vjvtgIhD4UkZDyrVsShW
XPjPLHAi/VENCnfsYXXfqA8wORC1HXtGMnKO3fnnvVbaQe9o0arH+Au3+88N/gvA
my6Ejo9naPdPumLPzXOQ+Pwj9e0aS3+vJTByWTHmybelCpcC+aSS9Y8+/xJyj7eK
dRxRa/7U0YBb4hS7mukfzF45n3QhqZ978YELqDMDRy8xe9SYvDkyvW48QIyN2yc5
4SWX76IDEcSCnNBtvHcGQZwBAAdMKozmcx8v+yTKpV0OL43rzPG9rpulnyP6Ts9c
531pQ2sw9CzTxCOBskvUHi9I5BANDz5iA5yh8ZX+uGfiOPcjoM6nK5FR1OyO4G4+
uN+nGlTB44LQw5iiP4SN38GlMYTs/Gu5K0WbYIctIwvwQWXJRXnTvxHj0ejNoBux
jWH3+IOv2wTvsLXZOM8JuvAKbTzlhAiNFNeTbvw7upSEIzpYptwbWJN2zDw/NBYv
aS8McS1NoUjxzZFk+ZLkIChOhyiCwV7iBtOCZceJnND6jZbCNhe7UHgdRboSy87C
QnxRFsffNJZuGRaiQRZ6Ez16RsofU+vTwXEXjW33oXk7nsqJDeGvl6J/XMyLdJ49
gtJF2cLgXGKPjVIgrV8iLU7IpVnH2D8IfuQQ61knHFWT4uE0PqHEZY0VC1UbyUHr
qcQW05Dx0gypd46pa4sHAwK8iDKBCjPz8MZSU3U+UA9AsoRFnpbp/SD67i4EfuaG
GG0iB8XJJxCOgsN1zEzVZpGtp0YYeDeUufkYKbDxju+KWcQZrbFNOcYs+xV4llZO
rzdOOK2WTJySpY8K4vrhW+JSXwEHU+fmqr+vnH8BEfFFhlWTNagGlt9TYN7PLtWQ
AcPc6jOU+gZH3vnuxG9dZc5ssbJHw2GxJb6btFgYegE1uXOUUaBCFH5Om0ACfpoy
Sjo8vr7bWz+KDFRFnVxA1PdCCVKtZaH/Emn/bYA7tENB96heWD+tRoiPuFP7qp8H
ixlNFpCJ3RwRtItxCi79XiEwQVtb7yf0wq8houC+SmJCOvXh90abm5JPVvAVKIhr
S4PPz1gpJqheQv3rPCjdeMkWBL5hi3tZS9xOaW+HVGzFgoYBaXjIZ9FRjNdcEMvd
xRb9LO0QhxFgWAaNQ+dABt4Me9eAFMvUMdPeUG/Sq0V0HMPd6b7s0DQWED4lQmWn
j8OmpoAK3leu5CRs1t4VBHRVG2ProgFZJMhCO2+hAj/E0c9id44HvuSkQgpTZkJQ
o75f7Ane9K1nsSTGfH7zpgxDTOKSbw4Zaat9oAbAHnkJMtAtlwHzSFrDQhugcbeR
yvJbKbJvRH7z+lpmWMwMtLxeO8ZG1dndoWS+4TIzbiRTWZopteNroS+qeA1EoY8C
oBA/8gHTwXPpThAwUpwvFh/O+syUHM/cYa1U1uZY5YMQYLyInwvsPwMC3wuAhPXz
bEpW1B95Aul3gxCsnVq1Xl7sTpCiKLLix5QnPpCIh74eSXAlfn/O+FPNN7quciva
MBcuPljQlmImqmy3kWqDHN/uh5kzklnPAgRYvUaMXUXNv+rHfUY3evPG3DB0UzRV
o/kXFt1WeyzxgSeRw2s6fVHyi+bpHJ6rvpG28lIdlaJI9ArnWCYTmyPrZynahF+U
A5ZEYMG700/b57CeQNKVthZ8P2M5U2fgbl4ha/xY62HRKcE3ncztA00Kr46McSbf
a31A+NoGecPE07mxzVnzr2RqF5fOsOr7IVRPfjN+FvcX+Z4ZLTp/Wfwctm1tPtZe
2h0wKFFdFVX4rRyHHGoALRQTAGQtZsbC/aJuSKP+2dJGJGj7Du8bRpTGlabUSRcR
nrXSSF+6lGnHrgPjrqfuXtLttOAdBsP+qABR5tR5z+Ygfnqx9646sQbX9SZZhVE9
Ml6AdcdlMyM0dLoIZksUQDnENjekH6B2ReI/uFXf6xL9w+80IwewhVByEaINxprs
Vc/kF1ctPEQhzSDb1hAMdasP53Uwk9SK5OLIbkaFQIxhaZjG+OQt9eK/ER14Rjkp
xjI9KukBvTlxlr4hp0pskXz4d4tBxmwrvwj0wPwwJlnrDQ5u6+gpLNjqhtLBv5HG
Ss234ZaiOV/muM4MFF2TAzJgAPY1SYGeFavthuFBVUtqaCjTpouxZZJZhiYXr3zd
JL3lPH7xxfsJaacMDkBOkUJ6BA3TmSBSkk3AARUWJPXDXM4dN+kLb6ELFIkqRrin
ckTZxioDJQiOW5ZTutkc0f/bnw0YhgGnopX84eVk689IpPK1rbwdwHsx9ix3EY4w
JE3vsGMZpMQPFw8JkpdR4pHrIjTZZdE3JpRACan5LG3UUy90T1usJPdMHP7nQO25
KQFxZDrzSxplhvCWmdYSMho4AUXiNgwawZ1wrG5pZhuuVfnyQIpp0PybM36vSiWO
6OqeHjZf/jSU6HZxWnyNrt/wm52nfs9veylKKnta3F71iTVRmPdSmCLO4paW+85N
7H0dav71eEwslgzgBcjdA7Dj0pPfAqfCiM2Dy7vtbb9xZabai/G+b10gzTbgJUmp
ouSqObzi0dHnXkWKT2hzYHtg0SEyEaptNbaykkceRfCYmjHdLxtVllrV2zOuOHOy
XdfOY5v6xXe7Z7ZQIKHssY+k5e4VEMnhQWUNjdqzRX5m+3jaJIVEtSzvvaYYVWpM
6kEWYgE/ZJFniVeNnC9q3qpEl8xHZuZh8RiH5OBCSa595AWIHqI4JurDyFo3eotw
dXDviZiN6kzSML06UrCSrQOUU8XGgu8Jm2IwtJ1SAoViOGL9YneIBY54yS5DSBXb
1u5tXZcYYcIESzk4zBOz7bHLBALPUAhw2QlzlxbR1MDOFKnsMEqypqEo5KToiaoy
OtewJH6PbltW6H9PkyI6NaApXumIOHTrk2kyCfLpFzieJ5Yg+O3ILqIDQdLReXdQ
CFiAkXz+f+NGZCtgG5XZBEi+hRimfwA43IctpUqC9F7t+BhP3tjWkQjPk2v1YCWU
zqgm6SeT5Egd5sy5xiWQUzATbYweCiF2Ifgv8Bx2dInD+TY9afF/QxPmGpc8YAc0
KOIHn9623R83/mdHjJpg//vwGKsFrvECIJ/ACrf+2y4cndJZLoheb0iqXL8ff/ep
yErOtzqylQdjA+Bhlud9o3s5HGbt5A2AQXDUixifpghm/ONh58zSIUw0rgi7g3+r
YEhaoNihPGXb0eOLXKTrsOqw6FjZITSZ1g0psZaYWYPMjvtS2Ln5FajzWiTTRhoM
W8reHMnC59QXU2RoLmI6gHxUrnVTAFKZfbg8mvhgODw9DqWTEAUnZwuH1IJqAx77
LXjbrXvt7xuhKLNYfIgioEO8Am6mM4crEPl3DQ/+2a7XqDsVjMLO7mvDobeoVPVw
7APZ+XxOH9IPfJoTK6QzU7gVPoKyUisa9tcBrugeaafh8DceNmoVi4GfGLYiadRj
KavaO/GpH9X2lpxpeNwMBtZUrzDsjKb/mkoEV/ZqFRsMvO7+F4pELmL7u79IKqNv
z9VBI6AHU7xGbTVxUoW9gczjjTZ6DTnjiJ0UNLtHN9HUGElVv9JRwK0E6KGsZwEP
VpBAeArOm/kZcfb4+gWV5X4C8GkOcc/AmzGSlHazk827B8v2MRvxlBJtuiBSBoXj
cNZaqDdmFOrfraKzzHLFdY2+gdujQ+9iWj3ZSNGe0b+9Lb3nJTS9bv8cqte6K4FG
h9NFC/pEny8+3jPdu22cwMQrQKEQ/rQ5eEFhSps8T80PhtVwYcsZGzMXqDYETWXE
3vttpS7R6GSNoMsECEPB3Uw3wEevvZLv1e7+DvYAG7josmsUFTCq12jO1ORGwCgO
cxT9dX6VK0XyAlT5DYirtNp1n+ERmMHBOV2ApSU1eBn7PkxX9LIA2xSHYOAMaxcx
ojNpAvqr/wRKMLi41XUFJKszZdMXHGjOpr12gnWkfmROyDTEO+wiZ5LlKw3oq9eJ
Y7YSni9PgB98dIYYmxvpVEmyN2aLj/2reBRD+sEgtelEdQNBVpoc8mh6hylIccJ6
Ai/uzevR3Qsa2n+im5har33pblVRXJfPunMfT8lOjyjbgC1zATZae0Xji4F5nKdH
Z0d5TRUbeKbZBz/AZ+Su2gl2h0vjETVeDHDaKt9knyYZZ+Xg4rbkmuCQF08HWE9h
7qV1a/t4biObsSTrKcddgOMC2WUQFwPzv4P6xJUd3y5Flek+nZzUJmbXNkURR/XI
Nj8YunCLRJtLFjnpm/9nHBtHXNX8YBdCC45+IXeZi9F+HZ/HtS1V57XoWClC03RZ
xsmtOOanuVWg/2Ass+cOQTuuoKRL4+4LzPq1wqVsIABJ7R5Zx+Gg1MDygS6vtG3x
JxF1ZqgwnkuNmwNs39c7wFFLdie4rKwohayM+ckZ/OyyI55emhDv884BAKNw26Uc
YDB9ES5csIlCDgdDPXjnXFwIQh25AvNYOP8pA+TKQu5aT6SO6lNhvbolmKZVe53k
EEELtXgLAzc+JxVFltfK36i5pFaTBrI1QxMnLxRf0rwXtjfv4+PFtjzzWZpjhUi9
HYZJAjlvQAfFw1q8AxlSsu0y86DbSeREgHoGcFNHl6HwJnvaCACfZf/qxSGEYoFV
9yfZsLkFlpCfx1+niOXy5kKCF5jnRao01jx+qc/Jgw5wm3YoyBJk7g2gZAkFh2lp
T9Peokk/CofdVEwYsAtYhR7zKlX84vpcUAEOPlnR3ZBFCLRnLJLbCnxwkRSC9Eq4
YjC17UkAPd6gRINpv/NGK+PmIYtGkbl4DXpjSiAZ1s2mAT8+jrJ3nolbGqOUjyZC
pcBsK7Bdzbup3uHCrhDu5VUeMS6cDG2JT02zBSMnPWcnENdql/UzCKwdfNGcjdfp
QMmZ4MFtcWGdJCrNICckElwXZoSR9t2lsdK03n3IFpe8IVfe6KkmPKLPcdpeFkhO
Y+XPlvB4rFc3SfqSjvZGJNWGpraA0nIqtoMlDzdhOFBTT8J8LqzDe+6/GQG64vSU
DH6UDqklAZMSKKPnx/5tfms5etvTb9gy/BPQ9mS6B6X9JZod3XSAELMGmnmENv3j
MZD23I4E4d62BVccXVFKAcE4X+YxMHFmvB/ujCkQgwZHXW6NQ852N7GcLGF69UYS
ViA7IO/1Ju52i8/AisZm77xSxx18bDr0tKWWNSF7+r/IvH09Qt6Ww6gC6W/fbLwt
LTneyu4LIMe7GTq8sQe/iLVZmZpa2U6LxhmlX/67uZagXIl7ZbwRb69lwPW/pnZn
JFXAYDZ8T7npFYJEXPezpibjgjjuBm0/cly5H6oZ9+wv3kIdpFbwWMakWX5uZWtP
GkF+zkDa+QBnlqYl9Cd832OWvXmhuMXqCHpmupiXBTOZqbXzPEjagjWWrF6Wkfxv
rHzvcPKbESYUDAF3T8mt4zpMBfaKsoG8jUAwqa6Q13q4a3S0GHttckt3v2Ocgr6e
TmrR8KXldIrkzEURpUdZ7kSC4wPoUi0UFsZmshtD3cg29uX1lOMQz4tJiWL6wruX
+9N42nwVX80zvkaC07y8xTR26C/P+BFqNAma1PyeneL9fQBifxZmEenc+pgnGP8z
LRnXeCah5elQ36ylN7ra508PI5XYhzJlWStvsDmGMKt61ytZiYmoZtMGCJwIMKY+
wb088LeAW1WqaQ9Z9c5sicXbsNrRkYbhSQQh9Dw/RAWtq+onImvo1spxZ+CBfEEo
INkdQOCETS8tYDXNf6Np8USjA4e7B0gH48OEYpGLT3Deyy6BCOHQcwnhLVZeam+J
ENuqnyFDI8liIs8BnJopaGIvHN2SAariLx0Fn6V0QYOb0wQFO+4fIp17ipnrCXqc
BRrx/2f8SCn8rGid/RbLmB4erLJqsQ/GeFFOSV71EEvriSagc8gc2H3ugg443koH
YUg1p0p3oC4+rmvaJ6rd96Cv2n0cIvDvW6nFibjQ8V2YQ2HP+l4oPUxjFLgpuoP4
UqFiqIolGUefKIEb5C/1wPepk5ZR/t8r1iqKn/v4QmifFko4mmlc4niRvqm0GkH6
VCEk85uibhY9anIBugtdNOKQDP43r0xnaBx8n1CeiPACf//Sqrhne9TZoXoSuotg
kuFNjFt+mlsXA3pUuxrKZycQqbyNLOJ0sOs6AfOxk2bmpEBmuggQGr+kiYAKqLuC
GTVQVWkEAxYk+U+58cNT+s76FFHtOmhwt4P0+n8Dj0JpQxNtQ4WDd+R+BRT7yAHO
hl6D7DKv981ucHY55WcYgQOj0SvJwAK0Zb5gHz3OlobmARrj4wg55RS2r8MYk9qk
N2OfJTUWogw3HlosFwVkymn/EoDIQ1UjacbCHcN+5v/WMtFhRH8H4mQtRDXFAcd/
wbvbPTsn932ngUpmy94H9ZpKmsgyCDBwM5pX51kKtWjS3j6umyGmhIwUiogQqRt4
/8oEhCf0dURSVfpE5+Hxt2mRf+vNhXcY/pawkgZpUe5ddG9A6y1KykVmJCshfVXP
PEKEhuFZ6eK6L/6FeVacy67ifBrIi2xvzy8UX4RLiJexnMazNHypoi32VMdSN71X
MNdcF6RbgR2GqugqS01Y/hdZ044E2uo+SFish/03NKv35fSpmUZu6eaE3KH2cZlr
pLhgn3IwbY85JDtOk/e4j4QhioCP6txnx8q1P8DxkmnA7krSdqE4YJuMkDQl+EWl
0MHMDg6FtjO+JfI0t6xOeqBj1c2gdgLHbKqd73/aExjx7QGHyXUxLa39UN+uyGZd
Em6+X5Bsi1A5VEGV21ifU5bkqr2YGgDEu25Pyby7YRIyrjRkf/cIRRXk4cHPuNqk
/gZC0fgVZbchNJhghLw1/Pw24CWn7Ynlds7IV/rpd0Q1Mr0kWerRVXHYeBtoSAtz
YWTBcsnCE/KFcmR3B4+jXGajJ8BTSyNKPPCxAETVY+ETSKjJ0U6HJSlYZDyRqBKJ
OzUyQpEHZOxxwUBTkIJl556z9hNZOy/cLA7E0nSx/fw2gCA0uWPibE7Iu4Xre6+2
2Dy1YhH272yX+ADf3VAG/ZIwB5prLXNVM4uy6Hm79q9yXIh3EUg6DHUdvXqBiRLJ
fzSJMu+DMx7XfV/S6vW0Duk/5UM5JOBBI20TqkY+suENmHiL2j7jIgqtOoy53LL2
ylrV9sg6E4weINr+jG8agdijc9jqgrBd1JPgfaOJvEqkwqZLhCuPay0MHuv+b/lu
srxScnp93voZpcJLeCQcybo47+obeSXNDTmN9qBMg+YMe4XxD0ijo8HCK6zaypnW
t8LXCHlyP+sPLdsR0OO3XmR9IxV8RJFOizUnvYxHAx7Avbu/gKSEaQRzC2hXYRyy
9wZmepuLF5S/R64gTlkq1kKAiZ9AToxlYki+RsJZqoumW/d0RnQTZs8dJoy6w+jk
gzJ6j9fbz3AhsU1F6iDFTYamzoisXu/5o9Qfw2PHslyy7CR/t8prB5vWAZO7mQVa
zcf4qDGF/HSe7MXXw6tgV1ezoiG6UDrCZNY/O20NfNMmHbwSglPt4nuNrJWZQUv/
42YkqYOVvX/huHz2uaXf08Yjwgexj/RUXLOsiu6roM23yKbMRDOOM8LZrGucD3Wh
dMtDDmuHtMTT09sD2q2teGgOl4t+Zkgv17ycd1AN3fNAi6pElAl6IoSGmC0FYNBy
AQTyFPQ2q8/sJFatcd38vjpXAut1yUyILZNIqCUYyeS2JVDT7UCjVpuz5PZTLbsG
dvtjFBYgVTfzegwFEvoIjYsBH9F5lMTY8FS9w9gcCsBdV8Kcz0+wiSO6bQATYK7l
hgc1YSNE9NF7ivFU4246gbwUS7OwgMgPWO7niQwM3kgMiBatHSKGQLiy0FErA8dn
vlBcFVl8lgGeqF7xNFyyTEBORWgQYWM4sT78EWjs/HHemhBa5MZ1ayZgx2zIXsuJ
JzQ04aJC+vh+WjrJnxbLgSMGXZDFf6r+Jyt3w/kYBNNaaVLoRMoOUX3A85oZXFDi
DZGING0ibUkQ7CBbFFSvNTZ5013ik7xQ/BGsJ5vv1XXvV7vnHKoiFQMC/01FwaKs
sRStiYWI8nMb+t0r3vudtKtb6FvJvSxSgPFbt5oazHBZr2I/Qs6NRes8ssXxOQ6h
g+orgJwGV6c7/TJu1via6pTqtqdq6DKokKYpborlwrZ9huF1HnGtNDROPgKwzZzl
6hVEKcFMwVAALz2MdSViSbsIUs0xHCcyuptfmdQ76CeC3KsQmoOhgMIQgMfkzow+
FTr1dd5Gwf7tAD8oJYm8hIsotvF/Zmbg+Qo0H5V7znUc42O65o6WyE8RY3YPSwVy
e5ZBcCG8hiKuDY8+fpIBR0j6KOCZI7gatky9vtUGJ0Iy0VRe6NQMHZ9IB0C6ZLTB
VpBGmYjA1P2F7G3GxL9YuwqVuwIpclflq+m66DWhhN9NFpe+yWrHMAH4Fw7WMnSX
rGUSIn6TNVdUWIuxKl5qPYeJLl9HmtjHFA07WlEUOhFL0DBxyjw7GgDcY1RqGQMr
KE7NuXwY9lvfTHbLmFo6w+p0c29mXqZQgd2cmeI47FXltq1IS0VcH/pgn+GX0XSG
gtsd5MzGL4q02b1r/IEqbdz0slAVpbJhsnbBRVz0QbWR+MSKjzKxifO8Dg3JQc9y
JgsCtpb27pYC5lPnV/K6wgAO6tsmLIKCh9DKAexXHZsAZ4DDC3+qHO4pPxpUqGHC
f8XRdG0cwntLJGXbbz31vLWPlKhD1wDr7JO9eRyPrdONS3UYIHaJsQaeccWat4O4
F4IG2CjJVcPEJwE0QjKPxxykC7HLViwNpSiTEq0Z9uYhKvSh10b2cBFD1+dAl7/c
cIYxekd9Hy/Gc8/de/epJP9T6YL+oUs1megp/CaLX+qLCbBK2G1NFGIkBCKTsmtD
6CX6ib4Yh+XJ9kU4c9/L/6Kuj57idZR4JskczkOD8uQD688XHO5f1HVSVviPVZjQ
6xz9JRwduX0UrgkedIO+qUDEH8o13isjR4d1C97FECH+ZRuBgCvNgtLjy5hG+9pP
V5h46ChDZJukTVMaCi9fkgQ5jIOxYP+EE/iVaJtmPMDe7uzG4SgyWyMLRshn4csw
ayj7GqMlGd3dV+mfIVZ+gvXoYQAxHgxmgmbgDThfJ6FMOmt6THWu9zn1furQcLnn
rQj9LiNyJaNph5NkxO6xUT8eqWn7vI54mWXg+dyQN7QgR17BreBS3DHhuHPKVixp
Esmzew5bec0Zo4tH4wGYJ/LBw+wLPsdLESnifmij8IXsPNzv6/Rzz2iXvWbsr4Wc
1gAuqVjdr8e3TMrMDa8BYDj1W5vWGr3yxHaPnqRiNwqCeDPN30talmaAVKvJpcSc
6Wk5e+4O5961Ty1gP8QGAiPkc3whs9S1rj7sZa2D8DeU6o4cz1K21IfinkmGO+Eu
4NE27150y7Zt6I/zZlqO1h7JxZtNMRTnHuyBlr3c9Fdl3ObzTBgfRD5t2LvUDHOO
/UFX3ljb+ytt6XHFNdqfwdDHHea2ISqGVEg3wrRlkIGQv5UHaECp9lpKk1Op2Sdn
8HTcrSbff3dN8HJlcLbX/Kz66XvjlgwHWGdQbq3e1eblhuD9TEOKEwvqZRX4Sb/r
S8j2Vq9uImj7DUiT4fY6EgVF6Kzu58NGW7lKRLt/WUNFYde9XJ/K6nrGegN+GA+q
xkix7w+8NGnj0uW9Y8AY29mnt5Ub0LaLvNhXfkBL9EAGANt29L39boh7LTkextP3
qiy0eVlHrRoGMStud27P+qqmgF24vYCR2CAGEprw+ISprY7x4CjIwq7pGzzrTpUK
IKeF/P2ZpiATt3SKnpVL17xL2zd23TXqz8BNseHxFYc0vn0wwCVkS0JF3D715MO3
eR6HUAEZ0laGrSQHZoO08ivpxIill3lruDYiOMmbTBORKNRvZCHDi3Eiq4DAL1qO
tTo47dYIfwuR1s5S5yNwNalHp4ted+WOOy0qqk5MvO+EoPXon+DQadLxIVA2zRu7
7djG2/r2PgFWl+lyg4aHYgyqDMd2EytTavVw/gNbz9UeHqVKglpdvKSuuS2SBXOd
XaKpoFppfa0mxGa5Lr5Fl29RtnRS3CAggF1/ZRElW7L4tKBsoHzCcW8jMn+Z6v6y
VA7i6VfN2Q534c/HFX5YhA0HA6kCQvQKAUrmZ+dkP5Z6jx2gLyb4vni7/S76Lk+U
S2z1lCckpW0JsBNy7Ax1+LJhr+f/hFWm+qoAglHoODfJPlwJFvPTgoMF9nvb+bU8
ruj7YptvxyW6tha05aJq07g8MMfJhqIA9udKYhzz2iX+JAJ3I4xlNToAljoDlNzE
fCpGc/nKDtBPpAez1H/gLfw15qII30Z3vTM1x7PlW3kUFZPH03hGiy9Ru4fHTDD3
pb4LxHOjpynLNa4x5e9iGuJ3IadNiIDbW2+NSKPF3LoMMy0mGgQrXqoEySUrbjDf
cfQWSnUUMaGlzblQEQljFoJ5wGUi3uwOPWFQQhCchy465fwIlFmRKnk5kvkl354Y
/MVByTFTAKbS/BwAB89Xy5nZJQzl6N72i+QrFS6GeJlTcItg54dVmHIFUKM+X4Id
NjzDW6YUSeb8M9HEF/vqoT6x4RDnqVCbiVVDbYgC4R3HWZ44lfA+E3i1HLUicr4p
WFdNKkOM5t4ScNjxE0ADjLOevrgYG6xEpe0ajfRmGk/Oczjlxu9ryzyTe+MD1d2t
bUur8iviyIc5AL4esmVjcORTKH8sM12knQM8i1Ysy/YHnp7c+rLZb8qdG6cFAAhY
BKceVU4q1sn1zgOyajSB//MErT+Zoxxqq1hMFCsl2LeiyxdbyA28dbw9b7Mj6OXS
lMR1l7+7UrX2UWf/e/XpyAv7DVFOxdZWdZwuLx51/qo3GsRRItyWhUSKXmQMt7il
+ecAHi3O3d0bt0E9XSVSKD0DNkJ88zg3q3d3rO4x6wVc5qGcz2K1HyiV1GAOXRwL
ShYZztzD9gdGZZ93sPTYkc8ODzU6PDQ0FquehIeb20UvZeaPGRRCrQpyalfQq0sB
MY0gqsr0tlEKOCvz03/LfaYvpAn1vuDV7MfEuZFafb8EQjaAI+tONtX+wbLtOX0k
MZZGprICJGJuR40KJSTN5TZLV7kYTzP15QeZ9MQK5D1gLGgerB5rAnUZyPfs0yU7
4Bb8eF6oMo77LHiXQVXuJfE4Z6jgG6nzviI4yWCEa0kDaetchJ0yffR4Opm9UEBX
r6Vq4fjsbOOleHzqE6XHLloEuH16NVIejYBala9dhTuXDWW+QwClJgPS5fBvWYw4
BhtXZXrhjVrOQeG2a+cEn6FXRPYJiI6pQgb2JmvTntI9IAVUij7i0WR71ltEAk3/
FeSfUuRmxmLgDJAvlebkBAeJD5Lqn72hzWbGsmp1jnYAy5e2HAGkMeCo28GoW5pS
kDIAkSqgZC0pe3V0tt2O5mtWiVO3d4Ew4M1GhEudBnShncYergiZg6ZUPYwQj7f7
1QeOnlTvIKP8/4MxzGtB8jycLp6hyKmdwAyxAZnNO/CXEzYyJkASqC/L2iPP8ol7
A/erB26Oaquvtuduam3DLutT6VfGAwwYeg+6aiM8TXCuY9yM3eg5v9CkIDfisnzQ
iuxuiQAyhT4AikZPVkgT5FMd4oD2RhlI+VZWvYZeGpyo3YV0xfvfnW8bvz1tXP4w
prbsR8kfwg65sA+p9XiHdbXA401kpcayZfYgvDmEHrnQ2/tonxsQXkxbhnrxjIIe
gQPMyhlmM0hdzFOhhMtlzhKjqQ3Z6I3EBg8vANSxNN1Z0sL084C+fbCpyGw/EjKJ
2UlBIPK3Ty3DgfdQDiCZ54DetyBPv6hSi9X55f+Qzjkokji6ZYdM0N78xpCdJF0Z
rVdJVV+v6WEZLbi/HjTAwAH9tqae4rWNJrt9M10E+aRYzaSV3Qn/4cqiiOdT4wqB
t20+fUE3Yy+kiQCUS1WJZO3kuhv5anUAlF7MzvYtrP3xCVKmEp0EoPYyqWK5LxTo
bHYYG6aLgEVz+JkoL3FiShB8wzPHCfSu52oPtlcXAi7EdA2QTCejPU2OgRaOT3Wh
5gSGGiSp2MrhRIwu4b8OPK3zacvidFH+T0kYMgnf+8um6rnanvp+TVhBWXVA35Oh
aDVHFGslthMS98NRRfa+NZ/8giNUE1w3yxXbbKYeh5QK9dgmTPxAdw3yvSZ1ib9y
9l3wzXHZtkgS3EA2znQB9Oo/F70TRp8itnN2DxqEbva4PNZ9/mXcKdx81i9Z2wXy
EbIytl8UoDaUdXsfirEHMU7hbiquaWmTP0W6PUE2t8yrMi/Wwcp99AzniNbZXGG7
nlQ64kpVFweEtFxiobCTZ7UPVSdzneWAxk5KiFLCgDvWNxh9qcYp+7wIuBT+tIMv
XdBvSHLJpbTcNtnsubR7IQav64okv4k0DG15+gG9B2eelGrl/FF4EO7uLbvqZCby
2eMCdU4EsXSXiaMhJexPsMSaPqXVpleuK1SG6QeG5quNP2OYPjg5mFL9rMJBK3ha
uZFYybu+X/JoPFBkwU0sVSbY1KkC5ZaYhAXc+3fbL40yhLU+RKm7K3XKurGnlOHm
6SE57G/gVTFbMaZOipWHEO4v5oZHyxeIiZRgUVLt813XcKrgDAESmlGEnZvlp4D+
exdaL/vPQF3MT6cgbXkRT+404jdutkx7YqWnBqyUfj8obowPqpWuAzFlO1/Zz3ow
Ctof7aD8kAbztQI8qET2Ityf0mitjBbUkYEL70uGNnunyiS9JUR6kQhMJ+QrRfqn
WJrJ52y9NtofiFs0yNMYzjA6L7jbRbfYbGAkDwUghz80LPMVriM9aqsvUWPreYW6
D93NQEceKMsoztF/N54+TZdMOrxL6tGtl9YZ9r1OqzP6DE661Cwv6VxkUyqBv5+3
oUSlrQIiIihEXFvPn6Mfj22k5wBcioevfRgagDkIQoCliEBF32QtLaMdRkYcjq1l
fuCF0DGwpK7Zf5yYOp2DPWX8rXtJBFeGlDuQ6Qs57PZwN9ueGf+1NZ9SRdMojfwF
vBj8a8PqaVhG92Oa9TEuFI+cQx2FTsgzgagZKUgIEY5wdSe19DA2v9c7XLmokgK4
sWgdFPDV5DWVdD1gD4fVxPd9TMAWkF673R0uhd342sxu1cdCCrVh4bgxhgICYJn2
nF9G1fnschVAlCkkRgG6GSgx3D9NdMaSofnv6vEfraWWxCwiQbL/063hJwrbgg+c
TcEXwvd3rTo4UFOLnyMGKNcBDINZYyz6YpMgFjkFfbCWGTMgBm09YQKOCqPVz9df
ODVaAcBM9E2DFSYsKNN2XoNitm0q04qPj+6yw9UaXKqXQSd30RRpbj9QZRRNizXl
lFUXffEtSXm3ItpA8tlq7IClB5ludJVi10MM1DoHv427ddOfyC/Zh+1iICRLF5oP
Pmbdp5wojBWyGKoEcqnLe0X5XQErAmw0/E7eDk8PuqP5yx/UgzCfTvkdAj0bfuHT
w2FtYF93KEy3KSPZ8CBsHzqXPLYC3FIF078aejANVgxurmYUq9pdYCWuEzWDVdeL
HmIh0eqYC7ghhO3V76AK1/QeuaqLUrkqL0+BT2jpAeGQfcPcZPtGHa6tYbfwUrKK
tp3v5fjzetI/h+KHYpwJSP9uPp4cbQjXKbRTDCaOVcBdNsPMgfuKtPSfvEdZAlvn
p/0rOWhI8+I7ehR2eFCUxIShjaORTtTbSJEPJUT0J8IOwTcI2hIw9f021QVbKNzh
V33KSlk5iZ8+qZ8uyJCfNX9ZzepfghpZ37Sno7PfYtestqhPfxElQkeH0aGfJZLr
aQ18VjbxulqsqrkxMRphlNjvGbmvxxMckmmXdRUIxACMHojYLXxBFLuKIeKWWD8N
2hblSOaKJlxYzX2dR1VOxPIY7Cep1qebk7UkM2dgDC/bfyo0zg0c8IpYugUSUfrH
puzmVayWjFe1wnfJmYqKYu4ZbzrwSlS/23izZb2omPG63utwAQvWaqlQEik2j6dI
xOEfLeHy+Eq4Nq8XmEoFJ8i6d033x34HI78Ejt+JAJAkDu/lf+xjbjb4AOL5r0LO
qEr3WtHIuCWK67QuXP8Ivuu4Uz9kddAy4VnYyN+TMIoEbfPaQCwBKboxrcWGBGHV
NJQgL8Y2tiShLWAeo5sHYxtQ4QF6zNA810vJjExeIBP7xwGyVvMzmzwzlxn+ZtSs
0947AOP7Tz1p4zCXkGwovXHEKGysaehEO2rarJEtHqHWN0SZk83IuDnZjwgPF6o0
CJ++Fn9ojaRGdCBO2cyh2Oty3lAIbYk9YGooEHv/eaJ+2pCeVcgtpfosOS9nS4wX
jeNsC28QXDZG8KwkM3drR7NrAhy2lvDnFVSkrtmv3x61ix0HVOWvDjEpWSfoqeRC
3W0fhrhOliM6ghDnT6H1FzsqZaDyj4/9jAmHTD81AIbn8WSy/EO+UPMRthqwccs4
+R+WmJETiInOTX9byGIqdtbjlFJO+48jwp3YlRUCawaNUgu0+CJ12tt8sa4w4MiQ
lWr5NIUlNk0QMa6JFhUtz8FFpco4QvQA11oF+Dkn58SW+T+Iv3kaIl5/LB3/qH0+
hD534g/78KHCGrlnvoHMzAS4YtxjPOXVchN294DhuB7gBJeLppM/ZOW9euSrwz94
TrTBfuMll0lC5rIWmSBwfmj5ck8SeGjPI2+aI/EQRzYoNuoxfZVu1zi800IxPuN9
pCFRrU8O0XeDV+aeJEG2LTdAvKuKO4k8qVddnIHiGQas8BNzbQ8GhPrVgBb//Ef4
AIuHw8vNVLmeV7Rg9oRIDwitwGObYK9L76kzGwDIl+tT3CEj/Et1VFOqGtb6p0/m
QKXS2gUYzgMoLpOBu9+UekFQtX4PkDCU0P7xP76C3i3lpXr0tp49R+WqyMD+cxpi
S61EWVaRyOPanqo79yHFwolPdVbfCXOQrCSNADxZAUEz033lY2pN/7+3o07IsTvg
TtZkphsMKDlMofHfrQbzEfCnHfcpJX/oxJTGZ0ZEn4T+51dyT6S9BEVm6jzwlcYY
TIx3o9iKaz8iDZqrpm2Oe4fI9mA1ES4cO8O3NhVmsqxNeqvQm6zjWyDHZYx0aCF3
OQ6mXTbVnLNgr5684cXIaUn0A7CHYCPXfF6/7qtzTOfTMt+RUXW/n5XFLlQbtMuW
ZMRMm8QOdMXryzEAijQT8BRB6UmuDAnJRM/0n+huvpG3yXVrt6WsGLO7n+24T0SG
tLe2t8b8epu7q/nN3dHhjD3FZ3PiM9mJc0YIkin8iGQFnntQjso95MUQ+6bTU7R6
u4c7P3nt7Zc7KSaxXRo6dDB4ldfrdJJG29MKjWg6kDbG2eOFxjVfOUxIa4sjOwft
3K49A/Z2bjVDuZR4yWHRb4Ak9RsYHFCT8DQ8YT8+BM8p7UOAo+/OwSDGJBxygDZi
/8qtjuZC7cwu4lo6umh63HmBYU7mcN8YRiP2p5BQqT8R5hvLHmWMC82XsO7G1HB5
7jOetJwImMgz4TLeB8EmVMt4pN0FXlIz22wsXiZ5FgcdlbirX/1vqHJe14/F+p77
z1/zIue6Y8j9qI6mMfBaXik3lupOAwraJeZ5RUUi3SdS2pemQkpOPF/vcMlaCNl1
rQ0g5PGB+8Dvh6H8o8T7khltOL8VTbM7mMQvDT98I/6lDXIIBTXQ9Pfe8WUm+73h
0jn0lxILEgrxvj+3+vxvRUBEwGqjaMKF722d5dffG1A+dDfL869XU5GWkz5QPib4
OjUtSIlcQAbkHQTIwV+iunR8sJJtKsBGSk9L6+zEm4ZXXMGf5B8FCtOT8y6nva3w
Lj+DqRdXhEwo9Ci+IQbBC4C6c1aTscSDHbIUL+rrEVnkrF1xVthPk6D9LNJh8aVV
HfZwfzfvqCFauMz6DIQfC6y2xLSkhbVpure36iaurABPDyKPYXITqEtG4iwx+uAX
1uQFBEuB6hMjHAleMcm9T4Z6OZTHE0op5kMkyOXNbX2gUTI6a3q2/7jp4V3DQwox
w6pgHGz+Fwm2T4t6MGqlxrRUjaCgwxCv7tu+NCF4xLVNAAskod/WvZO1UhE3SHtn
pjlPIo8DHAL/141FU+LIswqQM7ndEUA/U3zrXD4e/llaIV9T1SQ/swQ5tdeuFpue
W58/lZH+gCcGwEPE6M8RgkQCqFUAxxd+QTqPVpKxJJl5dDOmWhyxK4VTz4CgaJCu
uhc5vK2jv0gAp2yu9o+VCv+ND4Y1oQCeX4YYlcOFqbRaiVtUoLOeIFrRUNmgIRRb
9xSpYG/fbTHMBxD7V9kYJvRu6Nz9XgG+b9FHazTbDT/iT+/HgREet5RUZpMN9B0K
9rg09QgUVvSrkrzquAC9TjvcWyb53BuSs5fk69Vj+Hij0d2FHnE+Y+KmzqhasK4Z
hlHMsljOXYjltEPfC+PwhCLk05vrll4qnH2XeUnCCPW4d9gIIoAUorPW34fZb5os
1Q5IHArEHJohS1IyZanYV8sN2K5TkjicnQY0w0DZcBcQKi6GsRFgkbY2/B6JiBot
EmnB/Hf8y6qy3ZzWWtAUqJz7PQjcRkdm1YT74V5aPmF0t/cC8GZL9T6xFxBn4D3U
c9c0oyV8WzTDbMceEOPkvHtsLyWpTaeKh5J+3Pwip4QlDb/y9zSYbG7G1/W8totH
mraO8yzZ/pgUdOoL2yNbz4IgeaeMcebKuBOR0XHLlIFVhQgTSbACIXTloe2gE9AB
GvaSz8b0NMpTXtzKY8b51k+b6wMDgZFUu0HgVRKrEzc07Diogd8Ujg9DU0jSg7pT
3J99CEBCeZUzBiq+TNOPGnXMnVG98ELzis75LQU3lz5ItQQz7xF5tH068qw8f6eN
l4fyeJix8aTEgcoSXlNNPY6sOYSsdl0YcdBfzLsk7w0hr7wJZ1M/NTqlEPccKFPJ
wR5rQh9x1ljvPmqPibmZBk47cyQYdKZLbI96NYIV8zeeHnwXYBOBwlyvYIOErHvQ
ApZJVmJtjYbKFlk01CoMCIMRabLzxPwrvjDxAOQOEtGcGPyzpe722Qvyx7JXDAQx
U14gK9qBA0kSD6DBIr7WDjnk8+UswqE8dfE48hK+bEzLD/752QHKKel2R3cG2yth
vAxCJFbwvDEwoEvBNmm4gbUN45tpQLrnxqL9LhyNQtYUJh2zkP3M5MwXzgcPG3dp
3NH+fOY+y27nqzcLv5jF7lVof1wDdFgDmywzGpDZYNDndOoZdmzkA33a44bvnRRh
/0OOv92O6QLrXJLXI9xHVsllWf0bMMYxGYQ0SKcvKORo4bEwPiIDGBkpCB1sa8YB
+n2HxXp12K70H+lCwxhFMMnsp6ug/MjO0LI2J7wyh2KDCYpnqCGKs2KoG6qemUS9
G2iJJ9LhOcSPadNXWxsPwRlSoWgE03F6PO6Tb1DcBglB05wP4XD3a+yDgWhfDRGx
w/UdaCT8D0rVfmbIRH2Or9rb309N1U2VADEqAXiaux6yW8CI3kMmdLlcx5F6wHIL
GtlCcooz/O7n/d7NNLRknr2ucjWuy1YQ7jDCtx7ysvInALDXtndx32vGmTCFXy5q
iDQ5QWdvzWFkQBRDEulvMenIyoCODsB0cUijtwT2t47zMLVNc/EkTdyJpX1CV6PC
iAmn3qyBneuDbugP5lNcEgym447kuDb1sk7gIQx5Rz3VbBmEp8o9nqm7K2qlhSQc
HkGWLGQ9yTF+m8zBOooS9VX5FwQmoPSjzZmTQOY9Mf1IQrOGF0ljrU6MhOb++GuV
DXdhxx526H7f7vkDaOlM1A/OHQuwh/D5zr6887ykGDga9ZtpDRnkn8wwOkhV1R0m
8nulL+WuVySiauqvDRDP1zpB3W384lRvA8tb+NrY7EfUOWBXrYEBA8sgfT/UUTwL
q8rk2uoG4jEdLnf6n8i8mYDhVaLJsgMqsylWc6KwvKfq/P0BkLdaC3tfw8pDUA2F
pGTHctX34qvmAEL+P361yYh/iXct67/2BxB9dBii1+u+UMMYLA0xxUGBTOFHQnEH
0FFSRMkD5Ofu/iVCs4wkPqUbByZkvXyeJi9sVdGg10wOW8iTq1jD/6IRUVue5IVZ
1gn+9/wL7Bg/o9aIUUYymFeFeDuSf8MIsWm5fHU2cqpQpHK2S7HRMz0VScycfgVd
OPV/vXFucYbT0Sj8JO38zqrxWzg19GrmNXVUELR/u4L93cBH8ZV5J5p5qdcQldks
TLpILtKFdN5OaVrUyFXjZxnU73oQx9a5oXjos14I08mCsymMoyX/llP82ENO0k8W
HLCBMPx6UaoFbuziVNeo1fRoXGyBpgUumtij50+qQY6WG89Nn9crBsgYaZ4lIKDP
IhUjfGpj9xvj2LQGS0x72ayMC+hrUHXyrklx5k8ogUJrbo2sC/upUYpWVEDrFiBX
oWgeIfRVPLgMWZWtGj0B2M9oVvxSSa28DADA784fLCflyoz/TiLHA81L2Um9NLmO
+TzJ7j7mCiCvZnXq2tsXeEiDdVpXiysAwSnyvbJImECkDHcjsy22mZXGCMLFSFPP
5aJ1EK56lUbHa1S4FnNvdn0RqFSePNcqTD2jAfZig862T8+DR9gJ2MbIzQl872eq
vWj/ttL2lcF4CqV0w/NRfO/1DyrFc0wwHksfNaeRAgyTn+HVjoXjczUq8OVwNUyM
ktcugPV+0qHfK0abtChhbAtzdJQgp32SOaVlc4FdbEx3nAepZ29ap7F98NAlrr+K
XwAaE9/uN+m1gh9GdP1obR+V9W1a4kb7/CvkAz6mY6s46GhQJLnFubGDzD2kWI07
FH4B6mhzMfmMsSC7CtJV4guVfxekcV14WmwxaoTc0+jx5tufe7njsTrnGkwKVdWZ
zS9MNskHb+97bbe1T338NiirzMqQdsqxAvuGEG4GsZhOkVVYBfmAZ/S7ITFn9MoW
hqJi1/8XywbYdchy/CO+NAqTrjOJQO6py774BHlOYV31M2/MDXCkRcKjHVUFnmpL
h4FIbYGiGGoXqJEz7rXSPli041X24C78L0Vb58mPCRzzBPSGMnUMtI7/dKvFxHa/
GQTPV9anGH4GoU3rmTWkcqQsXTvVWNpS2R4AJ8FjRLH1XD+BeGNyXw2vY3aowpUF
U0VH9QDDml0iRhbpLhszpx2Nc9hMjSxeSFUa3YgrUJ81bLmuNdGxsLtlYUPmK968
VLkcw6vaGyyCaCwZTFdkt2TPDxWADpKzkvKarzYUXB3Bxzw9gwNoGihCOTRJgJIe
l/nKVyEur1lcolCd4b3a+an8uFnegOo37AMpLgrCM2xQvSLYI/xisCtxOX82/SBc
Ntg+bFDuwstWxn7nbEqh11iYwBvVdCbI6q37nHooL0yyPwD3gAPJxNfPN8/vvri1
i0pT4tpo0aIJrPCXBwirBcObbfGTc5kc/wpRaRWHQdYPr36Hhyw/SkNT9/HYl9uJ
dDGydqpuyX6Gr/2tzUdHJPiqrOLTL1as+NGzZZF82v8Op3KC/f05Xh0llWHRJVxb
iirBNFkc39c/TgbfHD4RIysWvwGObOAbNrz+mDmqo4GyuU29VqfCpIM8iiA/da03
SBo86MhPP4D5S+BAgkoPfO1MWT5Bu5aBl+EU2n2fkzhzSPN7LuJ1HzgWu7sOm4Q0
4sMrxEuiAZVoA5aAety0lRAZhw9jH6fy/CBLq1aX4SfpwCY1YXm4FH+HvO2aQAwR
4qSAyoHNSqgOoTd5gFVUJp3fALzNxYpjxH14f7SMqbK/f9ZCTh1c10lm6ekpySnI
IlZZyLheKyd8zP4JYN3pEkS2dpHppsxlg5ceH//zgVU39AuShmJnPvjuOxBuIgox
izSQ2/fPDIu2CCSMptKK9iI7YJBxG/GTUrCpN34dLGXeRp865eUth9PLifCtf0gt
6Doe8Q2zseaKtGBZrVW/yvDvNJ9MMcbUPR1vUn7K8zfoZqpNhbNU6RFA+g78s5Eq
u+kyCfDqNVgmg4xjK0GzCyV3Hq7RRAmkoSjGw6kzmic//9G+pg5uL6lAxP1P7Jiy
qX4ds2yBPAqzf9i4+plNZAGtB1vquLNRWO6ijgIrdFxfNWn6amjV/0X8wAnpUgRe
fVSFShl4jKRY+l+DHdyDM6xJKLa2O2DJBhSTYOh8AInGi0O4H21/P6KHrh31pTiO
DTqzRAamYf0dicpll//X5c28JaIC8w91LYDfhNQUitHmHSRqSlrKbHTte0menUNe
YGSKyRAr7Bvah++vbhqPa4a/Uj9EisXft/U17ct3MBcOtrODadePBkvFcu1O/fOA
wJ1DPJSYSssuIIMIH86KewWXg+cZmPxHfQ13wgHmbuOh2bRN8VE231hxGssoUlVe
lyQSf6Y117WO07MNvDIEnj5aO6dDWFoHF2riui4VkXIza12LkC+8qaGxyFT+jDPn
2rqaT+txW7krBLgUB5knrmbBthLo8/zohc/S8qn0jzv53BPavQroy/kBYwpJVmw4
pxkwxKTq4Ez/ykCYzpSNvWg1IzedsbNluwpUBaLoqZeLAhaRko2sXf0a+dYD4CJh
j2juO2USt1Z7BnMyY6q4f39AUYn7/putme3lusJyuyXHQq4OF1KFulrvU4/0wUWf
ZG5K7jLf6QGoblvrvBo4u2vzi3yLX+nqhK/uCF5rVDzDyIKhiDkZJdOAk0wYZvYX
AljZZ5FEYSu0swvaDS4zwozUvRQ/nde3JLgoPSYY5ZuAU8zslYOHwDDSQplggFfY
SzUI8WoP9AQ+px2t0KRVCDd8se/TU5v2280nlQU0Y6XimUcFGQu3gn3C0HaP6pvy
lWF8R8pssiGo9J2uPWlbPHqULmEE+kE1mYGMYsRcmqZD5Z7+EbJQOkDK7AipHjk0
wc8apJVrzll5IRSSh4J7HTSpi3dEeFnUR2vJuh1XOjUoX9fKTNcsehCXLVnCU2gP
aFwqYbpwy6HPVNO/KWsxkgCeKHi3hceosfRFc1evLVC4yhvNIwRwyi0ty2EUIB/G
XvweFNr0CXyUPOYqN27jBZ0ROJg19fGmo8GCpQYGEy6pV3Jau9qoaPVMD6/4Br/v
fKgZZhIVHtkwCn4h8+0g0DwQt8QILSUmuzcZ9bpaJGD2wEZlaGwV+BhSBJEh9WgM
pDgIjPPS/TuekqjRIXI4ERcuwIk/2h8TRUMf8ZRqte9RW/IwB8kcVKCkrCFdOKmg
Z1LkGinhQUXK8siEk+NRob2AxJboDm7apml15gypxKkLmyl6lCFQ5PKzsEGRrI/N
t5hKJLT0ec88U5empWFgc7vKlMVNMyCilkQBAK7VP5zA7+06lyjor5hA7R9CKMJQ
1XcS7pi8dt7QhDpAXsxJFcI0cFOcZQGrNsziJcyrj8SPX7hjTFqBeQo06M79NwEp
QASIDwNDo1Lq5fd6qPqfoOkJpWrZ8qhqjkLruHnLF2zO6600Bnk1ElZ1sfNSKo8E
y5IeKdtiDHl1cp6Mc5gQLXIT6Jeqtd5bDNsuA08vrGBPiljB1wZGaB8Ja1jvnVIg
/lnnRNL6BCCpRBy5Blg4J6J3vNenaqOfMUQSwH9IPnL8lHHN6yYwvcphDFcRL8RN
rgju06C5drTunJineykwbzk990HLVRpPcwIU5WaHvuMyLFNtaieFMMOK04BV0l+q
4f4QAJx1UfE60YAMDgkgZJCMT+g1hZknYJZu3Bemz7ix0aJFSkjxoIcR46wEPu8a
SsAx6zk8S97Sfk2TbtI2B0cGoAB5bEuAmmVTF3o/pysL/wu7S87Q14/A1VuyFxo6
XzTNS5K495Hvc0nKhfe1MSgIvbnKiQtPyhKmlXdDRJJ7alfRJkMXXUrOjfDM4v0Q
z4MgXvLbKAP+vsAtizebepIItKQRWKLDgYu8aH7L1bCubNHDzV/YJleJyalkBpj6
7NKQdmnUPXY3qZEoJ0H1WKPwGKhT1UMFBJuclKGTe1mpBtdW5hUlKpBmwLwgx2TJ
aXe7gj8uyXHFC2lemUW5DvJcl8h6TeW8qJ8LduiuJSAlMiFIT1FsrOjr1blsdGdw
EqeGizfl4D97EHG9dgbDTgyrxVavMZA9h7kf4cs6WmxwlbrdBAn6Ulg3FhqY9LnW
kcAlrCG1WmIxuYEmzA9LdMiynt0t9watFUM6Ghs4LRdBbNMF2GtAHevZx0jdkl+Z
3ZAQ4BgWf/P+tsRb0Zhy/W+LrtQx/lMvhX+AbyJruTh+mNyaBMoo1XDIvi6tdMqC
YOAkkRgy9MxecRPJettSl03oW/MbM71WwyLD7u39vDEhLTbMiuWz63ddnnfwmj92
eNRqdY4pRDolyaSBCPT+q6bIa13Ug8OHyftO43dGCBbZxTZj/YoIdOJd3xCjfz+c
WfLyTqpht2Tv9x4ne7vokhF35wXadRWe50YMKmQdBiC1YsxX1n/iJyOCqXRGtFuN
1WDbv7uUsbdoT9Tu2kwTTsPt+s7y2hxkedpf5p07/MCYNLV+2L0vrHo8X6RRbUuU
H/KlVcY0lp1bLOS6qru79YFUaN2jV8WDPQMdoXxHfHpDM9zNEwhYQ34ojXE6/rNg
7QOaIEuodm7n0XS3pSpM3G/1NTtPylb1Fwn4KdOvji543bxJG+Ajp+u5tgYkC4GJ
08JSrofy6GP8LPMx4EI57SxAVCEwA8XB8ICtjzTDWHn0naMoOB61saUElSsUBlAw
9shpJZOpcjRH5lJIcKSnhJbPdDuxNLLOA3SLBHYbwo0h7zrCY9sk+t144PYE5ej0
t9PkrkzDz7dFwSdwbKXe54OGdaDwllt2vhO6YAZzUV+eWzeVXBLNPb0TfpzdE+DW
qiPEVsQgSH66fOYckHbnfFsET0fv3jFQeZAOQsl+vlY7g9Z2hBpLjRCno69bE/0b
9A7yjgT+ON7B0R/TKD4eyZULC5GvmGbYguLeM1CuhaZwgB6eZBlCTqCmlXZvu54N
1CBwOmknfJ5e0eB1F4ZbYVFmZWuzEB35X/iSVzQNlMiXV70EjJfs2VEiMqL/AE9z
ryOAJwM5C8DsEGWfWX6UQJRgtOnC2AIQcOwOjN45Q98x6fzTFYYFPN/HE8bVGddf
BNCNnrb0EoBuUCfOLDrtbDVL1l+oACLsLNHKo/ieKaX9iccQ794sglRTN/w7aSa5
M93mbZv6v5zdExRxP4URzHcq453HE80MVZLwFVnzqCA4yom9WzZCOuOQOUTFeDsZ
Yq78apW3d3e1RpGbq4WYQo/xrlcfBPnaajLelY6n14itWAXhtj5//Z4ce4cI/zzo
NB+GnvRKMH00ugSrUi7QK1gq1sq1MgRK7mfRlV5puZDzQ6MiNSbSfNKdzRYT86MK
8j2Rp7UHbWC1c3WWQ1TBr/1wNIBEnzHQ5k5A+eNC/mapky1UsQO4lqGNcsmQ9Yti
SrhH5YPMgaFlcBpyxYjnBQtouX03eXAx2q7wM83VsRNs34WVfpjMIfx25XlnAAXb
y0ijWeJ87+YQofYSkcKyF9c0CGltV3be9Ac66bXu+n10Wy6GEIOLmPk0DLKOVQeM
kh90kEoBJuUiith0YPcorhd2+CB2cH9/XfL6P32/SVLfbhKesEo4/IV8UPdwmqEI
mX6ikOVZ2swim2sQyHyTjDDv6eWOcx5JSdNaZo68BkDcCiPwnTqKet+Qa/syRPY4
g/jFjPcCQ1w1cidPnMMH3swHyRP4v8ROv09fuZZt348TTmexvhYQIHwzYMRDQCIM
Msz4rnRmP0Uw2RvbVNcwkn/gg1dneHYAGj3ZXliKEB30Tx5yg49rA91mfIAHBmoi
2S+d2aNJmY4J2rJ0AdvoTntv83cR/oXi/9kL/KYEmeFhRn6eOfUww12ldBlbJjQg
vV9kbiPrlCramSqunVupvwNGJBnTpZ1EzGgjibkbPdk5bPkxoL/svBm+gXFmAvwm
GZayxh68/eZGQbPDsht4iG7dEp62K8Al3nL40hIJiZDOGRV5tOQsaOOMvwrISAAc
tsyNMqg3nxcCNrdkz1tKruutea2qa4mL5Oh4X+4v1tyZGVLuDwIM0n56v5e2VD2V
UHcdExIrkaHKsZp20J6ZjAkHSNLrffKcRG8BrQ9xii2kvRAqlH8df+0UamfLYXcc
TiTbQvD6u6P/ngW+Z1H3FkERjUccsPMWk4k4BPnviyIS4Lq490iaOZL9l2EIHkJw
SEZDYRjYETx9qgnIzd7jL2ExsyX3TC6IP+W+c8GKDi9WcJsSUBfNUE6ybZ86/ECQ
kVu5O1lWAyg3fczqHITHR9XeazRpOSnKnZCemu5XwLXsG//ulu7CJsexholYdbBt
4lFOE5oR0YM3FPJ3V/3Ym5O2PHtacSeKmyoqY40DHUWnajEJypfk40lt1fLNN9ld
vjysgM7mbUKZel6sQdctLESxFgP38yAIAj1KCAd1/B50w7OjP3WFzZobNFSRV79r
ipkT9PFG/iJt4tm2V+sLIKK1heCkm0SZzgd80X/zrLu1khcfSqGlIuvS6+mVnIYt
o93AcsTdWmGm1UxxRpWmrDkw+jJ/qVWkfaTZgDQEXswx3XvMM5tO39WlCUwCvMKz
pc+hvI0gRhvwSF8KVDaYrT8n3yfeuZ+sHqv0E29SNG+pWYOP6LEEiDiqJL4kjZGS
hey2z2pAAUGB/k5XvY89VWP6bcpoJDlTUNUNFkSnhVGE8Vevx7/cxqeL30RG5DQY
jqOTpszTKEAk5WB7jvw2G9DRbsLrCI9EVcCyfwrunP9uDbjbAy5u+oM3D0+wL7UP
XvLHO5I09JTy4lmbApKJhs6ihcfp6JiivFnajtzHLbXtzEw79YjDxbs7Hfj8Z5fH
Lq5t+nh5xoG3jq/CGpShLaBFiRhc+1Rd/uSBwCNPT/LwGjnf/g00/GB1ZoGtK6PV
dGDlCXJdVJjKKQKXrbiqg539QXFUdLfWalnX3RELiNIZJrtqRdU+Lhg0w0u3M3RU
Y9U9pO2VppoKzmLamjh1rZ2otSvv9S22uvmmhk7b0scnzlj8kfYR1vEkZkwUv6TC
zy1GevgovjNw+hL6A6ZFTUhUZ8O/LsIVJYuZMdK2pIjskRypq78Gj/oR42K2v6jq
DqmQJlvKRGMXE0b05iqB/09LByPMhlcXInLZemmvWoZhasRPyZxYcgt/A4Tghodw
9EYU0Vg0/Nq0blc6P1PaQ8ZiBs/q+KUtJHkqgfh1Mk01YB5mCPu5KTkEVhGehBdz
RZUtWNKtedQN76DgNfu6KMegjkstcC0/JPAszFOsYkVLmRmVppS9KzqzQ17QMqd3
LCSxlDLkv5+tsJ7SrzVwx0k5wRR7djyhcCeaoKqIQ7Jf/eE/fbGf63kO/H0cXw64
QLp0vyy4I0x9gYOks6cgjDvgUYxU3E/t6eaMt4XiDr+P0/lZ8DwNpuKvAE/CJZhK
OdlkiqIVyzlSrcHX5lxGQvkG+jkSHnj2/WwRKYferm5VgJscTKSceS0AodNiG27z
6tmhdGygkYqh9pwGrUQ23h/jT7GCt3QPpGY8ufYlLQA5Wj/vSF0BiZ4IHec6QWBi
oxhjl0shlowEYpAK4VAmjMxBCAj6FG2eHdX2hFkhVtuKPJLQd73dD8eh8ikwDYjE
pA7hmtMy+27WXFcpCN+YMO/7nFGw3dV754q5yQWle3q3/BxZrqc2mJvDLoEFbqk5
GW239sZpm5yAbDu1yyWsMn9BhmiFhu6IgvRZ02djT2LF0oRbWVsuChsZrsP/jnn1
qLZQLab5wDJSbYjKVtGML/oE17kcxJZplG+XfQDtYu0mRt+cS2RPm9Zts6ktsI/T
ZuswUzkYFbJd5oDrUYuU9G7Rw0bJHoRYtWhY6jgzth9l0X3U+fJ1XXUarcYKH49W
Ky2mgEgliEvYxI3XijjrMwbo5O6+PGVXWmibzjYVWClEcWzd00AD0LxMwL9T3Cuf
Sk0ec/qdxq3fKi8BPhUvefjxvR5BhF0RT91GRpvVtRX7Y21RL92/O64/bluXtiWl
WMLUl7ICTjZpJS4gLSYrxodrHYtKF7IJUH+XSu9MyS1dENMi9vS52ZEj60tdUMrY
0J+7xIrAQ5VunSPyEk1/ev19jSSolQ1Dzi5u36+Ccjzp1vv4UDGvN6bCI0Gqc75u
pA2WVuz+dmCi+4Me8cI6fjQIw+3vP2SuIu0UUVSP8Q9DazsNlXQg4rg44FOWeTO+
VS/XEp7stNJOwM10oGMEI3fGaPGc4vIaYZt81kbt5eOtFd6Ixb4h/1pvD81YrAQ9
KBNHztl+fG8sutw9gjY08SLovHXcRvOSK8yVWNqmCJ8tMljWArXONte848kVe67d
ykltCeHKFPs5WLAojrcXupXLvV4N/rwaGXO2s9v2Y/n8D8eHwZQz9Zs1nT7vN5lW
RohrchzNQaGWjo/lD8zvd8n+LgEJ5V7iTQJLDcy1d/gusXF8LVVkdrZi/HbCt67k
GpSPMU+AwhlBDwYC6dVHBSv94VWi+OlTMaHncRXGpVqFZOxIX09APiV+5lAQnzt+
H+xHep8FRUeWgVrhYKgDUI50GunVtIx070Pe5R/paBQSz/kp9CYrf82zcaNaTKIP
eyh9tU5D0Tvjg4KgdIVWe/dYftYnCpr/7D97G8TXM8jh1lJ+yGv8u81SOf3F/Cjj
6Qz3iCAMxg9MbHn56AVw40ce/LmA22/xCc3pWdq5JJ6JTAvVtCRnqVicSU3JdCSf
XAttv98LNCxM0Ql5L1ATukiQu0Pq7qteTSac/8tWMU5EuHaKT3DEcjtf0z1cfZsq
chJMyufbs7fOmwudoaDtu2mlhbMH9Igmw1FtfS90rgiTFFuv6MnSeRMlUdqp2beR
TUjR4VCAPpZWwkV7srR3Z0XHKmkhfm+glvVj8BAg5zY2VilxcTH5q+x6IQ5LnO2h
JmEmEAU85fZ17n4/pxddy7/1z7XIV1RSFrlwljeffgHEyL/2jZSMZsAX8kO4z5jH
68/mz7w4m/gr4DzFcdeVLaPbrvUtnz5mHdajOpO0CBhoXz5Hn8j01lch+GQijYfv
CoZWt178iRh/UiLImiDDqtZYYSGCsVP3TRW7uFnUC6ahDQJ/NwEeUmLyiZnnqWV9
/pDj6h3WGLrorm08KASUihZokBWOsTugob7W1lfiOQM/DNRx2DbPYQ7nqwZi3Ihs
wOukB4TrEKgq90BnPTqYzTL9J3zB/f0h+tun21pzK+qSHqFgBN4JG1anvU4CxGUH
NIszFfGHPvJOVKLkKUmQXAnEpxnFgVDGlIhtVNdHn7NR4UnMOLIybu9aAx6OiV+M
9oKHyxJm6T1ytyO7bnWGmxCnT+4Rc5rO9IBEFA4fHFgRgH8p6Yzpme/5xHePvMAs
3jT9WaHmEHEG0WuOn1laZDaYAZSgFOk8GpCDyjzPNtiWNTfQsJ5LvH+MWOAc3pqg
bBVr1AYxEEQdmadDIkGNFJMjYYszu7ZBDMDgb0SMyEuRZ7uUJ2cVkCzNRW8M0RwH
hrsMAeV3xnkx4+H/yQ8GggqKGS4SZWjTESajpqorI5ZKoI8nT4AFDIGBp5EgudGL
aR5Y/VeSzTf5QxTb6p8WQ7D4uJrWB4rueoasuGSm1WXFrp+xThfAOuTXGLOD3WKp
rzyG30I1GMO7SXJ+q/EVGgXjEz+rRx5YVNhzvC56V1K9JAf239u8Tv/i1/5eqnNx
DpjS/Y0qbIiZksWf/qYs91a+qa+TYrWkJlGPDmQkZmJsngpgu+7U5fm8JVuswhAs
9CNM3JiXMiTe8ZCPvj16srfh9eDP3hYt1f6s68EmaeN9D2JGKcFq+vvcIpUf5Doa
uamNyWznC0uDL2UY8a6cyXbvan74e3BUO2OhtIZXDHWinwB/Ga84Ks4pOTRCAMPS
lzNP30k8/s8+Wfop33PBjeDKqfbWrec7TH4if0OwRJ0Xk5RIPUC6aeLKM5EOhXA3
aj7UC08L6Ib9TV65E/QzYcC3en4Kg2bKgFQ0cEsz44TQhVug0yhgC7uZtAOt8GAL
ayKvBBFugR1KHKFh74uJTpnY7zeI05q7AEYqO9teBP6DHPtp6RPPV+bAwJn75PlK
I2EAhMU7P+gEKR5XiTw+Kz/vHmQTaHhwDNF7C8yGZFsPiWoHVftKz55M4CkOeO9f
Tje7lx6s1mqwFtxqALjdWi0Km/t1M8pWFK5f0c5Roy5dak4xbz3+5tPFYNXKH8t/
/85EZ1aFUULdjKbSch+7VprgE8PW3NxapNClAbJNgfSZBsEYvMw1e/r6343S/8wq
coEiZ4agYoR27HkgHPVizAVbT6uLIAwQB4shAzWpxdQmArbq1sRBN2T5Fnl9CElp
4HcY8P1rllN4YZ6DCfv2TsGUsWFMkcFBMGwy0v/noadB98ReF1uS+h6HJxepA9nO
n3fWxs2T027BHtyK5kEJtxNLRKH2c3apSkpwTKhPpxjVWHey+A6oIc3JgDPr2hek
4gLvTLRTkb2S7u3YUpPKd9ap1+4ZgRkUjmWs4jajb6uagBRa9KTaq7PGxt3Fh4j8
GEl7ZkMnJyPhK173Lswi9oss4Y2MPTmL9O3+DbrS8XyagHMbosZG020+i/s3o0qz
l7eN4Jeb5xA9WYXm7xSnFUfmJlaAFNvoFJVkJBnaOBL10Cx2kxoEg1ac7n/tDpMr
uILtXR8UKG1UaKmljKKTfh2FC6XPu8GfRGBEpufqpuSalzwtBVI7Fo8U2kqzBSPP
RgnDR6uu539+7SVvdTNXC4RPpldNqCGOZ+nSVwmFi+FhaHNC2TNDmyQN3N5ugqQW
r0bbkN36raq2ULPiusbvRumvHLEAnZUN275NVmyxMWIY3aJVP1OxMaKSsQXi+jOs
1w2BMKqKafSsD0FdCDGNcAWyjBxeoqDQ/WqOjTGEECXjHh0P1qb2MPmvx0fVKclN
jcXp00+TxpH3O2ZUp56V6FdMKlspnXgfM9sEww9KMJnMLAefTHLA6KSn5RDbWn5S
QEsaWPpLYvHNOf6mnweD/D01MJTn8jqHtk5bcUTy0hItGzanP52bzDPiiHCbOoz7
NIHLE/ZuGdyRRCy5KRq6HuxfJpieOSjRy5O/R1ZvxcI7rTQOwGHM02GCIfeo2lby
JWPQI4XK/BYlcW8b7gD6Gy6Sp1KpYcl9Su07bDGEgeQMq6gPDxhzfgCs3Ubt9ENb
XjrjNqHGYIre0ESgy7KIKohDyQEr7mq4+x3OKKaP6HkVMsM30bDvy8jt3JvRXy/7
OAFegmLMhqIT/GpCCryUielixqF6IUtRWTdsvXahLDjrVZ4cxEClBIT+ZdzDbn0v
J4JRLfbvFttfuP4gvxMvNl9teokRkNRwbvidmjGW2AQ/1kEpbOcSygtTa4js0sDu
g/71UOiMSkj3g3p323mkfG53SMyf86hPmoD1gnt5I+4i/etPGXKNaWVjcTWghTHe
ol98bfwORLhz00MC9gjwzXxeKIbhByPqUDWjcgOI9nWd3RU6bxxVehcJHRPcFIYK
JHE4mEZRpAzsDZfmExCQQsYotUJRb5uL7qEGIVqjD3bxU+93efud2i1xZ1/Q50cm
GdR3xWL9HMXBsXp3gueauY9yxx9Ah0oqNEy7JMHAJRS8CFbtIiKt26UvSc/JeqjD
2QPELTC4H0n95UPB/q3ypcb3Vm+268TXtdi0+I7/TFZzCYEjlvXQmrdScvB7atLj
dBGAOo/Fv3VA+13HNYdt32K3YAeRGcaX9QIkRIzG7cc8Lfuhq0LanRedggL+oYg5
5NYYmv5hUVOQBEtmxBzZliuWmLV0E2GfYhRL25YCMI/uSwt4awzdI6Qsk6HsL1JT
7Kx2y5T7TU82wplCSlnJ41q5AsgE6MaLWiv9Z7mddIn5hH5pOHkjZwt22wz4LUHY
zAUwRXyBVW7nwcPpTGhfLMWeqTPYaNcpTjDGAN8yGEX2pTn+awVWv8p5rmI/ht8S
80c+NN4TR5m/k+zSI32dByZRt3SkYKt8J0MqDkXZ3OcwrseYQQQ5Gp9TejyjsrW+
6Vrp0NQPtDuuxOhISOzliC4pcAs1S7Db1EqonwCeK8tzN1i5LhgdKtAsaT/NkgXh
kMpVXkBjFYDFCZJt5nXQkfPeZ5MFFd9JTqtL4kqLk0j5BkK322U3JSMw8MMytZ2d
KsuLeV9fRIyTZL+qtk0CtS4Ew87ljZJusxZTD6eBrlAtOFH1gNReW/tb8hVKRhwF
UPl8Byvv3gq0v7GCCzW927AOOOWU0zy24DM+yhWwmbJjSm427WJmpAyQ5TOuJ2cK
iwDFkmaQGJskvWzXfF5EHb4kpKKqimWOEqxN12ysdSf0vJnsajtcNXzbhO9d7J0L
PGXuoLus4aFtd3eFAasUUDf8r6anuvTVkLp8o/7IwucIzJXaE5YT7mmblzY97VVc
u+y52I8iXEvg6S/oc1d0RTR48EhcYTOgHiR+KgWMti1s+AseBIS3SJkuiRS2WjUv
SurfWzqBj15s5b3n6msDnyuwkbThlrs+IHV+qoyLhVvb4vhS9O/LHE305vOW8+jR
Vl3tawE6trm8/wRYdFMzZloVA3/5Th61MGhx1nTWz6U0/zG8vaD42AXTS3Ma0DXu
79vgs/Bz36p9ltFEQ/fvoxFQHVNV4RtShnrUT8d14w66APw+tDOMdOi0lJfWk/H5
+Gjy7+GraTNpd/BdmG//QSMA4USkfZqvl1eLCpkQyp3eReHPZvcR0QIOAe33Vfeu
5zDxdilyY4mTNI6VCuh+DVRNe7SML/mrLfx13GVx8S3dYfqJbSCdZuubg7dNSFOR
uJQdRjD0LJK4eXR5JxE/RyYHUphP6s45D1fahuo151SZuvRqroE77mPwNpk2RedS
PBHTuQkFoggu9cPqMUTwJSHHFkBYXGuFkNUZHsh9ZtgMHC2k6ugy2KbNtHfPdcOe
INzF0q25kQY3Z+Mo11MoLIZjhz1adlU0TMcTa1ZWvSHaZM14cMppvRntTwYF5eOe
RE7HqXJrdppKIwWbx/WiEXV7suWfCjfXO0A+J09JdgeNTpJFRA5GGvwhw/TUnkN4
7nGkSAh85tVF1AxKy8byhMn5GS8c13FuBmD0vJGFSq238iP6F/1g//SkWMPuc1l1
Yli/H2Sd4Uop6qMititqB/l14byMdFL7qUmBBlLvSZUyfEMd6KVDmiDy0kgTDdPq
NbXcRfdHFt+EyTH/t+pxOeP5+Jp8k6TF4irpIRrGsvYB+FqPAhZVUqX0sxMmZIHM
Q9d3KcaMjoE9k43zP6FENCFGGTea1ZIhLowcOQs4TQq+6qwPXToy6RPDP+/3ziZc
jM64D/vnqm9Zwg7K3rca5b7ohbrY6nUOv4BVKImnFZ8PwlPYqmJiCMCIeFDOcpsm
z0e5ue9nSJRs9j6PVDI8iCLbu0VjHv4RNmZuRMJNCVmguff7WPDW8suTGkDJ7Zy9
uVrRen0yld35qNC+PqJkbOdsq5lnCM5feo1W8iDilkVXVaKHD3Mr3fFe01gxUy6g
Vpd7mAvTuegYUmoX8CRLPhl2J4HwE77x0iOhEXVjKorLnpqIZshbyjvmt1ilvsUx
F1HXXRglU5Zt5YaTiGabSLDPBaTRJpet/E7z5Uwn/4uTTzymO2iVBpzmwUNnRkz+
dmYdtq5wcpYUGhXNXWcqg8LzEt+2XaizTM7G9yfO025qp8R6wIyrvWq8iIYR7Zee
iXxEduKochnR2n4CGmEWQXQZw6X7dBFktNNoWrA2WAH6ejJIqcXYwaYsD/ATSfFb
eGvmFc0W5S3Exp7Id3UOxGCgjTbfavBD0tJbf6gMfZopngnZziX6K2LVwI2mHWGz
9iT3CKKZ19/lNoiat66V4/BL9yt2w8JTprX6MZ9I8qN8ZWbxgHwMCX6E9zpFBu+f
otUJJUYlgutBqmS/iHHB80X0iT4U8NbCWCOqMaP+7TC2mXzVify3buO1od387Uqd
lwvuwfU+f0S9au3XRNgXKu5padT9y1yT1vfQkOSiETqjL4G3/V0p7CKYYOFLO4Gi
Nl7KXZDAGOnaMEF3BaL63kVjeBKIVb71kqUQJwwmh+ZkL54yVu10r3bOVni58UgQ
Di+Rak/hBDARVt4mxmYmAf3EUIVNUK2+9ehI9j6/0fHn2bhJ2xEXl43y1T/ZV3gG
Ocw1mCjymY/rqFP+syyXR+k9LI073S2Gh5Cm1LYFc4NgxzGjPDItfxYPcR508vcU
7IME+K+3Sl41PrZIMeh7UbGTsLGzDTPW/z5kaTo53EIEt00V7fH8I+Mgvzc0Hsgs
B4R6HULQpjHo5sRl1fuUgBfuJPd6YDPh+E63FstKaulDLmyUd3aiTzishS5Xr992
St/CY+nKQTAAsACzkJ17c1QiR7SftSE0resF11g2GXF5UYQeDZ+rhE9HXmLnACKr
NUwDUt6JE5qXTk2EplWIYCL/OPiO4/P2IruyvyAwcc2XKoiM1qIvYIzJHNSNhQaQ
fps2ZVQKgopY7UJgsSnWM3ZGjxAyU2RrqcdGsj3XddmMKOaEUWzM4u/Rqd6nCfGX
rocapZe4gKL4/+zhxLpM7Ce2MYHeyHVpAUJcbZOAbXotvGEpdtsWU5DyL6Vs7opT
8HHliAXjhW8FZNzGV9eK8qDA+8YYiLBc+wAATYoP8p6CFDASYgTDGQGJKT9kp+it
qF7yg1TnIogzZbFeXu2fqIqbXPpQmJckwOy7ZH87gkabVUTxcrJ/D/0wy604rfve
nSSBlhR7WQJtb8PyFkbIhiZiLdTHNBJks4jv88uTcfOHB13Q0P1qa768+zcdSGPZ
4hP5p1a485WUi8DbHvtRvFHJMet8pwZWyrC6/iLblwRJ2ZFAPLKKF+V5tgmZjbiV
P02VWTfJp17zxle2SSAIa0wLH7WYL3Os/oA4Qx7NJZUIl2soB55tpQ/EDBPHRj2j
Ktv5oy1rXuJQag7vHlHKuET4A9DiK2adopl+Rrj8Y4tLqDyYFFOE94fFtD3Jv8zH
bCTVum+cIuny2YJmeXSiZc5xmH5JCFWao0br2tyIZVcafdjbPNudTFX1HIolDWuN
WwWk/gqEScibjVJhZabqjsiQ6NVlSF0o2GV9RamXSiAAll1vBy9YJn7S2q2ZZ8i3
eZkrCBzeuzuGeyIXKpqgkxUEu0ClypCUrbrLl/bQArrfp2k4aamgzE4IO6yuHbJX
UlmHH6rSp7mE96HIWQgTlsvl7BwOxSqOARDfZG1q32bCqICeczp9Mqa06wCp79Is
WqHAiyqRLY+mrviuNYXZsa7r6TfMjdrJ/JT2g7hXwhrIbIErGCYH4NmCfarsQZT6
CSDLMz4SH/Qb10yEn79qiMAvv6/8DQFmz9DV+4KrNBPb/GUCJ9YRvTVkUVlhjRn5
Nbf/4thd82L8BWcFuiH0ffaN7mATvREdLro6Xf91C6cv/qjxu20VGNcZyU9nt4YR
gK0z/zRRJzhiqs90FK1O4aoW9Rw3EIydNWuVoeKOSW13xOagLQDcbiT6JOXJc8QT
Me2aZ6haTKPlg5W870e+qJmbUHiKb0u01Xy93W3MBw5QgZjLo6DEbn7nGpabjenQ
bze0TG8iQcGE80oj3hsR4A8GZ2DcG0RtJ899opbVm4vBWf3bB+Z++56ztfG76Cf4
1hP95XYls55hYWjEkCrWbDKLsT1II2sjzLg8857mUZbm38VRTXYyNX4Fcrq9lq3A
nEY01HagqzomzEIdPO/aWbI3G2hwDTFqD8LR5Gxj7GDImy/41GBExa8iDxoDm3l6
YdTQDn7G2VJ840qtE0P/laeQzfAKIKmSczh+V5NXgfN6ZkRG8ymx7Te6jl8n+Z48
6srvwYuJQ9FsPshUiXliQhrZGNAUkUBrfK9UN2QlkRZ2jm5t42uE7AF8k/dkMmoy
APXq7sRZWdS1J9215HEAQKTXawfiH4/vnZSFgyh9PMyqPNz60g1T9fHF3bfnLg1+
fFIXuQ/4p0cYfSf/1c30tU2M60VghDeT3SN8fX0fcM1tZvnWCX8DtX5sUQHpvWmY
Uoy6ZtroCTpqP9dI+uwLlWwsWrSeomOm3aqX94tzlASsXrOs+DRPJQMgUL819ycf
N54djrJH29wOwSzqi+/52tE+ifxgluTwTsf+t/S5bmcjVZI+1xDJAPn9Ocn+IzhI
Rw9rOGy1OGKuVk7ZTcIQNebu+J7Nafv4ViC8Gc3E2rLFnSkyXlykvvpq9I8HTgWv
DUBfqMT+drgD3w9duxa/tmBlFK9pDkPucVI4yzHPY+qYWcJHZYN+ZARYhUrud4VN
8qEcimjoGsCKharwx+QaWpZ/SW/59oygzyApqaKaKE9gzyjLC2bEhIMQzxKv8s9Y
ESvNZqfXnF0czSX23RfTazreWVvK0utjUcg7BRmKLn0if0eOc23uyJUbbgzd3jJX
yNo8IK/Iw+gAYUMZBr7S40WFZ4a21vUjuE2WzS5me5O2u1iNQ3/MwCSoKg0DBwlQ
0+Q6FJtve9/uvwiBiMCIqx5sEIYBfB5Ni7t91aok1k8GHSk4xn2Fbqz7xo9W4Ks6
bYaAnqfVTF+LCFt3TLB3A1v2aVsQ8wvuiTuj4BlVlir0SWuuGE0GnWqqgM0P4l5T
OUGELSx4iFq7LuKM0+/PRpE/+o7xnltiExqovHMq5x99eyUqwZARBDgsx7cqMWT7
AUqfRqH4GbZUc3kaVvvp2nzsKfLasJFQyktfNR3nt4FszobFnOqlA4jKCPttq7uh
J267+cpzS5/XeWxGbv5dc5iCQpta4bTm2WmRtwOOeCIt8BwsYGKGcNi6bqLiB0Q0
X+XfW++LplWSW8AgcIDKgjMpC79dE4aPhnotDfnPUMFzn+e0dxy1m0y4ba0TMCus
hd9p/jClcBBQ312RB8JgtELrqlm1H9mSqkvkmoWunuCE52uTzSdTyjbIYuSsmg7p
ZnY5a6XIYNuamn/K7ukYVszC+lMFeCXaKP/Tt/s7KwsQvZ9MnxSRPjKDKtBYEhAv
3XeyHWd7KIXLKkTkhKjq74Z6nv5dj/4GV9SE4oHgNta1ezqeS12bt8WEdWkYW35Y
TVaAB5Y2bm13XqZnyhvxqV/sJj2mQte+JA51ab5sBLGa6rgjg2m4a17qWfsCRnAI
NPFfAHHCSwGXHcf7kSyhCoNNl7BlDGO2nq/faKeoDkg4yXTkB0kH7i8QmEZe4Ot5
AfKfJw3VS84orWOcBFMUCsGahAsf884WViP2JC2wXj+pyGxyXA37hAY7wtqYSDYp
HtTaKrnU2l0bzD6qBVzgvrW1fHjXKOXUlNVZwnMJYulVCLsBZPyjLF8ErabVJpR/
hrEi4Vc0fg/iwwd7vs3yngZ9Vh+xejfRyZsUyysv/8Spn7iqrQGzDwy/4+BE2knc
53I+kUrdZXSYx69bYeKleMwWWKSptLu8SbSGh9gdKhdnod189CMqfGBl3/VytrfE
BYshD4RfOS9ycuZsh0mneMCVfk/2J7MshceQDR2n7b6USr908dPBvgMhzYQvQ4rK
bcNdxsExtYutHVVIvmwYtKQst+257UyQW/zntsDuRwHR0/NxZL5/ITqaUchDFowS
ZVIiMrTGlzfuva+MdP7Bb1qjx6Ajzy6BRV5cLdA5s+PjVvqyt74dJWEBInk6826P
mevh3WB126FcNlQTlD4/G1GrqaotXjtFx5ZnlX2SYWftFrXQYkWi2+dZNfImryCE
fi01FZ7rJCUv5bi2kdrpvZpaSBboFgLfxosPI+KhmVE0XxaleLAfHUQ2vPnO2Zxn
zOHyhfKmkc/CQ9nQ0qAxJ1zA1tRILLFRayNgsdGCJ7X3vPKLnTcppIhBZWvS2A7Z
S+fmbhgcapG/SLK37r/jnLiFq9IX0n/IZX8pTOTdLiKKPxp3f1qXtNnnVEGS8IfQ
p92WWh3Gum4B6vRSBUc0k8ztEOXprXoArX4z/mMP+F7aW6elRJfOMUa9YobWLmAy
8sE+a3Vo+1VqeAPL4G6cT8cP+gDazO4K+nxq8spJNMXThuQmrpfACGoiuWzj+tRY
oC7/e3rA5gf6Qwr0D4YiRCxcXW+nlrj3Kgn1MxKllIP7fxhVHqZfhSv0NaoO5f1H
8NfjPzZ+7XcBnhyjVRqABC1WAuILg7/ACu9gO4Ji3nu9AIYF6gYCdo0Zcpr2ypR2
wuK+BEdsEDy/s2bmdez5bJrbGswPLNsgvySzQWNAt7FOxXYbgMsa8gq1deWjROVI
YqNFihjM7TvmVUNnuM19LToMPrUwpaI8WfZ+301up1zJiot2k4+rf/6euDyc26ow
gv0w9S9Q8bxoG0P8YYJ5sJLhdANFk7MedsY117MzOjnFu2DFhXu0VzHUbI1+T0hC
xIN+sicQt30o+Qmm4H0QDAtkSDlY6AxAZTIu3L7oIReS8p3LbGy7pSr643mfSMQA
9B8ws8f7tqFI5zcK6lFWxcnC8M1FM6IMAWdVrDmEgpQX6qNaeV1jzqCukW0zotyx
0Q8ktU/cCIJ+ToAlYVz1YD2tG7sd1vdkFxGcFQqvmByLZaG8X3drw2h8CqGXD6Hd
G/vVnrOUUpZ3XdZ8xjndx+DmxxIH94ejsWsX2q/OBNpkgLPs1Y6Vua6rnOyTryXM
YNu8yIHhaaDPmH9Aeqg2DgAP91mj1uLwW4ayEOrO2xF18N95RJRKhTnhpu2UMmrr
lF5RrWf0EcWFmHl4SxQwBrM49G1Fkq6OIzaDAT2d8UA/WQlSpR3VZ7+Z4aoeHuHf
YcNLhXPphlP5CwEgS0y6o7CcLo3ty3OmvWKXEW7RB216o6wwExX+wiVZc2jg8Wl4
p8D9rSpjoYhCT92JFbuQniUxtarl5oOZVOLcVDdD5J54iuerMOGgPPk5JnoToGGb
tVYVrAggXkXSNp13DOUAOLBjM+j8yBtfRDWKd8UdBYnl/qnTAwmgdDK8/d/C4U58
hpQNKMDghkU/KyeE3zcCdvC+4RO9TqrKRwek0NQI5F53OEiLp97A3RrWN7BCmlSt
tOpsy4pVgITVq/3lkxx73lo4nqsGSdDL86/N5JVEW4LQgrm6z/0Hv01ksfK7P7sF
W8J13NBs96h8Tzp9u1GFqElGFo5Sx4+7lmVIkzWaOhGfb0hW1eiNwF1najYBafhT
ZNYlyMUY5HHxRVu/XrVbspZjCerLPcfrLFMKXPVEBVIGL6bdX1p95sZcafAzu9uh
hvfNF1Y3masqJEd+TIYEZ45aqdMlkP8PYHhLhMRsBuLYSI/jebXVqrc/922ndbiY
PiM0Sqjc0QOjF6dZNrn8D3kKwkdE9tTiqNiQdMyNmkq9M2NBNhSms6oT7nouWtPQ
pQJ32S6bLJLoG994v3lTiaid9Dm4pRng5EYUkmKtWrQmqNkrIv6JxzfnNYBKVRmD
lwWIylM13nLlb5nB6/2g2WEccmnn1T2k4+S/3C4+X5YhWYRh4OMZRVho0ed0ntty
pSMt8d6ufdLPMMQv6b6Obszu0o5qiht7XcGgs7jLqDydvxT8sLPq7xewc7HPWMgt
jApd+qyzIdMfTlW1nZ5c9yRBJa/o7yDkusMtsLoUFccoyJwQQ2cTecgkYl7TdXVR
9pzNEIkcTAPt2zdQoosWPwqW3JjfHuigzpjEg33W+nUP/dBwHkkGY07rFvVdvdAy
PwV3QXa7sk+65UT3IzvO6prNcn+Fe/cOgv0DB/cT/WZ/jCKG95XqpUwKjC4OOkLB
89GqYgJf3qKP/UjTwr0HQWCJLyy3fK0Ih/4ozwhg9mIi9VCu+f9Z4+xD1dSpi9WJ
/cG8G1fwYewQG1rGFzzM6xejs+Pdw4kFMaXvRDmbVAT4fRzf+UyY7n0ld8i6Kqp2
6kozqPP0dNZZZgVtX1tvJnQb55VM1TU4PaWrllK7HRc/SeppnLbSH+z5eH2KNE8U
dXJhlCk7/uHSJf32Or9JvBvSLlBbCACUUoDfBXwkf9N3OhI+6ZQ+Fq4QqKlU3+ev
tOPAiqemiTbmH9oKi2NSXk43qAMiJaSLCX9PAXgl+uwjHjmEgWF2UzxMvriv7R+C
cE4SGU2QETfhpM54zeQCL2eCgCBp0XD2NoFX4As3qx8IXOcM9StXlOLqP/9en4UX
DEDAbrRYgSgEoICLRix+zqjNCr1+vRu+I1LQtkJkIbr5k/WTc91M2U3R/SNOqPGV
ZGPdoCIRZeoz7SThFiLm86VNWZwisqUlve/cd3yoKZk=

`pragma protect end_protected

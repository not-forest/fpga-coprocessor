��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���X��f;��on�# ���5"0 �T�PL7T�0����Ǿ*�Յ�'x���!�����*��w���0`>���M�I��M���M�At�YY?��w�/��
��D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��Ěכ_��՛	�D
�T�da�]L7��~yR�����*̮A\�`q��*L����vh�P �W�%�ƣ�� 4V_'ķ�0i"4�qy��)����'P����7���X?FM ��	����Wa�5��O��2�R�ߨl؛�߆'(�}څwhe�[�H��~Ԙ��Q���fG��)6bO!K7�ޜ�I;�x ��P��%,6���~��D Q^�BS)&I����V+ж�Vp�ADP���(���w�+6>�����2X��ؖY��utxY #�)�Gj���PI.���w��{�E��I#+�LJ���DS�h0Fb����"\�{\q��=>G��c!�"G�2VS 2�?��[��Iכ��6I�{�(_��e�2����c�Ě ��sR^�����l������P1N޾��À����x�w�0��`!�-R�X�t8^*�����KQ�V"6w	��7���Q%:��6L(wx���h�[��ớ:r�+E�?����`�$�}#m��6�	6\�mh���	яzs��V�������>�KK�Pvg/�G35��>��/�{��O˸��^O����K*s=��n�-G-$L6�#�t��-L��'ƞC,bZ�*�r&zP��D��L���!���n)�п|����o5����U�\�a�(�#P�ꌄ�w�hIA��T m����>[;���[�j�H�7��O�uK�S.]o��r���+9?������<���;{�^���$�̧`�Lx������mSd��L/]����{!u&`2�������$�)�{��v���,�z��5	b+iv�6r����-�Ϩ=ڰ{��@f�(�2���<y����=�u�S�ĉ&����>��˽CE���䕧l�#?����o���e	+�<�UK<x?��YqB+��`f�/zPZԽϩ���3jJR?���9��h~F�Q���@��KJ` �M"4g�Is��z�Vy>�e<�֏��]m�4ʑU�==��>�BEゞ� r�,�������U������Y�xFౝ���2�{&��C�}ALH.ܶ`f����48[�,	���c|SJr|�c���&�B��D��䗠�Z��C)Z��F9ީ�Ԗ�ݞ��bԄ���'|%��ZY��)�����lv���=���E���Fo�Rw1dn��
Ʉ.O��gm�5��MPU�\��2�^��Z��0�<bWN6ח�R�;�'�S���� �Hx�m�����}�9���8e���n"� ��!$�
��u�H_�ݒ�U�o�r��Hi9U; ���;7�~��W��������P����� ��u^�ɏ���N��V������cExIY�sj����5���H0�~*H$H(+�eZ���F54�iI�ź}LB��q!��^��V疣�g�X�ЃҽEĮ���#����g#�j#
0�������	3?�Q�}����/�#蜾%Κ���B������N�͏edX  �_o�mj����ѪA��Rw�a�>q�7/G���Vs�O���Ob�.(C�a�八s���xv��[�En��J!}�������OyȨ�g��ц/��徆�n�r���^+��Q��6f�$l*����s߆�8�[�n��ݣp�w?��2���F6A�R-4K'��p��i��
&tt۪_�q�����]�e`LzI�Tp�Ҭ?�j�yYR����w�:I:�L~��^�=�{�[�&��y9}�B�eǆĄ\��-�B._Zz��[��%��"J��Q�n1�՘b
�d�!�������y*�DO��(� �@�� ���95|�J>�LR���
�a���	���xn8��Ʀ`��N�%`_˅tL ��P"Fr��	'��4p��A�K�4&3㮕G�L�Ǘ��n֥����8�n�ډ�q@���_7��t�j�y���)3�L)�x�b�W3��)�G�k�N�v������^Y��N�{z�-��� ����U3b�(��,6NN��SE�c��[s5�ș��W�3�g`x��YK���X�W R����D�~R�.�s�Y�9P�O�iE�
;���f��:mM�gC4x'�+m�n��l�FZlG���_ey�v��D>1X���o+ x}q��s�|�,�qǜϟi���
[S2�Ӭ�*Ȱ�n�@�T�xr#E�l��Aׇ��a8D�ʵ^W!�>�2�V��{}�p��J��Ӝ#F���������+ C��XXhY
���P?�N�`��lW�ov��ʔK�PXv��̙�b�4 �Es�=ʍ�`E)�s���	#@����Q� &�e�.��H/7���O�j�չ�uC�v2WK:�́K"��i��?�'�6��2й�W"p0"g�3�l?��u+�FO�5>����I�<����4T�ۙ��j�{����ʁ4�Y�#�'��X���=�{�����g�qR�x��&M)���q H_׋Y62ј,���q@�����[��7{5QD<�0D�&�`Mז��Y`�//Ɵ.�������d��ehws0*��$�6�W<'f����|�dlִì�� ���@��Oi�S�9����=��RؐM��Ϭ���pMqՀW�;���"���ݑ����}��愸[ȊA^�u�Jz�R��3�F����5�L�޾��}K�P����N|�1�1�q>�L�N3�Rh���Ԯd�$�����|DH+��yl�3:��u�i��[lN�y���Z�chVr�y�L<�]y!J��Z��~M���A�ce�g�y�0�b�s�#9�9��X�d W����pO2+֫�6@�+y!��Nl����?�$�w�w������J`���	a��KXHh_��6Gʅ���Ej2.�qDHP&��aP替�{��0ڷs�XU�2�ʺ\�a=���]@kR���u����h3���#h�8?����#̜�v��&�-E�m!�M?M�a�%Î×��홲s(nS����rDևc�ޡ���20X$���ؑ���"*�#���!2BU}�'OE�Ђ����g+�6��[b�9�A��׷��4��Ղ��ӳx;�ƌ�!��a !/I~E�yP���tfK��<�����8��y]F��6��h��e�ri�o���j��ȆG�5����g�0��Zwe6K�#}�ϞX�߰9�;�#)���������I)E�:��/8��h��̈́i �4�/��ʌג��Yc�	F�=@F�<�w����@O3�5m�x'r�<����9䨺6Q��|Tm�U��e A�=�$�˳ʳ��s����J��5��^-�uFV�=]����ӈ��b�f؉�P&�F�t��
�i�-kҘB4�6Y='�� -4&��;��tk�"$V�Ռn�C��Ġ�Q-8�=���m�H���E����#�r�lC@�jawwЗ[j��� XYt)�K+	��1�wBlLuK%�W���|������q(U�wn��!�ɤ�m[Nf�n�=����]F(����������ce�u�6�m� `�,���Y�����Vm��2�BM祗���;X�x�L�)^�}@_}����<���u`_�����=�MNT�b�b	b �/�}�a>�g��r���� ���*^K�^�|�qL����L�7�����Cq˓p�F�]��v�UIb��L��,���#� ���-��$#��{.���C`h���W�[�Z���������qē��B��q�rf�C]���_P%��}*#�D�p� ���W�"i�`ǋɛ�Ϛ%4���v9��Įy��i�el���Tɘ݋*���n���0&0���ݏ�<Y�P�^8�W6Y�&ʄи���wdg�?ju�p.&��hT��k��F�u"�q_/�>�7���ɾ�}Ȋ�+�ZO�Ӟ�P������:Lj�S����a��2��h/�?��$�V3�k��l\�H�#VH����*UDO�>�����!Q%�Z��K^��m�������S�h��tL���p�Rc���Nhz�^����/�JU1d�����Ǉ�!ń����9Iig�j�����,H���N�I#���H�y�vF������D6�N�Z1��WOe�x�﹕QU�|�����&Dl�����"_�SVk��l0��$aT�������1�<������nWy���a��r=Ͷ�y�`s�]B/�B�Ҵ�^�X%MD۸�f)�������h�K_�#�$Ŝ�NJ
E�6��ぜ
���+t�N�!��tAb�+�R��p괼Sُ�f?bPĖ�_i�(t�~��{2F'�}���(>a��%�	�9�4���D�K^	$ GB���y#���٦H�T'�O�p�-Ԓ�M�����2�WX�'ń�Ĕ����hTaº���_����;�չ>qU8��G(y���,Ӗ��N[0�5=�H<\G�q�.`;�㫞~:'쁈��r��Jx��u٦o�ذ��&CQ-���$��/{�-_�e����xy5+�*����Nт�ȷj�q����/L{@�lX�b���8Uqᕥ���tp&d��L} L���
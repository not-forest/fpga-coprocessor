// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
L+7praQwePH9Md56sR03Q1ALpN04tKTIPPrDeheXnZjx5wu8ubzMf2HZkhLlTjoT
D/8JJBnRlIjNfLQUd7ADwFUG+h9CjiEeoyDufa4NpsOheRoXc0jg86+++WxVVxRN
rVBNrMNx1Y/SiwxumqtWTd8suUdClMK4iJV8idgJsQk=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 8592 )
`pragma protect data_block
ooBe8S+3/Roe20cS73WvU3cRgB0vV8w/jMsYueHkdfmUidFafON8BqB9jNA+Gamp
lz0J3pLNEARgvut5SYxkn1Ft1/xzGLn9GdRQhgF4xXDJW7HS4phIW/KBwCLSvJxq
enbx2QDkk+bJi/0DTIGQJp4gTSIoTkKtBsQK54v/5bUozzM5dwb28l0p41W+nfvQ
CLvmgGJTmYh+TjqVP8qG8rYAFhNxt9frPf8+ZrT0cuSYbsbFR7uTeKOt4+Xe244C
NxURbWFutAaZNKc+R6dTtI/oYP0BAurgL8U9+esP88V5DNDKNsPZAc0OMgr9EVg3
Omo0Uh/4WKZAcLAIA7u/e1QRvvTRdsqx8qmeKwpdnPMz5cKlUDwouNX4VvjR/88o
jCSOum2Umx+1U584RZTqEYhbEGGcDh1MBpq4dJuFTUTwbMlAD+WArsb6y5ae1dZ0
ReqRvyshRKVyRWoVB+tDb4m2D1Cvo3RZKnd+/pC/HjWwWsrq3Q7iH/qEsT9Y/qBU
C6XGdJyjnFMSEf5Os8agOmVMOi9ORoyXH8uwNYAx1KoCu6G9vLdunNyT3mpHr0u6
/2n4Pm9E33Y9oKQ9Mj1uEp9vzbszR//2/dqEySw+pADVvveZQm06RjNKbn2aaY1P
YQC6kjeli0qzWHQk1UKTdGj8KFs+1YC2s6auNRWzkme/pp6EXijHvRzPS/H6eHkC
BrFNUT0QMRsIq6/ygeOnf4VRMZdThBHdg1hcNaj4FHn0nyBPQ0d+Dfjx2375yFXX
wtXlKJF8z0yt34RB10E8lRpLJDAuFtwQAE89aUvedITQtNYHdK02fpXGXolf3e/V
DOxeY4/xy2q5ihU7QdEnHVMfSVniyvL9EMAa3s3eCsq9AO2h1+g5Y1inXVOkqHI3
wJ2pPKRHs2Ym8xA37aWiF1ZblZo6h9VWR8lRRzo6bNXOaUHYQoIA/thyrpp4kftM
kpqJXQIJc33xYGCRMhS9leGvdthzApVN/2t4I3M8GyAguTEZgW9pFW2XRGKF05i8
lH+XhpmGIfDRtHqFebmofquS6mUnYQFr2pZCmzXYqvGv5X2ccjvXSm0QMk0Gh2f6
bFVSVpydY63jMzYQpgA0P9C5ipW9e9rdVVfu3/HFpguy2JJf3ElpWRSx3LYqIWJE
iRbhFW7BbhZjDnDnJaXtOxJ7sWEseG2sc0hNWfT4xXEjDu98N8RwOCaYDBjHZJiD
JOCQpMH0aHPTFxUPg5jmcuMWD/attnTb6IoSvxdrKKftFz9/q2kKKRI/0C3ofVRS
gtH+r5/tQC1ZxrjXUj/PXOjXn8DKjY0CYctO/XBDCpwRGZQ7mul5H3mCIOCl4FTx
tiFijGHRC6IHufC01AYerCO21D9REVO0daT/ufj9wIFCXRfaRSC040eqb8H3b5fh
SuNjmdL+Vz+db71mTbA43nGfvGpbIfZAsaL4ZNPpolZDJ7oqbh68y+oaKHoWL5Nw
SuaN/5UQLJ1da4pscvBylfz4VJ6Z/7GO/mhlApbbT2ru+as2SJfGB/wvW5Fghp/x
vrBrrMZokusOKeI45B+S7J6eNAVigi48U6I759AmGyYefVp+5UjP01ZA2+iOnAsf
8tCSeqdtzK0JmhgPDKs914hUuzg3wLyghFoGsOMb/xRSKnYnCl01wf9cdzgkVFP6
zVTvZkyOY/sxD27jhVNeR8+J93BMmVmHSc6Le9y19MaE2yPGIOL5srNK5yxiRUL9
dxGpt/SnzItmr1GM8gpYG8xyXOsBj0f2dhMF3Lus/WwZT+km0p1rIayXw+hDT6gp
vT3tVa3zuv9CjFSbOZ+Z/PxlRvY9kizas91G9sUe+S7VTIbr71K3W4XRYRNbQW75
gfxRoLZjrgvvbklQS4GDDquzuFpYhgXghxb4KyV4MICx9qAMMUrfFyyVIdJ4GozV
gcg9yMnhGR/KncoXESpiYMcd3XbdEzElKjlA1nCuN8Vu/uRFu3GSBfAkQa/bWyA2
FUzJ79Vxh/2twpM7GCJrwHdeAVZfgfEWiQwTm8j7SQdkaPcVwionz3cxKanmn3P8
ab7KgoutE0l8oiW7hcPCsGZqewWGIlYqD0dkgAHf/hAA8ONAuxi12XUBpJozpA7k
3e85HK20DZwd9+j0mdpF1Mu8E+5je7+Nu0MU7rqkK+cbQC6nD+E/gFzu3dOE6/HR
I2D5+f5aYCWTNeoQwg2b3+ZJuDk2NXWDv30oXoVMV1i48B4iczS13kzB8arB9qX6
+FvfzGC3Hz148IWmcxPLr7+NnN23Ckj71PHQaJ9j+60Bim7ePo/PFMZdIJ87dPsI
tpPLXztvcqTf2bDk/w2bdANKmjOtAwtPT563U3mH/cjXEBqM3k5TcN5xG+xim8lq
TYYkpaM3OXOrHWk2AGOK8nrBeV+agL4YAgKBvuAEA3MOloSt7hcdhPcMF/8IqnOq
TLYfAooVi8kdmx0hRIxh6sMrufrWOllYPdE/BcbG7XPgX3iwLzfKt9YvmjuospLO
FXFWwb9809gZHxR2zM73Ky6MnUWmDdyxLi5mmwNl5GrhYYekCaF5Wsdn+Et9xBeD
AfwSwSsnRdR/89njgtRpsdzkTIemvCNlF/ZSGBBEmnjRjHs9gbHNV/2mIYCF1sFD
HKV33I3QjDB5//TcapXpEiN/ZPw25KY4uyvls4fUi4QijTxl2rVsDB8F+Y39Fk0L
/lCWdyqKTywXpePAy+G3VxySkKl+mDf21AQULZMzUCEHfEn/3qEHCZWu5IFfjqAL
U1n398hNMR85ZtLPgscfYU+I89CLSf2skW0fKk1p1RYh/q7kNGOJjqIL6aeleTC0
SHhlUfPWJhh6mVVmUZZcug7OlsA4u1EMHRqfeybIMYmNzDDQh0qKOnf6s5MKuk9u
BLS01b+cxs4VM/daBNW2256yVfy7Nj2XqI960IGSaFcbrez/atc1d5u3hWZ8OmPb
krirRr6B8z9B9ike8OpyryrZl2W7ALN7EoYB21wt1NrlhKW0ITcj3fVdoJkHXkYw
eANtyXPRv5LmTQ8J7+WZfgP1AbRf4EygBEy8GMCTwAGJga84JwKbdDq0gYcN2wF3
pxpyPP9lE0o8jZLGRTdfGRHqmKY42tscNr4I2AtG0k8flz6X/4jwdmLuFs6CH36f
mI1LcKhaVAqpCfPwgUYvRRgI76MzoP2l8a6d+hVRJK8E4drj2b03S+BRd3EF1iY+
4j9NFmy0TXRFmY2FMPDRQjFD0dxCR6Fze2r7xAYVpFTabYuEHZpE246Efg/31sgv
fHdb+r7NjcxNhRfwOrGncAEfV1r9lYXPM+5tUChTltT1om+hjZQcUOLbJ5ct07vR
E5hLv2xna5t9sxvNTt2HZEwOeuZtNX2ETtFYyJbol8MSDQpH/YyfJE7M4d5gpq9R
pCoWrWj5jZHy9AZTWG1Az9dYoxRxq+Q5YfRGMZlBAM4RxYhRIgPXYWy8iikLtdpR
fLCooCuJbYVBtPmXrkquz40lnfs27V3njXSA3r5ik7OQi9X5NgvreFBPiYNeXLth
V6eraOQGmbh4dPAb7QXbCxVlP8vj0Cewrjnri2JczmFpk2lrE1RVLBrMhaJiBN2H
5nbb4J6XGV3CTZ/L/2Ownr7ifqLPC0WVYeGdvsswER97ocGSj8eiqg7rp+D9H66F
eFbeZM3GJRxX8Z/3w0at0jZnY/nak5GfKW/DmWmHtka8I4hYgbZ86VdlGFpSZrSe
u8cxmwWsbEKr9KT53Mkp/79o/PaxRdhM/MdoAmBeeOwzD3+P69n/DbYw/Y0Ftotp
4dxdOG/0mTPkCzscJjDJcIWGwUnnoHdsC8w4UQcOoT2DO4whwIag+dWAIBZNViRU
aEUh3ocbLuXFj5V3LEKYhiM4g/WN5Z6ZhgnaubLXgkchrA3aerkY8eH6H/qjRVlu
EYKnjAxYEl81z7Hd3tkjK1nL9UvXLYvOWVeqFohtQTgx/PYnCnUEKL9m9kNgfgcG
bK7rhQBbqJkOgSb6EctouOqkLCpmnWT4MBsNDqEJ8qW7Sq1Pqn7reKxMaQWDD3yX
B0uoTpwRDh8NXdLEbm+reqtzAhJJ+DUjeAqBMCFH+HgCM6YusevkZVQz8AFzWT/5
GLJ0/UWF3X8hz+xFUgdVZcm6xWfQq8aar/wAlq50WL3ZTUvsQEDADs9FmBTc/zZJ
6Ffw2fGzXsI7ye9eBnXMwYaUez3tyl6pu3/pyA69scYmUBlVOoEQrt+wXabL2Ig1
ztIWwyhbt/357VxfqIZfOCB8HRxvkuq4ABTFJOUsH4QEpsfdr+1rrsZRwoMxX/Nr
tqUty2lXJyaaQBTQ8ScD9Ugahn78ABeuHkYkTEGPVwkvmWpTpxikU3IuPNDuOass
BDnRWathn6qNYXed70lzY4ODMs7+7dlziYYAA6Jtn2Ytg9nYIchGfu6Z31j6OhB8
btx2btVAywIOQ9telkBpDF92EBzHerB8JzauuLsUvteoLXleOGEMvCh+q4bk8Bl/
JI8fF+wukX+XiXuMCh0OpDVCBf3ZNdt+lpS7NEYGrVyL4u/xbxMMNn14pwxPLlbF
GMjGphKjEZYMbGZenbYpamrw1rvs+65EP++a6D2kJSmP8AOMzuECSIwWcYmQNiRZ
sGNJzxlrKMQkfgga7rNiQONOuQO3g8trmGSuIspk9EFJ1AFe/YNszH35Ozt2pRM9
K2W3kl2g/JhPo8Ac8BKd4noFJdENFnCFIvuoi7abFMjiJzzba5senPfcznGckUOF
KBZA36LG9lt5RQtEQI5wB6Lis86578MF0PhUwqowuBAj0mTT/HS+WSLKAPC+mLPs
4vB2EERpJv1kokSKbAIY0GJ+Nm8YF4hr1S2BGzDu9UuOFGD4xgiyNeproFBYTE2Z
/cv6bXA7638flBOgSdPdvd4jrIBQ60BwMHxvD/syTqLV5p7uOorqMUUe/kGAc7y5
2S1gCYZhBMxoy+NMKEYbnf6jCDB6i6UTWdn9zwA+2UGCWJYA9wt38pe18b/qvzl7
zdCf0ofoPkWk1Hq9kiwkbjIb2gcStK+ZzEwtZDsFGOjTkIRQgZytSNcP9SkHnHsk
sIxX7WdgE+9yETZmKeMqtt6I2YnYUEGfO8tANHGlPwc8tArKuLeZVEkWFvqyp0lZ
ODkgJHrtcErdli+FOHJXZf+2+aBb7bUowZ1KnDa5Q4MtMCEDvx12UTm9CThu0UJG
QyVefX/Gsqqly+IcFwft7lgdOCyOrkPvo4lbpYSl156i3AUy03N348r+m8+eGhHM
B6xR7ZkPPRJ0ts9Tl14Q85/BsNzRb8dWz1n0ivEEvB55B4pZoPoxxeKGNznwc6LA
iIq7Q6x7ekrM4XKj3JYqlb+7y4kFMMhiJk4vibPmXH3gdAgmIujEUIBVDJ11F2Vm
j5Pp5Q883/QzC5t5CMXDopdd1ydpTTFeH9ObA/qiTlTCJviUdlUK0ThpiA/9qEJq
PUI6VhPwYdMa5ix8LdbSGpF0TSCdRO5GtAx6AV/gGTL586usndYsps0ZdLFc2bCl
ERbeYQjYRVNiB33cQB26BpCLM8G4CuTTvG7HysRdJgx4tUBhwSz9FgzmvW6fv+uQ
KyMWIGJ/3xy6TLcARgQxIk9K0Jm8mN/x+IFZtO9PY2h75QvlshV3W9Y3haqSLOTI
Lcx5PLLh2+vbTN1iP157FOohpuMuzjbdahtHj71JSbt3smULSEmr4A9pgcywgDxS
Yr6KEvR9cybTDkxWlMEcSzA77Ka+zKw4KnOsIoaV6LqEiaCoMb54z/reTGkyY1+o
ab2QJVgeNhLBx7Hnv/PC98+W5y1PBEtmw626nUsuJHvd2qTn1R0R3wsD+6JwF0pv
2DTkBPECfhpmDLY0Ma6NvTfV9YxXdOYiRXxeRDNRafBeXUckUCIgHXnRJ4wBfEAR
oAnXYLqmzuBgSppsFwseaGPrdLWfqvP3t7XIQB6AhH8UHK2g3bdu5HbnVw0EGYQS
1yh6Kujf4X0oSTH2b/EX7L17pKrvLR5CuF53roYsD03MDVo2qwi6qbjFdrmJ5hX9
YGBsp+KzZc+2pbXj2CXohODVuikNMjTR9bIkWROM6pBeuoMYCOhz2SUDnlPTCEGA
SoBM/VStqagF4KahcxYRAS5I4QqxbnB9DbH0RXudXNeZJ+4NnMb2mpF1kGMGBamE
G2BdTe41Jk4r9a1NipfbbKwPLY8V2+eLTd9ih46jvbE/eog+u4y7/ld24B3fb4Fg
5dGrGUCmsjjwkbs4GoLUikJf5w4AbYdOl01nhEr3cDgrhD2QzjnyJBzRUwxGlJ+c
yrmkFvXJqREOOd806F5cqo57xRnqeIqpNQ3M1R1kXtbfhVOnCGBGEPwikMFphFjd
Xx7SUwIL5RzEXplGBwQ32iQhDq0ui5hoTI1qkAZlCOcm6UfZ8o/E0MmOqWLUfi/k
5/SEz2lxdL0n2vTRVEMSpK96BYv7iBfRDVQxri2uUkLW+2LMcArgZHIij9TVEm9Q
EcO3ZDhyPbaG5so8/E/8jz1mRJhNyY2IuSA8bl2ylMfQ7odobeCPAX99ViE9KCF1
EMQp3tZhRiPX+CXqgu8Gc9PqzcYXLVxHkcrm45DzVJ2YlwldEyO1c9/d5gHJ0oyN
SSCUrVJpyjw8TMzbhKFXih/aGsngYmWbN1a1cicNsitI0quh3P9d2uYWGHVhusNV
XEoEEbMSBQyefPuS4mIXokSgID53bP23mpdiOg5ctoYmgBfZoncs4suM15tZ+aoJ
5G5l8ad+lDuwFYuKFXQoectxGaEfTv50swyeE/fmApZiDpJYkoP9cTZI8rbJ5LkC
Ma8yE8pm+6RzRcdgCV+iY4fe7zwrgGjk6hjdz+Nd0xTGy6OKKDsCmpcb3y2beX4d
lZTnP9xin3hQBjX0FcEBrbFsXFu88I8dW7jjf0i5RDtZae+FhX2t5HmyAhVWGsXb
mRDEs0oJlHO7CfvAWak/yPTEdMBDuiG+RUZ6ls6OudQReF8/uaXVeCV/uTdocmoF
3wkBcmYwJvrdKJuqG75nzaJsw6cW9AwFjZoilL6QjmzjjzDUokGXtZH/oz1hx0yE
1fGH02/WasBqxQEk+ojM7qRO5UKujS5hKNnSSDQLLwCeg7JGRgpEGe/9iq3NmzNI
XJQdhObf/6O0w0TlMgy6e5iEF9VIb8Ndp54G78HA8GKB1ScU66/smW2wQH+U8VbN
nWNJJQa/XxUPDwrNVyQC+40AphVIh7Btj7IyUJMLtFNiNJV/c1/yP4UcfIseB+1G
oqraJwqqBbPjZgPkU+aRaQuhwSU2PXu/sN8wkysXswX3XipAjdKIKLs3fD6D04l3
uM2g3xcPr6S+jc2Q4E0NjRADy/j5TuDMgkHJ4CxuBmpWUmYJmFIe39T6gtgi1Olt
LkwSed59//uXtDhXjAffgajTrGkwb949SDfTDlsboHYzexYLTeV57rYV7avRc5c4
35WkHwm/7Me0jrlzdAI4g0tQ0d1dAyRwVd3h9FPJhsMy4zXWHiKcLSkWtXI0SpAn
/rzqBVnVFI9F+vqkwb9Ad7SNSeZFtM87Of7McoEMCLhXfFy08m92eGq2jCP2BqLm
zZDf1n2WF5+4nhGiEm53W22G8qUSIgX7sV5B/3l1VWN5uLwmFw6eGhqXTQ+83/e6
5D0l1wlNhvk48Vhz4Wrnua79KF/rvk+9QXLob+SRHS+Y4tWdtFbmtP/G2cqp+wun
ZPMQecDHGn+1xGgI5+omyfA/+t8k5KYqVsq0qzq2KHfP06ZEnP7GiqHz3otSKfBo
jGku14Xs56O6er2ei2tQJ4E1qI9rk1M7BN6ssS5UDbxsDdXimVJxhQpqNcntquFL
t4FQXwDacyVQ4cLQiWTuxGca533sGEVY5NSBMBo/SIruxkziGNAuynLYVh90PVAR
alKPT5ygDftqQvMEV/alAZ0N0N6UcIFdmqnxWZHhvFBCNEl2hfWo7EN+k/m1bUs/
aUFaHxWeG4wDlORnWwf4sVDxyuljfNxB9pWmGGrQpjaeS6q1r2RxmB6YlF03Lf0o
d9eTBeJhBk1ETyLOtpl7fvhPsqUAAXb8l7eIbti8wT1hs+8gIBSNnGTQ4/q4XdoV
L10DZ3l1WE6Lu81ZSHNOmCNZJtqZ8vRL0pOvSyr19LH79IjLmGbUOcJVWf4ZwhPn
xZ+Y8QT8bGmCkv2WYcAzkwP0SRpoNIOV+jpTyKhrU3COf8dOtuQzDDSgCAQt6SX6
IBfHygn5lqIRWmRDy3cgyIUiFcTYik5E5IPUEEvvUZvbk1Xuwm7z0s4fcUsvzatb
wB6ev5yXieJN1bIKWUau39+cotlF8i3lK24PfRK+hbNW8P9pmXiPRPehPd0p4jAG
cJBSeJH9ULtjcGSzedqkS3jalPWxzgpwMopuxmEIsK/6XkeazQkcjVmf5lbQpNQM
OvD71iJYJwkfRny3AQpZzZKGgKxO9sr+kuO6edo0FAftRfHeb/r6FDUn2a7ShBuv
4PcYUTs2bbTs1/OuzHi7IBD2qkZn6Zeo0bF88zlPkfQT6iVSVyaS/i/Wa7grNg2w
43mLUG9MylWrC/I4nloQXCwj82xZc7gnyWUznBNte97zQrVwyGZvABLuRTKH+Qe6
/qcjBG51taLjDBBEhGEKeEqIyrQrb9cYTLKhBlP2WCk5IoeCKpayFomYdMxU1iq6
2wPXUWrgxgTf4FDqDu/FYuIDLHdHX1IVmXSn5cAnTrBXlqVV/23jO1gkRtnS39ou
fkvEKmcmFfehLjl3L0irvK8wot0XzOAplueHe3FVNzvrDmvQttu6pCFigBUoa+8C
YZczQ3xBXBUF0f9yZ+NYApXSpOxjDlqtPtmApDIJaJwMAv6ovfOh5YT0xupm3uhG
3HRdEoNYXmA4yHeprSq83Xa/ilaEhiz2OQst2ShsB/FzXMcshGCX0+J9SraonrPc
D+lC3jJkwy3GnCZjmL6sqHNtDBK69o4e5cC7BH3PR4lotl/7KmLGAZ74aoNvSzZ0
VPV5Bcz9wKATgQ01t2+3teotDshtCRU5ot2B2pqOUfwZZmqZEVlQrDHYcOscob7m
hwkbKJis6rRPX/pPc5k0HC3Cw9HT68dBIFaZGCWbFDR1TAxpgDTWy5nM5IG5HKp5
5tbRVVYoWS1+KZbgtWRxw4QHAULm29m4dZf2Ymv/kdmtnq48V3xFYbyLhoLdRaKg
Zf6PX34G4+2paSI1Ut5S9OxOt6384RBFVmTuDmzl1MDZ7fi+DYaNRpdMT3MYneMw
D0c3zpSqnWdQ/6TPgIrRggGj2k1nZB/d3NNpBKucsqJlrQtGXLN/dhG4q0LG+tYf
EoN70CUMJiJiCS8XbIyVJNRcXuB+jCkZLcv8XXR9jKRiXkDGVZ7K51TItns/MbrR
leUDGNRRYpj3FRrtk5ClmYzQz+ZS+2E4rZTYAyDwpMionl7rPaCexOwtG6BpxZfa
1XkXz7gZ6JjturKkAHg1iucKxgndKQYcKfXWP+ywCeXctDUUrizdA0PhcHQgVfZZ
ACxx1avXwRRqOgw3tukRSRIso73g/E5TepDptAMLNf73edZpLo5urSPKiIwGXyMl
A4tBvEWAlXKPtcQdv9WkyqD5E0bjKLuMD3CCgmJP6JeYS/VURfrNIvwr2epsSa+7
/f9KuYmhGZqP94e9lZ+xiIphYvCL/YfiXOoiFS0i13Q2qUSa384CedfUsGIm5lvz
yhoR1LMFUsW10XHsfA0xLr7cSbylBf9rsghTO7neqJpyEezKmraGX8xfUGESkr+R
INwHXrPZmGCcbVo5l4foafgzSJbUUTDmTmPHH21ygtDNMp98Ed7uSJQFuSEfv0w2
PC71C6ttyVChPWEwvK3rRAg2/f2jclWE7H+zVLCgcj8RaOfRcepEPuhDVjkhEPqk
fJ6bi2B9TC2NDDDOBwQYvShsNP8Z4Nqsax5Yc953hvoTzVySKPsBtC2SZAYEO7Y7
Btsk7yCISA5in0ffKo+KOnIj1XWWDpizAYvR8OgfzJVz7I31ik6NoDeZQ8UuvuvH
uMRN04WUg6jWklTmbSCbd0c45ASjBrlN1cMfCpqh5BbqzefcA5KNf4Lda4a0wWlx
BDSmvnAowJmmRqrgUkGo/hFp8Bj+f9piV41Iu/0b7Kk1qdDS+fVtMqKG0r8bKWOJ
x2d8I4BVJAr+Oh0joBllCWN5DOaGRnw57jjqBH70PLlgCOlJ2LRmvezsdhVJ4qZC
A54L4sNcDZvTSvnlTcULxBA1L7TM4kgnq7rm7KuH7J+5lRUsgJTrqk3lTVjqQGR6
cTPO/s2Q/9XBZ4o7on2ndFPL05LnAlY92rPdPhdPl4rFb/KQN+2QdMEmmrat2skE
RYzXihkZXg6H5Ft29GZTdJEhZBaqplO2gfQ6RwBALW+M7LbNRCLbiMqFuFCkMnM0
HmseD59KLHiLKPpMUyq5AJgYlJtmHN6JfnA0xn3MtvdMcIOKRBarm85sFhBLAKNN
eLX6N0JPncS2QMxxwY4W7n3ZFlZ03WZjzJOvQO+WkstolApSDkmfTBht0XYFt9PB
UZ9g9T58Iz0rihZ9eeU3HFR8Wt+grwKtCkP+t/6mH9G++JPJwXd8mXzA2lJVw2NN
vhoKCvgrgf23EW9uIXd36kOFIHluQZtUc4EyXyDSkgEmq9Qc9Zx44KtEdn5j7aLW
jxrhnRmg1tQigoUxSvqIlUgBanjqw79LpBgtLhl1JO09d7WLH4oaSaRHvbHxS1Ya
F1iiwb0S1ybKEQh+zWGWcW9U8jdYampRh1XHsSAT55Bc+sgWomvOXmrOyeZPYWJy
Al+FuiafShj2RX0ePbGCAgbGoSV1zFTcNd7JyATZOUqk+z1Th+uvPyJr/AeFs8x8
DZqgVyCuuFTPbeRS/j7FzX5tqpvGYhrSyKOJ7ID7suuDcc3vh3EZLKuatYwuMd3y
tpD8WkLWHLA0QAXZv2P+uclmc1xXnUGi2BDPvSSHPSm/lNam4On8IZpSSh6Vnqdf
wBrtFg5aCLaaOEBgtT02GhtaIpj8QoDIGszJD7+rALaG2Ed/xgDk2V4hHFFHpbk3
7MyPhq7VylPkJILuug1hT7UMWJ1bFeRAuCxSoHwlPrlVjq+RRn7Lu4albOLyklBE
cQhMMAfNgUUmr8YcCSzaVKEHZBI6F0ffVBSFAPSzgRR/vJL4oZFFsVjy5ALj/38l
xFy15dkkVjoTuRryMK+yx6HxYCoTyXXgmHoQhpSAqod6M3zumn6/HgTlECYI5uVj
uLxczdRLR2jtOo7m9MfzdP4cPeFikflcjtez3mWutWYZ/l47Vt7d0D+bpYNfCaLs
3RgpgYBFZn+/dsoMBuPtAtr3Tl8avRGLj0xGXdZ08QFkPOxwfQhCXYQzjFcvh2MJ
Hhl7Qz8mANeUFe4haYZA5OXe8N0lNPQcSYgdusFhkf8py6PS2hIQGLCcqdARxm9c
WKj+W1M43cWM/UulKWDcvR4VFfl2GPAgarJUshQkgByygheMfBQgMCpI8lMg/mIM

`pragma protect end_protected

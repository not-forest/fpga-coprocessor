// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
L94OLCXA/9jliuU9tqSlsqpbwkk2AFoWElN2rQx696zvD1pDbbuO/P1MbM2gOpVq
Ge9MAT1DRXpnkKsdy2qAi0zU1ZUq4bies9tSd7HumpKJo1NK78pseyD8FU4f82pd
lpQ7kJRmaLzwrSvnRYbNaRZw4gzmlfZmX3Qh8FTLIaTL9ifqColHPwwHpZ0HRrHi
XfyvUf8tDHB9bmgZkK2Q8s0lwZY+f0Sls1srjc5lMvons0+Hgr7VIQI07k/ZyaGD
vkVdnk4IqzDy2uQLvjuP5nspbb1QBcB900ebRtDGN8Bbswfkx4lGxT2DVOiC/qVL
v67V/afLI6eZMEZIb42P2A==
//pragma protect end_key_block
//pragma protect digest_block
InBgMuELCCI1ZXTbiFlTa02FCfU=
//pragma protect end_digest_block
//pragma protect data_block
iC704vCtDz0YO2BwfR7APV+Vm6nEHAHUAhgNu3EfTwPL6s/o9/IP5Pxa/RFLgv3N
NkIXQ2E3aL3TvXhI2jEZ75x7O51yIVcqgLdn3SMgOkZT9WmjgysA86DAW27Gc0sd
E5Hnc69YXPzTweit8/I86lN55L3Ivh4xc4ZY2n9ISdxXCoy51ObVlnuziumRURnV
AznBsgTZMvbnFKj5ci1nRZeEnRgCTZQ90LzvT4lzEVgWLwAmaJOvUy+crpqPDoSs
9aIGUYJiTFCoDbyhUXmFx1Wvvb4qTTq1fei7o4DhYSgDuhUYckOnsjSD0YpnZqFJ
CP4NTLy8QyWqK17M0+QuMAtNc3LzCy6p3ySKvXa980s6RntIyxx4fhuJuE3Uyutm
Pku4pLKQiipVWzeqs9pbIqJcoMuFW5SN3Dozdga7D7T96zeVpsnZ7+OqsMU9BUEr
lPOudeWpECOvnGWrJX9B7xfdNYEUbpKDG6Hppn4qA0WgVcsnGj6QSk5pQboUdyu0
GATwl0nJYxVlfqFP01d2wPlD0tLaR/e/JQwill+bMfuUKrx5aF8ZvlzJz8WjDmSK
kSL//JhPSQfsTj3nwBbIYuB86Qw9KFMscDMfY2OVLbfnk8ihdWjNXf7nkhiq5E+Q
/vi+TjY05J9ljWwbFSwxdv2x93/MBUcGv66mjG3O57sGhPfnr03OyeoN0/aFloht
JpMIEZl8XOJ8ZLrWzU0dK/J2Llqtx8T1/mIyhSkbcyz6jKdyo7d/Iyg6FGGfJOge
XHUJPOclisyg7ddNRNcashfP29ksSaAtRaiqju8ArS1pXnWkhEiidfznTS6FxieP
63XS1LZkrT35XFwGbrGoXSwKwB2WZ4kXLfemBpXXYW3IOHkWUY+KhdCjkIkltvcS
SZ3KNAx00v+TGUNohi/QsaYJoSSIUwc/gQgSC2oXdj5GrXhydrzwrEb4hbX/LLTQ
fnhPzr8oAWIy0N2tgGrHbi0+Z1jhp2aLnkgLNsDzglUc/2aHFpKNTN1SqJCHhELC
f0CofyOs9F0mU5lRwQLh4/Qwqa+pBtJE79kwgKRQtuj+tr+EvLyEWHeBPdEPUX6m
FLj7s85T/+V4lSTOsFIi15YFX1dBjjlifVZCdcgo8ZHQj4VUYc8HqAT1B6lvsqIc
+qXmzauD7eFNyXlh3S5QRqaBH56Ysu2X3ULkwRkD12Oq4w6UJzciSdHU2JQ4iE61
B6ZMst6rTHbDJ2FZy/jsJARwoEzYqgKNxdCN7UAYseLWrHv3UStmzqt+nkL5bsUT
5GaOAIHeEnJ4UgRMEwF3BrGRySgMv9xNAmdUhjDgstTvS6I8GbXweSlGsPLJBVsJ
w6MQkOf2izi3Axey9FPhzjjgeqoiWwZAJ/aE6Qqq119bMVjs+poLwKzanOa9IiA9
qkXOntJcHLCSQm0beH+I7lELQRaeRrcrmQNETW1kPtmYLOJ7jVKcOlUB8ZJZoHk6
qU/sja30K3aEK8no04bVm868cmzNMY80j8DXqWmEOXQxG9FxdRmyaYGcYbFe/tIi
8eCMQ/qG/JIG6VqH16DRLV0F7bAe/YXYBMhD32Z/TNssfCSnzg5tbvwKcleKjQa6
elBI6u9HRV8TeOvKboTYTsdgFH0oJsbmTexlkOi6WgH2ecgdR4l/gtQvvd9ejIdM
sGp0Om/ArnkwevFD5AMIeCEX3l+Fc9UZUfC0V4f29jCJvp3rrGrwnh+9ttQxd7fC
cF57CCoGcrvIhfTzTuFN5Z9xA7ANpCy+gnvpRCsCqU9gQRbJqXGCqccRunMbwu2B
nGJm1aEwULAMxcAKonluLxlFplD6K1wMqXVakEG2jq7ve4Jjsmwgg8E03+gGWr0g
c6Yh2NQZ197NHr/7qU8ROStcJttKDiY9jlXuN/MffdLIIwZtIQkz/uiGChc2RgTW
yR/zAL8qD5kk+SOE19/RQcT5ouAG9WgsZYYNLkWxEprGlch98qfiibKLul/q3mY/
Sqa5ATFtvWvTqMZSulOV9mQOcqEJP1pNAxsEt76tlLwjQU2qzYnnbpRK/7Sdm0+s
1fnRmhrB97tcOq/e9WpVWvTzNbcGOjYPA3brZXP3L1zX0+S0XK+Hivg88y3Xu9Zh
lPusuwz3PIQL9G3ZRHXYiuVDTGYzQP7Ms0z5/KgN5HLmNcHTWjJpww/qp9gCtLLB
IeEaT5L7WBrI99jepody8QZoLZQ5khIXZ4QVl8Wi9eNed7cWgvHXrCEX+/PM1wf7
+zEyCjs2WMrGKn0sXg69rB6j6zYqB6urNq4Op7FB51nIvs4Sm64oysXYXDm+i7pB
cAwKJXfEB3+CxDfbQZB4W6KNmFq8nMvNtRBnvj/DtZFn7LacjycB/LrQ7VR7GL6f
3yCPAfsosfdFLNwB2qhQWF3ESqdrgBRb06wlBXMIyGlOiwed+PuYICVj43tkJl/b
KIjCD13Ymwe/GzipiaCwDp6rF1rySQMV19s3arhBwsxMLIgPxnhqnC3jsf2d9EBI
Jw+5pZgQ9I9tTho3mhl1n2CuUy530FedYGoYbwKsONaRbzEqB0MRQyf+VS4Uwbtj
RsoVOYr1pCmbrxup9n/N4cCJZxThOSWkIbBeTlnyggLyr4itjXHE087lFl7YrQ4T
34xQbzHio4pdq7xlM9vjK391Lv6T5TMAUZLG/Qlf6sBkoTFdlGHw+mamyfVcHL5i
a9x0xUzSIZYVF/ecOnmI+HK47v4um2Jpu6jYzeZnKXEsqHvEurZVeqDABxHBW4EQ
JP3DKe9fv6NxIhiBLMAHrndoDOBgPF1Di/dXZTqLMQ3Y18FuoFNrsmAhc7R59/J+
AtO4yNALHaW7c4fiYocBj5zUg//sDc0rI5406ARdSDRzG4TbSZ4igrrPzkmjkhwz
cEP+s75T+ki0B+OnJ9H+g9P6CBziLbTb3RAyT82HWZ/4SYYFdQDpwEXGHA3VPWaZ
5Rjr/nmmUyoJNz8NPwD5Sj7GivugHpm4cmMR9yMV8oQyJU7XaOR82JRU5gCGjvU6
v1nDVxGiebr/VOFay7SU7507782uaGU0kCoqQn3fxg9CrfXgyemBegh4GEyhqrce
DaFnYqZJTOqcoi+rFsTguUdTYsweF5nhg9PZ7zKvJsWtlGM6FWQNWPxNOsrPM8MO
cLWIqyEiCQRmWdnxkolsWA+uPSW+hUYt8Gk+HnEap/WMzvOitKE1D3OPXPWcY3t7
eZW6o1OmqV3BnOhu8LqWq5r61HDKlwGq+OHsmZHE4mJ3jxeoHeVq2moTf/fEINg+
E8MHpjoMZPyg25nvKuOqi7ByCzkF2p2wDNgqbMDoYmDAyk/+WuqLjvUsPP5zIBr0
yLRB2EfgnoE8ChaPFI2I6Q1uCl+r+5xzeD2EgeVXWKkl3kBc+Qi+ZIkBefd9FEbp
xG4iOzPS1hpbdv+LGSlRKZJsEBE35HvIUvqsfgug41l8UEEk9u1OSiCR44Fw0cRj
zlRRBGf1fUErCxehmcKsvGb3ahHXiJffKb2dZ3c512tSErm73Poe7BJnFxNCGOAJ
2lRyduR4VCbyiRk6itccf5KfTyQ7hNC2UESp21B2HLgOhwMdXOQqXJ8I6kzSPTqa
hpRo+veqqVxKHwESPboooTvGwPpCIcf696cpUyxeFTQdngIpIuOmAiJbuQ1/OWC6
rN0C2pGwsfhM3ifx4mHf0EaVarEkpKvPuD/nLhXYRp3q8SbmNeuvl4XExiKb0aUH
jef/pS9gRJmFGrMqR3HEttaGcCAXGzmj+AMp+QuO8iVc0hfC0O8GahGFKDD76XM7
hAxtnc4RxzAGZZAbvkNKkJjM4C/hMxg5xDm8vH0HDUdGRB6GvrUfWXyMix0UDVak
RH36nG0jptrv0d0PZTj7mIMF9kOAqb3FjlQgpIR183Wl8Txu867KtbbODhlneSMQ
m/EF1xpU/8AUhP9nDQw4fXMguPyd1/tygfjKVSJ/6KqQ1RIOnYhTbEn34I3voX2D
ZK0XpBlt1zcaWyYpaPGIiBEpeJZjOMBOwM48GoaJaCR03YfYKMBUWHCa8yRiFQrK
jCtCgyMymairlz8itBH2Uyg6vJ1FResyrDlQ3rrjx6JCT81QRgIVpu1wFoxBlGhz
dbjzl+vC7gTgh6TGxVXndf2byF5nCoOyRHezc5jKS+vjwa31ZLiL/sTSMg7xA4Ic
0XUj9faC8RPIM35VsIe7f5xUGl8patkXntE/huykIHDaF5tWbkk4zATdT30tw3+w
69kjqijm/OWpo5jTc+4K915G5/ZpSRosrqkxcj5kYkVvkN1OrmTbPIiCflhQopAs
EqOjbkVjImaid2ORL0NAaWcdcRi4xgWqQ19K5tWty1PehLVETcHuzC/XnHeucC5N
tZxvvpNLcBUc6hZ/VHipO3AgpfwA1IEjpwvZ13usjk4VUAEHG8+dL3/NPGBcJ5Vz
nKWTnoP86UGqbQK6NqwwPxjpWN9F/i5xdhCa7HKI9yPfhOYGMq12TqfLaH/qVPG8
50YdquA2pIEOT5L05Yo5HSZBKnXOfBsaqdZ7aT547OG3LuTRWHCXHglvjBMV1GRZ
+0mtsWahIcilHPlnGiE10rKe0AjQd5prBVnIdtS3WlEcJgvNhOy7B7LaYjmI5xDg
by/vcuzzgnEtWkfmb80Y9RDP904SUyMgXdagMBoV3V3jv7YONVadV/cbS6ubk3++
O+efIO42YBsVyCNWyBh9eml/UCugkq6YqbyKCauCJWcMxp0Ixm3sEw2c8+fQ4ctx
DdEy1tO7UhHU/J3RlEVb8Jr68NHSaqqLsXrBhwwAE6OhRRe7OyY0jz6zNxc8SZQ0
0cfXz/uo3WY68Jo9/0Io35ZJv49NkHWKcJnzjZFXjq7X2/jjh7gdPbgxKgU54aDF
GPmMRPZJYuFg9vSWZIXofMBdf4oUc+++JIinCvIDym4i7dlFtDM0klcpQ7Of+xhi
jmXVN6Xl5x0Q/zkywOF0k2df4H8rJm2kL+tlOzqIfqXWRQcn7flUQ6Ew9tpMi4Bg
wqgfUr0bDF9NeGVWtadz9PvjDIZsCwno8ty+h7cy8Rrk5PwB2QkOcNrBkd/3khO2
AKK1CKp21syYJTdgrOvI3bJiq2KOeQe0FbpzPjbajaISgKV/ScYegqE/bpd37PbK
Plr3erPRgjQdBHNhnXloboKQAUw3j7h0Lxi5MTj2h8xrbIsC0e6lBLGxqSwe/D/e
4OaDcOV+I/m1rCUF3ut5dkxacqJZvJm5seGiaq6xSSGgOPWFtPiqOx4CExyMNcxF
iBxkHvPMiCxbBJnJ7KLpvVUljt3TEwchlMfLEV9Dva6Ua+lXTHaCRxDFXswZhlf6
Sh1aRGlfqxNGBdEk2MhUYOY/QpWEI5UvTpL1oYeVpHpaDzvN631jzMsPr9cI2nlN
AUdwAUNZ/0m6iKEXSUdMu2q+CReRpCNHEG0qAXom20EQjwBaIzDuZkDn5FucIkkf
TMUupmtwQI1fmB8xSyPGoD08+MxGWJnIcrQcV7XqUSSz0IGNfTmPlJeNmd7CtOEy
k5WZWIAAGctqXX6xs+EinFIw61RiTnyXm43FzrCKEEhS6x1jDPfEMzXqpuHliITJ
Zcmcl4M1orausNrYRiw5CkE2er2xIEcRc1U4kUoya4CJQHdKAgernluQw9AnIT+g
qitXQPI0sXQf7xzkY3Sndgn6IDBFgFSh1oK0tQl4mKKFPEGdzV5j4lh3xtL5RZpj
nlorY9xBRmK2/oL/MysmP0XZKBajmUaCGN2s2346vfmN/L7qAkMi7Lvlpk2C5W4/
b0MBtIOC4ZPE0fayVtlffsKT5K/JdL96yzW6kygmtbajIu5Iq+cvVispZvDedSki
H8/xjmtkFXD200TzNXhDBoB7tDt2tg8RBqodRrzydU0ogzO8kckqf1uwjVsb2sb/
ysb9tNrhBNIbUX8Fm776krL3MJ1vYQDt1zNaNmYs9EeSx/Uum8mUBoOciFXGnVsN
b4ww6+WLPPPDwOJNWGWrRBvqeKmXcy7Dp/ph10R8nJoRncIFQE+zX8hlC5//Pa3q
i/Y8EXEFDJYFto7tdmOPpClkHNSC4KhGYbI5MXICwPZwwi4cJurmbd+PmtT9Wrcw
lwKSUONsS0m+qJ4f3LBXxx3dvxIleWnHCOzuoqTiZyUUYlHxKMLx3yZJvggdNls9
N6nZdxOwTangUPMcWk1qgqx8l+N7Gfd3o1eBZSpsJXuKVZ32ZYSlX1J5xycFeSVy
QgeLEGUyw+eL98l1Zkgl5PHrADl9Uwxtd5/Zb1a7iOWT7HVFGCtBlz8VIv4Cib/D
wjc2Cp1k/GPOr+ShB3bSkjgrvO3Gy+gP1ZH4aSyIf5d4oFJMpgnD+1RfldbKmOj3
ef1V07kvklsFKRV37jttWyGoQv3LxP6qnW2TQ7+97WaPetPybaxmQ04JEivvItVk
A7OyjgwR31XMndQmDHaHZ8z5VQiBpr4UIWS1jeIzLqwWGfqaldYcWQjgPowtQ8fQ
p576s1YhK2a+8Iznrzyypx6To49iu1hc9x9sFpqj+75ONRWB/Q62lZXjsnr94mgq
F9hcSWnhpyGWwDPs52+Mc5nHpaFDMTZPPVQnqazTTgBuH13L1hIXSS2ieuVY9AhK
bJDs2vhbOvvexjf4fklSD+aCZTdQN1URLENmcE2alIFjMgUY4mv1befo9/dCmkjn
9lB6qjMfVVSp1E0ZMETakfv4p3sK8oKoHVSQ5dng/kdNEHW9Gv25f4uMGP2jtLEH
5EZr8ikpp+TDw4ix/3eU10HObVZs/LpgKIIwsupFW2OEndC7jhFzF30D+EDq4ePz
DbHnQUawRlYK+OXi1XzUsIE9CZZswa0aQXACwXlrafyB/O0GViwj+UYqVUao8tEL
L7FIZFwmTBtece7Oz9aCHkF0OE93wrWIlDMOUJRWSsQB9yzcAX+mpx4X2TqyoXtB
vcboqiOHV+92VpxFtClsc9uHyS2uU/a68fge1qm8b0U5EyKKZiX3CWGBZj7oi6yV
UIthygaFjixdj+K7Zb+GVp4bxdyZ69AiyWYwLnr4tGbW7zmfuvoH+DJmYYTvrQ7i
wLo87OGXT5Zcw+5WYfPHZpzR+Qs1pSapI7iNugOH8HIu6mtslrS8FcCnGf8ISkrU
99UmIJf9zTa5krhpFe9EWCn4eyUBRAsIkom+f6ZmRKM973znc5sYGMl3ij4SOeh3
Fcxk91nrO/NETOo0fM1bITQiIiYUwvOAU/qYFJV8GT0GlS+7rZoXYvMHYTEsT4hg
Ar1CWjIqDooaMbngjkV3ZYGgzghWqL8xmvSo6veLeEmE+dpUtIyt0qc3uJnI6GIC
LAFz01jZo+7/JtiISkx0yO8dEkaHVIF5A59mi4fwGdpW/VgBZRqdpPBiaFdV0YJn
KhwIBNifyQz++jW50HVUbjvOQRgqfZapAnfb2voHyScsRiprWjQ+9vYFqp6IoNuY
/HbCVJZPGtygnBF/F6yK11qC2vgQfHwiz/9Vtl/RiKxl16iuvN2Gh3RYtFL8q5yU
sv+ACUirD/CBa/mLvKAqsotfj6klcHMJSMS9tMw37p4zFXNy3efLyi6izSe79Obf
cXFoKf/YoLKilQYTNFeOXjEQs3R3hSYMaJFFlRRV4yNhV1NDBwMbbnJf29kCmZhn
5SnJ3WSXfqzeqbjmVhj4qemj93qBoLTCnSaNSzzSjpv0Ixy+8nVxsYNpVCbB++hA
Xb4olsMsE+lctehU1c8djBCQc6gHx9ZcQxswVOgWZpwYdNJG0NYot+xWLLY7Jfph
Iii/UzPCZvKGa1Glh07nCn+Nzf0h9Uh39odASn1MubqJrLMSKfbCD4n0baxDLIGY
bPX3ki/vUU4AtW/EgtyJ0sn4oNgZGMQWZ/IB3wijyPVKobxmsYc2PaVYCdXog9nZ
pDJx3p6KOuWqBvTaCj6E5EsZiCMu/NBDza7/dWScjRW97qRqIXGOtJIoRrX6jHEz
bpHPEvBgkqeqD2u0zAGh2ySzRN3SCMGmzd+icTGlvn6LJSMYZ0Oi13EnOd7rpq+8
3tUBQuYqqB/mRsAfIWOP/C3uiXdlUt02emQkmw7GhIXd1ISOXBXYaTIX5ksVVA4u
K5Olk1GTO/brxsvZwSuiyTXmkMWqv0WhTpUpeeXw4drfsF+J/NabwPhrehDZeLVf
ckGbg9TiZ46XFLIvuXcy8c7prY4JapAgdpWBmNp4hyOVolAlNdOYbeXkh3W3z9JK
Gj8P9b03LYxzrxpowUexqxwb/CohpGq9LEMIxzJM3UR/FB/6TdP3WR8AL536Cx8p
wOrvjPFdC3AEgCgjjivgQe5PgxnWQQCSVHOOnQaqccKnTn68XIj5Nw57mBis94fl
j7NsR7I/VJ2y1KtgUvhuhFcMPIKM0at8GlWJnRiVhSSC0aV/5aT3RV/S52yIqMtl
nq2hlUpqPFZ43Xs69IslwJloD3WMXMgDzg9VIJAy0z+kzIIJJ/r7IPvUk25CwdYw
eF1VKqqXwvdjs1VSUQNFWw3FPUlqVUQwEj9GdqxpEd5/2+7emvRtmPIZySSBf7aC
9+IuqvSmmnzJDA7tkWwtqPj/KgQZDptG07YbjgmhBa4X4YCo2fzOuRBhguEw/puO
I44QhIh2vA0GXaaNUPhHl4hRQr7OhmgrzGZSsI1BVhhy8/Cu41BLfMYThTbkhrtq
lddo3cn0/z1ecwYM0SPfYro9/PABKcn1tDlbGFZ2eIaojveG1TyVQeVfihfYWlfI
igE8pJS6DrPs6VyoD0DaN2TykfYijE/XPz0f4Ivx7FKj0cejOAZIgu2nVafZ2V71
px/eP5SBdf310lczN9ILjizFBvmfaDQrAfix6D16SaJpxvU5bCveaGUAgP75hplS
ZQ4h2hFg9w9oTL+CFTpHZNtW4NOMEhQQkwq4ibcqLhEjya0b+PdV0lM2vf+UArx5
8deG6aaj0csLrbq6b9hslSqrLnyV/V5HzRuzUy8tv/6MTVBCDLZf9qT36THQqjVW
84lOvBsBNJCf7dMmlHtxDTb0Fbuj0pThIgtt5+N+Ry2tmi8phyAeH8fJFJixxPVa
2H46I3O63XILLKR5XHT1fDIM70RVMbU6Hd3m3y7p9kqx/tr1jIQxkIdpA4ok7Olw
hNHvZJzd7d/4R6XfR1jA2bgu26ZQbri/nVtS1dXJMRvvTALbp4NjQdRSaSRBJDqB
5f5U9bi4cB8nV2N5wAwNxY9MGfXmguPjfeAELggso/wd8j7PMCrVPD+a/j27sJ/m
U9A9OP/Mqu5i0iU/VxMTPc8E+VjOqnwGnJY4VZzetafr104AfDYi2oQmPeTtCTGQ
1MnwJoxLI86UG/d2eq+zAYh7tYhJAFKc9MbDXjtAU5m/BILYZBNxDlNuRF92RWuz
nu4ML+P8zb8FUGDs290aOSFeOmg8q28bm9WncLNl8BzrPXq0VYKXg8Yb0JWnQBSH
J7EdbWcVo3d658yB8Z8vTU0VUfCX0TvH2ughdaKkO/ec+WALPnA4avJ3S8d0+5Jj
PI37Kp7ZAhwsPizH5C7LizTSLEGNrxbGfY3KMTCNeygKhqilpCFwRsPHA43uOkrS
LtFQFhiBRiZE3Y4lIUxqPVO6VZD6vPiUIqSx1BICov6XBfLzj/mjIR46GSjLdf6p
f/vwAVZmupDm+T9Okajno7Y0nPcxFlEjTBuDLuOtyJ+rj2vpRpGZFqJtibzYVJDX
bAE8qyPb3d1jTF8Vrl4WpQqABJm+FcknL/B+cFWRKie/BqIJbdHAXqx04j93fTAl
HPOsJaCUM/Kv0+QoQ3C0tynVLKybtOaLAMC7+XDFwqHZ3wZ4obPHXpTXBkM7GbY3
XuRzlUbv0Qh88ZfkXRFZyBQRh+3cLg2In0Abeh8LYUxRQ2IszFwKo1bsE7Dcyaxr
buVtjigbUK2CHZ1tDyz1JegO9uRQEb/IqDD83alZ8e7jzzeIkgDh0Evu874gw7Y0
AYZBNoHGX2vjvxVqnm6CFJt5H6lPvwQpc7ORMaiQMxvpHhuh9I3iAczPDUDkqt6g
IwPjsfYmlFZ2TIsEQ4Bhtrs7RIWMgPqdin5osLvoNSp5xv2ZiUw0LTk8VRgh/DVQ
m3cyT43l1T97l6OTPCDEaZ6IPXBsSjUkhnFKRhIrGyF6IquZ9LmsQwT1Skz3TL9o
KSXEa9198jKUK2CHO5B6D4AHozKM/339mlfXzvv3cCSV+mXgU9cLcW+laUrOITLK
13PLnmnuSw9j6iRoyANxOwUonZdQY53odpt47PUczoq5XQUtOkQ0mpCgi3yesPfH
zLZsDQZJpAmxQtbFsuYP38/m9dmkoOCohJ90qiBUcWoq5c+y8HaeUPQ/jR3j3tGm
SxAlyj1Cw8WtHz2wCn+d1g3F+OEwB2SNJYu9GFkcm5ZTbAC5xGvhpzn11aArrQB2
t3oLVzO+FqeWpIRTalZy80W+0xanQ0trv8fs+hXWb0wmBRNMsKxWcRKiloHex1Kw
UjsvV416OsEvRDzDtZxBo5DG71GBU+or7HqPzkqkP0NqxuuklAWVZKh4jp3aZ2Jv
zNd5VW5qAm6xzmrZ5OvHM0CLdMLqfoxrG2a9OCuRTKrT36i+DOFU3a2u2UzjNzS8
26u+unGXo0TMMLoDN1BW9RPocvrb/1NnGDg7C43gadv04Wwlw6MRVymSL2P+1DuY
M3JoQavE/gsIl1T4q6skLPYG205vjsLqWwaB7PvvboCv75OjgrDn/WsQu1pYatP7
r6Q4+72xU3xJmcfg+YFWM8FdRCs662OP6k3Ze/iORBDJ+FEmsadgJD9UQJqZkFrJ
m4SMXJZBlGzMwHUzR4iG8hw7N0NEszVRqkFfyvQPpfsTFuJEcW/9OUvNj9y8o25I
XeegQZ7IEi9ufi1YjqcE1MtFl1HL1IIiWCZaVUuZsL9iheFgu+qiF48sJKheSMYS
zIu98Lonh5R1gwvdAFq8BeGFxUQcD5iEZkkklE3V4N4vVx/JLKzQwGjdUtd5MYQr
/37z4z+DDl8glQkR7LBvVi7NxdyCy0KqaS1k5ISlQ7AXutR3wDJyIVeTAWTV7KKT
fMUB/F9WnDMHeYr7RlQ9BLgoKret+YdSBn8xFuuakPllLMx0eL4dVzQq5qqL0eiW
M+S/DGVXwvSdowp4fFCSNvcCFjkCHAxfvIJcY9tw8FsFKnNLxiWZVszgshxAtRoy
pRNWW2UkYPhEGDjCT77IpLDfl52/hKxcol6TB/YC0xVYaOdhVz+gMN6Miqn3+FN7
2B7DVEJdruJFF8qjn5LJ37sGjI0d67EB7bTPFjzrbUu+bnRNozSULTW8AmiARP5k
eBTDYq12EjC5MPBlv/nO9578RT3mhI1DKpZBbGzPe8/VBAD2hMkwq2IBEhtBeuPn
JNQJR6h25QVF+VYX0CfizXsT8XElt79EHfy11xHBqYclNmxCmNQU1t6Onb3VrJ8F
AFOMItInQLmCtKfodVwdvzIn5lQRNsFR2nQrHTj+7pKuPw0z4weObrqiQ2m3p+p3
DjlGCzXnJid3I/tyS1TGIIWd0rq1kVHv48KRlmVbgkSFrQo5J6wGZdaENxaytMBL
hLHGMFPZxQ6WtSdigp5OMmXR2y00/q21Te1c1/5blTsOjWvw2RAj294dy2H4ibdG
8PPf72zrTknKihdvLTaOsm9q+6T9XgM5hsBOG4keAKb/9U9MqUdrxIzNu0cnO8WL
ViLeb0dYMjsOb1lhs1LMcfL8sqkyoefQbF7eS4NIjxTgjsCb17Xko20MEM1+3P6Y
BSQEfDT4hU8sD6PNnDyiS/ZDZCvf8wjDfaa8Fg9Hbff8pQOCwQbhgjYpb0Yxthmf
4QF1NhLnwgJpse+E1n2o6w4qXHB9bfTwReeopXCjup0CUwM/DMPRXpmb9818nSJF
du9eFzDKPUHxuhYm/tM1ffm2XlxUHV9HH0LW9v5UM2v4Y67MWBqYJgvOmcNiizni
qPVUMFfYQhnxSScjiw30EgkBPyTj4aO3iZL8LJvPqc+Z0FU3G4F/DTIlIUIz6dY+
s3H/4mvgggyUAAXEwbHmxPHdxE7FmR/znA178YNblk5Soy7wXqlXZKiZUFksX5ex
6jXbo1Ur7mZ6ti0QNJ7XE7Qw7sONqoPcOmNZnGimHlzTwzHC+3hMpw6L+0aEs4HL
y3NyD0Ki2lj1y9+8jZZl1ZnR0N16G2gcgaxpgfi3OcwtY3sHcKbEd9EcBCZQHF64
pGHm4bVw3FbUElHfmnemJvX/+JHAEWV+hNvtffLN/TBUFBxeBlL7H7NX6qUsQRX/
IedolXL7iD0UPXtgKn30M0qtVO+IPib/rK3TXNIMk40Hpq4m8sNx3WC3iJNoIm7N
fsV/SA087b/PAWXHAswCzDpO1nr4xoTVar9iacyrERr1/Qty9SgYSUJt7LYF2bGo
qj8m/AD+7dUZwZd8/3pHJiRupmE76iEqkHUa+EWGbP76dnZxds2vcoYJ0mup8ALj
2Egwm4CFMCX5sNtq+1TyLS+mBvOeBs9/WMrnsLnRh4Yr3LLDUad587/uJU0eKjmC
rYVRQ+HmBhFiMKAjkLHeMijtXClMxHV5kPJkAfSCYtY+Q/ZWSyjW3OrfZLdKQzVc
lY6LyHcC+fUo+EXXMZVVHlc3sqX3Jzevc9xEqdPyPns/QQR50/3pqu8CN7e3C8IT
MAYk+QWlP3ZnS5oXG8LV01Ugs9PSW3jGkk3ugVcfNua5jvuJh5za8CquFDcq8R7K
sWo5hWh4PdfSxndGhFPu5f3F67A0aZzG4J7QmZ7aPk3OjDbRuD7VNHFCBeJdKOA9
fzXYvWz5Ar+i++lrnje1R8JLXNl8Ao4HAI7zseQE1WXqr0MXWEk82kJeZGB9Tvq7
VvJNcgZgjZhGYru/UqckgkbJ813RshOqEVJZWFhxTa76XjEpRxGK5uUguRL2tkT5
rHJ0nv3SyQBvknoBbI8kO+Oc2lnLY3jiEQfYwifjzetbZF8eNfnuLtvPpP+Hs/r/
YW8bTDaByY8QQtf1no1XoxDao5dVNKnfAHO5paOFpaGjQfGnrZ0ChXvkRyQ55HSv
qcnDndU9KY1aLBh5016fvMJ6MVnWPNkNjslzx4zKOupLGmsqeoz1u/EYhvvebgJs
bFtz19rKnVMvqK5a7sTHa/kzSt7Hpf6kbMjR8pwZ+kcGj2OTtxuL1UwF9CcrGW2d
/gEJYc8XmCrJNnDbvWkQQqFhL2vrtgsPucbWr8KYM6k8+TKch6n79Xm5ZzfpaiYw
K9LG614C/RfuCceKNijbYOuliwcXnUeIipVSLObHohdO1qYYEnmfSYL3IzVNm74V
wJzRJo1RcYnQL/zAuKhVQGliKx5WBe8SbTW5MimFM1lhYjzUS40FCtxJjXy+HBVV
SAJjTXh+VXJ6aqKdRZ9xPb6eompxIY4MGCeTpPDq2ToA0jNKzvhLVueHoaQrQGCH
HCJiyMn9RvlaUEB7xe1iVvjCbOMlo03c12omTmcprMgZTNiwgBvmlZ/syYQsvIEl
j90wbPSNyIQO2wPKMvL72kpwCVdVcsm4GTvW8J4a1H3ONpwqfJqE4cwJJ6RrrSNs
+anerBir30/P1Tlzg+/ClqvNyo6hYOpJOJ4gJrVwwKgwrr+7iLPtpUM6tjeoO/OL
OLQcONtxjfQdtoZofLNqWkij60vVodPnD+ixD5casdJFAv/xMJgld0ddYQVpB9QR
TABFCDOeEvFGswIx8rZXZ9QwMfUUlu7xSMtPDdt1qRBVjpxTfAwsE7Dr8O1Cht27
cb514YBPRLkr5IuEIHO8muEfrmNYTx602pC+o75xFtyW4qnMwu735wozwunMJlwX
zdOJIuOIjET1SH5NITkg6modmkR9iCCymEs3KWgqgah5jwqBCFMWCPXuuKnrmXq+
/D7XicpEQKXEjD4kr0gFxrGRlULGngw5tpB8K+Z/8BEOTo3U4+G1nKNDi1K4XWp5
jF03Bh/nmK7EEGW5fgln2OeYEeOr7+RUkWbBBS51rme3Cj4YFNCYjAYjvxtAOOhz
QrE0+rWmoCnL2cve5hmqk5+SE13dlyEID4dT31sRGNC6P/w9sbwXev0DkJwG8g7U
J5DrmOiXFlRqR2V5kGwi5BQjhFoxsoym44V4/vDWDcQTDwhvO7JULe88oR3rb0wR
Ac/izqH2nBdm5lW2ve96wPl78JK48cfZetiaVr0etWA4W2o10vvWSYrzh40hK+ue
cnsFAdZOKpMeQ6l6gdWq0/iVt//UEzB8M4yvQbYn+qLh3/Qet+lowN6gVf4RhGhL
SyZMTzzw/64fp8ItN11lRZtR82ufPPa6mLtnpGYXDGUq/yI7O3ONK/tH6HHqKCKz
nclTd76xNQ0LXM/Y3ueZVH2KdfgiceVV30Fh+9i89I9e/ciW8fI5XsRsMl9xPMmG
3DUYFPDLlEOqmNv3ixHBKMrjvkYh4/R9pRET//198ASGuxQ8o+uZLZO3as5PPtSl
s2pymEXqtA+u8YNjSGWunDlhAAa5QXHkxeq9iecg3W09tMKSCwVmsig4MvA4Q8zb
Fckqs/HQop1XH1B7eXn57nBXIf3+NzYDa8m53iW8hyt5CO3pSQqI5BjDzJXDf1fB
uz/wJODbkLd2ZDObwDLHtwd0vTWqVfjuFRBf4yVPlGVXVeV9u5jwCE830D1BMBn/
IO5koG9LBDvhLP1Cbvci+Z1txnTtUngAvNwxwPBSGvAWPo8BeVLezsLLmrp07y8B
dGMvsQmQzqQLlJ3+XXoIVBoUmS2OBysbBAHnbBrZQV+CCyz5dEfd8DdBfjT5SKYA
2pFsrGp26jsbuvxEE59WfNtecnK6LGwy72N7NfQ4yy+UEpcSOkgHGxqUNSZIW8Aq
LJkSPS9yIYkKVLHCWooHQA==
//pragma protect end_data_block
//pragma protect digest_block
C20JmWBOLxdcn9yzlMz4iouKRHc=
//pragma protect end_digest_block
//pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
rlBBv6MQ5cUyy+g2DiM3g1mUEkcBzYDX+Cm02/DIxCyE7ySX3OkhZlX4rJy+5sUE7jLVyzq1mG/+
Wx37qTweSAZGpjGvRY0cIT0XTLyYdxu2sEVz8C2c00NXPTvC3SyAB9GiBddgmfPfmqFCXUGYGp/B
gGWOhSLxVvk/oVeqFoXi9PsHK1ApqIgv6sDdeLJTK3LP0lH/Fet2AD02tCEBuhoItjLzsmD7NQxs
UIjJPLnnuE51JTLwKC60Qk8KAZA8vDe2fYaMhCKngmuzR59psgagYq19TOODGDrOU5JS32lQz0SB
NhQ9ToLDf+Ubx4dQKHEZTKTWbZAxpkgD1xvGjA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 3632)
JLsNwagfMaBP/CGBmuE+Mrx97agNfi9WhelhQ6khrPmSrf0KONr37fMEZM0z4PcXuqGS7KKHKqne
ieBsR6KmLmCs+4QFywzBad81bydwKe7sIN7+YeCfRNEMhhnRiEQHkaf7Q86OUnO+rtQkfH0snrVn
zX9TzwtTXmDjFJ1vSXfc6UO8n5lDVmH3yk96wiQjX38EFdkEhIyDl0MU8iXg98caW8rWc2y5J1Xq
3cE80tW/r0XlTsvo53pVLz1EaMjuhBBUVrhwe3cOfEAQsjM9CdCC/sLYJ2MnYG3ox5uqzUR6huj5
wEMiKOzimiP9y+SzO7rNgTqm5pYcj55NEOxN5xh0apAT3wmVXvp9KOzG/DwrLn3YqETVT2pnTjEt
zIiKQio0H9WAKqrPULmVOsmqsN04b1xA0QAaCNWLF9Jue5WqC1T8z4yoA5W1SWNv/Y/3I/xpv9Bb
/L671STWhrmuSjT2kpnELTa04PXbvWEZxbQoNbkmEWFbU8GSqwDU85QRZFw3QQgz7UfGSS0HEe/0
pF09GmfJykUTVUlHD572iz9KKMlX7FgReP6+ZCXaJ4lhhLAdtR+5Bc+Ao7JQ6mgUQLthgal+Xwsr
uCp3/BSIIvjwzY9VLoMrAr8yFz2hz+r42kojeyIKasI/cPK8ILcHqE8O5esptY0ZBsYgWv2Za/iq
nkaFoFVVEOe73gUb0+Iap+Gs6MVU9fhFD0/gIgu063tyNDSSzMNmzxqkjkY2eRV8yMmSP8PKHqE/
9eXn6Z2Dtu8JG4EFlW/FrnhsMoT4jjWGy7u7FfUMY1sfdtOibFtGuSszer/kEiU1/JivgT2hQv2V
7VGXwgxEp7m033lCd+ZplW5L1Yg3Q4Iuzdth6XG+k8CkoWs9a3yM8V8i2X3AL4HH3xC0IkCvXifh
Dw/8ghFXZdJWs8NF1gc4YTEwxLqi1/mjGV/A0nTQNJ5Vj7Pr+pAOy1t4auSRLDw9e8EVcGCI2jYY
kvVWWiMbl6kt0mcN53Q6o0B4fTF2QSpaNkSUespWQqOEjiIcpBxjTuERv3TbkhCJphfcljsJ591e
0I7H+QM88OHpMXTl0O+jB6fko5w7iFLCwHPzj6treq3XZaQ2i1Y+pfILWPj54xv45CrvQ87XI1cj
E3GYUhinrozIzpOlq2XCVbX1DmVAZOcWcMW+tlfpztLVwOvkoeg1Bl2Yt89OJ/pkA80JrvG3cqkJ
Gk8RAjgPLWn6km3tWzvh/Pwj7vh760Sy5JHuUSO98QmF6W+eoYM6SfFrl7aBDwRO84t5+aYKRqi+
bqdRR53frN9ceIrQY/mxAo5dds1YF+tErkjM/bn4sV2+22CSiEeZe/CxRSLFD1ZyiveO6qiYoCM3
Du+m3zFKAwOts/m6gzN1eqMtgs0NL0oIjsGIkXcYD7rO6AJSMIjHP+wgEFcnhH0geK6b7Kl4ZpmV
34GeH+jLtWLWtsOwbqycOxSGsFys/uV0sRXO2GL9m2T9UTGHpl7YslQjwGlZzlcWChgrNpmk6N4O
xxF/dEtRjwdjQOuxr1rREiR9suyljq3i+52TiNmobElRYuUWXzEmmJhdzUuyNm/dyR/F8TyUkRuv
Yy0KMJMpJhGpltXrALDrP6B9Xu+KHkhlBvzeIcXylg7XM9tPHsjkU53edgU3SpD1oRPgQ71ElDhu
mXFYLgFPG/g/yHXaXYS6sCP1t8/V7g9BVZvQ9EQl5Qrs5dqYPCTNmEYvGndfjtd3SLwhMiO41tqa
rrTcjDeYRgUUt/46txstZVq4jFaz3Z745ONbd1MmhKFap/DUPvYiRCgc0vyb5/XUmTqVkEDpDIgi
RGMgMxYnS3i5I5eIim5iBHOZb6RKShm+5T8/Wt3M+qh3uVgL5O8dJifaYcQ64MqJkjkruukYTdBq
tNyPr0cYdw3CMeQ5C1lDHUbgHpriOzE7WPOvVPVJsXholx8fHhwSC8bN3i5qOc1LvIrWYVwo51Ki
iP4q96zYCwSJLMd8G5ysVcyKcOvei/tCxpSzEgasF0hJcLR/esrrEWmjHJnzLfUFg3oMrC8jUz2F
ThgTs5VsRwF76q+JEVoO9XvnhkL84GQNetjYGyKZ/O6LDZx9sboPrhnu8Mh1WwByWcaxPYayXu19
QRLX73raHpb9u63DcypIZzYTgHZ9A2Ep/YW3Qv+33tJGKN1SYW9bMuesbchi+ciK0EfeMSIOJ5zP
Rc7r1SBFnMlTqEsWk8TV2b18Px4iGMmJkeCwBKG7Tw7csVZzYG9W98E3HUIYUAY0DQmm8PsamF9y
Dgi/EWMRfvrht4DpEpMSOlTzwNM6/MBfrcLliVbE/edtCXccJ528JVzf8lZho+AtroIHy4wGwuVF
t83oCs55+Bkug85/iG8NvXqlScSij52F6ogo+IBwkuT0DqyWPrULQjCQWZhYO9y/oT7I0PLwctAC
n1BECfmqUmt6tES7BsEtQ8hVY1oW0D0lJpbHh94Vl2hdWc2C8p18UcA9CR92pbnp2Dgqf1RgzxCd
QvwM+rVG3Ui+NQwotzEpHG1VigVAkp09ZacP0NQy4d3i+EaJggqvaWiU/Xan+7HriWTnKtC0B7oG
P+U6uZpsd2heljtVTFpBcr0vItdEAjaFWiZd2zKxBkmMYug5QhSObhV5Rb3NBQ/SXlKbGC9mNVKn
r0aRxrXPIUKnwwQckaZ0wzLaepca0aGIG//SiGnPXZvvoxYgiqSXF0dH+wTYG9IzjXTRt/bSD6fe
rjVdUF0WtK75BroB8U41xU0Lb7Ob8oQOKZvoLZuB35zNAQkRgO6jCTjNVfL1qe0cfBVC0uGJ3xjd
Tfw3f6v0eDg1bnzYaUbCRVyxudTvDFmMAOaYifusouJtKmzdizelfwQgVTRX4DEPpgHyLQh/w/s8
K4904Q8srhr6+GCpQwnW8DGYT6SyKmbVzKex4h/BW2CUCtVAsxGx3i+smQB+KI5tnC1UAVKiTsuG
wFp42p4oDRsSB5peRC9bhXVUgPnJnN7+aJsLJAqEqL53al4ldhs72Ic+D2ZWAg05ZvVW5Ev/XcLC
v864+3KTEdoPjoBzUfkjzdoB/a1mZo4y/5iHBZvgrQ0hZ2j1A4rxsD58hrBa99b7E1iMowkHKw7t
M8Qxyi2wmn7LfguV+yQ3PRcF67frZs8lOPZcAZopjgXrx8vV8UWH2BNzB5CK8KKtGrAaR8C8oqqv
nlHfsMZMMbo13S2JOLj1LHCITWEyKi/C2sM8cRCo8H33WkGv+aQOjrd0gu78S7iwDz2WzTwbll+Y
t2vyC99j8C2IhK+M4I3UE9yQFEMAuZ2upZkDfN9Yni5E7y/CZq/0Xd0pi9CqgHcAEPH8xpFXZwA/
G1lVOcL1QUOrkZ82+hdZ5kFqqr/FQ3KArZOMDYLPHm6g6fCna7UJbrZTcD0UYmZ4xTqzk4HcOgYz
1wOOXzXwBTad0tdqAKJsribm1NiK+SkahpxjaiK4Mfz6S+6lcpkF5u04IzR3au6IVoMuwUWB1bIP
8jFnUKuR1YtTIFrAvx8NgQOBZ7JPGZsznled4q0irlkg0dJIBdkUmr/lAf4se3GxkUaKLJ6S+rRX
hzpSAMQPhC++uzxYDK2f0WInjZIy1ieRZsBfh5WH896j2wl26BSIe8BHGiB+7RUnzdrpo5IG/4fN
BOVj6gR+uv9LNdb2vkR6FTc4ebddmMzFMuXka/mZzwuETCAYweLQTRE7gmISeYoL8fi9MtB8ghaF
yRW8didK/0GVpbZcg2zBZRb0T6incv2vyaKXARGO46acZkN94WXfrIuogcvsdNNPqVQ37YSe6SL5
wvus/ooYvcdRDaTCDtqmaDId8SueVrnt0XPn5gJ1zM/6lxIzxZAZ5gMJJj8zhgj3jB4ns66sMrKf
cG3JWwFYLbEGX5hd/6DuZIr7fF5JSkTsoCKFfdWHlUyCbyZcT9Lhs5KFLk1ondpU3Y7Vd8gSUTxo
dPqvNJPYicXU/XoPXV4XKcOOfdU3Yj7tDLNkcjsQSy07ptF9q3SOiiFU/CIZfX2YVypuD1zChr3U
Ye1aMuyTXcGird1TVXjirKJlUMf5+dbXbybhDzSjb+t8FuEQ6KZhHb/AnWONdNfgahmcFwDZLgSd
5P6QlQ+jrBUtxpER7NJccHCpr3++VHj6JXUzZ8lhZPU6ePCm1o81H4zu9Ojs82KCTHtWU/QrImY5
YU39sFi4H8k0uZJwluiXoAjjl23a7ZipFjHcLFzXhs62JQCDXBf72wep+ZMpDYCHP6o0yhg4Zu7I
8+XQv3Cakrhrd3wsR7DU5JnTm3EcVoCKEiyhkXa13CDpq3afEekjr1ZYIWyV5Q5is/0tQStIAjUE
NNRXiEVfsnf8wuxczJcL/YPgTM5gEcqZPaUQmr9VwV0e2dLe3iAmFzABMVWqos7XTKsIvZ5Bz7dL
xPryz92raJAj0ZoGdc55qYclzBAWp3ISUgXecBBbPE49sv26mJk5D0cNi2O443zu752SW7q0xQzH
6JnIFYCFs+6Kt1IjeWBWixHCIgdjzlE9CMW6WJoYVdb+y1e+hsWWfhi8S+C4SOAC7jz6faVqQng/
NGSTp8fR3odRgvtkkxtExD9cJotA8ebUCGIPr6dR3tLu9ygvk9Pvs2MtDXpVaP1rAD07kGdXcpD6
yC18b4WhYzo32oeNVCbzW3XG6bvpAWo0jyJMAxlbNw2n1nU0djBxRdbjVzxBPDvUBT3lrh/yXHOO
vSDG/hIhgdE+yifrEt7fysoXrKUD5ClmF0oj9Hb/1KctspskyQtYH7+D7kzMd7lik2i4qcD5+ouh
L6aObi80zE0uvf4Z7bZYle4fv0UXb3G+Yp5TVp302yp5FzrBP4CYyHQ=
`pragma protect end_protected

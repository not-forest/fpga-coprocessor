// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
AGvf8Xucbgh9eppGQILsd9shvUhYTfKgrQdT7vM0Xrr8lpkM3YlyR5GjhX8rqULoApS/1n0YTo94
ZdnD2vve7847i1SRfV1mR/WR9dJa7R8ACpRtyZTnmQGV1pq1I3D/wfm7PYGgcBGrwMKFUPZ05Yka
6ELtRnfTrialdRebtjdEkMvYsipDQmGoHBV74ZMB4YQlljrR8qKY3je+y0ts4MFdVVSDlH77HZCN
J6FJHMDMFiaFK8FHYfFzWDDQhjMbI7SjTFP4zv2UyWAoVrFmP2sn4NzFCJvpTOZ226rJG+xH3AX4
CEGp3jQ+rZpKpp8ubphj0SYVp6i5mFEmeKkIcg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 31296)
1HGXsk5qYaH9ZSd+Q57Ow9OfY1ozP4RcVW40HOpIDcCpx1v92VfbPhcHVcAWzjQIVdpAMwA2RzZF
qzItr0Fb3LZIFz32GDA7qhbCt0CzexB3t24B0g9AXnbjOk/C9rhJ5ciWNZLPx/YSJOpMF9b97Ip3
LDiq2HMZx9OQo2OF0szVspLNmzdXbOuweCVixvGHBgS38woZcdvmk5/qQDwZOjCB5K87RX9EWbG+
EIX3/hXlREtJ96D0nablq5Cb1yuVZLDjzRmtp1077leUymyXtiT/B79elzJFVchzPGAY5Ydpm+9l
miZXRXjTECtXZS5OM1xt0KM5f1uqc8XPM1FGNN+F1eMYLiXXdLMgEpDJYeKtbtOL1CvUWpEc/ovJ
bgqvce9/WkqcB5v2ETWeMRkWtREx0zv7icbb3Y25Ehi0zxUffw0O7gnTBQ/Woy/iQdhMvsieKzvw
J1Agy1YMt6uvMz2pJavRIKGsR8Zfzzh30mMzKuIHJajphE+VdTpO6VPzagkHxY2SaZO+HZeLWh8E
ZBNF9GO+SMLtg4QLb6LNuWq4+k7Py2FZzVaSmG6000mMjfIkBxJRhXJvhVt8HDUHHP3azoxMhAj7
PSSxUoPF9EeKd6sj2oBIXCQo3zUoUOxPNgKxf77d5/7goEeR48LMAri1NiekWBcEiDkCtOGS3+cG
Y32lKYLQ+75bp3jh7qw+0GmMatdbxYvmNqy8vhPZGm++r3E1Nwt7+PADZXk1Zta8+L2pJIVqV7gQ
+ZwAuiEGDYult2y7LznlhmeIqvznCbz/hc/+dpcu+nVbKYS9/aMGcDBikJKc8Brlb66PfVbH+x3h
ni7+EiZBixcLjTGgBdSkGhU0Tt+SFbeylinKQNPbmX/+LVPnC8D/TJz0HWDpmIRUf9cj21IQ1hMH
vHVV/cnp6TeMUD/n+6ZfAmJGrUrtsS2sfmG6rqQVr+UoOdPuRIt2tJXL6Y+idL2vfhLLna8SvF0r
JrHkRsvQdHv9sSCogWRDhoCTnktzbd0QwTLer3yfCRSqr6J4UDHd8i13Inj5sXct2VXXPgWJhwrO
CbUxyNtjK/SOQ+8NdlQAhOuK4BG0JWXMUICogsSDXTzzBFfhGLmFMd92uJp4BDMFab6YVoyBzH0q
BDBK89jwhpmTx8JUuoJz2kfSEXHcfdeuWuIzpLA8m6LCtVdHkKo63/dDxL1rOHDL6aFO0L8Dmzr4
Lvt/aCGhS6gjYb/0GrokR6aQmObSIRMz34O2kN/67qTKkNMXRkSoEH0AJ705K20VYaBSEia9fD+7
/SfgobEpAD1pY4x4FVKo5YZ3qf3RTduybJZm5Ih/eTxrNUK6yslyKNfBCuqRSyGsfLRu4BLZeCjR
/L+4FhPmxStDevuPWfsA4vBmVQnnY7tgp+vPgJLYqgIO6+CfQiJwGnqrNZPJkRCznUb4K61Z/ej1
sXU+9ssbNjXurnlLdHY9FeUXUwUbnZ1+SgOpJ7qPKMUmvQnAGY0S38CSvcBhGxtrX2Nu4JaToA5E
o5lDk3Maq7z+BUi5ljUr1W2ZMufr0vXE2MfYns0baufIJ1Ob2iPH0FDmdYgf9IcodiNQ6zLJC4gT
cWBLsbSTZpGZjmQMENKJE59Ein9+vfdMAcjUYsp6mA+9WpmD+HIuoH99NLPL0UFjQHdbraPOFVcI
toD6iBsTqKxI8ibS8cAw7iNwkbg/Rq841RnFny29Ybzo0eEF7LGCfaXCQ7MmPcgiamxiOnzf29i0
mJbmYybAzC43OH1XF23pVmdkxS7WtdeLI5xiYMTYutaDaYHNPI+/ysNq1wlfSJtcWMtuKNl63Lff
2AZe5aCRg6CR3XJaE3B+wa/W8NLPBSadaAng4MXPfNfayuep2z29ttvMFk8XEZXuQMnPMPtsMCU3
BmTVxsSDMrXX0weUFNWSHJV0r7Q8rRpipuhpl3p50TNNZPRMFZGPOSypTSVN5RCdSTpnkL5ACr9I
kJHtvo9eAEdvyKT7twZ2z5ID4mS6XKIC8XU67byYsn9WXAx8VfKkuxJBMuW3jElQiK0sIfKL7YS+
JmPpxV90Mu8Tl13QgniSUP3naX20Ko6LikbcN6iFDUiyROL4V6YpzU+JTYRv3ewx8nxcSTHxXklS
umPzHsIdBaSz+SWGTtQeHRK6jHXF2P6nxY7spZgF8kqY59edR+SuQwXoNIxGcjCSNriybcO5OKY6
jsFqyh06z4T30N0ZDPhu/N2MlDCiWC3F85CeU8YjO+6q86BfbqOZkpF1dK5qOf2OSYn0AjUTfPEy
fkuaXaYxwyzgcTbq8bEjPOfDoh0eKVGIWlLTvuczj4Bd05nj02RXU7qrC+z0PMXdETydhvc6dk4K
My6VbTNifpD4kZdpaR9z0n0YuYjwsVRC2M3/tB5JfUcCQFrQ5UQOUCIXAs33pf+TXPwOflCUGsuc
SYSpjxmk9IcyA/jiU62OExuVkd+41Xh4AuwX6PZAbo/b8Vk2lsbFoSaInahTa23xcBvUPDGhfm7n
ChV77E/Cip/PYmNB6lrjXCo6Tg0i0B880CDL+3499DfgLxZCICO5R+7xsvrQZvRus7JLpInDQFem
o8+ZXhl+GKJHWth9onsJvM2GOCxgenVHH+Aua2LjMqRbvq79DEavN3UGqq2NAfPXCsOSL7udPJlb
qyUxUdkshkxavOcOHtgvJSdZdUpzWoiay1Z2HqadV5V2pKCbnluMYm+AysWCBWSOqQImpoemd5u8
KHj1oTRlhgd3ix2kFhh/hFiXNAJZTYEwa7y+Kvy7xGRMiBSmFFLEgIC04XIuYps8Gn2q0XKS0GRO
FgtlpHo39p1M4dmvyiClIqzcf557w/NGUNAbe3oj5iDSKNRz/GZ2JR7AujzagiL0Z3APPOkvUHv7
DqGg3fseH2WEDjlyVRSTgK4ZInv10e9JBcDWptGSmoW1o3Dr5Mc6KvfxT+WHSUhrokodXn/M7ufQ
hA8S1J5lgerxV/Hfp5DYh7nixt/odjHoCW/2+TPaOtjeZggqZyvEJYw+D6lGkXqcC1MWv9FjXGba
xf7XrULa1D/j6fG7DnC0UjtLsK2DEnyGMj0oZJyVje9Kq4udq1/PRGuMswbX2tOabPJkUVijIyMr
PStQkQK8ow5O7yYuRm01fXvA+iBOE8f8uNY+nl4ktdV14P/K+aXtO8UDdJt/+mDKuUoRQrSmuvso
1+fvkdOp/sv5BWJfJFTV0Bcs209z/0wrjoaU8/wL/Bs7w3WzDepv0ZX5bkoqfUVGI1JWyTv+mm9O
8YGDfirYmtuvbUl6KaxV9yFubxeH8p4VxwgdMvfjv/GJysocXU4ymLObwbBpbKj3loe9U40rKiIW
oc5wmJ6SjfkFVLhYVyrICXEq+QSTQBzP6EJWnbempfoFJSJmqivSie4xmH4C/UXMlCJ7VN/+Iki9
9lugskjJnnoC4xdKgXTHB1fua3iR+Zpk6/n+34fL2fcJ/+oEQqPaSO7FFYJuzL86p+ek0IsaGgYB
596FNgrXwltdlpYDD3nRgsINES/T4V6OFRA4zP3P1t8igvUrEXWyPNqQdf57rupIfZjyRBlzKHR8
oUlpgx20XkwfDF0oGVMm3QByAZZ0Rm+xelEUuQd5egL6aj1nFAS3wEF/GBlZpoLZdvu/ms8iomve
LMo7KCBif3LfU0sqDjc7QohiUYE6tpCAH10cgvf10ru967Yk88h0kPNJ8asM3PgdEUJh5ITNJYxS
gtRDGZIr3NxkmWJ5HC030wBLREL0SqlUjeNU+ZuRuHi08IbienaM6tf3bLWICoYibnP/+qH9Khsr
PI1JJ6PvHW7KWq0NTmy0SEPiprcrK2Cn1Pekb8tVZ7imHQ91yrh40HS9jjLJCIMlHK78//iJPjJk
4ZazgdRnK4UYFrkQKW7/JkOo3UOebM4S6DEnDAYe+wowXCOsXoUKuu3ODevmF8fsnU32vWbBMHoi
ucl3kd4UBdKNQNVJb83mkurPhJ894WR4tjoWDKuCqHPXAIhm4gf0NNLhNvcbb5PAg9sdY85QkbN6
+Nvf0cYVboPGQUtWyodhyDhbhSQwRAXXIh9qACScC3pPaIZgNaBli6rncDxGRnz7HfQTxQ/ub3jo
qlGBisKkwLU8tehppHvSaL/W3KiDw/Ot/Uc4c5jil4Qxukc38220sPsa6p2HQPkV2Tnai0qGhf1h
VrmtJLkvdyo5kuDsTwmCEtZGA7oIB5CEeG711DgwKte2miOPXPzVM8CFthnqd8RCIsoSXzMTpyvx
Ge6XttCGuLqY9GZCPtSWKPeqCvY38SP4FdRldLTutrEaiz00N/45vDEK+k7dvsWWTjMaAmYhr7Uw
ftrvsNaUOQAsomRrnKH++WM1mZNBNFoF1g5fvJ4N8waXPQ6sEoGLL1HLXM4USbRwSAxz9zLl8nGk
cl9ELOfj1hF2JgsBZwvDrmPk5sJAGVjqhMbkNqwW5wLWCePczQr7SGsPWFIj2JWAVJkxoW6K5vf0
5scPrctDSeUY5wBqbqxrJyzqzxMRDmFZRbXp1oq7ww26VMrDGC/0wNW3XBwSSbPKdQTAcJ7qPBVM
lQXu9uHu5tzqdF4MJeT22EBs0zLmnUXBDyXlCffn1YtG9b0DP1+UQLuG2cmze1wIywUzcar98M4f
5xBVXKXsEs+dO0WOdN0uvtOT5AfYxlwgy8uRq0xgBzS3+8eblaAsyd4Jyr368Hq7C8V634R+HT0b
U2xdxxL0hm+9T8ajZxIalr4AM56GbKPtN54QOge4Ben2VjVXeiIt52y01DeDyV8D7JAhA1htu/wB
vK23ioSycyyCPE69SbfZiDath81RVrViCQcGEnt9gA0L3dU2/7REtlV4LFJERBmZK8xW1F7esx9g
mjALDLfsTSFj2B2zPbEm5BbaDiPUsZanxMemFcvw/8ehCu9dlmXBAbCoqESoAVro38Gk1jFwIlWu
DPN6TyWQ5Hm8Ro/am6PUKrBcKbs/IRKTG6QnGG7S3cMd9oiuPr94QKHiqO4/pkZuyTSn/knno4q8
NciQQlX/tc1XjgeY/DTxQvwnf6k8CTZD62bT+0uZd+FdZhbRho11qZP6ceH6UGP5v1Gc8MB9NjdQ
FukKf9GAuWFRhjxaxv6z0k9QYekdQRgKRAnphpAgHtDyGHsuU4vQzxZuM0pBMmRhAjlKsWUm6nwt
03udTSGf9ZKS5FnbBgldaJy88yKbHUZOtrPnrc6+oYG7hFrvpQf+k43bE5yAuIPgXkhkGHAx6NEL
o+ZiigJYDgY2Lo9hAwBRKZn5cbTBlzWRHxP3gEDB6s+P9vrSW9p1HoDnsw4C+Gk1rGsy0L1KhyDs
xa16p1BD6A3QlvIAck422d3IoJCccVsLuye3S9CECSSJInZVM1ruHuXL/FauvGUcQ+jy2ULsqt4r
YHxnkVjOeUALnT/XNEGsph3wMoihmsGTjXRpzxo/c1tp5elEU4ARxHIibw6gnbQVG/APpJW9EIe+
hIu0RTaNjq31UV/7470M1eM1F5NTO4gA5AK8RDoyyz9hXecPOI7eEs/POxfiwao5AEixzdckhV8G
8iXOxZJtC+REEv06vihXpN3I/oojdNTtgP5WxT1xrWUbtq6LAX/4lO704JReN3nDMKPHGGCfj91Z
+i2EgJhKpNynAU8ir20mveVbCS4dmqpxlPIekuR8ibwMwpOxQZ9OgeV2By6MP+Op2iFzER/a+80g
vcfa2qukQsVmCJVF6PlLPzbdanaBg5e2XKbCK6DG48nCvlkv33cEXdad4Y2DguzsWKTgMORcYBet
gqYJXBAl+ovJtB7jD+QEKiEKzQwXpicvJZ2g6Azv1Ll9Pyqbp8eZyckfh49kBVmUt3wz3ZO0f+CJ
EEgX2XBQ5kjrBVNIwDoh/rrT6sHa4sh7mJor5M6P2DS4S2Q1MgSseaZYtAmlYWho+jvFK+d1JyvV
yeEt7sZ3tqj2Fq3vf0i0Bm/ICL024pxt1TSPlYD6fX1+Uj0KeLPDrkOK1pVSWTEfGxjp0MZYYXST
8esWj7+mQ6gc3wGYNok2DJdq1MwI46Lc1+O2C3XuLlh2CEK6MVMaXc1YJGBI4V5HkB8twa9AFWc9
DW/BPTv0JuAAAnrJZjreTK20dCDCMlabYf6gpl/T81uyg6zF0kJXfDOsK/NtqYgLC0q+Ix7BRMdb
VrONQ4afPxq9DWs4uAsAq1CaSR4JYsPFEidvi6CYuP3gnyZvreDCFBy4xGMZ7/zMCwvhhMwUBOU7
MF1d+DXs46axcpZyT2w6BIGuW5Iq3Gvm9Vkf9adFHhY7osFSiIHTQoF7E9H5HKWNVLauQ+owi3C7
xgwJ39RIWoAmJHI4jfb3ZX/+LXTIXoABpbONskEIPE/QWnsGiIEag8DJFpg4cQkvOPHvSXuNPFl4
lSsWs9YaPBb1AVwF/fhCnD7V4qCw9TNicRTODbg0TWVNRwlecKhIvp72L++GJmc6VFu5sxpfCrUS
VPRbYqBIlTqC7QDFgNdUsW0FeeuVtJnXRdw9R8j84OMD8/wuJD1HIlEroyQd9PlNnrD0cTMr+12w
u8cYaBLTz+VLStxZVKRuYb4n4JgI7gHT7Tjde4wdCVpO+3k110zwEArvH1xSFrez2FJZs0F5xS9C
OfdXHPWEe6RrWvcwN82kI58YE3y2FAvGUG4MZRq4r2JsmEtf/BrzqLIsjMiIQ67gVxqzcn7ip/BL
9139luWEMi98ScycNK//rgwGpMxaw76lm1lRLzksqQof22+JGYy+ZvF4PJBh5ugJduEkxoxZdiTF
rlUkxPa2hCBgHCIwRRGdXrMPf/MbEUJtm4eorSKlzKJvrLJX2mqU5LyONbLbyvEK6BV0Klst0Mq4
ngc9uBjtf6gYSwbwDTTRBaWAr1v4dFLtIiuqHXzvjZV8KM6/uHMW35GCa3WiTWJ/QkFWHQ4jbFDS
opnB7AfNelA6iseTqEEpyZ2LyQj1KzheYQUKYOPApao6R/I5Kr/6mEApOnUIUxq6MwDso4K4sC5N
noNCoLhVt8jeXNnAhIhuKSDLOZ2pMf8Rh4kmEXZyMHRqQT3AW3RzIh4RuQpTbxHEBFClpDZCXq2n
r8kD9+TkXTrinK8MOKOkgHjXBzppiZFbjEIsvXu3NDNabqERx9iX/+uAtm32NH6Sqd8ERl1ChVob
A1G6yUVIs4rtvNrUGz9PBfk0D/GL97YSeHxQGeJBWYiYItaP+l+f/fEBePPPrbFWe6wdFcD+rLUB
T9XpggYi4KurJksE4r9eSa0jSt85Q7hk09ssOU1GAp/nhv5GwMVdiSoD6AUKgIulzsyVpObRhYXF
Beyb0SOsmreEzeWKDvrK6WHqxVWN5kveR6XS9JLbnvtFuggRFgFqcySccBbcmVDAEA4aA38KqJxJ
SIO61t3don+uoZGpSzznPUp606OqPkF05hzUP7ca1zjmK9VXbwVLc5m4brhAXJ7QjEB7jD1DI4A4
+2zJwF4NdOoI+YJ3wGyFEjaeZy34CYE+6eLa+olPkZhOKeaXzGgVIMuxsTqjb5MzHXLtsJYnPUjR
E8TGp48K7F1yZpI8gZa+FLDmIM4s3ZjLTyVJoOhShhUYZ0mWwiiK7/LCGq8N2sV92BM696HNIJdR
56Jc+IGe1MMas3e54MMiy0uNNOwuSHL0GIdbgMu5MgjaedCuhJQO1bf1PN1mGZ+PrZPbbcdiRgeH
bidujwhTHeTRzojmYiak4oaRwTn1Aw+T92NtOxM0FMdRhZaYWvqPaE+cpIe7IqZ1EcGnoW7CZZaP
97W4+U+vhG5z+ZYBacR5EGgcY/Ihqx4u9a2LtISUtO5cqAJ9L5H30dA2fL7FumnR9u7L/1ZCGWnL
29oGmqgMLsmwxg8fgw+P3HSwQCK+5lHeuHdoxAqqC2S2M5AViK9L1Essi5eTi5v7FUR+Pgeq38DN
9VH5fjP8i90tQcgWeoMXWX2Mruf9H21b14ZCUkDhZwXPokAG7N0YYrTj02l8PeasSv1HSRptKmX8
coxvPpIYHZ+TIp0Y7WNBsUH2ZKiv69naOAqnCZPfOasFQ+3W3XSlcZg31UV++4clYbitUPUlr1jd
akSt84ZFl5TzOK7tiTpgNlhWWF1j8t6nI+PWYNhhYyKfWjeW4uHNAiWhFqV8R1CqUSbWAoBbm750
bb9mkoadJ2wKepIAIBakZEVoEBN4cfrJIkE8w65zYFDnH7Wl/O7dxkTyhF2cIdGWiBXTSIqqOvD9
MgNTs0M1LllMa9mhbGuMoCYwX9L9xoSO3ZXaK2hGOpSvYs1oNh7e10xdJmDrK/O8Ntr5MyZSjymb
ahvNTqaG9WmXwnSutjBq6M5CFuNCuNbmCbHvlqT1wZHKbc4z5d7EoFoIFmXhGxUdM12u4fHId/Xd
RtDNIcsVaVCrjZHyj6595nMRbSWTw/4LyVRe9mV6+wF5mUhIgWp5zYc5nyl21Ik5/16vv+/+RxiO
cuPFkcqbOGuM34t/UnU1PGF8ngjKFSb1h2P84ctsXJqLMAEUtcHeu7xP1bQ2qhwKOKOVvwdEUnT0
YUKhCp1L+ViN9WyxXukWY2OeP2ddbaAhfJOBLIMuua3WwoChcS+dWhXH558h0uqNnvCDR3yq9uPi
KDO6t6wC+PaAzi/7lY2poj2gVaFVUp5QXOMfwBkPihLflP+5kWUj1wDA0xRjKVjLnGykY8QKg8YW
cEhJ4bYxeDW9t087BnwsUPMmbh0dUZYazyxEgtRYJ1BeMFS/dr5EmCWmMBGukHs11y97cQF3uTyy
5iWx2L9jVqqa8dz2vUK3ZdNyKh3fO4zse1GV69YAnN5knlPFmtHBg3XPo1bHGN8oPJfDiIq4a6K+
M4yC19jOmdpMFopaONzYQxvg1DcNCH2H9SzHPvVTJ3w7/ydVVMNZFgTSijMN9xv8vpX/NN2KDUKT
WhKp3sMLmW7D1v/pvQthA7erPBvRdIdz/jeMhII0HRgS5LsbIhgGT1j0rxT7Wel1sR2G7aapKXbH
MbNntE+dC9+lfK02My47XkpmWDqVe2BkLs6dhJpzqt4gZ6oHoQkzbGRziIZcaTZT21NIRZ9XzUgD
9xljj7BqVIc0yDzutVJmsgsK//M/JPLNu1wbZN0qX217DSlOD9kgDZ/mPZGJX9SiTq2OVlMGDG1I
XbNoNBUiqX9gRbd/3mS0kF7jZ3IhVlGjt/ApUYMQbQ2DoBF31dHaCwa62Ssgac+za+2dbYUTm1/I
JJo4R6SUVL06hDKOoIA6/dG0OMwpjBu+hUCJ4Q4SrVudTpCqtv8j1dbYXNq3szdF8Hjq+ccLEpbI
Ftx0cEwSNKTrF85P+vE1NVFMTFS1YMVUDxEVGKOBhT/QrKItWB6x8Jmoqsa5rMdgqEoYyge81HP6
EX8p0HMRskmeL/QOmeRzdVeKmUq5fPqUbCVdhd8SVZ9D5OjdaCWOyAyptvetPydJu1omCga19pue
oZhl73ymsYIlofntMMdqFcrNWcCZ7U+wZIHwJiMsvPOl/KapMOtQI5uGQ6/TAEsfnzaOdtrG4xZX
f33LqAUX300UtbQfuqi+ylfLoZn9o1aimnamuFa3UKRY1ELqxwQIUUtWQ6AhTE0sNjpwXcFSj+ou
IcrO0B6AUnZb8+db7lf56fyPa8YH2yzTFoMovc5kTmtcfp/DDJy8VWC/65/mkeh7ZJq1+ZuWiOjq
7cxe4JULcDSTUGb/A3RKrQh/gFKIQieugyyED90JZbvWCmCBdhbOv5yG8mQ7qxe029n/nP6f/tcG
4wrjo8qM9CbkSj5IwyIQ0a2OXHJoCGX81kS1r07UVQBaB8Lfu/o2SBReVPtQl0xoGVp3fHlI+S4L
BVY2YvFvXKbCZAU7YxALCepihERFN9iAuQt4tyCiKEFlEaVTO9Jxt+anZmAJOfVTdG5VmqQQjrDs
FO3HUQE/P5rMtKKbcT96k81QlwBKzNKaiLFeDhDHPq2jdC1dKiF8wrPjlo1wQ/Ng16TDnuaNXzg3
I3rCMB3BpOftCeYJdDCtKoKD25uqLo0IPA/nOmVUapEjCbhR/heblnL43OJupMjZ+RNnhDCbEqaP
5nx7nFj8ohyEgiJMuzIEXVdYZp64ZT5fyc9BHLAZqyosqUp7m7pIdnWcdLS2hR0w/YX7FsJIgUF9
mTzznMjhH+ZtsdxiVnnaVL8EW219HNy0VbimhAYnF+WGnEcW17eACNLSFIKecaGoYlBjlUxvJYqb
CvY4sZuU3IZzRNLssOWm9Wi0Abl7EKJg/fnNMsjPEh1wTOl2eqQZyu20YLaT6FXRvYfUzszijx9I
RMkRNleSDUGRRre0Ah3XavKGWuRj7zZqBNtEYSYfUWrt2A/DCET9hpohEH/m7UM9w9WQjgW+cQPZ
QfTKjl4JX3HEoYJOLtCM8wYdr+Taofc1l8W1AgfGqFIE0oJjH/8oToF0DJBBjfU5WOoLYv+WAfJb
r1MKp37N7kfhrLBFn9JGkE3rVztNo+ZKIYU04ofoDm7W+nK1+OBA6r0HCC8ke4weFHTfS1m2YArN
K0q/g7DMlNs+syH0qBo2VfTo198e6hl0ft1h58zNXfdhDv4s2HF6790652QXT/8de0pH1gz0KdvN
0BWOqc3lQPDGxtu0n+gfD7ii776PdrZaLpJYZhfB/xE8O6N7aVuDEBz2y1ZV8q++Vu97bFRELxSg
1Isph3Fn4SrU5Z3CKJFoz7LGiUfZs0FYJSx2dD9HswpW615ibSPrdvsUntX05q6OJm1yL0Ot8p0k
wagW1T9pbZpt8MFIfxuIjjUgUwTuAtY6pmc0+r+ZjDy/7ncSdkwt4mrhsfiIhZDafSOA4J3G9KSC
v3m1iB5N1hTIpliKaRtoiJ1M2cX+Cb5U4g9zsXvMdjF9FOIVBuUI41E1sqxG7vhnCfGR9OZRkcU1
rb4LeSriNZy/B1qPPtmo1nBLvP5cU2NweSd0uELsgNohTqN7LhBLRtSU2OYKHs/V1bOykLkrWJjo
fkIo+0y/zmC+QxmBHXTbhBSPdTFu448aN4rFDj/RzrlSzOpckErX1otYiNknR3KLhtM2/nI0pFjR
VQT8DL2ClUPYAnEf9AAH1TF/bOsU/h7rSOst9HWhl+XEK2/Vtc3+enyRqvTrlByyyNnV8xeMq8la
cv0+9IpanQ/5JYPs1ZzT8h6CBscKIkTeNXdQOinVKKd0FcfF6ShVgw2wUTZY6oreUGIwzKodTz9j
jd6+4idJLjCDWfk8nHbVOfLFGcRSfd+V2MnTtSY6BXzikQ0NDF/+TM3vTQer54/TytX3AMS3WVSC
PnY5DdPSQ82kAU4zAGKvU34De27ueihvHfoW9xVivWT5iu/kpIlvFYwakDxcmXWnVmrTWKpBLiBr
4KwFnP0H8KanmGlxY1dXl2pAzqx1CaRZSSHfvdzf1SFHEiPT/6e03DKEv3MvkwzSU5XqnT9aN/Oa
tWcwyC6SjIeT0rLuQTDqeqvQ88fTKNTp9knADgscM+Bhcjvj29lzuV609mIm1wThUp9OR6c+jT63
44AwGK3UiIIKtbOM6fkFresNlJS2hETV8sTYmkHUA4G3d4s4halALPqBuRfrMvodN6/z81i9WRxU
JwMxuwktUyHFmI/VUswMnrLrwGqey3F7BNrabyI9/z4qKFSKsezO5AxqRwRp8syzW02yMWV1MmmP
Dt5EYAfKp2+AQil8qnaNA6UXiJ/Zl/clP5ykzLKaRSZ4wH2nk13QsWUbN0O6Pbra6YUH7ngo3JtW
rMGp0AFrDGCnnbmB/qCofSvsvQ+oUxXvLYA21MrPs78zlIzwAm98ycZaqkaQPPzRre+fmlwl96xM
H6D5VG6i0pnW2hbXeULLeW/w5tRjhi0DzVC8aluua/EzRc0uLDbB6lKeR/4lolEVcYqYXaCokOnW
7PnU5KEhEz+mhPAzm2eNMBdCWbMzG8d6ZpPbtFTHhkxgADg3reYRvBHBx1tO5nMewV74asCQ6vAx
1cBcziGXc0vn4ZWQDN0zseosseLMNjTyA5XBM0VSNtFR635jLFy+4XrOcqn3OIBJHJvaNs9XGV7d
ycQ4o8/8bDU3e7Dl22+v2lAKAWwh+g44eo7vmYvx84zqiNrDFJXPw/wVA/+jHYseUl5ck+5NpsbI
MaIy5wSEGhxoTFL4RSh7gwHXN2ma8QNHYsPvwLeIYGdCJig1EQ9zQs81gg6YFnGe6UPZmIkAklK7
QjMqvtutG1dM9OCCMRNvGvZDU4Ofd8/wbbrVBcZiF6tiMbHR6OQWDX2E+qceR6ELP7OjtXR8/p+/
ZPLA/x2jnqVmfJUYp4htgRprwJcNVyNqvhv21HgYnno/or+F+vrNBB3qpVAHf2IgfhDLza6IcNOu
QbkcYnQAsGtulQrjxMNnJbgGz68nugorYb7qvklYzMRWk/f/BZjnu2YFwyyBP6Lz5+7TwnXQ9IzY
sdrmYI1Yj6xAbypqv80I75Q1YckSv1dLhunDCeakqL6rRsASfAmn2Xy4oGG+HLk2yqG+bAzGo+uB
Y7QOmvxK5ycXznjFhE3ZukcHA5vANbThKtzUJ/XzOsUMhaa8iy6XvKkQW/LdVs+S75pGekstZy6p
eTQbRw0u/SFYcEaEgmrK/wSuQzLxBqoB7tLhne3p4OeXOWL18fwimcxcgcT5H8CbyP2pzwldPIfG
qva+dttHo3tHPrYJQQIBHSSphRCpgjGjJKE555TDUe0X0aPXS+MtXwvv297rxadvHgEf2VuEhHO7
OP2HqBPFv7bJT0jYNYXQ/QbRTWIzZn6iRYyzawXu/uHsdy73W042QLTZnID2LHfFEww43hCDEAIq
n4DNJ5OHYqtBzqpM5Q5+XCBP236rM0eqBu0I/hifZ7ie30LDDAGZYmJgRnciaE43oesty8vntclb
s+cbokCB5lfNN4HeC432HRrPVxeIdsb1vtFlXQ59JWIlAGFxXi4xYF5clFNpTnE0WLiPwDBtBR3K
JocesBjA6KsuTmDvfAthmI1QXW8V2WZ0sNycTaVKNTej6Nwjwn1C3Rp3QyahplCsnbCL92SxWsZ8
ogC5Dd6hWjAd+a/NsRuoPO4HjGj81OYHc6G1WM3bzcmBmS/mtBq/HNuqSv9YDo1TPWzAq6L++Ej3
Lrn65I2cep8YbdJBvCKCTwyT6jyKP4rUJZqq68D7iZoY18TraPBGvWwjX6gRMnxCihjmrEEEP4td
e71mqd2p+1XIwxsDD7KC5cBf5a4e4/ZGb2kpQ3F9wzLVKJiyqU5yFo+A4yS8LZT6FkafmQQt5B69
5GLhcLcEbU8VAJcgQEeuMYmdgLjsSiz3RGGOplJs0AzgK3Dy/5iVbkUo25K4yUHfmt6kD77B6VO1
yi0un2aPw0C1chBZUBmK+ptn5mR/rrZjZ29D9xQo4hNfHRCg764zeGmuAWBcGXvYnLcX7tXbRgAf
A/IQOJwG8QVQsFZ9LZ27UwxETTr18QdNB6iDySLHuFH14l+K9yYRLv9ymRLY/kP6XRL7Y5nH8pbR
FkbVAFoqh5hoSYTIYUDv/H1fQfnRsz8pCkYPCM60Kc5pGDNtUOjl5rM08siAW/3ljGjNvZami24B
x7i+PFKNn+WXXdESOuM3UV/l6YIl/AyL9Xvm17hqZW+ujuPKY6y4W6TRDviYrYZ4RYhzVpUVFKyi
8bpOrLb0Bj0a+FGhNIi9/aXgTkx8HXb0bS0aeBeGPAraxa+qb4hfZCPeyuCtZT5arJFK5nKYe19N
bpUO8X5a5z5OwhxepXBfkqj14QLwdrgooO9cRu/c9J4fqn8dozzqEJ6C0f6AZWr89reQ6uOosDEf
CBJ14YY4OqjntCHnPO3F8hvzzpoSMqw73tCWUgGceJxVpxvtZcF7WoXk9UAG8x5UUN/l3B7bRDw8
63KAXLMyM7kn/XRbeW6olUezhy4loCOUCYTKkmlyr9Je9pjMFd743QmgT5sxIFJXDK1n1y+Z0fqf
ZJL3FnyCrGq4xUDH2Y538jQcULWtiFB5TqKFiazXLgs9P7zt/oTNq7u27f27ZyMfW2vOAMBB6DEW
gk0sOcE/0tuvQmoV2hbFBYlcYWa4Az6yz4mzsqUFnyvgI+JQNqKcr+zTwP+mbPd6dIgtoPo1PXq9
IiyMPK8wVMPCKxxzIDC20YMhlkhVIowgFniGY6940Lpw7YeLZxl8FpZP/orGKAaIuq0H3pa47Rlj
/DyMLkRghv0kJZfG87wqZE2KmVlEQ0DsBIcZdFiEa+NlaD0oUcZjuhzdZUKIOnIB+vnf8N+SZVAG
o2SNUfro/cCP5NDrliyMS3OD3l+oDKjT6rqYmXbWox/I7QJuphIjDfh6yPRwqA8SqOyVAVGjOxBC
92Dau9rNUlDY/lEwH83l6YbiRefbBcpMt6tG8I0p3K4fmrB0SNyMr7zAH2sRZvLIuStsSIJpVKoF
EREqmtJ6mpbx2EMSUoj9kBbBtcHsINoq9RA7LPvVRwgz1FLBN5bOU68JMw0FLnvhtJy221Zzf96T
EBiYXGpWTSJbGHrHOL14WkYRX7cJlhG6EaKITE5nyS7/pWn1/K4Di7Px3QESOs3Y/+ihYAU0JSEb
A7wTmqK3EGR68fC6f+ey8vO/jZMrHTKoESGyLXxRh4eoerNfCTaZVCZevJvBlyzuIPUWNfMA1hR9
bt2Gm14m6OnAZ5Ve6ZnoikVEyIRNjCtLwQHA7Xvac4Z+5igpIObRSfggOk/BglGWL8BNZPzRm8Ca
i+PMNGKylf+mheSiyNfXeNq//DOmvDsB8cDcRNvOBLA8DK8Ilz60hVsI4MjXvQrgHu16viIyCL3V
NVIp4WguyGHrgi0hnCKRL8UTQG6atwXAgxTcB+SGAv9uj8AcDWdTVYmuiMu37XBjm2XHF4NxcXxQ
/JSUG6aHN8c5YTYunzp8+FYcB4vcbsOA3MysasNGgIstqBnEACcd2YRymxe/OzMQoGTNqJaEL8p1
xovJeoCPOOkubp3istzf+O9w1HNXnFp7a1COHllbdu71EcMG0SgPPhYK82gIGLmCQMh4MrKeyQQn
ffjgI+/qXLUAohYgqjAz1vd3sABDmzt7x3YxhS71CQwGaJQRtVN23MXxlqyLJZ1L3zqJE1fHcVK3
4L/25Me4XLiknH0K9+8ZMHxbmaHtFvv/6oD2gwYBorxLvPxUGjDABYaiyZPU182ztPLApu9ALmSf
rMdtfd3GEyORGkVNeWt4+Yw/a8JLEbiKgONi+pXZJaYRlRV2cfy2uIwU2woNA1c8bJYT4u2chgvH
aB1vJxjfem7HV05WZcIQjNvfcaDMVJT3i/UPiFnAx+S0TfSX2AbHC6LvM0ZnA5nYCL5sFeqLT0I1
KK0+ZOAORjTneerLCq4hPozKK/F7xW34xzXy+zCJ5czGS0oOcrYBLpSOL3Z7bKbBx5Xkp5EqJck2
lwhUcbC1Bj7AXQ65i0l8x661ssxTrK1PSrzX67Zkwr/BOD97pEwSKAk1vQc2oCzM86pHHcqrs4Zt
osOwJZiyJxYJpf180Gb4n9UvcQEV9ra98VUaSYRgvlRf/vG03J4Ze/69I67zOXvfx/TFLW/s2A9Z
SS44WIDfhVfp3LwPdTPpmfdGaAU8TKNKS+SgbaVHZJ5ngqgvwksuU/8LxSqflY0Ym3CqOL/P1/Iy
xtYdHGgqD8r/OiubzyBE5KkGa60nR1h+ddKFHmgMXut/Bk7Ltnkr5MGekhQue0jQOgKYxbUnXSM/
+gBNl2ZSDpI4F6Sh1juxueS2YyVytYB7NU113IL/vqoiLjVLZSLyO//Vq00bjgJNqzVvQEN5zbHQ
CRs2DrPILq2OxZ2E2wuYxoCp+TiiRTuLA2zgcBOgKv2ZkFk0Pkx5bsuYmyp3Axq9eEM2UfPsSMvJ
XjEOS/v+IeR3VMlw+MD2vli9sPC68qZ8xDQjCk/zcrzCZCBGqp+w8DAT9Ar9JcwqiRrzgcNQTYje
oXUUVVZXXh79g6rkpY1D1hG/ibQn5ppf8Bwy8zhjxN+5ZWLaUkM/saR07ANdEby7iqB1TtPGowzp
WPK2KqA8TGZBztCnzOf3YITfzZvqFmymTTUono6IulEhmCcJL79xhtuEd8QGweuf3ETunzOk1DwA
I5hFa9TD6ZglaP6IYsV9jYZO4/g+WHcB7UsoVG+CNyEnAhKeBNdlE26TAbj0xFO7FDHYh1zxmSCG
1FXdIltjkerKeVCYeOknGhB++I2ZSX2nJ/5cOZnOta0AuHhyGKjdBkgvMwYwF+CpXeA7v5wBDbBJ
hG9+Tu0Id8nF5xMsfgo+EWCjbhxDEst7xORYXDZQTZngvpaVzhpK9hGdMDuZRYsZopm9rITKgq4L
Fd8uttf3eyc5Ai7rFCeq1CIKZ3eBaB4ZR0yEo9YxptsFUcOUyWTd2ZaTRTxYeA/9HHiw/k3xZyQk
OKXWv2EPfKbBF5f6D9cCIsQadWDtWrM8Oosd0/atNvaRh0FvvGFIsgV5wXxhej7pB5sgr608igHv
fFYn3/bFC3gi9iefxrWi+Xgq4K7DEc+ixX1Sc2JVmbu6xpNYow8DaSaSsOGOvPoHlcdhgiEDb5n/
OFdP8JoQ6brtfNjVgkWMMZbQN174Mjt3wDWro5rojUyx1wxAR4prvvH3h1142CXxIPJitOWHY8aC
k6QfkozWATvN+1JPAGBvusX0yNJv4BH7W5yEyOyTw3q7rN3wkyuJUxLjhZGUqoJDVKXLClS/SJvJ
Jvt36SvwhIQMqtwWnvne4LsAOBH1kiNr9w4pvgkX3IPYHWel/DEaYT9Zh0c6KA1qMpYU2kZR3ITz
+/Ied4QuMtex2sIV5UvA2dCWkpk7qOugxfb7rqQmL/yoRU/6aWeHMCusI4ocqQ3DXEk0qBiTsNKM
Ku2s5ojqMJE8I7hwJwcMWl/6UYcSAxL8pj1/O1q+jU9ulaTZ9L1ZL1eJ8rC2dO52+7KoVuh8T+c5
TFPE2uc7fXlAiZAgBCDMvIHK7wjpJiho/NAObbXhQVZPS6z0uBUhtsvqp+bGn1wPwscvqxGMuCRl
RsPi+ocFrlhcXA6SA5qjTLr46sNCjtl4L9tbjBgMFmU/XV5ZToDyH1hjh4KmsCQK7DoSQAhbZBUw
p+OoBu386OBTRn/N6N45FFuqYKOAR7CLFaUPIxqhUNzakaqB7jFI3CMxp42WndUcTYEK2jFzloxS
cL4KYTfM80AVBw1VmGBZG9A2d+lYYITcGrjNEAdqqHXYR1FOriiBmNZ5+RyyTr6BRodDSJuwJMby
rT7uSmfwudbAEQoWqi+vuMZZuQyhqMIYUxXb6kNxaOLb7C+Pwt1nU5nKqEiamH87hdAdHM3yQq0S
U13+ebyJsuRNR5fVyn57HtjEvxlgXln1KwvtK5Sq92VrM36w0RCBEv3QE3bq3okzGdL6MNC2Qgmg
HOi3bIcjatfD8o0VrBkRyzDAXM17XTjPwPvUxlYS1m234oh9TQihbeSBUmmq3WVwFxjCAqE82Myu
EoP3PhCg8KhYSL/0o51RNCtjhoIwD9oBRcDE9QcBKOI0PJEEsTimlHVZFAqvLMaMLsuXJClH/NbG
QGD3d2mOy6KNT4XHym10N/EZ7mJ50RS2JBFSffv5eHGXVZZv6r/pu+5VPqdNQLHBnVvbHz2JT3Nb
inlKjPNnG9kJfzbz9hjtrnbjHN3TV9P85QtoiqGO/L1lIIV4bvlNx+NvYB2TSN/4bFAsdJbQatbf
1W0Ejap0K7ZBDXWGUY9kOmWGwGIocqwW5+LjxOGrbqXRcYwhaZM6jXo0zzuQw4WWPq0O5nWJM8Ig
eWkRCk44DPZ0b+w2oshzc3+Kgxf6mL9apHUJQvYiJGlC9uASW2lpkiER8HQAJhYLCEt3/EQfq8aI
I1gkfJpUGWmQxSekZVz6UGPVbMAMg/ONNxR4lLBKSfVTR6jzc9NJ4TBmZjMwjvvsppHjAuPqolsk
QNYXktGT9rxrMAnPweMPfkcAkRqllNIi7wpKcPqEq0UccRQZPlWL98/Q1EG62d1lEN16GSWqwRy7
7HXxj0wF2bQyyraO9fjQecY366CS1zPt4LgdpCiJ/z3NDZHwmMohct1uVMg8+lSyvq7A0OOGLBFz
gD8mcZGl4gVuhjGj857VI2jmb0psnuNietUwVBvOMi4fyIvxJb4LhVcdSCzrlAV6ivPxp3FiEVfy
lOGBtlfLU1mWTMPLj+AsWV5w0ycVnZM8J4GC+pgSC2SWR4EfCqT4jwtA57kY0dmEwk3D3bSIn+XU
NqvAfhcTgHJO9CtqKw8xdntk4jryIRvuR7TzXpRo66ocXHpGJPMCgmCdtn+fa+zdurX2bLf6JFTQ
nPU8N7JtjSUQtefZQMXJFynd9aG30oyU3jwgAeQ8CZVvo6i+Bqau96Uvlznd3u0ZumJsj4XOQBcZ
VtSuIN/kQRb2rOQMoPTAvw6d4L3SFRCnKKymBUjMa+/+BGKjYmB1G0fP1c8L9NYoZZixLVtN69K3
QF8l5FxuAw8fIKj1mHWLfs4lIMph0WMWgpsIXwZ3VxqdfgKlYdcoD/qG6aTJybndB00/z2Be0/jK
mpu/tJOm+1+2+sZejSDN37aVp6LVq8ZPtV/aAFSXcJza7nIgh/BJka4bSf+6ZY6enBTJUnRlgCkE
CZNoG4H1ZTZWx+8B3kVUXFC+xBlyngO30rjlYoc0VILgAtOe++Fcfdt4lVQobPzLKCDtX6rZoIot
wIXHTEoxL3UH1NtKHLtZlCLFggqOIKUaCfxvONehFTGe1wuPWG7IYQRNIAdRAS4SPKRTOKVqzn5y
MXzGC/WPuzvl1mpbKMXV7oPLIc1ZNOQV/r9HhfyFSa82PkVkyFJJe0VFgl0diwd9Pi+y02++JusG
1gKaoYoNfTDANEDSHKiZieLFEuC/tOWzd7Te0WQkbWifS8Fl9gCgCsWoA2H6YZ8hwX5ZfCAGRlUF
DLbMucASCeWKhNa2K5XjrEMGPuRExrqQYpLU1bnEnxo+Qsw47vy9gzr+8fRCuZV2DqnOeTMKhkK5
l6/uLJWRw4D8Ac2HJb3SZnVWW6SctT9tH/7OaGFAcohUkHXQKIyYemC6OJX5uLXZD/1Cd8Rs/Y5M
nFWfJdzWoAMANzF48OC/8zQmnzm3CPQR6gSUuhiFzBpcFqa0Y3soRPaExoOgHLSgpQgxz0D2UvOh
SGZUD4hivf9hLU0gExg1R5m6sgXTyktE5Du6HWE4C52Jj3jVzg3bPMEgSaGvG2+vwVIRkLWjC8JE
3SD4eKdULlXTm15xHVEzhj7Az6uNw2HPAxSK+rt3ictUCfSY6X8JHoK9wpZLX9fDRqdagqJuDqaw
G7WZYAwqp45n2ED/bQmbp+fdEHvVPaup53u3zqEg2JJhPzlNlyGEqrC7HnHT/pnfchmzLCwqG5kW
1dYW3nnpEP2Y0mzgDuP7ZbIVjYMqfqgY/mtC5X23e0xkyqx7jahZiepGWTJ7HORolU/3KmEaLwWD
rssHYmpeEi8imAjI68+ACX7Pf669xDmk9haaU/rnI87fJb3CUuQcvGNG2kLSGqGwoGARsvHj2jii
g2ueHzLoB3e9EllSNftT5zsW9ctvqSCdALWnu/mAtKAcD/a8PnTEiHlDRbll+etthdYTX2glM+OF
9xMRRA3gkUnq6ZXF6MrN9ERl6mVzYa+rSIN5Eb6N/PBlZMUGjzGjyRpQkwh76PNuaIL71OBWvKp7
c1W/DygY6aF4AQKSslMDjhMVCB02OE7w+1XTsNvcHldru8dZQcadjvoLXi1rchvEy4ZKP75pj3pH
fsGbOXYjA/KN/I4XfxskNLyimdKFAkZ7PeS2zzuKSOHk3qFskLXtMmsERj6P7+N6hx05mhSz8NzL
ja3yBqinSeboabbi6+Qkla3pD7oZE4VY6teHehM4Y1EfnSoaSg+KcTgUJyT/YnZvAQNu6N4e+PDH
u15epqT9soBedgTVRCEe9SmQXOXYp63NtKwgVW+VsMQdCl4ulZMIAar58SfjtDBXj5s6DUXHd0e3
LRxhs57HbVTGlGzOYZ7iXVWV82ffjKPNc048VxQpfZnHSxIYPnX7VnxntIrSvostLgMq1I7NsZyR
qA/Td+M3n4y2oD+njFzL9MTAXdbBKsYZSx8uY4RPb7aFhcTVL2GvDFM77iM0eq7MOkzmVq8M7cv/
TeEw3V2KMObh/hjXZCn5S0qOnLy0s2xeFJGHGqrxD6RWSY5lGrU9YOtBWVnjP0xmsy7tE17kkPzv
ZsvuggNgi4G/WLpqlLScFFC0tyy9uGI/rF+nt09bdUT8SR+ooWTeQ0SZzYyw4dLboeQ/WBnvpw1B
6ad2RBpVm3IOr0EQawir4ygpkc6+ZKPEVAMFYSA7M/dngcJSB3qsxYAwbLNGAmdXDcrQKikm5W/o
VvPMgABQoy+qynJBgqJm6r+uNvqiVZYsUCojaa6Kt8mmBgj/zBo4zNHaN4qkA6RCEaVC+320iNOE
9nf/4vVk++Wi3nvk8+7/riFZTpJhssypTWC7MaMX1wV7LIavSuSPT5jwVBEMN9SB2+I6fcgZVvvU
5NKHE2wIJqvMCJvcEO386cUGpBKh6+euxFC4+bDHVTKJaLnSjxSCWG4sd2D9kv7wrIPM6X47y/NV
Nl/yQgQcNn0d6Rp0m//YDT/4cXt32p5OxbrnEdDCIeFK2O6EPyTHfXdpljIByLh2WloauAK5zaD6
7pbLVTCKweyU8qIEh6rSSvmlCS2kRcGJRafsm4A1t+zz0ip5zSKYunxYqDEZjR+uRc4FG8rfjnsH
6fAiVGGlbeNcvBDBVjNqPm0hEFSNHiOr7kxXN8QuZVm5CE7D80swxPInWA7VIpBDHr4Wd2wNCDx/
DSVnkRSX6NOnESJ5ltAy6aXdkZzyk7OfQGM7TqF/DtlUeAhxji8MoxBJyIUUg7CmtEsxrjZj1fo+
2QcAlZ8Bvntnv89yOnJoZCaQH4BXU1tM/+xzueFrqL6rWFKs0AFB6SxGSb9qY9qH+xO3AhRRzaty
EFXFLuApC26ymdoTFekJLQh5MKFQaSMJVth2vTyIjAJNYrAtKyC6pWQneTVNs0RsWWh2zTXovbqb
DIiSmxbmhKwxgeAnl0VB6AGDX+26axk1xiAxhGV+7vYhsqXUNH7l2D6s6mwcPvkqSqXJ6iA8fOGG
1pmRH0Gr/P4rynX4iDzz8l2cVstZuxTCmjqHXymGtHVhHuguL9pr8BLtSwdx0CEHUQdrFZNB6Nba
89F9vtWYErJPXUWSISaLcojgGY3PZBapxMwQ+uZhRsP4+kPD9ceNT6+Jz7bJYYDx0DC7yyIykPjY
DHsCUNnejFLSGcc60a+xO3RoILInT/5k64cW2v6rAdpjooe38Kx3MAesFPq2T1lrdYSTPQVF7TKc
jJmG3KnOFF7CbG+RoojMnXRY5ihJhHNRvugD3E1g5gP/HZm/KJjIvZvJCrm3d1S1B8u6rJEAQo2U
J64L4JGNk+9m2yGNyXTcY3HdKbMXCgnS3Cvct156qV1zG0J9lp+cRTC/xLWYNZGwupFnNqvq7LQU
cQWqruqiAcBOKIy4pbMbswnMLq5JzA+vKoFelEkb5U918wiq/XQBGEaR2BRaNSjiUBvKr/8Z3jR+
J/pXD/SZmYEWn/rkuPb5+WdaSnrJ8MAU3x/Q7doQAdxmzEJvF68iyi+VsIqgJhBVgwfAcE+a3xub
q+rRyL3jk3dDuiWR1gaMrctN4f98my32WcUsH5U2JnTs2w7ZEU6TOHA/laUj+clXpsv3xr8pYMAv
B8Gj2Dynxl4GM4XZi91Z0x5dVA30dClttynrfqiIH3J+73MBSz/1Y5VIRmFs374BRe0KqK1WppPQ
wEqn7Yn7LTzfF2WWwlTQ1ZdEXq9kguMbhdXna0BjnGdMa9R/BYWvYAAJ5zqC6zIkL29PoUVDvY3o
cYR2vllrO3kJc+bVS1TQI4XroUPh9h1WM8+9YxENrsIPwgjOlaWVH5nRVRieLjwCIra+7Te7bH8D
qVxSt8JBZFb9pwZkEAkDwfPmtygzd9ebPf4dHkpDYuC8uBxnXPGmfOSe5nQRnhKGvHyTtQJel7Th
RL3YQ5BxOBBrFA6fdaBJKVhnKSSCnqmQm2NyaVRsRiCdihygbTHApBZjPIFtp3l2IqeH+YzjxiXr
2rdIZa7iTnWLFZhiPE1waIqsm203+/ZLgZuutPsKUO4wVy1zF+X3/4CcfXquy6N5Csqym/J8RL8I
7uRce6a+vtYhnA9VU3ePQBPw9Pkh5V+siQoUNXEyV6HyqsES9JzeDDwjGN0gYdGDX6zHbCOUFNWB
2xpGWhpbdYWi2+SgZtV1l6UKx5JY/y3XZprX8U8veJh75f2D4qj14GTlw8K1QCbYHoGJCa7kLnis
p+ouBe6W2c9Wz7O8OLz0lsfmAOuAlQlr6+FAGgJWEIB3NaBGMdjp5p0zvqFF3eGbAYOvc6X8Ho6K
GvItQ5QPEpg0B6hQxtgAin70iVQNxEJ3D6tjQeL9IJL6Vlk+P0ni4yb6XMVmTENS4DnPEK6VPrW8
1egKtDDhfd6Ox1d+caQzVszbRPkzHn50VTy3269u0XmcrhFp87yGRgVUABzLSYVCymbYTha6bTbv
KVy+OdnEJmoPOCxRugensaX95iZMYMO1gib4tAQv8HIarDLHdN7fBZhARj5M+lMOhosGsnHZsFFr
0fYqSZ+Esno1Yydm8EmgzH3vThKzvgOhBZjkKk/URSkqWRJVWwc6GRJ3iEPITelHxOKhoigPW7T6
1OoOMeG2/X/j0V0jzhnvc0SP7N1KRw9AFr4PeK/hFN0CvrjTBSLFFFmc5zQHIwKGGtTHMWRCtnM3
CvuRVG3hxl/rgQNZp3ftJ0MUDZhziCN28FRaZlqrSZMnYG0Zj1rod8uZSeWDaxDoj7h+MjsL+Y2/
BusHnXedb19L+AvNMZjG1WppQaHb9Rm8m+08iSj5BfXabD7ejg/ej0UbV8nCh9HK2oPwcHGB8OIB
jJiFf0LAObJlJKXHYvzk9cowoTYB8jGMH2ZcGV6/sxZ3Np07swoSlhyewgFWAJLgpoV5IoSlbcPL
rxU5m0fGBCf36kVfmqYOb/rcqswb28w9IAg6XslJN87Tt4obQIKB4WLmqYzRSvqmChvAukQdyXi8
vaQiKrKcNIWCiCDr1TXPv6rMSTdSXOYVNsWLNiRvI8AOy7+GjY+cK2EAatF+A41uNAULATZwKjln
/QcvYOcDXPkdsFrTgoPqiVl+RXU5srzei8ggsUKxAqiQ1sg0bN58VAI2N7vKwqbg57FK/Nxy1BWE
zVHxO9Y2t2f644F0EY93H/Isx7/pXvl92iFP0Y3KZIN5rhoHF2CXuUOyGpNh83qsM0V0SPSbQUNB
HyJ821CeKY8Zoe0DHlJ5WDe3KiWI3DHSfk4RqeYWZECH4PjwqwaYS5fLik4NssxlLNIKTD2VAsEw
SEsOvnAxNpvFKKyQX/tktyoWtgS8Sjq9sXnOFLWgMWu55cIur0Ew3NnNuR/v3s4uNyhaxntTh+8J
37KQLJ0htibtdNn31L0i4BN6da/6HOTzdDQXfKgGUWuzB37WVBFnuV50ed8gpW6EajOQ+husTKFS
Ig8Th/ZTvbAiUEV8PRpwBFVLshW1eYTC2PtlBGWTsdjbrb03P+sUmeqTddllyu1rlDmlm5NqedR2
qhRu45ZjIIgCAWNxNw3Zz5ts707mLRnqkUgGfUFBWRhgBKu3dv+NnYVeUyvLmeu8zE+b738HJPIp
bmP5woNUrOZ1lMkkG2A43ERBXSv9tH1/EK+huETT2n8YW7RYXrsNcNfI4GckRGbGV5Au+g9XXi9q
ssWxpKPEA6RpwvZzRB7W7oUssP7KuefpjmhpbHfrk6vhDLHN54mrNPT70ZZtGXRz7AaPYhbREtv0
V1BPN/haxk+BQGsjZcpWywIPCVlF09hpcx2uEyLyy005XzVcvkqKMs7zf4ri/iWAW5Nz8AqWtv+2
MU02fm+1jsa3FNJFS1gb0by0SR35y+Rrznjk5bLvzt0dRLsc8u1aZO4t9ApcFbcT5F4WKgd7trXs
GQZbKrhJBvzlbbHjTl9h3id63NjZqGdKiA+JHJ93hoXJA3KwQcnX0JVzdycCbyLOQsM7YWEqgZIV
f3WP+Ew2LxI6mzvbWyBQfIv/Oa4stjXbzTNE3JtkvqGCZ922d0B5fFgOx4j8kijmVGZy4AUhU4Ux
xk2rWAlunnz6KUbTsMUs4WpIur8zjczyfVh2KZV+gxtx7iUcjtmlJIZPAv5EZFvIs9l357G/PcUd
OKXkGqZM7KMco5SSFrsBScPhlxyu8k+Sn1hkvqtWUndoOUjEjnQVNSVFd5yXBK08/cGM86FXRg3/
lj6w2CTZlHr+P2azSaNQmtRNPYo/ObsCtG3A/HxA79iBoI0080NRw8MG2UYy+KsXh/5fMn1998aH
2mZ+IaHoKcRtcMrrvlovzVJIZe98xRx633Ai9yZSfWY8OmVOWsC8k3K2iLjRRhPZKG2fnq/YeiB9
Y9RayqQ1rjS2Vh73r6EM1gA6JVO3RwmKQ2BkrGJlvLZnorW+rejYAq9MXkSvtG7n9w4NbhztG5Zx
8G5plWhnDQ2IKir0hnx/48oMn/May5HV9SDrbrkzu4QTwNDnZIs2qiUJp1rNm6oWQufRQU9EPBF9
Dt7KQjy56cSpjvxe11BUfdF+iKXfxSvUqFcEAqgCsLIqCJE1G9UFzl7B199V3Bp46e4Jz8kRmPwA
cl+oJUsWrSFPumQ99JX2rtZBsm1iDrhDm+rk0YluSdTeDy8CFi0+hMu0NNUfdHdFbkVJbyZhJp8p
DS3kuoZevK1dcWMNosG+OtyStKXgM+XgfGHG9Su1IxPxH0yvuWVQvIl4pWruFJd6hVLVT0vARlMl
U1opTLNevaPS968cZqbeDAJpgTdylLqHM3Bod5yQY0QAp/PNwo/UvHPXVC2qxBfaO0bqJuKwzI8Y
n8LdRL4bU3EKPNl37lnE90egz2GTcwSFvCkVPskswzeFCxLJFjUeWlhNWi08zkJ6jvRyYgItmO64
TlDuwTGQewregNJpET6gOUOfcwx0aQHnvQ7HiAJskhqt6n8C9NmxH0Styxh8w82R8G7kJJdB0Rtk
LBwpkRYwZMeLl6vzTywPx0mYbzXZmqvlFcmza9LMJXlrLWy/gn00eJGzcDDQ9/ue+/9z8lTaMwr9
5B7BATDlLyubEhMy3yyuWMTqTsPr/EZ73yAN3VE1srGnKxZe/Ll7xXv+AWWxfJydklaBTxsG8+7f
pyLl3wGVwt0Mt6oGmGk2igRLmaeezyFb2cFXUwlogJtUCykcTnAxP0ndVl+aJobMk9ejAHNUpYZV
O4BQsI0/Hk6E5vByAMAu51BA1YtzjaMvSM3zwR4mzhEVA361y+8HDTPlWFjhY/RDZB0h4fvcFYXt
rvxYdtcFyXpzbkFbVfSg0jupq4bJkYwJlMo+/pv8aPX2CD5rl1ZvUBj/+QmNOCyQdouLoDh56yAC
XnFrBgykiDfg2NdA9fA+kqnnyJlGUBr48UZVk2YpNgPIVNmiMM3NcPU24eXxIWu8ir1SZyVmR2lS
IfTzesvaHYE8vmAu/Cg85X3nucZc7HcNHQeLBpn1guA6fX9Vi7N9rFC0dGX4OUrE5lWD/lWgTBgB
vcLe53fbbF4r/3SgZkOvHrxvfjds26nyQ7LXxcI3CLI3gekcdfeT0QhPXq9XQ+2Fk95VR93wDrOi
B8x4+VVECWnjRMVM+7p2wrHtrsaLdEBUBpmv4kVXzKLahn5gXP5nn3gdFVKvbNrcMS5ChNMVEPnw
nBGFjqVwPF1GNN4++7CVlFlj5YNRX9Wl13sGQwUMB8yuKUI9ivwlu/wgM4FrxvxqiYaBbxxUdS6z
sCMk0fceV94gRojuaeDPcpjzeMV+Y8ykfKE6KYIZxtkflWYr+MflgrI/vfi5apzknTMI/sBtVDN4
+7/+R4Po+dbkMGxgxB5cuDS0w7cdI0RcaErogDa3JZ5wxw9B5CTr4cBXZNijV/D054ggHyimJPvE
YYZ4RbzknE58K+Xeg70g7B6uc+S967srL+7LcTl1RQLjOPOQJhflc4uuaHyDMHPCHfziT4nXzdio
K1mO3gxbAqAsh+4ZZSx2sSeTwErW3ClVmdGAayOzwexMeKhcaFLiFrlfpLWCyxOpZcGorS/TDZ+h
aNQ7pykwxYneHwr5ih2OX8vF68szI6taYmY3x836OjsmUgByOGkASEWs4D1kNVwmAaEsBkRXDprs
uScs14cA/KRXK8Cwur8+eb6AMx5C1mD3S46C7kZbCL83H+wh0lWjtOfjW5FgtmDdSL8HDYyibWx9
pDXhNz74Mfuml4uZ8zAyy6z9KdLDUw/cu7Cj/vE7MXNudKbOxudzu/uaSwxjLDL8N6LxBcun0q1N
CXOf9+Ir9/QYYMzldTTd2efYb/ZZB0IXFs/WUOzbN7FpJqddiLnmA+8znLvOr1Pt7RJojzpTcopq
RPfpAneO47PvU4qZcazHHLQxJW+Bzl6Jo/+mBXvzgBtiwLvdEmD8t3tw758NDzyrN3ksh4905AUf
ClsMBY1v6WW/iGKiiqd7gKrhzDV12CR7HzZEPSjoW2NQ7EObT+bVMxaNGh+qG51hOMgsNluFbVrh
mnLDoHIV6NtDjetSgkKOjJAw01sxOzSNMbJ/iBKA7Ea8ELGC137WpYXXUk46awPAJlF9qjZhjXIJ
FWvdnDtmQZKqwrgvvvOVvyjq6QtiLJY4mVI2gq3qfb9KABkEPZej3I4X6IIH5wEK+nvWEtdADE3e
i+BBkvPYCWkvausuGuXoDpXgvVAbwnQVfjFMnzBw57jMHImsqJRjoMxldynn1xCYDnQijtgxRSLI
cz1f0J62XfUWOtGqR0vIuaVXiGyzvx1mwyy9XGybvtJqR2P0Oql1r0p7e3HRBdnJbn7MDZiuCR1u
qq6SEdmYqU3aGj5nz4ZlZ76rUop3nVCkZbIx03Hc3aMUMJC0WFYDFCaNCz6tF189kKBy7qL7rACK
k4n7B022n7LSobCqQyMOnE7rPKgxLGtxQWwYWg4GFYUP345K4z9JHUGHiwMIZIbpLrP+ovsXw1R8
XUtg0dXrWjA/gyNgdb07PkXXb7NmZFfzxtf8ocSkaDE/nf7Cu/ioa6SP6tTVowguG8hgq0tFtbYC
j7LaT002ez4dmdGBXiQFZNfhYORjpMM9g6hnlPapl7mpEtJpkfsx/pK2JIUnXMSQrvTQLfaAWzRa
w0qHLwrdpsUnDXSZjmP68+whzphieyolDFMfugKFK6kdWHFVfvSnOo7mP7uqTPh4idFiFhMaFa6o
8CoiJlSfKQpZxnIrA56qHZaGzCsgoJxoAifOKULL+uMnj+165ml+/yBLs2Vh6z0VJI/T47Pjb283
l5ofrzNEUcitR2SBfOlZle63bZH2DgCGLTkCbbGDwWI2dmw0F8yTj1OMY+q42ACuhxLtA8uHWH90
naRGyux7UoAbIlJOjjuigx5YjQul/2fPbgeAfdYgs7HI0z/rwTDUux4Wr7g5X8Xss8Iw/fciXvJL
r6FyEBlo42FxuEdfFD/v07vxM0fbesYacK4yRMzh+6u7MpvAlJp+ku3TT6LqbOUiNOl4ldGeLNU/
DbXuSH+aQscJ+zBxrL7I2swhNp+8CSTzB3QsrQ8cMYfKx8cfqqXbDaHlY2B998rbqcXtpaqLqxTv
iG5lbh3EbLTKRVs1buX14HDQPeAMXUC7kz4Y9H1mCdYqJy6JCbLvPGLOQ70B4GcwAKbp4eZ60Tkl
NBfBE90wb21etETI6QP1560+nVHMbWAvSH1QgzuVhrDdW6TIEePGVpWQ1toR/sMJ766ofhHwMPUF
m5lvc223M92fcNkPuXHFBBjHHIefy4GNWIr2O1anLceFTNI9Q+4X3GkdzZ762EZV+Swd5QVHaw9A
TkClw3Q3JBCHUTK6FOjIyWod6n7zrXYrGMCHLVNTIFvWi4JAnLfuoc3+PoA18rqfcVjeWpbjtq4W
ekfKhmA5DsziyVJQjJhAzNNU9iU6iLCsts2A975oxMASnXuJW4kOxsIRbAv9zR3yj6nj/Wmg98N2
CiLoKHwVIqNT/LVade0O9StI6IjX/W2UxxmtOKE3lwNpsPTGRBRbq7tSrSsdLpsxBQvmPJ7LJ/C8
fhaFh0W7gsZbEJIKFhiTeBuBmH0qsWrhNLzMv+6HHY0eq5a2Uidb/DRJbEZBXcst4b81EW2zvwXN
vN2l1EflhNsdgCYpimKuGx9FMMUdIUFXX0XtPPPlvUN82kOtT46WR0jThDObslOyiMi6Uu4xn1kK
/iAWQTnG2JwRzgE+kZQfASjwo+56qG/CqiKIvsTagB/SOXGt8x1XkH+bKU9vtPukk15o0rU3hco+
DXVpRpF/wPYyzQSgiZAJnX265TuWcMF6D/c/4+BJknlsIO6QKz3q/BN1wxthC89s8E74anmOivjT
Ro/8HIaTajb+M1GuiM/fEaJJWnjpD1u1eHpneE+0JfbcYIzgWMp04bg+ShddYlcyNA2mrmgKTd2H
ETmCexoMeRoD2oA1Hkrt08oS+bWGnHBIeQFhbnTqi9VqfDXm6HLaqdXhBr03IuqF1oR+ysY5IYlY
1PbcZE/dtm0foJF8krzrWbZkW/4rD3dWV1saP2xoytXJiO/YGmVtR7MUFyFmGS0WC1pHVRo2vcEQ
i+jT3DPJk/XDUSPF3+gtXjrAN5274IIQBkLRlM7NfE7u9mxfxg09OsgTUBSgmQmxhWgh1KLEmo+z
M25okw3v1HPLKqETeHPUDVLkZb0jb1nbxa3dnb5moes1tfn99bhO50TqDy2fIXnlOLd2HalV2dzX
hkKb+qxnGbFSduhCUOmH3YJaG6sJh/SvT0uzKF+dj98mbQRaYTJtvrNdDV/zW+3LBaXCzylDRZTw
mavlXj9oSV4VDdKKYUKedUUlUd/NvI9pYMH6Pds2uHrE+/pAfWJ7YBguYEBlVF1M+3e/aORiiwgl
CsjUhNI1OpUImLltDz0ppXHZjPSJ/UJFsX1ARrK1VW6A0u8p2DZcl43v+ZJFylixnoww6LkuMGpV
9eiyDClJZm65n7iDo+RKTu5yVmywcXRrApe3tyIlRAx7sujQmuPlOd+JG4mwrReKlgJAMhrdw95h
qH5/CWlGKFeiFnGuTh67qZzAEKbP/ewBSWFHhUF74HaHB73rgAcBlSh6nm3/qHMsO7pCPIbQ1bv7
oTxf1xKcBa9A74S0M6KQLDgusJzTrIURXqxZhUZDk4nUYO6JOCZ61SsYvnbq8jwWK0sKQm8/D9Rq
WvbOg/JDT/uuc1zVI9pzGu5CulpcF5hfyhvSTiPiOd+lv4RTF8CTxsqhXQaiAwq5XlouZ6Cqm6x6
86xmXNipQOz5mRAMAh4o1UVKBbl5NAjJygfcnInuLp/TzUoaVPO2nv755RkAJVbJg2YNBWjLIgEl
HyU1AgnIdb0PTcRyAD0k52Dx0F01YgPHvbd4NLKsanjMOtaG3unfnBzrkw8VVYPK1vtu06oinCMP
7C0FxvUTbTjhsRHu+hAwoB5EFceyFlrdG6lnEgQ2zNfUkukG6MOAyhhA5YEksDtGDbzwEcG+W+1c
pfplk55gJ89nb6NAPZ0m9uJDTzcvSi/2n/AC1rgkrnz7QQZRKvwr/KuuyG5RwyO7TD4UnSQ58DsV
diWgALNm9MUpe10KJHIaBYmw6q/ld/EjYfLJMHF3mpibwRN6Ce/TI3rGR5cNn1qN0Xk8Yea5VRGb
Bp9KWHk+C0gA/NtfbByZuLUL9AA4Ntv4dY2sHUkHMLnZAhB6BewZDTq7ZXSIZwgnjNzLJi+8p0cm
+Bje9To2UDNYSODfPn19pBw8tsQcbe8AjKINlPZxC1X3MRBmN2xiKh1uk9WTOpXSA0Nxpehml2Ux
EE0M14nEP8gLeOPHY5jujtkmEVwdS/8ne3PKEM4VqXYrFPkGCdrw8DnE32E0qwHvkL5tku7BiQB7
3tvij9oLJdRe5b5FVHefge3lLciSPZgZXkAAt/UhZXZvwWhKgc4G2a6j++ME9Crg311a32sHoBVq
5FvEt5HNxElDbRF9nwge0YtqVmDctYNNIwVOHOdCZivfXriMYVzaUMm5heAW7JPx5Ul+h2sYsDm+
EJebIn8Iuzoi+hqFY45JYqS4LdiGRWXmFlNNQgnp4ESYxe0YmhAZD6xvOvgYeLOY8GzWr+tW/XaQ
dVqY5u1/gwmjf3WpnwcQIYFJS6FU0gbzkQIgGIM4mRKgqUvFvqVzg05EAAK7ntz5OiGp+4IRxj/2
ckDGyDl1LqsFyqYUQq87kFeMVBdlpWEWFrCHjqNTCV397GK8/DuAeWerA1mlBK+a63qJe95g2tNt
5h4WxKMQ77akahx5NNxYUQcD2Y448DAQRICAAdcXCtDVQcSUkoEREF8VvaYrzT3sjULg+70AIQ5j
jlIj1rofyEucxd51FsO96fY1SSo5mUtiPcoQ9UsPinNeMtjdSqMWMVUZrlcT1/ENgx+Lt9M+WrbC
Ni3pGR15+5TmO8/7RVC8JI4USIwOcS5s2w3B5Jj7BCwjR3KXKnA9z4Es/HBsPKS2En0ndVshwDeE
Bn8xVlv8UtC00aqsSRC55EAjMEbBw+YRX9yaCLr0/6QrF25KLBoR4wDnvgseIhgMMlLdgVi3vEOA
sWDL3hW4mCAA2nIimoizWzeu49c47Ev0za6Uyf2n11Fxl94a+NyIgmlj0rzB15SWWvpSg390i8XG
LhgpL0MqJ8CuSQa1JoG/mTApTXoqbla1yWSNSjjisjLlpfQMOjZzslg0Kf7JjfDV3+lgzYyqpSwG
zi5SX2p60mqGlgm27NAYuORGl1SZx1P2n6RqnsRJj0GXxJ8EAnMOE2h4G60TXKEUO4WcUt32E6+7
YUPTuG7mYwZU/qZkbnH9sGAM+EeUBreu6Z9/A4yrYYj/4nSKQBz+wcUGHYdL9SEaB4KAkL3eun2q
eyrwRHTmIACZa+teE1icH5ML6KJu47gQsFhwDop74MgVGIEkiKyFca6swkRw8RADw0LqlI0T9HLr
lucqfLw69WSxdMtkLHjNU9DNe+eakmle2uVQqL5f9jXcIW4SOVj93glS6ChHVpIGOMbyh3Crhv89
OmXOlRyL1M9UqWmH1e7qNJjTyQjKLb+4H4WjGn8DVuOwUcoEaCFqe4BLvNMyBEFQIDPTx2DqoXc4
2rAwdleBboWM18HhkadYRO6nTVM/BWsQNPhZdS88kZuHKe0WVWRdESLbCUvikUeGhlRwFDK3auov
bBR8BYFhC8mcYpes9YGiRZS1cuXD0Jz+gY0UvmKoVMHTY8oTTQDbQLlQL17vKdJMhis9DEGOHRZU
+WkO7zmKf/Aq3lS5B7AY/uEBYcQvg8bok4CNWgUxns5MJAz5/K2DiDrPyVgKv97SOHsCwAkLR2vY
PwLJHSlwfSCwjOTUu1oD3br7XP5CXK022OEWTm/tK41CN8g4vUwv50xvGJLuZtrZVN0z1gyv0ofr
8JyysHTJQzmRcZTNmynfQhCT1bl5xPkFbxPjJyDboRDNCC1JGWh/FsXkbqFzQc7f5D7wqGv9lSWs
tORvSnu0SdJW7fTTQQ/FJPVf8IuEB7rm+nB2sQu+NHd23GQ5Nye7pGhbA3MH7lrUIaO6mqWx5xvF
umdWCfk0U5SSAS4e/0/TA9l2RR6au8KSSecHMKW4aTkyIOJi2R2WXxwgBGzdYQVU2ts15SnpyXip
MGLi3wLefTojQM0zy1B93A5MgYPpXQZgb4OOw3whtGuOtp/c52cR6V6HsHLez9LPhTZcLlb+TodQ
AaKJQ8DIfluF2pLnN53ozQozpUou6Hozu/QkNiipZplZHUNCBDJhxrXAvrdEmWvMJ0j8DhykHB6U
WeiTwkCG2LYhv8qRXDupvua0P2YM24PICZlF3fEdNayIBl6aHzMGybn0a6YTMlrbxwGNZ6aCr7KG
UFRyJIFINWLiEHeTmNReRq+UE8VQOjOiGjZbSu40LzNc3eh3tPorMV9rnI8LcGoZX+u9Wydi4FGv
SVTjwEj+TzJ8Za/tD5JlbG8WCO+6zU+R9kmeazx/KodtAD7SVU3e0I0er7XY9/fEK/kc/V2d5pYj
WkoRMn63auW12edCLtcmoqZTBUArfeIquYt6YUBjmt+qBi907EVTw26vNEQ13qekbmzfrLwigAut
bBP7LwvnzGozfb/QqsnjH/w/w/OSmSykFB7Mw8orh5XiedaCubhzQqQ9OUqyiNoIy9wEaaI4a/f5
suQ1yYfQu0oIjfPbXyn7YpB5oe+ALP0ti3V5xnjeVuZYk75jV0KNM6iXYP7hoQ9QVmpL/wWuM8Cd
J5G0GrIy57zrHVsR9UZiaveTZrQrLy/lTVsVMHw3DF9Ce0aXx+MxpH4mkYiFFa0IA8b+hi7jJN67
0zn+VgVPubukLsjQgJ7Jw+arRwcwqAcxTdvbvqs6mue5hREuGgyc7zTeOF8JDVS0MMYvjshYBVq8
zavl9jf71qpFovfIDJdeP0gOZN++5YFjs6t/4kO9jzZrD9k6F3bibOzizjsGMmBEgIqWtJtUCkqF
qPtCka8h5FP/4nRNMpy4iI03Hl46VeFNYuemsDuxuc2IUR7w+Q53ygnAea9V0Y1KKikFJ4rP/ePQ
X0kQN1OYFfGpVpF1Zz14KLgAfqHOz9jRJy+TSBCUzj2a0TMAqYpyRifxIXQEPHlVi6JB6aWvmLuw
QALfNROJlJdatKbSzujTDcOtiRvf6JYTMrE/RX78xybiIOj2zfpM27kH6UNLuhnMkBDU7wo4E4Iw
3c7aVtKRwVVTgrnQUQIrhkmEBx4pbEOFY50CZll2/myl57+bi0/zak3M4TheX9Nl9+G0VJW9WwNE
RVCQW3VsDjfqYmlNthds6SLaWUXFaF+MGGcN2iNGlIuyf5U/DAD9fToMRpNRJBS3aFenQrWcoDQK
BWrw1tSVsivVN/rcPmjfuVZFkq+UgqRN7Qd3yNWSe/cL9wh0wzCEgkygfegcheokOia5qDE0p3qd
0YxnJOvlKq4o4s0gpHaqzf881aX3iNEUhnTZElqukBRMtYothAfZVHsYiABHI1lbIuanAesLM1ef
D+A+CBuzRioLZgcrySfVksB+FcXdXRDfA+iqJ7Aw87senjO96oHgNQ9BMyib48xL2Lc9A3l5F554
rGtvjOaBXhgRBVRO10KNPhRHSfYmmorI7mUZUveBWHXQxNuiFyjiOI1aTPrTlEmve1yGYZC3h5JN
sHysUuaDnZa3q8JXjs0Adad1HE77UQ5vzbPjzsvGZEGZ1gJeV4E1jVGX2hXVBdvSD91axu7zrT8J
Y9RPilbgYVUAC6Ua7dV60y5w1/EImaL6daCKpQ0mKJenSH4lnHRTbix+Cre2H4dpiKDoKRILHeEG
LYkw26R9k73j+5ETeuc0joWivUDzg5Wm8VUOj7DyZRiYIP0k9UoC0BzHJGIClp7nl/qqX7di5cA1
snszaP2+PCq8gII8SnUmmq+5t3UiSKUXyWwFmatqyZ8SK4BcR8wlwMPh4Oy+OB2H/dcShf2Y5I1j
vcyKSVkqkA+qDcpk3YNzgprySVKG9E8PxvTptSrOjBB0k+MnDb62/ZHPmTK7gj1fPX/LjcEbDTT8
vIHCHtcitENedJg8CtCFkZYYpnUgAgLrJwM8NbBNJFYdNmmWfk34iIS/gLTIWgwafaj2Z1TmcDLd
5jlrmcxGgm3OWM0Ow4ctiA9PvhdEL44I5AjNClbR31pdGkRZxgP8uVE66QDCR2nEcVq7cBTAG6/z
2cE8E5jUZO399pPHrDfNcVfy3oGbTTh+XAI9OGUw+0OJJcqDRQrhlUH8dt/odBm1g4ZyyOZOfwdj
Q3ecjJ5RRQjzOZAzW1bGbCrkS89zFpFrkw2bol66uc2dtZCQpry5pHAIikZF3Y0HeadnVkdaHQYI
VHgnJqZzRC9UwquIYEMfMAu9V8NbAgwAXn4piekA2XjyRVdwj2/hFKEG2vcphsuK5noviZxuUze1
kZB6tol3MfYNH6uT1ROimfM7iRxX9SqZ/OU6GvfffWAiAtViGKWdX8EU2eXzb/PYrE9a2WQTQXgQ
2ghEvCtwNh7/9pHaxlLbvUGuFoRBdLxgitbLTvZ2ZZD8/+j3APNmUfLzFiJHGjNXwu+I3eGbX1Ph
vKI90CAsHV8WyMXQWcT0cyU7fhHZ9CUPFIoflgtJk8FVFR1e4QtFKCBnYny7YeeY5QABEWuJFKzJ
9EFGIVtmwCb+VVBfjAM2cZOV+sIGRrH9eQvlda3/6WQQsVpjXsFZh0+OvgM1MnCYm4GyB2OwtrIf
dPvFQaDmJMO+6C3MtIOwdkcP/xRlsBYC5HNwCKvLqRobrqMOcIf4F8yaBSAaS0CJIm7/OXhA0kgH
pFuT05M29/jGJxTy5+muWhfQg7SqArycsdwqb/c7bx3gix3cFpMvwiwa5UYKeyZjFyl5lkgLqKhu
/jJR+HW6wnLUWv5rzvTXithK717WPBepQgg2XMmUTqGkuPqN0kOvXuop+d26no4kJ2d81QRIUeh/
O25zZwZ+jR8QL/MivGBJ9NgYHZN5D4GLktQvQYmpGRGaE93ghFbpCbFiYbr+1Lth5KOm1GwYef17
p74JVfS5/QQ1Q6+lwsyYeOAciJaFO49AgUAUpItWEt+RwlqIQCwegOq/wvK+BAm6TZRu664Ofnnj
1mWYfpS/uRH9ddwnS+G4DqWyiFMBeQZLBIptf1O9vV14X01JQuSmmaD7NCK/WL27ToCAEQnjp1NN
v30yaXowZhS4jJT4l7XDrSs+/Iu7Y64tchstoJoKip0csBMculYKVQ3QI/HWnvWH7kYhWVZEGGex
ufQthzaSl9NgaYPkMtK1QFgA4bUx5p8Rg5w1+vXBPEgtX1ZGDBplalcM6v6L3K7cZSgMom3BshBl
Uu6iepWAflnPmAS+wAgDACHugv0Y7Cj2r5hTuSQk6pUDRvHlOLJKGb38eO8K20NVP4q3N6pdgbiW
BKxBtcuHh7b/0Bz8+LcwL3F3YqGNuvUKhSjMePZiPUHtUejNB+5UwsSQaBUbrW1IbWh+qdG40+Zx
q+sGn6qyY4IE17whsijzFHDc0xAl06Rr97PqFud0H/faoT9A4aHTCWOZS+AolXXenMsmYwwn6gIo
C7yFg1BGzngPsIyoCIeGdjUx+2g7e5y80nznb9RRxknruUSXYsWUb4CkkhLU8BwsS+KnTwNO92y5
ymcxpuvIwFPQje5pAVnFQp3n0LmhBu3yWQeIZcRZToeqXp9LK95OPaSLBTh7sjeBUNkees2Kuv+S
hpBybXd4VbhqhC0QH9y2xSr2xcSJzjBL6H3MLqZoDrvYXmpTvGUFpeyCen17UAcELi209cyAhuWy
4fxiDpS1ydcHvKvZUnPmCZcaaNMMZx8OffDm0GFkJ4O+0INeJRKcG9zdfIAJsPtigAlmoqzjTgzt
75+3064Y+ioMbIrLqqXB70YEQm/Mek0JShi/vb26xt0DYBQZIrT/Wr26jKK8gRUA88SZ0G3f9UNF
Ys/8Zd3WFXB0HsN9peBIC2iBUEe/FMBH2w9l0qIfzI1/KvJdYpWhAg/XsR1+IbPzfHsjzxutY5Qv
30JGGeiuyiwlHCJbg9h26elbMk8dvlzsJasbXWYBd/xKUfqOTKXIWrMm+kkgCwHB24wtDivnGndn
TNA+ZIyMg1GhAWyYBY65Y8fF4k4H4sNnk3z3Hv6DqhWRQduv5tE/z0TA7QrVpJarahEssigkF+wB
jHgrPCw0H0N5zJ/5pXtogbs2uDcFm5NjtGOgGFIUz7LcacW+wzpLXsemzLbJIaf7v6XJ4akrb0uY
JMJkSkBDpPR9MMc2s/KXOt+wUAznWJoC3BjsBmpgZDkB1KdnZCREbTQlsQc8HFROFgL90Al0AgDm
L2Za17xGq2avcj94E8ZrG//bneuHUghgyyyEWITGtH/HAr/aBvCh9WBoiuy0vX8XVfZH/KQz85MU
BNiUdWD9tEbZXlq0QIabOU1QUn1jhfjWwzqQmYyHrFGTtYKdrO6lc39lVM/csRMTv1gGCKGtOnEA
wtSOpOLEZJ99ort06pyLDeopnvMDw/2Z4zzvNOl52AfQYGEMdzb1TlYgM3NYjR0VommFan09tmia
Mk4QkkyThwms7duiwne5t4CgrEDtQSD8HDGzHihz3UgIYUPDjhSHfqh9VfnU4/CNQl9sP6+qeu7Z
T8yl9ZGky90gOmRBpE9AlEXf2usU366dXokL6TkEcSxbL4lgnb47ybX0S2g4MNjtPH6KWgozOBNm
eYL1GayIHeU7qdc5RlQCPThAE5wXMCQTAhf/MWwe93F31egOTAkjSRwTPbeMnVSdiWQbDT2fQ2pN
jWWS5DRyTi3lSvaQu/9sY7tEzIGdKrf2F+b11ZwZniRyDd4VO6BO3B2LdpzpL7oFUlouKxdECVYZ
BKN75H6OUjfbOVguui31S1XCDR1De5ga3bsjY4Qe5CoSABmg6zZ9JOaBnJ0jx/uITMVjO/8Ihlro
IvmzsMQMUoRu1v/V/XyT80Us0xqzFcAmj/J75glK5oFFht/gxoR/DSZr68pLaqaBrjc4+iQGxDRi
4RQlsJvs1Yy4qPPycrmfvGiD5Dh2nx1ddrm2SJMb3Be3jiA94n5t/Idti5fvGhh3LCei16kuGE4R
v72z5c0/43Hjpn+/6QsOxD33V5tK5kz/AA8oDXeDfTOiKqNVQS6iMX6zqy6oPfHpQ+7J699clj3l
hCQfoGBge5dg4yUnLUSXtIKQMrpPbkksEwqpaT+6x1uNO6jZJuXQt92rByLikdeFHYguAXI3y0Jf
CEyjc7pJIZoEpxJzvq7xIvmPQk6DJe3/c1Xw0cDircl3//2VwQIUsGZQ5jpVNSocUwBNfWaWx0qX
ORoggUuUvwO4eFdCE0AkPVaj2TPoofR4GofOdnoYga/HvKKRonKJ4ldVa9VHr45tBtHAZ0ufbNHG
6pu6M7kWM9Fnn2bOR4QfUudFpqjl81x5FI+96/Nd9moNrc467y77U5SY4DeaImemqSZ8sBBAKMem
yMdu0J9hfA9pKtJW1LLFYRnWIYSrddyDeVMX+GDEzMfS6BoXbMIl3A8S5dKl+LtQk7TC7L/lzROG
5C+1BZWksAy9w8ZGiQRyi+nPztmxY46e3lGI367GAfo74TWiWLMCiC8QXR6mvDOpYbhSHPeNwvTt
pNJi74V2kbvR7x3fDZlFp3RHN9u97lhQPLzgkNIRQigK/FJ8PP+zG9Lr+XKezZF4V2P5vPfczjVj
z/2jHbbwktKJ93lEeD582hQ2aZpZIeq+DWA5GseY1jqtsk0dlTYnzC9YswUJHFd2aPmQ6vPxylKS
k4rZBn0B5fmjpZDipcTlRVDIMIBmwS9O8peGKkhkZenuK/IW2rKEID7oT9gNSQgWHmd1P+H3mGk1
Tcu5k6BT3MbGpH/b3LPmtJYsqqNzYrTpUcThCyvsGGUhOSzv5wWbi5vUXP7d58aNRc/CQ3jGeHRh
h1OjcXoc7J8Q6WNPFmq+JNtGjyaWpPOfsaBvFsNjQJtBIuoAhg2rtMeHTj4FN5Ck0bi1LMMxiApU
WFXWd0ZO4J4Q/vJW7BNg2jxDFWJzqCVw9qXtUxhIByNAykMlIUN5i/smsPk7GYZKU/Kr+P/NYa5f
0QyGV1yJeZWtvrge+2qFVubAz4uwC24dUtb89sJAaiZvlzoqUs5cOKhF1EJQPojSfzHBm+P/+Dpm
ObxUTPhiJt3SBf5jFRfKIBeMeoPXy7CAsr3SedW/2kjRiVld8JLbFdw20TMItuGsUq2RQg7Y+Q40
8Rf02yWrz2s0Wal3vtZ0knN4N8eW8JwgQb1Bk8u3sQZf47p4UQQ1pR2JTt/yyDuebwfTxP1UXgv/
EBZLaGLKO/8XZL3X7DYChJQGI8fb1ahEp8JS9uenylN/cbizhXdfqQjexmQl1wxM/Y3arNo0w4ER
yPnO/rknyvGw6nVYKf4krisQ1eiFJaXOR49Y8WhW2wNv56qe/tpOWmSy6/nvM2ZsPMv4LjVTJp0C
FnT+TguiXRYxagPAWNJTO6HMeq18KYfGAIyAqeyRcgnGdjJWWpy8jPevecfFzxGjuZIrtr+IAMYi
TGA1Vp5yXOF5QdLWwDR7Nsz6XUYwmxi896J6Lupvw2/5Ow9Whm+RK0nYPN05HfAi+ZFmiqgmUKNp
Ea7Ws3z40PBMCkSDDL9KjGKW0IUTtehbb+ZNHjipNg6hCVK29M7zaSi3eQdcc2/lDHBTs0mvVTzs
2/wkPdk6/+T8ACMNxp/tSpv+EkYEbPA4LC5Dt/YhduPK6p90k4BLQRab0c4D3gnvofDW4+d2BagJ
dASr3hLPtQOCfYm2B7kn/R6Ejw8ubLygT8nugOe+VqdB6MkHBjRgAGiBVTCVUqvrc+fq1RY743tC
BrtLBFZyt65eoaG++Dj/yjbI2Wzl2tGpKXD8Lf7X+jhz0/Hgi2fuccIFQt6bimkhmUaqMd7gAyHN
eTN6Y7V+QeWPXISm947wp/3YtzLO1EwPZVKiybzgfphHwwUj0sWpAZh8bhhlBSxpAGMC+AQc8vnk
2UDDN9987XJN0VndCInF0WgchsIlQdx1fgaSra18Oql25MqgEAvVDw7Jl2Vovsrz3v7wLoLk1cEw
wgde+WG2cwAiKf8P7/JCCVWcK8LeCC7ZitFeBsfa+THu5G6CmtBtQFssTLsjCUhoyBQQ73GqCYFg
LAokwU6khMg8QlMJEKa7X+9sOTkswjkNHUbM45ilWt1msRiMZS2Ljl+xJ9eUDilOAJ38Y1Xi5Pai
wSUcroiVxp6gVZEWGoNv+t8QUNLPnvuPpAs6/0cyFWk+K1Edx/xe3oB2Ff9wA/g3c7uS0V5hc4ob
TEMT45Cms1yiSHCrPIMSWu/YJJNM+/R3efIR1gwkE2xt7X5NaUYIFXYSC1lkfY3kmjwXskzxTAH5
gjsLwqZAxd6dGw4ccX0N/sUKx4NjCTzGJvYVl/YNpKjuZJsoNLxwxNEUJ2o64alEIREsFdLrDrdz
JHPELZ1KPsw+qjGfeJ9wlafW73OY8ITm/JA0L63v5D3GPrLNDQWMsTK2OuVHSSj2wOuPrvk7Jvbr
GQonvBabuLzd/UzfU6Sr2ydmAtg4NpHOxnYkaY3dtXsrNouLuiz7QLBf1TJ/tBKa86zn1sPFlE5B
EGV5KNDn4RhJU7MpVffZSctdHt6jE5N50aJrukitABbwpUHyLXtp94d5DgO1Z6B4bx27xqrVTC+j
Z1I2nsAM0gptt4BhUyY1wbq7fkR2N3mo2jklDAO6fL4m3J30EOAuYdyH80WBY4KxflCZ+X9+RE/c
OdQWU8XTAMT2qNJxHdkhBPiyJUTGMUli5LH1+a4VM5cGGuBHUQEnv24XhZeOQO+IHpX/bPzH6+Hj
bg7kSKxsdLqFnQotzkxVJ0FI9b8fZoGJSK+tac5Adiz02keectB+ms8cQxq82+j+hkpqS9YguzeL
dgbJeWMtEZ5L9QNGGVQ8JLNj8b/E9yUIo9WM0ICWjqt5WoTBfSu8m8nicrzXxqcmOuXbFl72YfB8
y5c1MdQfd83aQHIHxwMmoAgVH4s28cuK1EbnEDkeGZnFyqS4EGbjO2pDAVcScLfSHSyfl11da4O/
yo3+JN56rmg5jsWSdvnu/siB0tLgEMwCoIZZKJXBIvKZ6qFh4btn+wc7xrqpGfJByL+oE1uzBu/w
pCN5ZdpHVhtriq7EWN2kIoPk5wT74E5aiFS5ek7ma1QxHQZgl5L8ahuebpcj42sMhNWKu2eVQklN
0FOOH9hcu3B1siT3F5BkwK4FjjgBvIhY/BWnCtIkweBRpjQZoHqwzavzi6gGDWrbSo36dR6rxbRm
Ob7FQWYTZh9/jAgZl50QdV9TOIkt29VrcmWsLEyY+TMsNRutM1y0j+pxvj1NQqt5bc4aPfKf28a5
FbI9VEH5er2dmq1F3btOwlVTLv59Hd9H47e8I5Ub3BzwirwtuAo4SuYE84yj2az7hlj7TAoBBoLg
PMH9ulqSRmy263PajfV9Yq8LhhyMofK21bBz/u4VNpUeabfQxdz+QpQ2tRtEPP/dhgRouORZWIaf
19WEYGCkp+4cvzoy3NCuPInxaiTaVWGsoIZ/8FPeoG97ouL3BSoJ0mFgMwrl6ebFbFUXuv5F8kkC
aTTQWdax2dxCaLQkbEJW2kyGlB9mBSQj9XphxduFenq9N7HSvQmcYawDTJHmqyh4luuU/MtwIL9m
SJ+94/N5AXZO9m9bgoxvpDbXmtmhTBixBQrx2CJYi+A53arXvdZC4myOBnCp5m2GDB2WorjNbj//
5MLakOLgPL9Gw821sf8VnErNNUOpZ90xFvDG5Nw+YAUljMgsVV1SDG73ER90Hv7/s2VCFhzZCwKE
g1L7uoZ7phNDC/n3l1f5ts2ApejVlRaMz/+acH0pT+gaP6BobHjnDdZkfNt23+awz5O4lxp2ODKL
uiEoeyJ1r3hg5+OW2Wz4+CzJMKKeJKPV1ip6HLeVJUvkE4KxT+j/G2Hben6WC9lbQySLQEgI2bVt
CcQjUJW5NbfUVomaxrYe8vw+1qLx01XOVamiQEOIUPotTSJZhAc2s+al1r+47oIubRwGVYJd3Yn0
xFb8hgey7h/1aSRjtuJPqE/typ09s9v9yy52F0H43AlkezYy07GcbpzYINUCjO3QPPmz3oB+uD/+
2c8WA/rXVeg8Ege8XLqwVmzMC5e7OzvnE7+zovCDmVaRuL67FhdYexq/p5cQqJqDBU3uxMbpHHgH
W65FNkz55ollzkK0DMVsZd5W3W2WFWoucw7SkLWkIo9EQDLZDCyaH9OZOMUq2hIcr+nmeqsUmaXy
6ObaTKTnnK6+pT1m6Nuo0WfI/0TCLDegd6OJZFtw9zgVjHsx9sDb9bMf7HtpWFxj4ATHj6/etqs1
Rk1P8qouWjbyci+hTb37ijKhOQPKOZ0PfokHLrecahlGHrHYwdaivWTF7enliySD+SsoqjXgY2VZ
xg3xofuPfgbhq1tluzzXBdFW+PVMD04qOjqoQ+PDxJ3tmrBe0+b4dMxMrdT9cWZlfio42X7cmsMJ
yF1uyxFN3Qi/pTcaYMMFq2GAY6mSkJB7kVSOWcaZB0kmw4hf4I4Kt1hj2n1l1jYTJKLBdixiBnsQ
t/SgMM9HgUZDGI+QvdtmlBlspemfFkpFskLIBEafndExwGdnuRzSgHIpKpr2SidxpOdR3VJ4zfN8
s0FziQGBRmO2/X+/Up1Z6s7V33qlstWxleZg9uuFRTrXTPT503dF1bNnX8mBtUzBit+hMsvS+S37
beLpKmHe/s+VORZNFmhndbzo2gi92tLhkUSkGQ58gvmPPvKZySQDCNhHuYbOzVWZFWQuP4lvKZzg
voVLlmtZFy8veVlhjkHJ5Z6KVTLvBDx0h0ktOJPc31oOuuZmhR3vSnrrKdGlEymhKD9AUub3/qrP
qAigmLvG5tKTJ/u6p0atuS4tZ3tMOqNcHJaT0Ke0CZq3+9Q30QMTuQI+s/G0GsqFtFxMxorVufYt
dCk+KT2MFxL/KAKWcN4HHcLYhEmBCjiNcYCiX543Bl5og+/AxDwlKEg0tzBZMwPT9n53TuZRqBVI
uuEACXBX0n31XoKy82bSDUU8oI3oKElGrdHlkidXcP+fkOJRXB8ZEFxzFYcxJguqLLEzYKGep6f7
iiETl9sbyRiC/QPgkAiyhvFE46+gV5UMcTWfs+3+ubT9PxHtw8NWbi/mc9LJXldUHpdpNNbFMjp+
vrvJylE9NKlbcb1DOAA0KXyM76/AjvL40F7n15OVWoCZu+REbBFbJzYyI4GU3cc4enOaQj5KZtDW
r1Ad
`pragma protect end_protected

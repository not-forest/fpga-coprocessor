// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Ud9vz1hUkKH2+1gUeLudqjyiqZrAizl5mSsE0xzNTpuSc1AAou2ObbluCSzpJHe9Nyj7fHIthPbF
O0vv9cF9Xkmh+3+QBHLytOOJcfGymjsEi9+76VItH9nC8Eji8uyg9Cijwaz02cqW4ZtxUVn0gjSq
wfsF1IDev+MTR+eIW4jUkzVsI9SzYUzvvu63IEOZyYw74xa22lOSh8e3NlutA7hNDyhg0FdcQXuu
OK55Op8WDehoLqN5hmWXZ9pW9boCMBLT9mOrT9xv9+9NyXG0uLHTD/+XYnCa4kTpeJhZBXtb6Dk0
o0lHru0+k5A2TrcQKhDeBWfco426Wx8JWCj8/A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 13840)
nteOUTbcFV/BtEPDxhoidHxs3Ql7FCB0wJu8TPg0bc5Zgya7COgjuZB++JOOQ5GdZRnvuS/FGsH9
bmMMHc0MZoPSs09yc+Ea0l/jRyOSXhdT068vwpddN9RaaYU2Zaw4HaQehVY6HNLEUGviXavpoMLd
wfvB3AY0/JuxUDhl18fQLBZXkrYnxsnjAvw2ZZysPB4c2pJt5yfYb7xyEZ0uvEJb2tPIFkQJ9gIl
jqB2SKsKzxDeu1E6aePCZGL/o6Y6XYbuyp8iaRmBcZv2x5W7V5+281EtjlCseFSGWYjud8QyM9uN
Irzlz8FyAFq1Eiabg99goB8ev7d7lUEctCZL7Rwxp8dJOMwZz2dzdJokhnymqUsrJ0Wnr+TpHzEO
NHC3h5kXnlNlfyxMs5d9yrAnlsVBeLIj9dApOshOKOesGYixCzKWGEuDeqXSBDT74NEl8SaaHr/r
KANm5Grs/5mpJiZeGUCCX8eVwih5HIhdDJiJpHZfSYAPv7v1iZx2vaKmRAsv2sOiVQeba1GvwKQN
J5f3JIWMCwpBqluIlEbvdNYbMlAMPIdYJu6OTHNTqCSIxORNgexUu+z2y0XFWZaHQUWOvJbZwjCl
opGr/60HuQLhXVtDTAOW8wS8gIG7ZQpu++z8fH6NEsB5vk1wZFETcBXyswJ66k9OmTpv0agReb7t
DMDi7Voxf7okvmQFd/oAMkcfe0IZzcxjMEW+0PbEq6sgcB3ryQBnIVm5eqVq6KNCxdAvPgDSiU+/
6X0AkB7BXdmnrdrAUdxFf4R3zp3mKLiUAUuyl9ctpQUq17qgabvmO4pV5QIIGmCR6VTPZW756wr8
Iiza1qlr7x/Q5IwqkdWYIyCx8jHtNqurcXDFwllbxc6Rpn7xG94FO5/ouQlrcxnZYil47JFVn4y2
7ttihliloyPx1vhiIF+6gEk53Fy3KvLBOY/PlH6I8As2tJDTvj7TlTUnSE9fD5mY4WAFjeAr4tm6
vr7h7m96SR8tfKhTmp2gUVUk/ucaOUMfYlEWtZD6HnfCcX5aS788uBqRs9J2lJ3pJpCucHGFfnqB
/5zgM3QtrBwfWOrxfgcjAcdYl/QtqNQWbNjAKp9QOQMmvyfzpD6C45FTVqOxOWCdBbjgPkHcwkjO
ktOSpHeEa/3FNq2bJJRah6TCVxCL/yk5rLHMAPv8Hjt0hZOVucUO7lXoY3WDyNHiUK5XKM8FwPbd
VUF+1kDMJFQNUyXaKL7nwJow7vkX+sWUOIdfWIM81L+cy/mMWbsCZNGJDl8bcOzXR/lvTY4+LsNI
1LtjhQTDrjdi3eGDpGKxEEKUWdoMylCeNFcEl3WiFQhyuxaXjGsSQaym2Uzpi1wINZtHAY2/PMtj
N7koojp0S8qYqdzumf05ax9NsHsDYB1hZoS8LAqTroOCZ7FzsBGtYcNudzQXkqFW2IlZOo/XmTEk
DlbuWf6g1/ZiBMBoSuRN/jpZLi7LAhqSyTcAyT09q8CLDMDs4KmmKVewLGXGqVduYXpWjbEi4YVz
YRzHJ4tliwTzkguJ5BlLYXu9bHSHMDGmNHWFcEk7x63nnndb0kSdbCNs+jGFRLhPlx9slH48oXUG
yqxF+mzNpdDR3a8vCmD2iOMg2e2pkTQcKTRyu2J8m+Ke9iiuOfcgHKkkLuerApIpmZCNyS87mhWY
jjSrmZNmpRz5bd3ahKJ7rEOLPCSJCKHSwrdd/17yd/lROuP2QPCla8gg5yXmXsa/v9y16SUgYIbN
hf0X4LwbZMWA+K81oiawQJc5G+Tk2AcxXkV5X2CVVEGQT+zvmo5alOU0qFzyrUTyjQ0W/olzGxQF
WreP9GLmiBCyfAtkFSrqGf+s7t6E1lXdMzywiPZLvqksMt4YskO+GDYNJtKOgHlzoD2Xq5tVIuyZ
gUO5jwhMv21etrIDMfsCaFXf79ILv+9gqrzhRukC+9Nr2pI+RYRHrw/mA6XLikeILLGZ61xS1oDQ
IJDPOkBsQlwI7jFU9IHE0vdWWDUPLfme5adPqesDOiwory1OJ3dCz1rUX/tVkTBXssNocNM7oSNy
D2eM2Qj+dV2INiCS8r6MWRUdTVP5vZ81FmiQoaLVZzBzNPju6VVbtriIUeWvRiTtwK4oSOzk+/Qg
UZWq74EHmxE2w0sHQOzNSot5kL9cDXPdNcS7U5l3J0xoPuHZJmvNrCzzn/07W/PB4fvdi3rgSZqA
9NVIqzDj4XHZaVZklr8XQp0fj01Ltdn4T7K24Ri117RWbhnBgKT5/Om5q0x3M3TeuVW2qSxTSBqG
pvl7lcv1tMMxQ+4mf5h/gqVLyAK9Qp4eKVQAcjTJNgCcFj7rEYw25Amo+JbIfG/qemfUxmQJxqJ2
ZofGF2ABv9VrOyT+sjS9LG92DrlzfFmKfEXtRCklTBzDYXXcxE3TCIO8O+2lf9MM4PL045ipbziw
4p10gG1J00R/pJGikoDELYwwxnH4O1YP6vKcHF8/gh2lhr5M+65KAqTXiR+uTkrUjTMoKY+04Nyt
EVgDlsPgyl5Xt3OaeDduTm+pPYZdGbHVxlxQZGjR83MkSimf3yTvJ6Rt/ZHK1YKFDnZcev1blV0e
O/+pJNifXK6Z+L2w56uLAJ+QYOq7ZYLqPGs0MNKL5uOYpO85yCTPA7H2Zvv4MhvCKR5DBVZf7mf8
OkOOBIQ5Nt491RO8f8AXzw5feI4iq4tZ/Va+Z+qjatqpZkSDNyzYLkI0ggPVLVBP/z2Wdt4g5mbG
MgOoLdXJ19ZsIU2fovkIJYtpxmkoxxPr/3Bf/0B3bcjb1zqnBhdtnW0CBPGnnJLvFIId58eb8rWd
vHJv+TnAJNnHU92UeoxsKEOfdve+n1BpOfIEhX6nsJoRJVLpo9PhzqX4xP1/jIXKhxpNJDhx2UoR
9W0Ln9tGPB29WGTXBlauIf8gtLIQ16mMS5DdcAnlffdEzxwmGla5WiDBas8lwt4zpo1fGP8GB2Oc
/RFU23mXlGDhtl3MOLGtCqXliyF5tMaJoWtkxb1V2c7fYOM9/My27glvcORQobhAeaVXwprB0DC8
ZXngrVnxwVNFtbM4PII5dVS2aNUGB75D5Jr6euHtxaV7uCkqRAkM7iAFrr7aVhxoHZzlJIb19DwC
WiThA3TugLxMgBKfPbozcUNmJDhe9818T+fnNhcQ/N2O06gzdMc6SgD03A3trrQX56y9ESvMGMAv
mchDSI63WTjaJ1tNPim+qs+LcgwFviDCTNAu5bUFMzFhKbQA8AjSbfz73qvg26x1n28aCpqlf0iS
hzMq54KcTs8SaMZC3ShFb4IqdLhJLL66MtiPNQ28srD0KWmdnGCN9HZXBo4+xreGkpwx0vJ5iuK4
1Hd28G/W4qLP+d2Y9mgeeCfSpPwaoL/eqVFiN6+jw5Q/J+VWt+e1rahoTJzUzrZ7rdC3NgLYMTHG
ol0Bezs6xownVh+EmpuOyUa4RiN8wlfLRnXP3t1/xX2yebKgfSPNhsj1W766w3FxNsmyY/gDYxfE
OEdYyMdxUfjBKWlAztsKz3M87SoJMgH6JfqVGfiNV2E6PFr68Am4u1Tfdr/y8w09gaQ9d8O36z/1
vud3Bj+M5uVLcOBExHVaYqRifwg73P2EogbGqGmev94HUDU0po/M6FklIhn/lIC3bgwu9y2ManRS
rW9+cRR7V4DBPqGcpkprLVhUvIl2sjNkZsyfnx3jG3HsQT7Leu5rkxPPs++RaewESaYRuMP+c+Gj
wl01U6JT3qWDU/ul2ar+6OvJfxIqC/hNOEOP6YqzIqwkTpAxSw8IueSHLr29AoAdF4NedvU/Omkp
MmgxZ9k9+MTh92BQsEcH1LR0ljwdBudRMCeRlHs12NZ5Ue6o3F9tDvBlO1/NpOFbFMZnujiKHX8h
4jw/jPkfaI5b9IKRxbtyV92CQtYwL8hQ+2hvRtiZgZ2vNeeQCDwZoeBYT3DyCBhhAKFZE+Oy2DdN
79mZK+v2Fv2/SQ28CJNylo6wkd3nhl52qn+OuPQg597mugFWp2cPlihKNNI2mNYQ3dSTUZFqcv5i
KJxyFbve0+nOT9tRcA4uHPBQ39AZzRcM3+Sb/L6kYBJOFVVa97pmaXP7lEZr0WZ0GWPmm0DW5mW0
xIBAyE1TwiX6SIznF8ElD+0VA5Blx3YIPEH1VBN0OtJFJ69qLmRkBij7f2Cc4yvnv1BPsvpBPqUI
SPyHl/3EJcFrbbSZiF3X2M4X/ym+lL3puTI/Hyj6J0OflqMKo5Rcp7XV9C/LwOdBsAOp+QQPsbkK
joJAXAcU/7wzmlWmC951JboEY95J7/n6BLXgbPLF9z+yfLrijQoRU6b1v9thNsk10em/OmrXkBgp
WihF/JOMNGTZV9J8MRm0M3rjc8x+6pw/lnibmVCHAjYFTw96pJgyzDBdRcbJWPFPPgXCfH+us/xo
D8IxH76VX1BcpmjynU53f8vONxvFCl7w13V491HGLgoKbCTamjaQEQdzcwO3k1s4t6KBufdZMdBs
HN2D6M6c4gwTML1NSu8Hg7DpF7tHQTVdoqC3Mj2XPeLkwsgPEM5urtLHWl9j6LIdhA35bDCt9KPb
mkXd2JZzKxTl47cNbXlz/W2XCEbFXWAyBQqhzglGqoKc6C3RmvaotDfouN5ewUxG7l9Ikefkc6xe
tkKuVs9bpsP3BxwKVftJWYRo5jf8ol6xQfB/WCI/DwNjR3YUGiscFXJ6+HJ+8nvM/QFeWeOxh4BE
w81YaAgDBZOZ+1Gb1U/jDeLFJ3TGn/L+GN41qa0cBGGD+My2DHkCSSEOye9krqKAWEtBcZThAsix
Yzc/g4ctPaGKTMqkKVMZBTImxRBT6OkEaE0VQuSQk7qw4IhlO91pwB8fiFmABXhY/UF+it4flGAK
QTJuNRk3W9ke9NqSFpsIVrt0Haf5sKKEaVgaAUZi+9c6UEbDiIFIZ+ACIIoe2OHCDWYCZt95uhhe
E6DW9cwhKmGyMvQ+fVBY6fVB8rPnOX+k04sKAA43p8kMDxg/qKkD27hIcLQMkupoYHYMu5//zRt7
b3IO5ZIAsVs3AGvGoBq6sSFir9ysNmEFRnhzeOaDkICrKflI5x2iUzSl94kjnSPNz0Ps5HmEQzW1
SvboaH6TshSGmFXkGvkKA9UqQE3endn2CNqKm3Tf13dgH5g4dS0LtLHRA0fAagSAxH3kC4nHnxn/
8qN6LpX0JXbESS0N7QseanpFR3HV9/stNM0XaDiH2c2DP9VKy4TyvHFOAs34iZ+VcJ7SZnz/diS+
iyJO8wJlibop8yl7Q3Bfq+CvrFOmwmISWEVrsCRqBYHqiTGUiY86a9+R4/agLKZlg5EKIk8xvkNd
Jb2n1J77CS4S8NxU8+MAT6otS+Wkeq9c0L/4KzqnQ82owJavyIgsW12N4XisBQPCY4IUHQeXMQgn
lIBjq8yEOD464uJ0+L78RqNTf4XtREaqo0+PCmA/tezx026MRfbs2gWiUiWgOS/8SOQaECZVmX56
DjlLP92zHzOm32u9zv2qSN0FuybV3UQvLTv2OEy1yUukTWCamAO1L0/UMCuX4I4P2ymVk0L4AJj+
q3vm2OLxVnp3ddh1uoj99GC0z9S6MLf58/AofZsZuVNQCfHh5gSv95sl6C+GAg22gXBJFfrAJ2BR
2vSCydY8SWwzeEMS6NQdlOkGqkW4Bv/qx05psU/FAjfOzo8SjYD0OMskue0UJuRtarZFUunrFay1
2BRgSBDnyxcZHeL858Ara5syjQy7lcd5SyMXxCNhdcyJodl6MI6zAgUsxWzQjkSnWtbPMCCAqGbr
giJptBIe8XGUXEpdIJNyj45Mugt1OuMygmlSsCRQIld9bua2Y6bFd7JTjNpPzZMN6KFoUmvhAl6C
3Gsqh2G4FiwOkSh7sMxy2/WFwArjBw6IUVsJsEyKZ3SdM88G4hYP+yTkalE3Ih1h8IVO8D6j7wzE
wrjVZME71wRNfgYOIyBPH2mgKEWBuCu5ouJEK/noOt5tdGyDJb3dAbLV492yxUaYXPnaKNr2XP36
0CSntR7bn1Dk1+H3mThLeBNytUk6rQbnW7/EgweEii8zJ2F0NcNFc6Ylw0OuT4CnsbqgfdMoNVoC
b7LSMW/Fm1fNUNAj4qCp46yszxdxbnNLSbBEPG8P8Q2SmiPrWUXdgOESNRv2fQyBjWnBHrpQz2mh
cjgIAENKbsLOtRGosLEeCxRl/X/jtq/jjc8WyJ0S0zxI0cSGo14xAHAbo5d0vAvQ8Iwq+kGy0Qi4
uszDBWzAaWUlEaobC+YeB0c7Zsih9eXJmCkntPq9MmwUdoAqueJ6yAShqOpGDVzwSpT6vRct4HDb
VWsD/yit6TJiTyZkE4QjSBecDz0mEuQwy+C1EYpKNs8DqDibC2KD56JpXqqculQZ8TUAvX49lFgC
QUTICrsLQgx0QXgbsb/WMw3xtMymv+rfo2FBk6neXZVPkde79HjkBcnV7GEiJohoLw2PyNrZfvl5
Gda9cVZvJ1Y0bZbrYrw8iHAxqTYNRMjoWGwB/VJrHKufvRG8DIJZIFVSiyTxhXXBQXKqExgw0/2V
QDczA6wWOpCBbbLL6OjTqPJaA90/eA2Jf3JZXTMU4nSQsFnJmwIPCipgV3gaN7iRQqJyeclv816N
CSCFqkLYykG8t9XKEacA4FDD0z20pkqN6wi6lJm/xo6joLx00y2rexMNaaYFDMAHUtUg8ZIpifb7
U6QlkzB45cdroXX+Ey2rE9HhiZ1IV8qd1IJCHmObX7dSn0MRLRkJ/zGNFze2AHpiBH5rojilLhDX
VS4A9l82SzOtwNpNbZ59u73k4Ot/CASGQC9hYHwDFfBS9qRGh4uNxmmhofn7gYyFEaoR2p0fK3hP
o/8LppEByP+VSDjam5rZMXxXtLxArnJWfNRtnOtAIbXBDeJjFilpUbUj6OyOtHKqcCbNd4FQ4PBq
Fi7kkW6p1ydkoE+d7QYxDEqozgY/Snz0COKJMXGmN4+qdHamdi95/4wuKlGjQAD75pAOsglfo6DF
AVZnyceEibW94/sfhC3u47geUG1pYhsRP99MMBcjdkcTvXJpQN5Drjb3DXIblRr2YvkoNw7VMJFF
13twjM9PFn5TOm9qlw0V3PnXpwnRSYRAo0ax6ji/Q2wOZfasDxCUQURLWAbbMtPI645XugQCQ0r3
EWdIOXKOJbXeWvk/AMp8ROg7JLrrxvKr+R6SEbdsmMRHU+KhMHSQUO3/8UJ4TBnX9uoZ+QG/Rq79
pMWBdHkJmdxpqC5pMaO/dPEkgRSVvkBCOOB+8JFV159BMkrasFf1yIVSGzYvimwPWbkJw1lmEZo0
rTzw6sFpvu12sHBwU14TcJNqKDzKC/psdYPo/ipOZzMY0/pOXjWbBQzQUnV9MtI4++V4TXLpahZG
QMckNDf2wfkyqHwQJtxP3ze33iTM+2DN/4o6D4Dwu2yzPL85Dcf9VqID1nYgQtn+OQtifPCNodiN
Q6Bru5OmR1G6xY1MSGi5czFFP5O7JrWvbsOOYjfWrL7UxQzJm+aNwoi7z0geNOJMyt6efTkOfnDu
RfIH7YG4Gf15KLqnFQQDaO90adB5G2go0WoQamDRBc8TyKtyLTU10WPNVhgf6vIsOLYuiVov/U1t
g2SxhXgw3gDLAf9fVQ3zhAqFuRaImFZrsJ9ezKUGOxl48iurMojB84RGfuTTTYentwbGSfb8Uda1
H3o/rUhasfMp7Lg2D/tSgkouqhGGlbXOCzW9FZ/3tvg8/tuaNO4alaEq90uX2gQMmiefhxQ/kTJk
wKvo703ctEdMbCgXJyWEg8ezXDcqCqiaLPDVDUyQI6w6BwY4aSAwSGQhh8mIaFD+n8eEoWmXKT/g
Ky6YljNVYU1nMvHkMu1a0aJRP6SsJ1DK74zVyZK3g8lJ1RApRYj7IWJF8FJp4HdwxyE6DuC/UUnd
9TO7Pln69rjPGestCpb2EpelPht79z/XSFtyFyTlcVO0BOg826VP50j/hrltjUKvVh4Do5HYPSz0
ihAOvRT/IUZjTaf3CGQZwMTPBItZ7xMm+kaCnssuzXC+WOrHJ+5snOg3Qqr3zz6H6s0E7PMiYYQU
hD6ZEyXf0P4Ti+IFScRJ7lrSG6n2Q5t6GrzLh8gFQzfscdrW0Si0cqWCfqipNQnHL1thb4+q/mt1
2F+BfstctK4LMZu/hB5q8yqYK6oi7ewrELXIhWl6eC7y1t5VTHv3UJcuXF0SUZpREPmJmwdUHzi8
CylFoSdcTyj3eM2vx+Dp+CWjumq5sp339YNui3t4yI0ZptUvpeGH57l9BT9JwBdnrG5H8MGcKEi7
aCEJT1dldT5kpGNwI+0xsh+Kh3ibDgZQDxFiAcbnhmfSumpgrf9eQvk+qhYScJfBVroVT6MoX800
On14/BfJaEixt9ldhJb416FQPxbxb5GHHBtU/jXvGneS/rZ2owb9dAO9amCRA7oFRs4XCvtMefEz
Aw5CahPsf4Sy3zOusLhIHCNaX+PXDLpXys4ncE5r9tIg6qVFtLmKXZVVaOEWp4JS74kFtsw55+Gf
X4o+Runs+c5gLiyslQ5uzSvNQjXMDB35DUq8Vq7NWbmfnnU0aM+eHeiTO+xw1LsAWz8cQEScqDMO
atlMWXUYCj7cv9Ziz9RHBTASBYUdMubu1LdGGBsHplZ65fG4hMuwA/byc//bKSPZmunbyWw+cnAv
0JpvqxUrNo1uUIJoP+OjHEk92d6Mvvb3FDPmFQaF0VwDr/vuovqo61ofQ6rgw1izwOV3SllDWlgv
Ody4/pctURngqRPvyVinMlxOi2huOToob+GbWeHz6ekznbOn3+Zx2GaVDz1fNAYPs7dxCv9B/jmD
NQg1i2Nrsehpy9aTadjUW6B4daUqUCQFMPto4vxQBpq0NZc0FZ88ltsGMcTQe0WQJE5GECpcib7U
mGkUQPbO4lcQ10WMcBoU/L+D4lj/ZXWRAqT8oRapuulnnur0wu+1GvO/uD0roG+43fuTTUewq1IU
AVRcIMLV8dkwTIGDNnEN6GfyZdqJt9sHKc6xc4XM65hbo5Dcz4WY48O13HTYV2LPyWrDiAEBnMXp
2UkPLSvdPhhONAotD/SQMS85J/cMG0uvx6nE4MfcyicvY6i9Az2JE+6TI3zf9+Inj3bE84qoSymF
NRAlmu79gUgeN6f1IP71MmKjaKtn4eBDJUY4/XVwZzU3DKrfo3NGzBBfykRr9GVZKwAd7vfcj6Qk
AZksRLMPls5bqqwNc/OiY0GKXrjrOzl5iPysi8ACWkenT9AYVhGfbM3ulANhrvRceYjoPE5Rxc/t
eVUmXO81aOSUorDOjshjNibMmmn9eOusAlYu4xTQ+tanRrDedeLKfH+Ah2jHay+ymyLzYCLpPqJr
aiQYLcsLVZcxUtaRsh5mUhvCK++nqMGoKihsqnlLQm647tjfMJZJMokME7Wdpfxv/1skf8uiafbE
5Q4ug4nyFXKa3ol9sdvWM63p+gSr18c78AfJM7dVS2Fb8CO0Sr7ngoARW2GKqVV079S1wOOFZZik
RQHYkgey48Y44+RSxWFUrO9/vKukfmykiI9yMWt1cx29vkfGaSRO9gpQsPYxzR2MlHQMh9HWfkeZ
g//52Vb/+nXXDWyPjtWCUSOso6CAmjW2AU/X8ZSoEislr54HQXVlE+pOCEGN6rvByp5DrlYGBE4b
6Tc6hWYx8Pa2KnYKaR5ArFLbXflG2jomguaxqD9XpfvN8cnIiw2HdwYvsXf2gN6nOs9A0ld2rZGI
l1h7ubNhKUVscdTH/IopVmlSN39bvoRJD0ntR64Hq9TX2I2OtQ56HsQuDNPNfRO1QaSTxd1pFpF5
ztT+q96WRctKEWWG5KXGGm52CfvfQG7Km66WOl/aKqxAOfGusS4Mzo68jF7SU4vraA1LHwW8++HV
Ez3jquQQ60T6aA4mnyNG83A1IgL9m+s23Dh2nVUTyh8kcqa90PMhcX+dGrmZelaSBQbvXDZUXv26
CTSlHmWsee/bMeL2k8OtgF+EYCmM21f/YKol8BCIV0dzwJrXNr6VfjKHKSOrO6E0dcVH0Jlimdt+
zhQ2izv2c4XEtKEhTxjsnOo5Ajuepj2ynzr36dG8nPSDEW3eImuBLb6jvZgrlbYmpUg9tlU/YfWO
1HUGybczOYboyXMul9cjQBZ1Fd6sVLiQzTNHSWBTZgtrFIF1zWM7NqtMaATQUv18b5UU03+fRLHy
wIuwWoxku1HywlDib0iel9EK2+c8PfRGUgwaHDKhGbuYIhBvwmzqwCW3uXWwY7dWV/N1xS2SJKKu
YrFdQXNUKSCdDFf0dXsmS3rO/VueWDIBnW5bl6R8+icH68qL1rRYGOBqdCCWooQ5UvLiKrN2KDph
BYKWzq7IJuD4DOEXxGabd4FPh1tZTS7E5cy8JMYckzGw3nXYim087xcU7vz3/CcdvFrXU+EiDVsk
uJx3X9w5ZUixlrqtxRpdVj+sr2/6v9u9m2kh6tiZmLOUVdYtoMfBaieDS/HRdW5Fz9ciBIDp+z2d
/+ZeEJGr2jxuNjmpWoSI4gzF7FCqc1G3gRWEJf7W/tctuygTAVCg/+YNrC8YS2YhLE3kr8CbXCF0
Zog+UIYsMk5aOaDIx9xcjyfzN6bp/Rt94KVczKZshva8JzBKgTuH7M10/DOsaFXANflHBH/Xlw9y
XZRsZny+PpymkdJp/DFXcXM/2afvRpX0O5ICbWpLZXCyNeiMx48BO+oCpddlplEUE+Cgif6E92J3
/Di7E5fa/nU7exLp1MCHHzZJUfpVQYKHCQWJaXn6WE42lvx5tZ/oE1pmK7vMROvQiDqB6LHUFBcp
J+hUzhwEG4RvDtdcuzb4IrRb3txyY2zRUXtOWweI6PLAehwLn22akfF7wT/MsSCrTq1qJU0AvLT9
/Z8+2G0ylac0+Cf9zr9qPIApyQeVYvQzDBVuihi1n/1eL7KzfhHNk93BKeQDgdNIGK2wxCTIjqnX
4/8fV6D+ufedIb9tLJBS8C1tg7fk26kaqhGaaof0k9XJsH25PTSi9oNRa7UQTp1rMLdabRF5tu5D
gE7pLf9naLbHUvsWhKOPqISP0r8p5gmuR1qKqqGkNDuB0fOZqRVGsebRmK0fZ58ovyeR7VrKNH9C
oH90ymUx/tXcgkdxWlV1dzu+CsAUpHbX6xC19X6uAI0Q+QJvmC+GTxzmJzRwnPQJUPiqfbEhd5zO
+OaJJDdb8XZEv8yPaelq+j9S2+1hqiaUL5DDrI4p62UdbG+3Poi5kHdkdzC5QXX9Yb/U9b+4aetg
+HBrf4TwoNVDGc2uZRl5CyPsp5Eg+O5ijcUtbDFVw1DoHSZJ24AY+b/Kr6R/1BzLyZ5Dn/8Soxmv
x9dqKa8t2htaPuV7bK9IVGvHnzAQ26bzZJbrzIa60UL7uEb0V+i0l/NXjpDL8MWZpaRss7nxp0yk
lBXDDgrQU7Q3HSm0O/Gt+xQzg+wpk3AO5DiVRjELftUPUs5pPVQXuVoLdHTUwPR6JIHfB+cVSy+d
+/RRgt2R69HHi6+NYZRhTueEdqxheba/rpEw05rnX6NlShfYpJGhQAro4YBlbm6sce6WeoCIxHuM
TpMrK83v1qRXwyUGQ6FQtBzzQ07bahB+xwbjUzzkMYk6J1iIQT7EswgwtndpPMRnBiVIJo26QCl8
L12awGU1tfgi8bAsxyOOKIqd37FxE1xItgPcdNTsOSj/VJpw/mPZ0/vXG8T+eSdOLw6rfnREltKE
rRQxvRFRHCqfqqwxWH7CDILwkf+LI7u66KnnezYRLuncXpgjfJkybBbi9jtIiy/4OB9ohAjK7xVE
dXOOOVRB13uGaB9mx6combPqRIsnONq2teLor7Lzv9oG0a8c/zhx9Y6BXd/NUbKS5syO3VDMBYSc
1YRtqm+8+t5hE61CFyftSWNQnWKkov8B1z8o5svFOMjFYqiVbghUmc3JWnpufLRMfCO0t2ePi4gd
pXthBXPCrPmu8BM9QfgItCBW4yljsXWU6rZQrC+iX1Hz4VcXlAXpoZuNh5Ag3QqDe6WKvkPEgPT0
C/TabMd7uYnTmzgaOB/PWAjQ6WcADIyb37CuhrWSeg49qWVG+pkU85TqsBdVqg8PZpda2T+zVVFr
IqcteAvn0KGHGnr2346spEpthdcpeL45Son0Li73e3Pbb27gTtiWdykJlLVe2fyGTtP5R25U7AV+
aGozPJbW5fhLsk1vITB2hw5mui26AJLjIkM1zqu1m2wC+NcSn46Ebn3gLeCrzHKjbYNl5GAsc577
81e9Es28DNC6yfz2F1RRiefRC3oom0cyoygNU0IUMCZD7x2kh5lU4e9lYvE2XI2urlhW0kDxOsnE
a6GKlrXTp4tsDaHPTzk3TGwGIfALV8fRI0l4iMDa7+73Md+9VO2cLbFBPNjJuqSGMBQJ1d7YjQK3
hBS4BHKtD2AfRV8aI3G0U5BjUE2thwUkgaRXuKY0Gt5N0p+odySXrNw6EnYuGPfTPYGgMMN7VH+y
+kHSjazfWGPrirxHNMe70Ng4OOxV1vdXY3yj3PnvCzZgUbvipKoagBW3UdQP2/ZiiYMfCLGaDQXm
qE6LmbDo+LwDtokVGVhmzHD5d7GjmMOtQBPfGqJ/EH8iXguvZdZNGN/MILP6c2GsygYTAQOk4Zo4
eCz1/lgczLa4ymn284X4EpwmSXcyjz9og7aUNo5OuEivi0CpeszTs4EylX2qHgWXZ7aeF+UP+iYl
KH040AM9RUQstO2J8zHZGZNu4bwUQ9OaEGKPjH22PVE3QE8A3+7Gtp5hxK3vqDlZaSmW6wPjkTuk
jkVoBS16bLlkIgaQKk55jGXrqoZ89byY6QRLKwsgD1A9WloTtUdMVPov09M+goOls20hBtjZTNQM
Sm66vz1EBsJwb5IfUgBxPhtVXOnAZSy+/2LZzdN7u+SiFI05HZdrXppJGivsyEoCxXGBwN0ApgQw
eSv1njyoaEq+ABTjDoOTUY2GcAlLgvz5zTb4vv/WbPuh9UO1axRayzuiT1pYOo7BvAbIQkjIUE2b
48O75pqvYQvQoeJdiKSV8NYR0PNGGzyOfFfDbBUtUhL2OL3c5kJoKjZDxK0Qqkk5cdrJn3OEU3bZ
E6BLywnNtkjk0kIxP+sCdxeXqQIrNQaJdDYKQ+UuKAMjNXmgZqBta/8UC7DcZ/2wa7/FXRWvyWDu
e6nD1c0tH5RHY5G7RgK3la66xdIrL4lWAw4XlW/Eeajc7HEIoPC1jLGSwlrxY/swx3lpp4tcwi1B
wcIwzqVE28ESje5ImR0cclmU+Yk1se6nUKhKFXuvJyELI+2F83zViCF/0BXLJ42FY7Hl3WVUc69r
3v88HFhZYPTsJAaWkeXQxdHv1G6jNSyq+ttTVWBx+PNhZg7lNtESOdyKN6vEU8QT8mgh+eyIpe7r
gQ0LrCZG4VwQLQJPOqa5JuKlD04Tngah+IThNMIA7pkwUjTnzgJSWES/N38X+1wsOC9WdgQez127
lwqNJ9qn6tAWcqJAzvfPll8pXi9NP+uzzHaVXREg7lQZj7j1jc2jbrtV+M+0/VsBgYu+oPb7mCBF
LKnymJ1jZn925gMN74ENrWPbnCDL3SHxXuZYXx/FXoVRm57qC4srwJE8ZudNXqCgMblIuu2WIeoY
5zVtLV1A4/+cYfmHsDX+jZTpBxMz/Jp+Nsb4DauKj0Zirl7aaVllDPvpl5kjfE87d2CTzzA4Cf8n
YqLspJNH42fpNVmJ9NiGDvBZkCROU+VwWIYU7mk1hGlwz15ctLERpaXqnQoy4Ax+Tc+tfM0r4s7W
J0FDhpQNppKc2ZpAHKsBA7uKqOFvveipHkZM8dAKsK3JO39kqwaxOk2UYwpqnsZzdX4QdwaQYGqk
8ig+wgQpPcieHJeuxZ2rAoGrAQZKEy87ywqwi/kENpKUEszrn06L1NufDXrb9daEMbSREPX951AA
8WCVYgvVx374lJxSmI99w7Wy9yPGcuZJzr8Xu7NbsiWcDyZ6EvAWViFD01O/ry2P3ejDJ3HI1vhI
HgZbRq5IljchKBwnlSL7Defrz4Q2B6Cztp1o7gjYu4iyHjdKMKnxo25dYw/+Q9i0+JbDH6LfsQUO
jCXJR+i9VNuX7B19zQzpVhDW9cau3fpsIcVh4YelNtqLug/xpj7V9xdk8ij+EWNyfcSFIW6nT8of
uApsKS4YCzjh4jkHhm1kBijNtWNUtAFqLev7co0zf4E+/z8xCwqBvC0y+Zv0+RI7dX9S7SHb1Yx7
ngeioEEDRPlg5298/DPL1iuMCBRgvcCyREjaLBQrQC48MJx5fPXNRI+h78+YAyLbsmFZ2zes7k9d
kVWItzc+HTbbIJE98TYBxzkO1MJr4x13HTYkahvbBy5vqEjrcqgOJSMUxlY6mR4lyzw0BWNu3tmG
DYYDH2rWVyGLSck2ULN2wCYp5okaHNuEINlL6sqKdMvzvA8c95sZv30ncKE16lQXyIjWQb4/f8r7
okHZ6BTR8EY8+sEiNZXCgKywfJBYjvSJ+sBhHN/iyfJkOiDVgLTqIa3J4pAAbzT3upB0Ema+0eJR
tOLMpnbCKo7CrMUHOeQuxuD/3GYoAUM/ziwqv8XTBUL55D+YZqbk3trUm4xNq4POyorKRotekOdF
MrdTdoeKmnh6USdi8POmRq74AGwVUI3IXebJExcaDG6l4xo0wCqedZAPd1yfF34zv+jhYIS3V7ZK
UyhnBHrcZglV2pT5AO4hNKMmLWEd4/ZG0BSDxMfDwR/ReXi/pC0jtxABvailMwYRhAxjezySDOmh
hxJBv8pS2xZy5gR8ipQQ11T1MQBh8HRD6uvVPmlV0kk0DjSFScetzEKKP9hTyw4Ukeig5HQ1+TTP
5AzxhTUFUtW+3AKwByg7lB3r1R2IPtSYtP5jENnNccOySyPIM5XBltCtoUulaI3SOkzGWBQcrUv2
endBEFd5wXz+bKFSgsaAX6NS5hAHko6wbQoQaP+q//cvU+3vp61gLWUSXpxXOK1XhGJ6dmLxp0R4
1PoWptECJ+u1Q/QmXZol7spBdWmRnWhgaXjR/jq/5+/B2rB0bjeHbBibZeU5Sw20Q1hFIjHiY6NL
AqaCfutxT0/lEmoLPD+F6gVqtcu7yyEQ+3nQl7q0PIlPSEBoe2Qz0f0sWx5zMvzsJ/vKUn0dwwLB
ws1K558wZP72vthodCrpaV+TQ/gAz33x1yZR2j9rWRvL7BSk15FtYR1Fj2QCZHNzLUThE9ia+ob1
g0aZg8ORsSKQYE0Jj3eTJ39v9nSEylHv3870Dmw3Ul/myU3l+NxXaEX1vUv7huE9GWrhYJzOQNg5
TcvjNKU/mILjINTJCc1zfLMi20Qs/+FZphm1MMTocv9gzFM58ciOB0czyAUrgCsv+NpawmU/Wtpz
FndDik9W3LJrlmn3VvFK6zkzJLvZh92SuwJHY9hM6gSozUCdX/wSsSwNWJfSzV+1y4wZALw0FGSa
rVjOX99RlYpE4OXad+PFVuVYCK/nMYQ/3MfEiftNDyUJxGfH5PQLmat37CU+CEoidS2Ztch/MJmA
hflSWqW7hi/RNW671XKnoJmpl3DRL84M8LXWANkNzRUkNV+ZV/Eq3iaNu4dZ528rQXqPkyfL9HBb
qcW1RpXTS6k+8zjye1fgaNfTxKoNNd26fugFWi6wOAn5beRN2YYfAwkg9IPIsqaDZVw8e7ZYF4UQ
750nGylC7LjSRv38y3tqzQJscTWcN4ypVBiR2vJNKvYbuUCVrlf5wTGV+LRqedAqXQPlboJVpcCc
baUAGgcLWsJ52D9YjgAwAGHvwzYc73ZmmV3CY4ijTTvJdJKf8gJpKEcDG2IQCA/imUfIQ3DAl+Q4
RVWlMaR22TjzhGp+InV+45nKfeQWpdGIadInoNsVE6QqAgywl7td6NyJbkUaNi6f8ArhcdeS4nFG
UgVgty5AE/dytdigXA20IQD4MsyMO4J3wO2MyuKwM0LzgV1F49ltHf86ourDiME4XOFUcRpk/mCL
G+sFIJv47Gsuk5CUAPb/x9A4NrjajAJObau7YOrJf8+u04KezzhNxmbdPMDG2E0mmsUvV9XrlXuQ
4OSt8cZgGvxrVKMsaVH+QDaxhegBD2FopsAuISfIypZ39i7d80hyMfQomMdn1TDUOvZRKfK+xtsV
ZnOLWt0Xgo32ZTRC+iFnlCEFvro9rBRlmKZbPUoJHkTAHWQACXl0l5F5sGixkdk6UDG4RMJ/oHsZ
zQJCFLKaP8oTqSb6ONqFhaVNwMKren1zaC/UQnqsBwsIxk1HbnL2NufpjnkpCxnIwbJASE3gk1S7
6/ng55yjTKJlaZz9XlCGVUY2XfJjY3ebXHqrUHY3JVmPZIvwxqDbNOKn1xK2rd/M38YLk0fAJyIA
rA4mrBARMG0YTpwNWlbvARGkSI8Cy4maNVxH7IzRaMom4riGr4Ap/aqyAJSg4CNYGNr0H0qlGPV2
W+WLXM4fpZf/0qep8PuD4PvMMe+wqcqOIvf3fJ/MenFYGP7b1s11xmSds1XQKf7iiVSlw0rGejW7
F6dHfbojvQeYTSGpakfwypsX7XCaQ3X/sV1LNd+OJn2afvZO2tDuixzgKrEs5Sa9TaIiEP1VCAoQ
j4OuJPyAJmrBCkfRgtVpNUGAfvr400Rmi0AsePTQJHuig57CaCGbO844jwy4L4FSkXJfcNwsyHMU
qYAI4FKQQtorTkzBpXbXiliKhQ2SozKpZC4SSA+4dH0WfjiBPzWcW7wLa3OnGM7Y+chiQvist52p
+9H8CH1ALzuiQ80pGLtRBxB9obLtLMfmm8FO2e/nwT6EOW2jad/xQkYRRSeVeQoDP1zVvg9EgScW
AmVyB09q1EBu+EoFdCzzPu9snp1DYze4CpOxQ3mfjXfi4jfPeTPo5p/l6l+W889PZPvkf4gJjLHV
YzLdMof5CTxcVOhLSEJbqyfBAQsnd5zFwez/FFrdUyHd19J7iQ1OJ/8Ruoolbjs5vHtLoFfMlY60
wvU2GQayeuFzTZbzCFBBVFE6Qk2KrVWv+zHTSr8VJKEW+aKniSGf0WgG2zaL2FsOLcB7u4cpHa8d
B0rVBDxbWUGdtHZHxk4a680JXDZl/82oB34+v7KeceppDus/IpPm3QQ0feJEV8d0gDm7Ad7b//ih
uwRJzx4wZzmC9WAqvtHRgRH0ooA6QkzzS86OfbNPQz7j+KuYhmjbEkrg0EsfFSxL5NpEDjx+5BMN
J8O/d5MMf/SzhWA/0NkIk8gmRVHT+sEcbEQrDSHaXwFy6DdD/WFpNG6qigEt2gUcuqylS1A82lAk
mHj8sAIxbad7DlS2cIaj49jR8B8Jva/MHgbMQMmshcKbjE2AtZqwLaxHeECSo6aMbZBNdNMUYOXI
YCA4oqwAY8LjT1xaM0Nj+FVaGp5U0uic+NZCIhmgt5g0yfOwWlsBgr4Oi7nfTxb+OMM6zmWwNDyy
i+4psGal3mgSOF3acXNdU541JlmlmRCGo9wGI4K0DMrbOCxZJWp3/jKOygTXYcg4MiaKIDvlKe2M
9JVNrjyngTWEGdKRQ+HB6tc46REfpNrxSpxgZ2pY4Ytx0Bsb3zFDP75DTkq52kAiz/mvQHyYhiki
yXhDDtRYGql9TNPV9p3ScmeKllyJlpav+SfhXg7hYaIrQOYK1ak8lhVRrmTv2eANvQ40Xm/2oZ+L
BpWx5FEmuu8lcujqWobZlTAn22cQgvx4tbqKmaSslyF6dcn+CjkTJZrGpB1S079bHLH8xl3Ah9QY
KG74yKeMHqQIfY8bOB/TAlcv+aIMOSQScYEBPAnFla5zFSN+HlHrR/6hlmN2GoN8rNOh3a/ggzc4
0Sbax/YobpIsDqS4yg7+MX9F+wD37oGCXUwO9S84xVMPwolyHW0U1E9JhD+PpKbZaTxFhUhd03KF
TvLmTctvsgsseInesxj+is9tgyG/ud3DJEynhRR05WObS9jC3ivg/PnsgyFQeOFzk5xiEAxslOvo
hm+YFyHbnYIG5wvf+/ZgdxH4S3BUcAtmOXlCm76AepJbF3Kq8Plbxi7FpoiMJeuD08kd6Cjd5N6/
Os6pi5z0mXO48nTOwGpUaAYp/FCo+9isHYvZ2ZFdcrdEDeDF9ZmyTsCveGbgW4fCtFbxfPFjlVQ0
BByXT5YiRC/8w3GCJfv8bt147ge3rEwFsZvtCk1DwsaO4XQER+20so2fs52pg6I0QUbuJ2oIoFuC
+1pLtLL5FbGyGxI1rknlXXf7jbyIGVCu+AlHEsTuH2gUfYHwIlHhZlBtifz3JiQ6ejfemkyd82g+
gwhzoK2C0gsWeqJRO6APy9i0qzHgxZteBKtgceAcwjFA8Lox4zxjQ9WYLaEBNkeZ36z5oh2afWs/
W2g/Niyv6rdsWzSmMFLsfMAU4pUXYEG5nXRSEH9h6cDpeqccX4EzzoJBkqqcf7Rj0FcsfJHAZt+W
/XDVkY9+HBKwkDTFPi8gQxho/kLi8cHKRARSPpffRFjVJofmNsD6qHNCm5euoQ==
`pragma protect end_protected

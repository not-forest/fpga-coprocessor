// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
GitFu/fKHAlgCJeZqUh7kX7mCoHFGJ3hZe3rpxl9rTzZ5Vp+GHnGwdJ7eDemCbz5
d7fO19fq1frQ/Gx4ADpZpOz2XKTjKSUx3h3qQnJPrR/XVPb8X6ZwfPJPQziBW9WS
dutxSRpbH51ec2dn1gjen5cEXhjLzZR1jjxNa7OFRnx2FURfzmjMdfpsV5yTKr2C
e/s7taa3V+1N6vWmQFFpJ4UynmqJAdDLUfWSK+nnm8RBbYuDzErx3gMY+2bGBxVy
uat91BbwARPZql5UYQwOkoUEeSXm2vcsz2ukRcXb55Jw8qG6QFrx3LB9KE9xa2tZ
eakHOhpS/5+dANGLIgxxGA==
//pragma protect end_key_block
//pragma protect digest_block
Ny2Ci+ZUMYBPtv+AOBasJ8E32OQ=
//pragma protect end_digest_block
//pragma protect data_block
CB+b5hmc7Y8URZ6sEQVSDQyXpfPCZj+3dRABQFXxDJlw7LnOezIOC2nWtz7wLf75
p9FFx0cRBwnf7hdoG6Hk+6cV5xb5FiUI6BQrvRCDSX/oXYB9cUffaLWuixG58Ch9
nVwvfznjrX5Lld3/sDHwK49qCkss5lDx3wnf+3I8lqmD5dFeElr5MHxYBLxcJL74
L3mg3l3cRnR4EIuZ1HXQWgQ2KSt7HvXumE2NPS2gp1cHRiT4feiwopm4uNs7C0K0
PsQWaKeUgGCXUw5Myc5dnavYUJsxLCWOj9GsKGaViF0N+ZoFfSB752l4FNkwwax7
5AsRP3w40mOgVT7wg+GYnz9VNk//PhGJmF6SMr7ZQTwDddqXoRrYE5ZgvnEguICy
U3H+jXYvusw3ruH4zbm91bCEF/6GHw7tVtwooVz11lyKGwAefUYyYlHvkETOpoRE
ZgQEpVaT0aT2FZUFIJDFFO1YFlZUzkyF+zOU94goPPYZ4p0JDGtF2I5iv5VOGZRj
fi5peYQQeJce87bkqdHYutt5Nlj+wXWbp3tDzhJHHUzQOf7A8YKj6UC+5bjOmmeh
C1vgIcbWv3GBNX9zjiYkjQ4ggMxfRgj/llhNbqWsXDLUyigBTXwBZY8UYl8XJhvl
aWqAp0TaVijAvVCKo+rRfA+XyhiTVoH7Xh3YWjOz4r0l4V9f0fFyRflLvUMxRvTd
9rQ9NOcdJGmakj8LqPusAIKPirBlFkVQglBcBGaBPHkJXhMuf218bDUL2Qjz+Qmz
LrzZccdODezsWzdis5C5zHLD1vmqTBFHR8TFSl3Vk8mfOH9fe23Re6sBc987lSi0
S/5/lgV1hABx+4CmoeTdGkAQ0GYJyE0gndqjJU84RgJRkU5tcpKB34ift0AQ9lMj
cjWGi9/SfXUpbwh/XNZpmOD0XcMtd3rFyrVON1yL9bzYtyfeweYPUbL85MTwDcNs
3HZt8xISBApD+Eq4kVjTC4W+6furiFreXB5hyC2iPKIoY2usD6d3vc5xrpdyNqmr
08dDw0umv4zOfe5FS4Z78y17f8jeGcSxmuq7bn3wX3YTN3EiuCWg+pDn4oxKqdFA
TZCFC8OYmb+D7146QIIgUUPyfjtvJO94v1qM4guP2sKTgmjVQMtWZWnJcxk20Yt9
/kp3sEiRyy1fOgtSF/qb4As80S9O1VWm2AaMxx50oAZDDKsic3EWbOViLJ00Lgrr
/zYY3gb1ksel2PKlJoUgV/ZEBwDwqmjEK6uEURGvwkDDOWil67+1lKn00uH1E+sE
Li/EyLWvysBh+itOouuOLJvHSQm9V78er5tqEc+vefWPaTdkGFJhhltVrxkZ3Gq0
20d76ITmtdgwiNFUAV9/TKDHyQzWaS+tWKapMf5WXRPkdwGHhux5Or29b8HDDaa0
hr/vYIHbg+ZAuflrYnMZGSwHoxcI8Fxn0HREm3mTLxd+3OW0/NWFHbeU3g/NcPgC
XE2MQQKA64a6Wrl4iXduDL2jFoB6Cw3m5e/oR2uWUCF988Xeq6lZyDXxzOJmPoRE
msyk9qi5QzKr3vd8yQAuvZ2nAUN2KH+svgpksMHFwJDzu2DwWjegDCJaci8ndRcx
4SKOMXe3UkpD/TupKD5BrEs4R+do2ga35Tq8u+YExg8IUNqTaskdlYFP98RDi4+Z
QcVlzkNVcAPtERLgZVvFCZxVFEE3YN9Af5FPjoAfBAMITpAUJe4aM9b1NFAUJ+hw
ZgzBQf9/k5FzekVTkQ8RWH1adHDLSNMjw06TGCN4tcY1PsJzfh9hAA0EqdtlvMxN
q/JT7v1qpcujkqz1i/l2+4DaTvpBiDNhzpre+XHXYeR7Vv6mpGu/vZ4InFtTBJIi
MedJ2yMXkibWJUos2KMe2Vleu8pNpRNiDio2w57JTk7hadiHt8yJdOuKasAttEY+
ZPpLFrHTTju8u6ktLHwiWigN/b4eAuooZLZCHTSS2DXoXz0uanyxS4i5OWGdqrxf
ENzqGanqy3coSIZjqpQS6ARbvGqsHd78cja34+mmZXEsnto944+dAmtCtqXC2xPu
6LqxoI2u6BosK7YEmJu92KflUsftpADb3SXGxur6KLlhO1gCDH7sSYa6PTrU9Pfn
K1vF0uRUPaf7eEkWpFmB7y3XKOMy+6dF+eK68EQj411hTXr2wC4y/0EP2W+X4590
y9iXuykaM75nqZUdxPWw/Y+0OezFAglWqSxXDmIJX+PUNHnUVBM0TiUV1AflLr2U
uF+XsIEAbD0QkcdlOfBMdckQKJDH0PzNbphD0iWMHexJnzd57aPmxzEKLODbBzvP
6TptRTU6q8qZyCg0tO5uVeIf3kuictTsjZ7fwlI+vlbJ9JyVMWWowIB4inv2AjWH
5URnAcA9p7m28UB8ufOYffkVcPtEtJZqUMD2BpGl6v4yC8qo5wvKbpmHnfaWRMU9
nArzezdh32UZKjoUCtRq6SYe7uXNsyq+jATXL4s9htgxq/AO1746jGqQmW3zDt5Y
/PEDPOE18mUZqwE1pa+ZLpYWTqsee7lsaGcXaMSioi61DiX2C23lDgnZC6LQib5c
LA9LsTjDYb58Zy4NwGFMcUu6s1MrLRYkmlIdTvcGA6060bmQAbyutr0wtZzEXZCD
bt6vmvsMV7U3XGvFf0warQ6RfPenFsui+vrWU+KgsL77dtMpBU7vxB8anh+jh0OH
bWK6t3l5611c4QXrxvR2Es/XPtlThP4BCKOKAYIMrZDOV1PpqHNwjkkKMlRJNE2T
14avTD2HGoHHS01M3+gnaZf4A8BqtKUGX4bJ7JAIefezD5O6li5JuanScRCx16Sf
j7JAWxaMgM1GNasXz5XFnUtFPz6fL09ktli7mpGb3hP5TCKMlw0n+Ul8UhDfGjpj
4M2/pi6tIJbb5PWgFEZNPxF9oqZFfC0NVIRa1op811vbgGYHCj7DzbqgbJj3PVPi
HYiBxCsqKlA52MBRoNE9CCTioMQuFCIr0YXiGmh0YoYaHtoAHXe/wHmwXO24m4OE
Li5d2t2hT0wgCOB+CyfdyuNu5RV8YyhJ9kM7/aN4fu+eRHmIZTyZMkkWEQJJbJJR
DOIGjAZXLibBoQLV2nffbaby6QZzeS3JZQxgCVRdmnyqjP/ywWGV16gzryZrev//
8HKzZNCV6ddzgG6mGAnon4G80QAuxjO8bL5mYSnJePVvAW9mdg5f1nHTvmq1jukF
H3ZS3Uk36IcLWjg6cBalpnssln63kQAdbr6c+9lEqFpDKL8oOnjNDrVoOazKMAtH
ZPr4x3sKUGTUsT2g1/ha1hmAjksfmtVElr1JZjwnVY0b9WViAle2WqWnbhCDSZ2M
veQ153rTwUU4/kATu4Tr1qxzGH4D/YenZ1YZXpf1UxkaDE6cJ2xa3WvB0aY+yRS0
mPCRJBz5ea8VGrj3KpPeou7K43W/lrT+hHYqSh/HBEIAraD7Rd3NCi8/vInNUZI3
Y08pvlHE/9QGGpDD0XGaf68a2PVKWWD5c2N0o1ePo5s2KlV7SaB4P3Ngr872FTgX
L5skpBNg71xHcLyDcLiKDmp6gnc5WNSpfGfDaKh0HVqJTqW6A73AzNeL44y+CEFO
WodldtwtFTWA761Omic3V23sTc9v6C2vfJsEkKHG0NlVQYmj9AQUVShCAq9EdK4V
nIWHwIKDfH0EhEpex8gNB53qOX78lot/edj3B3e8fxsorrrDvGpCXEyht+gdfFq+
jQcDY36oxSg/w3R5S7Cw2Gk9DsKiKHACFB37tXWanKUljV3M/DiFJuDIZk5jrgxj
HhXrY0zyX7HmZA/1IiRFRoTD7uK8Vr70Y3glfIMMuPQ/aiZ9+U13CwPGje8XWKxA
g5P1byTMVQfdKZ/w3qtZHZhNjHnEDO72+ca7CzI/2GF4qbYmSQbGwsZ385aLfbwT
e2VQ8Q64oDTDwq13YYmeGO9ZDoxD/bUZ02qoVkDNFeTEpujAa48u3KvrsaM/a5RJ
jK84UnJv6lnlPPQRmsE4B3spEbA0p3nUFn1SSyDy0P/gk7tUDfD9O2DoC0hHMUPD
5WLmFQPUt1SXYyW/UFC/dwD+o5UwkxswSLXSwNjEaeb9EAAuqwGGnn5foIzriMtu
E3D2FRf/6gQKJjtYkIHTn2vN//d23vYvIJExjuqG5n1wCJf5yrS8KO0NQKR3rU9l
Pu+9mEOTsLEhpWgJYQ30MnyIw3NWMmV47aH9vnOUSsu8BTf9GOOrN8pZxGQeD41D
eQA7hnomGA72DzihuQ1MD6uOOHNK795s6Tj7qm/xCj8tDoEc5sVKAKC7y9fj7tL4
+iQsY3xxoKyY2TZvHsrMjE7mzKBUHD2cszntNStEkzRG66gQUllP+EjxmubUNE3w
e2+qGLm/vlFbGDVzvPuXsw36aoSVBwIwAAoiNwBw29qkZOliwwEiZnO7NdnWN+p8
ShAOmmvtYfm7+0eMXOcPaVMY6mJqmmxn5DIxzPpog4fe25hF1/gDLYiyG+f4S3EA
RvwqE20tyTrHu3o6AAR0F8m/8u28V0i3wGr8v/WgOPeT/jFDM/aDp20uxmNQ3CGn
tkmgssp/bT2V1rK0uRso1SjJ95ZEWJAG/HFEYC3eVUKTub/n0fjiiTNFOqOF02c+
SxlISjR3Ah1PT9srw2A22bd6RThyYnnDTiXAwlIG4173ptFlCQuXw2t/NJlv3p6l
UUMBBuJA2Ux6ImQwzBp/M/jI6PKLWfW1LuUsOLIHkc+OTKk40p8O73tNTRQRuhTF
cnyBGQa9XD7zR/wrAZqwmw/lNUzz4kvIYT1dnonhXRsqYPn78PkwHH3ZWLz8qhDa
vZZ/gw/SR41tVDZ+/F8W8BK52kKy49eU42NhF/AqPDG9B5G778q9LUjY5JH17BJL
vq0ZjOOWy0J0wo2KDiW/4+Y1lqwGWgiDrw6e1WKnj1AArngx1a8wn6fGP76uJsrc
qtQLBWjf6sm0y7dqrpKchQ7n6Rmvo9kPee+rasSlotGzq/YEMa0p+t92hcEqziI1
kP11NNpQcZZZLxaWEnxI5wz4OPYT1UW5kvRKLDjXTKf2UCjBPC3Cr/JamYhtkcbE
BelXSVFEfFIz5SO3KIepYJvoh+BODuTaymlYvMHBGL9FY6ewRbvNCO9Yc6RITgCQ
lStsT4Uz+/zQyUPKE71LltQf6dc7v5Q8L7OVl5UuFESSixPMiHDHGEJvrAZRGPmq
fR6HMLUNV1jhkB4KMH15ODN2rG0zvnrSbjqhUOLSy6eL4vEf1ZeoJnA3IWQbciRR
89rA244BXlcZoIQX6FSaxThFtlcCncbhgicMX5jIV8GBXjswHA2bC39dztXiMgnn
JR04GVKf++25EgtufnEZokaZ46wKSSATYomCaK9NcGdvNIkI0QCBjB8gsnZuyEVq
CXA3UZ3fPkHSaEkFNjp8ODtwqCoCk8RGGSeOptARlH+yC/Qs6+Sdv7oxu5XDEBHB
SDEPFLhMtDdv0hipRC25jsobmJXCT/iMdbyM645ngUV00bTSvqcyGWLyK12J1d9/
jU3V/tKeXlb5uHlglg95uG5b8TLJ5fSwxrEQGnV9/VT4zei1bduzsMFk9/Olokcf
NkuE8jXyMuXTv13WRErgHySx48XyzHu3sqj29LBAASoh/uGDs/54gkvmcX5yQPro
hBTzQn4jWi1183PNLszq+9c8xDDUZwtfcPSpFrJTElRJiYEwuZMZFWmpQf8sD1ee
TjUBWMd41s+FNVBegaR19bpXJFEyAfOMZBRXeyV3W6XFcQ7wjUrgGs+wMb6dnsRC
ptJOrZ9CALw+4vDaG39SGyPtIvnkLNdLqGpajo5jYJdZCOmmfo7YQWoB3nYGnOxU
vNjI8w8gv450KoOu7nQL3MNYIhoSWqigxzawWMMkySvVG+kYLavMqXMnouwWZUPl
GssYwrc81qKKbxCHduLAy0cO4J4jwhRcfE7RnQZ/JNmTK85EOoRQ+aO7adfspXUD
HTDAncTs3lPIfoXa254STrz4asQitI5VjSKHLjT18wtjkoUQrmouFHUaJ88hpVWR
2lwJA8KH4NSznD8E1Qh8QZQyrPoXxnBGSS5BpzvYE6pvjw7Q6xe+JzOfCrpliZy5
PU/NZ/c1EFdSDxmFFIv7nwwM8+ADOJQtjPtD74FR95q7hqHEa5vVUV3Y6HI8iZDn
p70ZmNZGlin1ZTIHRLY7uPYaCkn6y6D1l65qGqDU37K5fEPXlkTNvHuUHyWtPrFB
VOoafgOnOTw3e6u0EKnyrVST56ZxLWRs5S4FYuBEeYV+McDmZy/E09tafA6Y987S
cX3g9HnMbQy4JvCnRtQfDr80TuJIV/1ZGS53tbcSK7yW9fZAzN5TY88wF6yiweNY
W/gTx6VXGVcwM4tHZEXV5fwsSHxmOupIqkUwAu+H0TXje6Bmx3igmgg2lhg5y/D6
GsdqvbrVLQyG3CUtbpb6VpnsXBXZsgKt023qvj7LDL0HT5bsgSJ0IYLmIRe+xTrH
3WZx2SZo8tADl+otlPP83QSWWMmsJGtDddgcM/kiEKRPJg55KnUkz5ZXDYy2MWDP
S5IUQJaWqHhPX56FlU0Po4umUev6y343W5+AQYEsaMlTmEhJ7uLP5HyHXfdvEp+l
1kzfmR9if54A47l7bDtXf6Vercpz0/0XmB3hCxNkwHi4y5rUR+jmABcULvRmubSP
+8AXPLJZtYMr8Z88tEnXENghWWiYelQAynJvVdFdSDDIaDEN+X3RE2gz+UKXn4+B
K0pKCE+PDxu4AIdE2lqsSH052B4iYBO1X3iROViMy3w3oqEdcRTdfZ/NUiuOOq7X
RBFBF3mXcK+GnOnQLOmpSa95t0p6SzQe5NOo4FQWi24FI3SQfwC8h8xLTGyJvTg6
t4n8cbhBSskn3L/vzne6jrs7KXmPuYpVEYDaXsIF59HOTRUnKPGC6fa8OunqNNQg
VNgMgOqtuwNigu+Sq1AsiJMuA1KsTM4tRNfJnBzUo96I16NRZj6BMr3e29NBwCE8
4XK0WOASFKfesWOKAi1Y7Tkobfqi+s/5NrAaHwLvakjXeNbZvBmVxknAxdaidFAt
kWmFBahShFn+hvvOQadGuQ3nqPX7waLRSFnVy+moaZrxACXHpNLQTk5DJIM/rA/D
Ekc7gTTuNVKLtMrs1KbthohCoWGDuQ6l6NznMjr3CcHZSXOUZh9KxMV620kiEyug
rhav0nPkvXQzqPObVZobdNhY7EfQMTwtUJUCdFEwl6QPTNjRBgIMgZVPZ1I6Yrs7
JOQo1dEDZSlVSaCywU9ftMBYVyW9riWZiPMU1L5FUViKebzKwqQ1FqEN0CiZld5v
DvJuQAjy/kvzftYKYIAI8qkNWXyXBMtgoG2K5GtCLOqRiJKPLaV3iokM9ZD8pEMm
tnzKp5NjFGh+u4DPX4PAjaSwX/0MYNN+n0tET6sjGlvgcXeH6ofa+r2/DZMbLy0W
Bnoi6mbWJ+T6AR4TVSo5aDYDWKvhM9f6Kbj8yphKp5zMMt9gaVekEfctOVPjnOwc
6dUUdw1C3lDbvsV6BEJChhJz9Nrm86FAnZLSAlqp7MHQB3TOuLhPRqLOQ2zy3dqN
I61IU4DjXgnRsFI608ZX+XEUGT5iYkGti2tTcy9Eq4F0l1jhUQdEPMxvY5Ci+pEV
va0Y7ZqrY/sNjY4/ewOjkU5tZmA4SlHsiuYAzyRJQihQRz2uiYdYn+x4ohf14RLB
Yq7XvpPtZGMDzcEAfG/4UvDb7T7ygkWj2P7SgdqAEybIYFAQEZZJ4KjNE+1c8wR9
UgENMZcubG9jjqGHHvlpftu402bNz/TucEz/+pWXrOo65PQEWjPzIugOx73v4r5f
X395ns/93G2b6RtibowqhlCL7iO861dSrKqmBixjY49ixgI3A/M2gX9xGjW1YGQi
3G1V22r4QklG3m3yfmQlrT2wdX1G2owH+wuJDTyahRqU2cltBXNXOAG2HHa/TeZw
NnRtDsJTmoTzi1WSBODIUkMySmNKcfsxbeIaBdgOHMM58yqkslsB+j4eYcCmfSP9
BcV6GgP8kfn/4vohx5Xjzc4oiqcMeFPP8iBMzh7VVDjoqsFZr1S1JEL09ttzUdze
7wo52nhh01z85F/73JLe0zRzDDV9aAUBzJlEo55MGjJciqKH/0IkZXi7Y+5uSNpc
gPiONnNW9eeQutEwd1Wpsn7tetCt/OWDMahoMZm/Idg7X71AhGc+ZviBiCPfvsKa
4fnAdYZ/gGccd7drH1+3bHZS0A2+Z2izy0n86ENB10Qccm6WpKqvvkH/tYNYF6T4
W6VyOWWz/kwiBdYw/FePSnRsL+rj1JURrMyL/zgLsQISnAHVitq7/BTVRMI5alX1
ncWgMvBDXCg51uVlofg0o24f0M/xR69tRnN0I4FqYaJipGuWXR2ne8PogIbIRaVi
YkXVKgtS+9I+DGTiTBac1IazAS2fqtApp+JeDYxdub+2Ge2D2lomyuN2430c78a3
xOpXQwbcbXj8aouZkFeQnEKPog0CXw1Y0nVIXU43H/arqYqVs+4xULh+fq1tD6p2
+fuZkhbD4jpZtdr3Ept4FayVhHmQTG8XovcgxB3tFlCk9NHIUu/t1nCqiX12pI2+
f/lxeoZWAzFOy6HHI9ycoyZh78bfSnozKVSJ7ntpIaa85H2/oP5EnA+dT1YOg/OS
No8yAkEb/Y85vduFNJ6EXwsN6B/OP7uz/1tRoaAh9YtSYPk7lRN7OFIPaOP1Q98d
MtuswOqhXLL1VpbbDpQSQ4/+SZir6XKXqaTTiyBym53IMpcfR1dNf7lO3yOCE+qm
NZ1AqcG/gSYuGG6eIXzu0yKhCUHSiZA2rCx6yaS54jB2WTA2NAK7kxB4Dq/3LuR8
Sb71sO+1OH68YRLPWWGxbiky/qAQ6TYNf4QrDDpev8uOe8690tBXpxrh2Y9fZE3k
GofZLlvec9QC/0O7YvmHf1vo/0WQoSBG2OtopgsolLKc1VLq9SDlURI0hvE9P8dm
xkaX0ZhhExXK1oEXn3ZYVx3fvGvnDysMpfRm7k1ChVsuW5jZqlioqfIxRjKtqxWf
lg0kr54KoA30BNoZEF4N/F760CQ9oHgDJ8SI+nRmWJVbIiTJNJP0G6ciwYU3ydp5
YDgfu5qHB6tcaYXWDRnhBAxq3e9JjiaVeuygpcL5tq1PkbNNejbMDOJvrDX9TAmL
p8Fr7plTGf4i4cYC3625dRoIIwhcJDv085JflHW6Yw0azl2asQorKZXP6UkQCCDk
I+VqvlPqc8igTujCuDtaG1XNXYWw2sU5qBppWT442tyKYailzxXpTXVV7R3fBZyL
qKy28FmgcA2EhHHO5zInIfwk76cD4Yh68GhvfyafqYAPLnHRUuTiQ/7JsyC7L8/E
zbClwnWuIUlHIXPfxF7Ba1pAhzqy9/y9rpGOku+2jC9W81yqvspIBgdW/+cv0f7U
qJvNna5TBRFRJ6mhI3jHQzuGi3g8Zp9BdCCbTzYbxMTX6FJH1xgE5iTkTzZqg0j3
4qQJSf721Yt2CJUtf5taRqtZQXLZzIesWZw2ZHmgLbITFT5WRCMVPcVA+dFXWTXl
nvvE55UJkgDTEEcxiew9hzAJmkR7d5JwR72QX+ubKMDD7EEG7GbhbYlzyWEQfiXm
xi5tP5Z5mPJ/xy8Al+Tl+vVQN2SPDgEZkv8zMSKHzQvd0Las3zisydLAhlamaXTm
1JzzqwTbfnmlXypYteY2wg==
//pragma protect end_data_block
//pragma protect digest_block
+Rzt3rKlYDfXP842vWRiXGPP694=
//pragma protect end_digest_block
//pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
VQK440ubw8m79pyf1CmeYo/25xy5yuCWHuy+hph9KQ1q/q5ce5kBs0lGbITRfXQBnMinFvRD+7oj
07bfLvmqRMhP/UgzRQmuIlaHKGvpSeshIXee4V56MdamhncqUF0hgWHgIBoM1BxfH/6LzRt9wtem
rSHtN4E1VIwvcCRNkN7tejSJeSHV5KRUwML0dwJMIB3MLthVA3yP+wb8sd1GSSV3hDE4EOxHY3hU
YXuwjQTEJX+DwEvzTZuOjf8MOLgip0RttmakN28Ze2LeKiwZb/CGrch0ygslJRCqbz6bRPE4vxqZ
9Db5IU3k2BPpcqzL1aaTsEECXM8kENR4O9uAnw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 67568)
8jiMwaX137iFwLpACaqq32Uwx0Kr+5XUBj0XhShpnjG27m98Fn2HIjRRl3I9BHFUFZYkc2ynvP53
lHv3gpmQPgf+xUGiHE9Co17ogIF2uS8TAv35NZvTaLN1JetmrB3ZYQZNzYh81y//rgP6M7jWRFQV
NXexS318HEz8Xulm4+zZBsv48S2yDN3wJG7GIl+uxVDjRpCJh4sm9oW6zLdO1H/hNdrSA9PIN9XK
/CE/3OQltBNx/emp26xH59CjZsaSN7w1mZnglq5XGFpoFtkdhX9Cn3XmXVBzylxXgJw7yCVtBw5t
q0Wf7HKd/Kd1cQUHWfxTsoUbmnPTKvmdd5hZL6MuQCPbCNEDZa3xvALKJJXZWts+pvvnm+oEu7PC
Aj0EbQMiYyY3Dy2VvrTvOuAVtPYeEMNc6zO0q7ydTuEakW5Vg8hLxixB2JDB6R0E7sgdC+29Ux7p
VYJH3/HggfGWhd0ndyVI0kKoA4NN2nnj1XKd/O0H5P+0uo+lNx3nZItZ4KTZVV8HeB4CM8fTYhvV
lKCHJGsYTfqE/+1QOzluoej4daLNON0em9AgLIcWOpr9pGeZoO/lNFajLBPczBIX2q5Z28/GUz6U
jQs1Q3tz2HWVEtXvt62L2zBFecx6L9W3HgPeIpLoGJ3LQnn2B8HFNB2g/lodIscJ6LDBUdqUPdG9
l+9KIc6d8CAW0pV3XjWy5bqQWgrHGotPgOQtxZovLOaTpF3DgJrqt6D9q+uS0LKgRfhBQ1D4Qd1A
Vy5rULklZQTGrJEmwnBUkO3soXuisduIPDlIyQzMyFXbhiRLYgCtc9P9v8TqHAk86PY8CwdKLomu
Mqkql3RrTvtyV30yHXcM8gT6s/Fp4ONso0IbVJwO9jxlEK/o8Y5elBhCYp2cSDXpmH83Y7acSgtZ
E/yFQyi2jCWB8xH/joTwse1H/1koM6ELHro7ZUKA3GVq+GsReU+Knz6KTNCr9iXY5LXz1j/QHZNx
G2n6/Ykx1t5H8FV86dxEwi37bPj0fmxpGW9VXpdIu0QNOKZCQcsYKy0fXM4doeM8dksh1S2966gf
XxkWrH9VskPwt/qS4GIMoGkR1GwLd8UIkMMu0uJWd/rFlGbzwFxbOGh/n8POleCLMi9LQR9icToQ
WxwzTHLHL/8sNoFyuN86CNnqFYbFtdfIt99rFbR3YmojAwBTb0CciTJfmNwBSo/5cQzyKrksf90k
1kaIlBQtZ52TF0BQJqvIkcC1rnhVYBkywUZB1AIUmUiohsqJYNqkFDpTS9Uo7ZBSFkEHn/Gk4Jnj
+K0i36moD5rE+fZUTAmXgKtxO5h7/7BonuOJMo0oSq16YZbMVaD+bNA9Yk5EUQ1Xlz+V7jv2aNUd
jJ1CIbP/H0PXUo3zNfY2bKQfCwSQJgh2RkaBbxITy4Lnr1WUdx7FSx6FknYPDScg/gwdCpn/mZ75
Dcel2lEKEX09FHP8p1kihY/YuPBpcWfMrOccKRfTfR+IiLY1z31zfOBnz5kT6hsJ6poHtRZEtRww
MAPGFB7ux+yvpzj42eWfwu+3pA071F+Z7XlYZuWaTQVc9IwMCOlvheIruS3KfQemDqlB+TnmPu0B
ZTa/M4mzha1v+KHxQp/DHKadosLjKJ5LkyPLtmtv6hlhRQK6RFU/YZC2auJSpkkHAypMMXH54Po+
mjbAyaOZhWvUe5ljMMLA84qd/ahnZTiSjAn5rlQBcRAmm/77kmIZYyXEGfIAdzBxcbFkibQlxeiA
SnjwkEzi6WqDlQVDuRVQh1ip6FvMfo9VRToZJLdEKRYkK/jMJc+I+n6ddQ/rYzW/m/eytcgE1prq
E/6RR6en6tk40f3EbeEPXasSm9nsYNmc6cRSqurmTobeWQPT7B+ihyGWIesZ0/LkRDb14Gv7iKPi
WFW9CbSGoa6u+8NMIxCM0JEWzja9YJ0tKh2s0Oa0wIFhWs601zHkFqWfCCiIopyhDF5JVx2aXAOJ
qfKYx5gJukog7IGV00tFlk5ttlGrDpoXqkDER7WGUVNWK89g6Wq5Q0htttI3MVH+DOAgk5wwRAKR
C6pAOqXbDR/+cgJnqf8SDwlglUubik81iXV/Fq73eKNGSjTpcGWlRgH7zeOQzv71STGd3S++Cnf2
dHpxoF/Vrygo04pMzSsHRFs/20F36lACLJVlzO3OoHjqwEohrup2hHwvaOn8BM6QuwQtNyegCRt1
5iFq+W7VU3g7F84S9YuuMdsDpDwTustG2vlU3dRmM+1zsHb2Z5J2ly6B0lzJWk7sRWBShY13QJMb
lGjeNuY8K+We3w1mamIAN1YeIge0jLuXepcFggc2CRkm4RxdkI+CqwYcb8jRY2YYRGX4XQbCiWQs
6L7O7IMTvWE85jqECQMxqHLXZLpJIzvrtMniOUim8CY7tZwYbXlaM4YVHCJnGlUn4xln8iZ1VW6F
s33RaWcwUEWUrBN7/8oUNUn1agragjOtqzHW3DQL41ThCnJYKCOvv7YqpsgT+IRUDEsPry5B/828
0EJ66M2PmW9MGm4fGW+yR3CGibESP4wI2LFwXKzES+2mj5ZYp6ueevFbaWRSalMmsnqz/z80wKql
vLvsuCg2dzbFH+XcXpvLzzXy+phwF9zgY8B2/PZhcU6Rstn0J6H3+7OX7OIPoTHv4lv+A+l5+uOg
ZkpzErgbHzHbC30oq2YdDQKxQqMqVzaAWQEF9ddADWZDTIT9998i+chE8K+IGUs1yPC69Xz39V2q
s7bIg1Sw7QGWMtnLS/y+EAYuFSiLCaN6u0CqT070kmfuSkk0sRcq2SKcZURK1/85ahuiHH1R7NSF
mVN3AWJfVvxkEOdVd1YAti6YywrS/0pmZJr6sPpDfdlzGlu0pX3tiT4OJo/S6PB/kzIHsiwVUXbk
HHJSCQSaZ/fwGXhOKZZRF0Ze4k62HBSonOh46j58DDgXCU+jcmArg2SdG7FZ61VqfPWdyzyX4nr1
9yX+3rKjz7r33MrzLYHIsOX8mh2RVP54tewiTxXkYgFGZlHK72bRDWz9lI+bFweogWgY1UChxS7h
S6SbbtdfYdWlIyxlyMO4XL1ResuILGnar6tQMfP1IflJFaAAkb2tEgrDvVT5Zg/8xP+IT1BDOOfv
tRXEHV5qx8yNxfEqvm4xT28GnWqUdpzC5w+HXEe9bgqd38xMCoVv5xFmi5xn4POtAMCY1foqGITQ
RPD7MessPw0xcX+fgJZboJBo/aflEfhq9s1mVfqZ2m/uZvmO5VIJdXxQMSuXtpt4pBxQRbtBY768
9FR6jvlJBXvb+HWXQQYZ9F/QNC80x8Wan9DbwZWke57o8OsOHHh6PL9r4wnx20Fc9ChoPb46X/su
CyCqFMkTdzgs4AUT41dtOPvyhnZ/YvEJ5rEY5p2k0Wz1yDZw8XflkjuBa2pDOn8ByNYANxfQgzVX
6dkg7965K+9QurP1saiDCLfHj9bMlTPk0PPC1+IFINrVb7XgWctZoN6DE2nF+mh7WfoekrlEJwmK
kSmt6zaFSZMntzKcZjcCxrtDQWC5FU8fcLSyVUMajWDBxOkRFwQYwOhPFfBjQGKmP81iOm3rQ3Ff
4oXOktKcM71D6/tuYOCnq9YacLh+xWNeHyVo94QxJcv1e6uWCjAZBi7LQC6U6UJ/B0L8dmmttkF/
DHAmwCNHfDa+iNLt8DeO9BKLDCgVb1m18erHUNc2LnGy53bsCP+kAUplbuz/qWsaTwGaxM0mInpt
qvADjLd1WaClfnUn3Ogdj/Hzod8kRMuv9IMm7i6O9RH2HQwI5Uke9++lPkLLzwtfpxZw6gNq5eWW
4ccnKa6S/oImvx7uXpK1H1Z9vClzZGZ/lfzYABFknWG8agc86eF43QF4HNhnfZXbL0HM9ariUEEc
ugvOgZQFtMK16FlXG0ppZzSl3TanudoPXqiar80n/bgL5zJZw8a5jpacnkonLUHQ6/0LNJUTyX2Y
rXQvWIQulX5BrHxIYn4zZdbKZZsfeAEuatwRaCU19NirJhworRzL7azcYaOWppA8ZAwpYrn4QzR/
8IdNe5xyd3Yq4m0JXohbY558mK1xlQUBayFXL28t7EG26Dn5uAzvbLqIoGwne0/lx6WlqKohuIWb
G8YyF+qKqmMR5wcICRj1ZYcqHks0w7qoK+7BxDmfVeCjZl9CnwO06t7D2PkK9r+Mx/gxyKXIMr/F
nZncHsReO46rGEWAeWu6Y7IVsCuLy2k+8K2cFHSUX7VMcbeqP1unnTnQKwzyM/OQHpm2/EioPkA5
GkbM1lqtJM/R3Yma0pbddnm/gsKMecFcAN70gCqouSTIvtOC8RN4hUUaQp7dCgqtX6iD22HCKpLI
mM51mTlmCregxiUIh2EZEDKSrBKi4aNcmGGMFY893zsKemLumxIMVcesqADJfwADJiwh+nUEDs2G
8cA8G7F6bJYjUOC8RWu/SuLUD+MWurb2+YPGPyn62lJanFl3qNkaRfTOoF9+7ydFdBAdBtchK4ZW
CgrGnOF9o1kQAOKiKf8st8bHAl63R3OEo5OCVa1f4G/3SCSTw11/DzmcHgQh7aMdkoDKwZ/y1/Xd
NklbCmF9se+YSymrZEEOurNjWTok6oUUCennkxxUS/rUsQzrNDIUIv2PiJB8smbu6CawpHkzi0/I
9KNXTCg4hxefQCRDUXEhfl4lNp87Vzb9GwXeCPREzbR8SdjvESUBKpWS7rjO06F/WedBpRLxBy+Z
l0h3pUvyJEiB6abeWYqbasnWs+LiDSx4lECWQP9uTv0eXO2L5LOYWwvE81Bj4YzE9L20BZcKjIMN
szuYUuY2iD0zg2IhNlXXNfdb8eAH3cTl3JI/z1VdEre2lDZh+AEnxrEe7yrayyJjiuWXSC9yth5J
l51nbD2U3lSIhL8swZ2zuawYfjW9Q2pBJxx41aoj3mPKb0SEk0NP3OMf7f0pHjvYospo0EwBMCaP
+v3mab+mfukRTmr0a/1V1TPMDoDPwRuvmrgDPc3vH1uXYts/LdVAE4/a1U8wLMdAgtGo6T7uxn3c
X+CSC6ZI6z7JLfCJ6lheCN6XLM7Yk6RB80y2iplIliwEoSC237QJeSvLcUV3tfgLBgYzM/8owcct
kOD7Y8+0/4bA3P5zW0SnPhsfFkArKji9N83HEbIAx4Ri/Ix/SoXo4UKtSAIPFKtOnck4JGp9JYWs
DRsvDD3WdAqaDQBkSGxiiZExLuPpF/byt5AbO9VY/RtXYJNhKNPSP1Jw3mghrBOEmvmnPM5XsxP8
+5/yxpjdlQbxdymXIjLzPH5ikjLCxsNHmKt3U0cqUPmAcUNh/nRZUJ66ZMT+1BbBZcjAREUvddoA
s7IRkXpqow8P3TGwO1gIxP475caiUUjnL0hdKbprdIOPpXJKzbq//JL+qEqQdmuFwW0lQSkffZTf
SEc/8n59wywf7evG/jG9vziTZOrFHHKPh0kbpCuzYr2yjBl44VyWeAy13KPMEDz5BDsAd3xh7HEN
tdz9aT/gs3iMl9aEkst3RnFH+LOATtphylyWDRsEFeodQh0vinHj8flZwrpooQ/6SfmKfluczv8u
QF4EFE2GHDkTQ97NXmbOnnMokoYSwKfRFDMuz94vfJTRQUPyW8rqVhOvdcjOFEdF1sOp6tCaGToW
yolWUhUr0DAKuCpJijwY359DFUTexOYgeT4gf4u/3+P9F/WlkNPWep4g4B5UlK7a4xkq5C6a1QoR
FfpJE4bhAOU21CtRbZSQoPMkDq9q4jX/i4pAGS1HlYCkOOk04Wf7kQrcMEgOW22+G8dmqh3XM111
DxrEi18Cu5sANzFByH8Ir2nmGILFcbgDSLzjp37Io6b7cYnrpFt0vSx8EFQ+6PAOFV2W6dpVADFL
4KHI4eZn2QWe1na1JIAES3vp0T36FWtHHs+vOdZwD0vl1a5U35jjxRjCIrswvM3m2Gv8J8scjY2N
5d+xu6YAF7NY798KAGKQuUZTlTCkktT1wmuXEkNy2C7uvHAwnD1VUnDkuiVBmMSVAMjtBoAwkN4N
xo3SW+j/eG43oN7ahzW8+4RE34V/ZMrfMkX5sB/aigZjaHLELf/9rT11lMPs3yb5oJYojya1r/lJ
rJFN4uv4Jz3x4eozpz8GCiT2Jx5mwEMZa15o3Amen05FvL55NClppsUJkXYDkXmgVXWDN5V9AXlA
6003zY3Ben1+tsB8rr7kyayIj3zH9mnuzLIqimKopLZ7eVBhe6F1a+xzQQaKNe8jGPxUIog8KsTU
joAMjDZQJW9ZWO6zts9Y78VJPr+/TLO28zEgJdnr84OrJSnpPCp64Inh2JQVdpOg8sd54Ph1Vpqf
1LfbBjSJwRIUhQc63r8O5HTXFENCRgPx2Luc2V0xLNNGszGSt3LbISjx2GfCeZinj+jXQeDink0q
Gzf/Pp3iicmo8vsCYsYsfNm2+YKn/jFmoKe2CsTW3oqlNY8hUw49Pr4MnMpof+znLQJpEpS5bFUd
0vF/ElXNv8g/s6hUgpkb7dyKrIiwX43zt5FuKQVq88ZfSR1C6jAZnk5foFEk1laX0ie1RwCnOyDr
QyulxDnjzFAH9g5UiXLWCMU1Za6rwhh2JGgfuvhWCmL5i4X9CvmAmkz/897clKvOUttJM1u5y5oP
T1noW66lFoerDGrTUpC4tVs0uMVN9N5GRTufq0PtzZ09/8o00nrPt7qXPhZZi9igFCKrz5o6G8is
6RomK+jTb3YIk/RA+noyNlHLASYg+GdXmGvpeld/w7lRpUom46dl9t/VHv2wYUjvaLSUvWA0n1AF
qDWACPb7WQuwlO44JKrl3jTr1blrfb13cdNXU9SozAulFhcPIHD7/LF12P0XMZQOYFAcJGBliRDg
p+ZtVyQnwO2qMxTQ+P6VktPMHJUV9fQrvEbzXm7C/BbBu7wx09fL6/yPQmyecid+cdWGTlMHaYWO
a1haKrrvJJ72K06s/tXxLRLbV9NLxKSbo1VcaTSsJefWE8U/cikan+2UsTZeCErHo0aS/h9bEgz3
W6V8nk7hapvhsAUD0vGRLswAVyT3zGVH37A1tcm0On3l2ADoj84UXxIP36Ise5vTjda7Rz8t+8+X
qdEb1nXMVScbyUgSHUY5XRP0+eBTp1NUP5QUwQzZGBY9yNYzZGdwFhoUSNJ6l1KlyuUwwbi6C0A4
LaR+sRWhgo//Lwq8ae3y9NO7ivY3AQZFKnFhBahEBBNKJrt7c09Is0jLuyIypJsLvqi4g9++Hdde
ieEiJ5YV4ZJEh+p0GEoJCGA/qdLjK33L85d6osnY8KMBDvYX9MLaVYYJHVUJrdOYhdpWgQg29C3S
zko8vjCpruZ1u2bVee0jEN9k70CyvSoFUvh0dPA98smBFThz678aoBNqDOac+Uayciof8RdH70N4
QjBaVoZTNBXsst3i+BODWYlBauj4x6fhKDMA5bPZwOIhs2c85fckQNrNJ4zEl9zeqWjjWGJKY7eb
6kG2Lc/zV8n1Bycol4cKdIox80r+skSWBIESnjhNezgg7etgT9eXNQ9TfgSbJVe4XtY2XpLas510
DgJC0QWBP+dFy8wdDcWw3toQy+nMNWn6dH0S5llJVx0rFrBM6fi57rkba+Jv4sq/ze5Sm/yY5ze1
7WKvH69QTDVKgAyn442kwKHKjKMJzUg56WktjndvSaDWxklyoAOR1efddNqLDHHJ3wXPagOO2YMx
l0+HZtL32nKTEWhqwIj+/SK7WrLD2Y4tSgrWuXY5IEg/uql3fFlDUkoGsx0tQhj4BYKAcZfdHk3P
3aGpCjybWzPuCiD/VxPBF8S3Cm33TeH/ZWUPJxEuAkGF96EanIgYJhYJiz43eCqJ+9DZJRbtbave
3RbxpHYK+c0H2weGL1efsJuKYCN9zETTGHhT2SgjrrevtXr7uiWTOvI1TmqPnD9dGZvH4PtoHwv7
A5jeknZnsWYC0Vd02CCFo0La3eJ//cdvFV2V5ea+3Khpk3ur7JEQEYimi4N0HcL4kG+hMZKPOtjR
2maVimAgO4JRoSWuxXgxKgc0QQvDV9mXjstM2gtB7BijqWn9RiPds6dfr5djkfSRuBozMwyz4zgS
Q4EZ6Iel6YZHqHv56qHL80w6NQXuOZ6gkAO8i4H/1ZauXBvA4TJsi82b6Cxj9TlXXLiw/J11TrRB
MwEy5fpxlfjO+RNNWzE190OngCJZ0SZFFze1aV4gNhDdRgH9dU0NEjIuU2mXOTk+W3HxstOPhC6G
0NG291uIWcFJL7c0LyCHidObTPgG0//MuTS7ZvoTm0mp1TYllVYAaGaLlmmG2I4/JxyT7Jq63Dpd
PximMg5n+54YDhCDYBa9dGigMLWSrRZpstfEDgH1/cp4DhxdrExiUxzzvxg5M2H7GJfRPyUhthm3
E1884x6pIyYcYtaaUidsq8TNWK7vSeY4pmrUTDm5KTQ68RFUdRSqNnqLQVO2+S7J1qv0SsoqtekZ
GZhH98vJCooohJ3381awBKEKPJ/ci79MjBQebHUZOdFLw1MwrSF1O2R9vpW9CEMK/IMiur65aa04
IZ4/cDv8RGFEct7S8wqu6qHnvZNqGEZlXRwVv2reXuzpJsYExUY3r25B/VMdEeowDv+dCBCbdn0I
ZNhHTn+MaqWTfjHc9/Pyr21tImpMVhK10yxV3qY9fEGw0bhT7KsRSKHwp4zFUYRXlJAQqsjf9Ksp
VqZuOnHO20ObNwfVWszxBADBAatrzHEjIHgFlaBwr5zw1MEciVeb2dZIPXBt1XWLv/irhQ6Xx3vl
26Mwqtp9Pq9uxHDVatJJ5WLuD9NCwMrdhF8VVJq+KGpi70m4j8KBsfN46FtFmLR8hYvL8v/d85W+
Phglj80DjCqqPVDAW1EyprSTH/NlAPNdwKY7Fvrh7RQhLzu78sZhY8un+WIRa1IozMtzndVCR5IB
FW1b7EaxhZOwCfgMPv8VGRd0BoskEYk4EAukcq2uJJ02xjUqfaVYMaHSbA81FStjB6p1dJl6MEeA
JzfcNsU6BMGywMqng64YZgBmaXPgMJLqGym4nsc8MWnFWxkKb5H95Du4b6dus74Rg/qg1evGriLt
9cEL3TcHgKVbr9M3kL5Mhs/KyDvE4FBoUAeErGXIzT6dQhUxfN0eNCMI15/FIfa3BSmsKq7hjCU4
JB0JxLauzB9Q+FjePdIm7Yf0llK8n0CNAOEfwA/UyFrcapw2eyt3tGG5g4iqvh3h6gqYkBdZHvM8
VV8IPpVq+MWS5iFsGCLJv0soGUodqIFMITkgsiMGZmCeoX1TL8Osb48XFE+ctzdNOye0+xyuMJGE
lQuDdnOjV6WVqsorqLM57TdqnhKdiaZA+fHL+92LD2bzcln9o7cCI/QJi694G3Ehd0BDE3t/Wyi+
HLUHIwU9eGsk9T8IZo1x+Xen4nz81uYyhSmBaulRzlTHAdGb6UwhV/FJSy7Pa5+nSEUdDXXgRbvC
OUiE2ISP3ZvERY/++3exH0wR3MoI3O9QF4/LPDGIe8Ss4rwtC3V0K2Sm47pH4GcRw1n2fGjmMRIZ
IObMjZMFTFHMN3KPGeRvsuxWPWX4X4Kb/6feCxEckx7hiPN2Wnlnwi8+nJ0gMX7ncWLwxTXa4z+R
ZDdUyFxmAfEfOo7cXK12wqVKfESlKMKJo3145RizjCWY/qZho5vnEJyY3qPnrarGOKNtuLlXD10C
90VpAOWmUXIGQnbgfUuk0dVAb81dkNpWsWGKoIKH6wUSMaq1DJe/Z+yMmts49HGCeKjza5iUO6RK
8a6LvNF1+ABtM9FzwdUPoiuuVx5hSB/QONm7IggshemnRmAQPKCOgfk6XLWhO2uKo9o99inW5TVO
XJjA8MI1ZaJlefSoYGXWm0IJX6PkuIc6gpQlEua32saoCHztgEdZqR77B5/zDgVxYHKcA3V9Sz0U
IOEk72c6Y1dyrQ5V8crGRYEv+8aBaUzscUTA6r72n8NWVe0Tj4Fw3TXgmW71weMr8+LZg2A2NvSg
/kQOTfXoDUy3XO4d+0DxIcJDlYkuh7e7Gp6f41Ig1Gz1qgYmQvMOCwJHp1kioorbVXD/j+OtCXFc
/51iK8G93a+9UicorYygjhEMa3sMBkHedPeYEOMP9biQtaFCEixDosAJzF9sAjNiOUOJ6+7M/SP5
GAxMZkXLM3oh2sG7HWiC8FB7ZmgBtNQEUPWAtIuOTkemc2/dJzDcKmmsGEs277wsKt3d5bsmpbNB
SZDSXyuV4bEGlhUNKkToe93pb9wNBZJjHgf1lVfEWm8lSYoPFI0VKNUiu8kL05tWqVWtyjDT5OSb
3uS7nqp0IMHwfE4eK574kbWHq/UlQBWxysZKz5WH4viC1GIAecLC/oBvD9381xKtM8g2q4/eHM9Y
BB+0jvqZA7MBQr/3DJ3gZCau1InyOQgbAja/fdX7XUF965rTTkVVwsiQLnpSqmoSM8WGLsn5LnPC
ADTk/pWHOgLOeHAZ/spThxTh+1ra8Z68aHcrR5XdUTh2aB14o32ENhvBYAHHxLyvd1uJs7rP7IH7
jGjkAeLU8ns5UMlGAyXRGXZMxuLwBPfcvCftoCHDp9ATYq92Mg0YEN4UfLiarzezzgtvgCHpiB9Q
7n0jWhZ92oKRcLHsaOyeuvG9fN9fZqMKOAKiFgNv5Sa0ZsWvz3fQpQ9mbRcrEwHsBtUF08FNdPiS
uauWqwBz3VcIJTJ2zYN0nCPO2aqut7lI+4a3l0Pfe+vvFMHJn3hOGFHx1VVA+fAXEDqBnBwThl6n
2UVh0dIuazHTVn/ip8URwQ1SLxrURJueCoM1aINccXsZ/pjur7EmZ2wQQk3QWEMAVmXuYKwI5Ciy
Vq99qzfvvY5fLs+/5GUhbzbk7ZR2M39s2AH10mEqmA4F+TYNEhsYcdajHhj4LZilc314uN96lvTj
cn9XUy5NUHcJJBSP6JUinnSUYcxhDgeGSXEJBdouRIxgoPe9MK/9ZN5L1mGZTFuLIEwCaAQrnxVS
UTS8cf3g3MBVKJ3qAz6L+bSvgR3Qrvi24tAuiOYrGGc3kyIQdM36HqXEZ0phS0j6AEs6GICepUqR
xkoRvTSS2GFYs8jda8kN7CqErg05nft/WPzrDUPBOpE+7ngnZwvevuMXjrPpaVX5gcq+DPIaux5E
ImVOkcHzZzKeI70241Bplt5zuDZimRdh3premO2LJgwF2F5+FSpJT5TvdNJNKs7tlr0xqn1jc2Ua
Ub/cysIhlBmeuknHC7Dj+Mmn/jfQDhLyivvWTvYFm4wgJeKGc9N/J6U9DssAmIWkze0mJ0KaQZda
AXIPP5CXvR0iAa7ijxzCLAAvNX0ybEMtxhDX6WurrRn4/7Q3Kob6c6qWPnap104VjD26ujm5DoAY
bVB5rnUDpEZkKoVDJhBwrcR6uCX/lLjr1h2aqWZK8WFYG7E1Y5yUPkVRmkSGUPw58pkaCpiFkZgr
fMx3b4Nzo0GzkSD6lVh2EB5mCJdUtf6tXrEALewZFZfkLKNAzTapKwnejL2ZBmtYfXvCzNKb3Rpm
kWbZ500tQEO8hAyvfnAlbr7DK6R0pOGTD56TEuuTuHifjcIrSh4zGnpos9sn+BEj8ls4XWha6Xsw
r041CLMVJ++hB/nP1+P0bVlpRpnEmJG7veQOh/aAcawLfCnUDiN9M7bkcPWzwAmXDezYlFGizEPS
dQeK+UtEfpdJ3cDb8xQnDc9KsHAfzo1wFWfP0h2Q1+Yono/WZd5rtuKJeM9N3rSURqWSWsu4NvBW
n+D0f+t0dJzNVUiNP/gEzVcV4xh9XcDJLeljd+OQAO4lM7EHsjPfyoFLC7xXK0on28Rpdc5ycAVD
FO7qtuqfXzeWLlhsW/lCJovKOqsPD+q5cNt43xe3Y0SAke0AXk9f8FtpxhfWN/uauW+pwrSV+sGm
aJJjRljrTXS193+RG9fa1+N1g2Wz8Mf4IsPe4xpzXOmsB14GvA2mymUgsTu+d8dDzIT0MSVq3PYV
3wwK3CZn8S6LMN5cio5ZnTgd7PHRbn9gP4ikjPc3Qcvixq3amit7QQU3eBiFILjuWSj3gSzfxGuD
AiI7gK2IC4/ioZ2mYZJ6W8xJzw0xGmSkekWruDp5tOlR6jJIX4KiLKnxIuFuj6MmSGiub+LHuuAm
HsIeHD471E+PiPZo9dljoJWth/MumVnx5BKPjPHDLrSH4+bPktqhf8DmLVKF74rj5b0aOENtW4sr
ukC4jeIuIRFcwAnePHQyC6tmEphG0c1MYxjkEMYdR/BJjxNpnGm9P/58cbJdCEqaFY20S6OFB628
QM1s8Pl93JqJGNw/CuG9qpPNsbp+F5K9SWZ5k9Jw6ICtE6kOOEFq/P1L/IdePgU689KfMGoTooe+
GwZrKS/07zaXZYNSas9hproff0rJxF9XZuXMI3rEt7b4Qp4gdLxH5VaGAEDTxA0PXCjVm+1FQkRg
mWTKaLDpbgous27hgUAXaGuDZt2s3zr1Pt3IOv3zdcBSe7Nlx4MRJb0vCn1Y9UKDlHFW2rE0w5lD
JPfeJ2S0VtFElBFVL6s9ResYzSubqefWzF9x8E4vaLExO18SHO+PuLGQcHWUPCo2dtbpkWnz8y88
+Hfpcj856ngCQzN+5FDAHj/4dxM+Qo478dPoMprulhWvPITWCe/89OA2oJgU7NaeHgOKp3QRMGN9
5locffJSJhMnlr6fWHo8hnIAclGPPK4Fhs5tXmGypkMq5fvML5lrYj+QlkZIBeJQyWk45t1cJzZ1
8F++Eau5dzy2YjsENRIspz5yZvnYQx66Ei/yV4lH6CEK+mvAdCCKOfEtBs6S/MSlzK0EPak023MN
Q2dCcLk7tyJMurleaNuC8OeJl/ack2Du+SaY47ArfZnvoTnoztJf2oBzwDXyXDsK2tn+fMR8Q+Su
2bGpqGuHCResONIuyeDxz9Xe74+1wVPpnzJyL6ln2DRVRMURsQXRlTY6JKA4d6O6Gn6CqlMb8mas
lL2v6IDdu0nGUX46HeiWVIwirVgozOu3ZTQ90UQB6Yk/7bHP8mZZpccOLwG5qO2S7jUnH2RNu6VN
DMhnMkV3TZMEXnXIE9o/2OYs9JzrTQivI61/itPfqHnEOcKZYb5H1RbphPvZ+bGkBExJtJdxS4vO
W5EI3ij2Yf1jeOQh6ob21jBhMaL7vMWOBFKytFtlNV/PCQrOHU4xPjWParl1NBE/49yoLFud3+cG
Xa+jVOzcdqfkISf8eZ72NGDOUxU62GMa7mcSkptZclahkVEFiLy3snxgjNGyl/qkVXtKoucErf7O
5DVJ4EYixWWGHWwEx0/SLqS+H0Be2Lsqum/hhX5oAdUcZQFXJnzw+H9hPQzDHXuq7WzJnQ2mOaj6
wjKRhIZZ5s86MqwE2TNzCJi/PfCHdt1Ayt//dTWy8H2EXXyRyM0lCaKEKyYfsI155bv2ET1VjcOh
5kzwFbiAHFwKibQRFpSQAJ8fECI9iL3E/uJFCc91P3L2NdAupFTKaWMdrVNmJHwANzdMYmUndRkc
Kc/T7jeaSG+HK4TbftMriVh7Z6WaBQjc8RWVpCKaWdqAZ3AAWCsMFIu1o+N7UNN+dEZ+oaN+60OT
SAh8oDkLHdlC7JZoycMKn+JO13VYeId2CldIC9CLU7g26z4lAwm5bEEsrX5Vghvkyc2/ke8kGjVd
6vXg4VXF39AzDJ6FJVJKVfjX2PSLeHIkqLYU6OT4wY9enIwBIyVO8MXHTNEPbvJqOgcOdqFXiqdO
WxR0+g+2xdioEOHvma8kGI6LBsbiXLHH8SXDTvHtW97v6ce2feT7PNOkPrkEN0rH0T2aPRJYWj2B
lCT9uhuVERooPy9ZPMl3GZhUMHa1M4nZLgbCe/8Ko3+R8gvSs9IFzjEE1J3w94zGMip00kuyltgD
ImlNH5phqHc7/tTPjw2M2AZVxh2lXNZ41jqK7FrnPuEDvVM5HOmmh8ZUsHZ+D8XPX8cFiSsa/YGq
eBfHZGKTpPkAl78BtyEp6L6ww/Xdf8BovPcXW4PZqnh0A/JKi6Oo1UFFEqB0AW65VGXk0zqHhPXv
UIzkHhvpOUiD+PdeTrH1t0iQelWbIQAyn53evbnSGOpYfuAqOT7PTOueCewdL7sP7kHzWabpZCT1
UqX2ijnsU9lIh2FUn5rFoYfR9Sqd3Rncu2pfPT7Z0Aokk804u8mCQ1pEdKJ45UqX+S2v4AY/b4im
NAacCs087xUZ39ABEswOlYThpd3Xtopu51IVpGGVgF5lH8aAsSvSb0SlZmiDISzqyotXXrtjvc0r
5fg9hb3bzpadcDtNxo40sMAnqgM2E8xZCEz9tQwkYAnUg/7wqZ+D/TymI7HYeIhO2oW+waRdbHLE
qu2ZIu1pOqHRyvmkdvjunzxYkMaMG62CXQrrn7RkAmqea/onMq950h6nywnubSsn6aNQ/FxsCian
jdL/pSyDRceaaQ7ph0ggCqAqXJz4KF5wsz5ny9FIpjNS8d84qcBvoyZ2/yt3j80oljOBG0AR1e77
QoXsIxzUjwhK4YY/eIp4b+3o2Ma1024NmeVyyfxyLvDh1/o1yzm8dlfPkjuldnoJS0N9K1cN4wi/
8ql+qze5C7FglLO5aSmX1L6I6pJSPUCyEP+8enoAhIltvGqc5L8FQAB5DKGavXBaDoALiVboa2kT
oxSuJTDJPo9I86n1e6J2wDrWT5PHIg4TC4FrWZGsl6rYm/TBEU3gLmdCpJBwLdFN2K6QinAitp2P
2ICFjeHKj37XFGIbiyHz6FVTza0KTJxVs2hp8ZQ/mZvxIuge7hQ0/PwACzN1qOKxM4ckXIU/1Shm
IdhYjoQpv+CHMwyljkJZXAvk4rwzIqh+VqodBAKedrj1BbWNdkFv0U5HtYvssgNby7oJP6QCAqbV
1++7X4nRC3t2CWmLtoXd/inoC0qdIotsVHajsgViRbJX1szxmbkD5gg1IPQPbcNDeWYAppfc2/Sm
PM4J4OIeLUmgE4aCFSPfpybXhggb0DF4xGdm97dGFCMpdHT9S22wqK0OytXSuqZqfmhrQ7eOydAV
lOxFv6EYGai7X00rjbVk9Gt7vRo4D8UgQs/L1Ch/Ljsgl7r966yVCMyD21BBkYobPng1Zx4LwSAG
uNLGtAFS6FRImqSqpXRsY2TD4QcdX2zMSJLtwDqOaOHAEdxPmAAgD9MmVVxfVsBiEa6FwmuYRG9U
31fHIf9mGYrY0AYtGs+E1FVS9GPCy54AE953x2OdPajMqQyyYLXaXDW0nyPkMZtUPJUQwR2qBz5/
VyvG/1dj9RF85obopzk3QFwf/q/j/N7bymtsfwnBqFKoKkfZQqtpg5eqr2BKGlZna8dHNIG6FMZv
8J9OgylJ73hJy0oBeBCbRXJpAAnB617VlzZQ37eZ+DFqyqQ5FNj3H6pOUaZP94IAauB+u86KiXNh
Rvnlbn5HFyMbbA3rCcsJ+F61Ewy8EheiQ4v85WDVpO90tGMsTgNrxlIvR9ZU8nv9199wrm4BB9Oh
P4VVpj+5tAMZrDNL6WwdRxhwWPv5JVFvoZ1RvC1pM1cjPPBnu4KiAajDZQ/cvzWXR4kRR1VuvzgG
iUE/xhXk3EPUIcVXz8FWUB9EgHsFo4xWGvSgImQtjd5OMFDjDQFEfiNDgfWJIr6ZdAvoMWhT697y
DYiKkaojtGYNC+5aFOvIiPJdRWrREkon+l8ayjB09FixtVCHPvHFuocwPTqUq2YuOZolxoexO37c
v9fBvMZQy/fRM+mFzDfWbsACnMsWPUAKGHkU3Yf+BbmNiNQoT1tgA98nKs+SnfuN+aQcN4gm1vIm
17OmxK/2Y+kLyCIGw9pgIi/3Sq9O3r59Vq7hv//w53kq1PfK2NH2GOK4kG5pSzwJe5DBHCikzsyF
Mdq1z/uIRBNRNl+IHFwQjsw4/T/5Qi38bcE0opGFOvWdxCYMipagRsUXrFZjhVRw5x9xnvFgSEEY
/zqH9wGRjsQBxTb4lZ5XxTfiDbhwAyRgXdenOtzVj/ZX0AU4jrC+/m9t8DbVe9ECo7VZXTU2nzm7
wWCCvZF2qjVaOEkP2JRruAgeCT8fw+rLS0Kh96IBFNetsKIt4DAeNDnRtIwF2+YpV9WJhqGOMVrE
sMxhKtuQq5xFfOQHHsVIsbmNlIcEueoc3/2xaFv493CsOZkeiPNMeHCLHDoi8SE4BwraVjWpoaWV
QeVB60ZeZMT3/Yz8ArZ4GwYJOjCoWmY+/q3A8t5W1ju4cu/D101BVgUUKkgAHZ1O8YivtJbMrWT8
Vpp+dbG56bGPvwzes9eMz/0/79TiO5pqQf0NAxQGof75EGEc/GVMkWQX2a0b/932usfgp9KksagA
qKi5oUv1uav8MRG6yLBaaIcDdh5PmiZOSposFnnSex7Cunr3H03tUKRrTM+xOZ9gU4RzpE3hmL8H
1HKcARrQ+sd4AvG9yvuGUZB2ZHQBzE+weNqJ8UAu7jBx2P2fy+1M9WsIcy4lsO4BVRas0uGkAAUX
yvt+nscC1g39FZZN88tbnWik7K2s/ecL4P8uHquXYxNZoLRtdBLNdUayTY573JBAWUIE1ibS1nb1
aOoC/hkXJwQBVIM188bRk/9URM8tILQZvor348ynKlQyBqdFYLh5a/ohgubEqW2n+wMxK7gQNt7r
6vbcy5LbeuRzsdvr+fc3spz0JrpYqi3x5/qt3FCmEQShR95oujunh2j47gyFoP1L/fgG3f/ybf0h
Hbczr0jEYcN0P9Xq2878DS8GgTcAlmrhi+IGvjJbOWlAutMuh79ssXD1FjWjfbCkdYKppk36lqX0
GyxKBNduDj4Kf8C+wwenN8RUDYuK7XzPcVW8nmPf82AuUGH2FrUmIjZ4T6S+9nyX/tXSG6um4Qgj
T8xgYoQZq4qExYv6Nbv0UU0Tb8vEUYYXOGAOacGplozDxYv7GwBJ2d84N2o3CZNUSE4NpuUIYEx7
aeA9N3/MIGSi8x7HxjKSMqXpE95HqqP6jhsIc42/Rs6H210u7brmZW6aPeyCxdcya39nf9uj9QM/
BW08HZ1oz8K0Z0LWh79+shT2wFCzT07xGMZtJkCbG8cGc49VciLNBK0asHrF1M4LPBG0i3Ylh+B3
cPM9NukEWMMm0qH30AjiMNNdA+V4gtEyAUwfq3IZFaqJEo1/FliVwrmzAZB3cIMtLVgLOUs+Q1An
3lMTGQUUqmuZmS8KmVL5ZDGhHgnd2WmGgEoOXCQWl3PWECBsaqni6HNBwt19rChzVPlOQbWpg1XO
NMdBkKVIq4GR3t6IVcpSPIsUh4zm0glcIQDiDpgZLhzDgXxko6i7Gk0sn7uTOo8sVI5kuPos2Buj
0PUNufJqNujJUBkGEJZDfDEgRRAcfYR1FP8MOHVgW9YOJHkUYnPEq+KrEPK5MaYssI0cR0onsvbm
yXBl9dRt13FlHTRBcJ9NL1sa/BF79XMKPKQ2rFvzLA4f24JNqbhyRTOEbLCejJrrLvS1/p1ks0Hg
TlvYiyYBW/Cj8pJcA0ogogySkofm6G7gpkeUCgMX2DODvYDcJi8/qMItXV1//ihZJ23fePrWTpQP
Lv2rMUT6IqecnlEattz9IPVC97mL77pA9nM79WH0oTaooohVvMDjaNmCa/TQyLLXXpLdgZZNB+j0
4IalZ648Sht3XTYcK+OrTNErqHKq0BpeEfMTdyhmZA//fuMFFd+BP7nzKEUVda+rBZRo8Ir5OfCR
r/jllLu0SEdqgoFD97JRBen+da2UhGPaRsvntvHiK31L4jHXcfqCWqcwKuKc9DxqxGUSgksbS4Fo
aNds5GnrKu2+4ILAfS/AzjtvD/Wojhj0/QmBriEQp3nxgtPIHElmlkZQHqVA7RMJ+QkpyBdcqybs
Z7Fv+TrHiey4++8DdKW8v9nVmKQT/IIACcod14JYqazTU0hNVgy1y7k44SHkGjL1uDgnh305ct8K
KCANo+hQZ7N19tRyDgTg/pI4VrjWFjNXJe15suc6NVJDtducA+HzQVfNkdf5V7Uyv8Ny+wxFMC+U
/6mP/yrlDF5GIwDkxEO+iJXZguiRy+iJiMwbrFWXq8XahA1mtekAC+DySEVE+MvoHVTyhh9ZlGsE
XoaoES88gdPACszFuqnAAIvKiRDWisj2Yc7ai47cJg/c9lq/lb5QnqaDwKdwfBDFbjx3k+FMD0sA
rjokKpU2T1U1TIJyi+X1tIpZYd951PLZDEeLFhXwf8KHI854HWbbEgRkEk/Hxq2q2GhFC04h80s5
e4dzwfcO+LM7oDYGyWMdeanJR7odLEq3M2eCsJNQ34Ug0vXO4F3q+Jkhw8RMy5HiG7x20a1RudRV
VnXpd8z20+lUdCIJQYnDbOSel3p04yqcW+gcq/WyjGF8XCURzDW8eausPu+Mjy3TmjQMAO4f8PtY
vUf/TR5GdBj0G9KUQvrWEh0y2bK7Yr4js5Cqwnr/u/oN4Yk+WJ68in+XsyzVmOtxuDBRRzHqUagC
aIPSW8Uu1fO03aqnq2dG8RVdqd2toSIntHkolGAV1SVHVtUHMbAhnMNS8I5SL+VesxTywWMTUEj3
1K/dSmNQAslMGYNrleoLUCgT8ALWSUfLXaH7o0kPXUBK670H2HSqp/co1g89peMopV0JVyIUszkI
azLp4yRspySsorqmYXZU3QMdF54MtJFdcN0ivNeS8wXE3IgjjFSpXfk3WM0goYPi5+2Oh8ytLsN8
AYlOg7eWF5QJZagmKS7prAe6BgJ4pSsJvBfbYiNQUnFuFwWLfIDSrJRA8+Hz6suiIpmQrXKqIVNc
A8f4uO65/AidZxR9Bjk3qMRl+CMiHKXZbBuOyc2mSy2IEd2fjAO6UMFOijlfXJriWichCO14fkHu
KPn+b4xYOaWrUjAlvq+sdRKEMTgL3DofSRPyittnSjeVy04wygkKZ22FRPofFhMLluB+hLXWqrdI
nk+TSX1coxFNHoKqlUW7d52m2EYd7WgExTbPjR29wRSC0BAgzqyWihXY/G+nNDF0kH29hzbLQcxp
NKtFG4lO2bCQoL2iWFgApjQohEyQxfUGQfyqN1iVfmz3ePmqox4UajP8xgs1d1YIDcm8HtMnIdPy
hA8RkVtMNRiTNq8wX7KVZ+bltIgosOAx7mfklq4TCzumWwGheXt4+8ZcSEat75wjlXIylosroOZv
hEJve8PPGNMAlkRJQF+dyKXJ+Vrr3Krt0R5UXyI9dsKar0MPQTvQ6OzXcyYkHvx8azeE0dxKq1n/
I2iFrFZew/6lGUROihXr8ssQgtgms5CEjjk7RI0punPk2hgSpcZKuvwUR3Ph6Z3vIcpGUdMvgabH
J/gFd1WLZIAYuEnrba8kY6fkFtea93lvFVHyknZDX9FCQPD99iMqsfnlTDNWtr8gJlPOUD8vQ30D
/81x+1KO9jAGH0d7n5W4p77ITDN4dqAWVO7PkdUFaMfJV8QBspF1z/KeMxCV645e4fFal7aYS70n
GAFB1UJWjNYffLIpmlQ1lgf2kEXSynOlda5rde/2YWmqYzGWPd/pjEVvFvdVz4ieFqei3mlz5kfQ
UuXHtAerO8QbVP1ysaSzdb1dDJCTG1DAQu8cfdE/2rMaauqRXPWG9RSmHuk01tDv7Lf3ArjsN9gx
XrgXEjpp07QRQlZ4OAOMD4TDCglYr3v0py4Yej77isRRGUonTq8oXIJp15Yjreq2ZnbhL8TstRe5
GgPMHsggoLxwhpzKGSVAxjguXJUP19AKC5M4eo9BybbGGwp4A0klD6xrPwLYOzRiuEH+IQPcS9W5
fl7cBHJppte23riMZ/Fv3I3BsTkWiDMnC8wuIJ5keeuq1W2pW49MNaVlpEkHmAMS6IBtv/bU0urG
0nc6XK17hX6A5jfO+8uf988/oyiBk2ej1f2nVenx/gIFU02ng2881a/bJzAOS78uQztP2s8pTKWt
QeWrt00Q/rH6VB7CvLTpeD1iAGSfJnCc1MYW8mxY5ylBGHavefAGXA8SD6kLEnL/rZ4zjA3CDz+I
OwU2LKTzCO8LcsZ+Tvyd5uRf8qix486IlmZOwHl4vc2hva0leKEI3/aGWZEYbOA5mTm76wu4ovkX
S5kPTTqewyve5lxivLf3Zd9APxeR7j7Hjx5uFZbCttfEh9Tv52IVmsil5ExtKcuI4g4XOXthqbS6
D4zfH8HS517siQf5GVS5Um5KNavVF7MedIcBEC9C8LhUk39UyZi8V7go46sTSDwy8yBpJkubCUQW
j9eeaz2uZd3qCY9i3CjYWxDIoXglySZZve7mTdLGvh3LSOR7Hlz3zgrSNN/C/Q0Rm4suzOCl1Cy2
EBrL0ti7oWaGoL+8z1kNZ5DQo57MHAndC/kgz6MGrpxjqpMFn4uKt44eM64XvQw+AFdqur6Vi1ky
5YdlTHRGg2cUVYx0bWMHU3mjZuMmFsqpy/L7m/Bk9RgOp2wE63sumRcDZ0QLWXoKtab0yBZRZuVx
b7vgtJM+fdVnPgIogE3I/mCY7kKu/mCb/TnDzUflbaFTbWGYluN1p1uzG9EqPhuAgejq461baPRf
HTBIV79od53VPuSQdY78Dpqyhj5WXMmmWWpoIlEsPFF1ALITXqiGnGY73jfMBLl44Zj1Vvk8GVVD
JplZBPJOkTw7v638QcVg1I/1dsS9MdMM21sbAIPiRg7tCDEjsWPsCYXZskXVX94kuZVsGjnmUgCu
67zRereeXJ2JCGTsjzhyj9sPzmTk71e5eoXqwiFIQK6trhPxeJv5e705ITC4DOpLHcTkAZ2ibfdY
PzltfWUoW/NcUKKV/an7FMjNPXu17+vjXm/NTQ7AvhTiK39y7Lvhb0fDrRLmR+HAYA+EjAFO1rY3
CpQtANaZz1DoJEMEP6XEvm7hiyZ6ctdNaM8mCatRBESkIbDW2WGmNwQ84GdT4OtjIyl+l7T7cOI6
849bnI/1G4JThmyki/hAp80+DmVPxKkb3sHSYXr2Csy9CsiWGakMk64gIXqWdiaTivHG2Huk1goW
TGkE0mE9Dn8LIEvFzBc+fr6UJR6zO55u+w0zE7zFyxfctO5bQs/BV4fvci4YaT27ebjK4jPqCUz1
swDeTFmA9a1hawmsWWwvslE1HqOO44mRWeZRH/wFYcEha9cuURrWnkkG0ZBsW/wNNvapglINGaB5
q1/rOcVfWwKEytdzU19BXXpRGRqktR8Wzu4ZDseHZLfrRSPECvdfR9TjB/aOJmfiVA/fEAkA3lwK
fz7No1celfPdv/5DYLIPGyPBoZk93I/uMsOQdi9UgOaxkbltUj/Jv1zn4LYQgcFSo7ytjGs+JqoF
uSN7SCchBej5bSDdq98uU6qc/YAMIslVvdMEW4z4NZwGzqw0S4ZZTgsDg4MMnUGrwAyz8sjLU7k3
nVRYY1ACr+OeCEFOMoqVgyaZ4NLdn86LfznPs7yQxqdCXpVoG5ncBPadAZlOuRSUqqDgN5ke/Rbu
EjYHv3PZtPTt3AQ6X1bLk0QNATAv9YsPLO6SBivjSLdRcMN8UrWoTneVUcAyGRe2fKYtDNmRJs+q
NQX+h/UfVS9BSN9t9/HDb9mK5aIKdBNSqeoOmmCQo0j5bWkPlmUpl0YtBwFao/XmjS0X/vieFZX+
3BN9fl8OBub56KGGfmBf4XiarerqmpyiJ16LmktAmMRrf8GRM1Z326Ta/Kfxe5dbbdVMga3r3N/2
p8z/pe5QyUrJiGym++D+FcXizzP7xe2/XF9Bcu/yj9WJ6LZeVCGKiPc0WRjA67FPHFeHgJxnfMgR
MoKpCEFgyvQYLM8/+jB8mhKf5G4gEaciJBSps1pL6yb9aAV0w541Dn5QDTh0kSuVYOFO2KnTOCIW
nKlpltFsR6BaOOvvz924JTamfmVcwqn5bR8krf0yxDeEgyAO7wZkgawtw+nBKZcjjdwNvB/65VhC
fpcQEE7xaePHtuzhH1fxLUbo4TzpagToUL/mI5rem7Fsf4nruLjCSWvl5ET12sLMzBfPx7mrWW7+
lwRsFRYmX5pfW5nIb5oDv7RvlISJlbFb0MrLSg3ni9vliE1ZI5hlHUx+jgm/tklkUZLjHg+NT47z
FNgsBqLWj9I2MGfU+pk9KNwzmAHizkQApLW+haGAb8PvGIBjbJTbIORoQq5P5DvPq9EkDG1ArGHA
7xSTRcID2GFE/WMGh0Yn4WlW1fJyiUFwrUqc58+gI5hl6vb/CG2zaqDQ/a2x7iwZo7LpuCJw4R42
wSZXdaG0dxYA/V29Yt8mbMlUfFVb+0RBPN/mTeDls2yYIcD4W+1HoIvvwB6q8amIb08SQBK1kLJd
2ohMNe6P9HC/oycW3lYv1lctllF3LZibUnd5ln79hJnGUXzb4nHxtbbIimbXbLt2mDMOYsznoD7w
zXSY5z7tUfIzba9drRvw46aoNJ4g14Na+ThWSRpr+HWBJA+c5Heqnks0Y7RpBwQscbEhx0YnzJT8
lLGBwj+QpncVCPwJgU1HIXBslGWEDMd2IXOIWkV8MK4G6msbcOj8OwrAfEcDmwyT0B3nS9m0mKjc
CqaRF/nf6Kj3M36S+HtU2/7ZM7FbECUyf4YmHtqnfXoHZFkoBBYzWzml+uEenvYm4zyRi9lQ8abN
lpCHvzPBUKHYAnQS21boj+zWEPPkRYV23YtK6/vhV3yFpJhdUhXC1wHu5OsReb1Wpo/7uoO4QTaf
+JCqZ69zPEKRRl/UvWlsgEgaM4YmBA+ExgTi/HG7Rrlwp9gzi5/IPpGRcgALG+/GCQjg045eRyD7
3hTFI7+8ZyT0gGfA6gd7yUS03dfSCmcINpJEQL1q2VkW3L4Ch6Z0aBXhk0RBLQHT1B6HxcSZZL5G
7uiEh+ag+NfkprpJt+ABTFC+k3W4k/tMU4cbTHlxbJz8Dr82gyLYK7MhhOgdMT0VI33JXvKbOPQQ
VuK2fZzXU8H53ZdYOTq4AnvYV0pDmNhrRW4fUzqUi+nvoh5TDy7hfh+uJ5L4dhnhzJRgEONRhMcw
vpqMwLGIsvAuav9XY4xSpXAoUsGr4yAV7bamr3C1PVhBIQbQCGYOyCCGvp67zIZGg2wa6y17aT6y
Cy3eoFnInAgNzADez7PULMbCUN4/cDs+lQZyX0NmqsoZIHFf9h4LxfO1mSEUSTc6692JGmK5SSCp
sr8haJqlL+KJciZSWnp9i+ZPtt1M7TT1HtlnXSZK6gJt5l/FNiO7HzHImDaRrhdwR2ywynkX7s8I
nIpUhnUB/oZ+ICxImYUBncxRs1UkhO5iluV5OS/cBhO2Y+XQDCSQzcIEXcH6DDPiJQFAI04x2jwX
W5KvU3NJqIrqxMszx24l5x5EzJxdcXand4DnzrfKpMT4Z7JSGq8y3IQeD5meD5F0EWiOax3ox7Jg
Ol+y9eJDEIpNQtfdD3sUkps85JqLAH1K98oLeWJk3Yn9pM2fmVuz0wFakRdCOrMrXVg8n6Rcn4A9
TPaBlI2u50RzTHSDPDlLf7T1hy5ScsfKwL0fDB3USx9dNiD8rb+bZl5YFJLXg4yNGeYVDc9GFDN3
/H5GT+F8P0MPaCHsM24B2lncBP1DYrRL15sFgmv5E6HYeDfAaFi1muVmsYTXi16NsVV53a1RIGcE
WczuekWdU4Ywo94wxJ14BhAb3wRyOf5o3NRbt4Ne37hvKPMgkd5y0kuKszGo+Dl599nNYBtDg1eC
NcRMHtvvdYqJYRL0uYz5rCbfkIvJeAVI1kJ2uKqh+RlXlajbsQUoUghLlDW1PRkFkzPsZ7fWgDaK
363CIpfvtSeTc0kkGVxtTroZm+WTF29WZNktOf0YNTepwh1//FE+brxa9kTymb1DId6B74NtLnn3
nzZPWph+U4xQ4S9RXTrCX20H8ErgMsH/f6klSzP9SfNkQdNSBivksDt1x9pQxtaViWOS7ieFwYEr
yKakv3CPEf4A6lvmRzhDaAV9xcnRJ/VIb68tLCLc/AqWCwYTKpk9h7Q7HtCtXgYw46sqi0W4C9o4
IVw8ULAow+v7MSv5fl657B13p3tZSDphRq5m5bjWBqQ89TDJmR4McKM6ceA8TUAOCPbvo4Ylx76M
qDCCNW0i5txtxmfU6EZjO2fIrzsZb4gobMIatpf5tyDo1pU7s2JRSYS85aiGTiTZHEHW+5+UZaqn
/k7pTJ3dDNjnlNuJCYJ39CAl+69Krn9UuM5f+nkJ5RRc/2ORmfP2cMRMg2noIP29IMp6hZDOowUZ
M23q0MPqOcBWumxnLPZi2kf4iTfFtwDNEdV3JHb/0u1EKOAJbbPJH5OUzckgL3ce7vFfFJK20R6l
SqxTKXIR6l3kOnSXCkpT4tDJpyxqhf2u5cQFNTy2LFRlvGkdAfoJKDou529Dm/AWJZvQORLp9AJq
xmKjisTTNNybFAA/pe3F9CWkq8FfLVsQaIUd0HfP+ZXBGDlQQ0cPvR+RGsXhV74qFHcBhw7ZqFrM
L2Lu7a+/b46FSUucUL4WPkiq9Q7Q73zdrAPNLiy0t76zDOjs+zcp9XFXwBG3dv1UawZBqv8xCtZg
MIrpZhebx32P0D6EDely2w5jqAXpm5U1fd2LtnKvkPaI/B0IICzxm5qf1Rs4RBei/eADUYS+HkEl
tpjZH/WkuYmps/s65WdWVdruCWAkyY51LZg6wQzuR5VshyjUkLDNK5OKwJKIZBMogTqFFTKxIQb4
cvpyr3sE3mPpNZ1OXLwxCfGEZ2sXbZU4kqaA70knQH9B1SVJsx9Ec/e/p7afiDU86ZJblbe5LXUP
CkAhPCm/qimJRhg/YL6/Qh46g8k7p734Xy5l1n1+NhUhT5VMIhZvn4H0a+8ad2apE6N4ZaWujgQd
5KmdbXg+2ECfscEwZlM6PQUQwmAL6pB6g6lLPd2jaIOWDOX8rVM/pOcnL6q0tIP5dYAUWV95V1wv
62LR/qMHeTn24z3BtCfv6578mE1drZnFO/QLlSgaIWDNC1VViyqw9wIHr+wLd7LCjMRsHZemyJeb
0uJVwZxPwVUcZV2DOTuXzXZfLCk/uL9kMY/zHDEBxqOCtFCus78QVAB5ClSTLUisctUGdAOGsWFF
9z+RubdzNDrc2uV7s842b9j/0Xg0BuG6zmcSH7+V3SVflXI/9NGusnioMva4rgjhncKhEUGfBKvD
uK78BkTekrfPTFZ5RqXu7DTX9RLbP37BkcWjsiBOyApagf4HpnDvVM8uE4Uow6qlExx/qACBFYVt
PB23MdnbA/4AKk3mJJRilBsbIloeik5NpH++0SV+Tc3dD1NNmQhadWx/xWZsjH8Y7TVAYo2uQ+if
9BRATYWScuotKS0eACYJ9yZeeiVvAfblvwgqZh6nl9s/o8+DlcPv4eCpOHJxc4oiT4G5SnkH0RqB
eP3JMUffJ55217GxYUWRhWIq4/ptEzOudizhUrt/yUXQZePlRMX6403vHD4Zjbp/GLLUgA7L+Q6V
ddK3M2LT/Ux6BDR9k8bcohuj9kAeLSj8GBEnceJ0nJO6Qo3RXHukBn1VMbIHeuHY/qYf+DZtHEBy
0sweXTgafGBW876Z+sEdCw1fqoo9i0BaO9ouEp38DKN1DTwtYlOVom+iNPQNByYXOWDtRUgBXHn6
PjGrTJLPhs8PVU4VzO0cPlWgwHA8Gzwpi3fNQt+nHKZHPGWk+BNTQzNfyKw4ncSPqSJWs8grgh57
HSBzS7c8uX7yMldG8rHVY07siVubu8rZQxsTW+gFtmBDT5SRuhL96Q66uUVr6I9usLR+Fh4YeWn9
e4nNSH+I+0gNMDwjy6L3NnlvRKYH60PH7Oxu8Ku+wBJjyBZ2iHz5UHVQ1hUNcMfkXQOfSwLAh8+z
ZWC1Y/3a+55JGXIgNLyBpJUJypWjP32E2BY6xCPVqL8VLO+Bxgyxec/Tkqnxol/uiMyXOrhtCaMy
LmZvo4R7tbTdjSLdbu6l/ukXlY2EcOVLYas29OTYxaZ2d/CwycLryq3zv9L7gRjFtP7l3bPMZoZn
S2kenkKwPJWXkB+ZaZTiB1TmODd1Tqg22dGo/HasPqexFLF0HfP2RD5cSx8Tp7y/o+BGrCeyDlI+
C8wa3QoMpSrT4wv94MCgjUM5g39wLTCkcDefT0Oz88cuw8vGmDyYfQvOehlWZZIog0BkpZ5Ij+Jt
jdAeGgUUHKz9ngoILrowdLUN/79fBsRYT6QyP1jIiL1eDAL/erlfWxDlwbqGWRXWy/jCBe1krFmC
SDd6RgX8JwTBoMtPQgk444zauZcqT0MJrLf+fXYZv1cxtR9eHMVOBnqbZuX1StFjYrf1OvmJKXtr
SXf3Pfvjp0idy6Ja4rgkay+VDxax0fUbQvmk7YkVfYY40eiL8HclDzyDRiBCgXb1UCZazbvIBXX9
8xAYaUWLcRYgQBddYhEAHybD8t5XD616m5Z4q9/FTrIY/u9KNxh1J4y+pZqUOBAnWApwQu5sVnyE
p1MQic72i1kGZ6wFQcK6eIaxoJcOvble62NCACY3XVqTU+O9HoIXHQTm7fawhMKVH5fTB8rFMRq+
s2yzRh2+1jU7yjDgVr9e6k0SZOtPxC9+FfKSMNadeDuew4BJX3fvhMui48cH8sOm8/f/SCAsLbwZ
+1Xrk4qyuwOA/gKvql75suCvSPfwNeYQlwvZoCxRYQzhrJg8dSDD6NRmHzv6oeK/1W0uUKInHxE7
pW3i4VLrvVnV//c12zL1ULLnSLcJsrf7xyuSEwLZMAP32OQ401cvWCa35MNV9EM9ls1erq+21qgM
tHw75Wd/WCOLtZ3fN0weZ0T1D/VWmJ6aGea3WafxFtFF3jQZ3tOV/tPfpxKUl0LvyQqDssO7ZWT/
I1LxrgGMmhZdDgjCjhzLxDy/Cqt8q//3mkvAj/dbpqOdR875E0wYlqWi2YkRA+xb37yivppqRRp9
dN/kHNxoSTPe7AbVuYWA6WDZo6WXQgTxUFs3WPVuaBkyLoVRbUxjLDizB4vjVstd0fU+HFcEPO4Q
HKUkJgxxHzyF4ZJcDIAIot3ZXj0JzlyV9BFaua4H1tpeTV1n2I1CEahnooXUqjLTa2EqJj+MaiHB
0n5mr5NCCpNWtjdYBdKKDC7l51SSGakmfqShNnOhcZv1Dc5VgC1IZYaOzt7KKGbzgR5z/iD7T6H4
loBvbd5feSwOkQUKoj1rY92WOpORNImQAKQ9Q2pUn09D3d1ce9SJmU8Y9e0+TetKgW+y2AICHDCf
YH+jwZjD9Mltm21WzJnzMp0RRJEvhhqhZhuoD3ArzWjevXN8tv4un5W52orz+K9/IcR9smugcVGw
jPGbtADH5FZK713dLA1NjI/Ca9dZAvEdFp1iz4enMrsbuHOyKWyJ/elA0KkTkq1CI2Nzj+TFzMU9
+ClCtrzTVyiaoSte7dCExpuC1Zj4P9HksHmCc/bK4H2KDb7MlVKbReviBoYlCQS/5GMn8/KPxqSM
TLx5UW8J8kGWCn+llDduRSMqUU4fymtLd9xUzSzgcbR1GieFai4oRdMucxWel4iHLS2GhR1A6scE
E3/EYdz4+OAQ/c24t9ZPVGrUR1Jz6TJFaozWnMn7ez8kH5Xa3hRZGlpjho9rPMClrBnBYAeK4lCp
geTuYCAeVIWcxjz3cL9lntquI8+4SHGSPs5SYJhhVz57PgGMOSlLrdHN9rTx4mJIOazhd7tIxJ2+
RxI5JnTu8F0ABSwTqrnIfJF7aEKzH6djIbZspeA2YOhKZHbx+pg6mVr1A6CcvONgaOuMXiQU8oxf
q6/TocJsoW4fyJAwcu8FHFXWor/BPdXe34uNBe9feFVRMrm0l6Y3cBmKmw40BZyoAeK2n35vbYt0
kIb3LpvQU/UaXcmAm8ID5pTKdMZoZgzes16FurErHzFOsrWMmYIdSAeyvMPLQdLraz127CXVL3Wc
D1fJ0/99ZhASN0nKDvN1RiDBdoEUapk1WvY6WbYBPym+xpXRs9Osd9JWT5AQDoLp5bCDAl7xJvHQ
Ceu3Wju9D0TsIr9wY8kpxk73FZec0Te8uxAd/jwv8Pai8JgEQAzlrpS4OMyHeviuBQ5GSlYE4C8S
FFzxVyWsqVcslLqrP0cfLPr7sBN3bIwHZ87CcFp7V2H8i+xWgyFFphuoIhYIben2onTEnfBJxQ3b
PqLTf1MwNEH/QboG/SUeGaHy0Y3+t+qgvuENX1ntKCUp8fy0z8g9kSRDyTU5cPwkpQnMgdl/14cj
xgazLJ7YQFQqx38N/pD9IlLnyiIYUHMognLuxyp10TuGbl4KmwoeUNLz8QC2eog2jmkoDkK33txu
o+pp+NItoQWJLXIajUf+uygpZDzHC39iPhmuz77qZs4MBF8HDl8VMs83jK+mxq4huC9zY8c4R6Tv
v34BsZFGi3efIcPyBjin9JEkYCfcGofkf71Bfac4YuS/2P6A9/WIBHHCuLfJwqaay5QGWjhPt6D0
7w6WPtGcnn/Tn29vNLDrDn/HKGWZ6ekV4jA6Tbi4NXTOjIh0tjZHsm7WnJ1twYbiB+niSC/ag27O
WMKcyfwf4m/G+SxO/DrR9kuVOPlLwclMgTk/OV6qFSZHqPuO9g6BRrdanSBDjFxT7JQ8qiAVhs/Y
WPgjbpntVSBxCG+kXaBcqEcgZqKmSUn5+f89/b4NIwg/+8+XhsTPxePvaXHd6Z1xGA/S+PJW4y/F
QSXBuzZadAZMgClP3Q5QwQDrC3S9M54gq4pce+F1IFoci7SAosXxMKxYqGAOqgIUzcEGoiz2xf6Y
ITSpPTrhbiTmgrawH+1vn1u/9RoeeYfsJPPF8v71IV2MpEg0xuAaorMz+sD9tk+etcWsh6Ux5bZy
Wj2z7vZXhrofM1P+j3fmFNuWblxu7XfTov59NZmVtpktuL2Q46LEnsZxjLdZD9VE5ZOueiNW7IAE
K91CBnP2d2XI83U1FUhzhmBorZU/nApk6YP/0RZnEaSvJN25J1A/UJDzZD49pJKAhuxHOQ3qA4pv
z8DMnelIcq8mshgjCzeXrJEpChm1D9ejyuV+LB9DhyHgWjVkiH8cPkaiy4FqsWDL9Twvp9hMYjzJ
j5Sdrxu4sbdJTjdW+Fdl1z6DuKUoVI56C3znz0usx5qHKCo/5cXIAZYwY9c9oIpVeEUuDz9F0nIH
2/H/a0JrsX0A27IHhu4Hwp7G+1Ati9oQ7YMTvlwXZZiJ2rpAMsq32//DuD1t3wOvW3VLtht4lEW4
HvlZiY2Y8IAivNVas8zADxfC75BBPfJ28GvHsf0Q1RzQOaXDJWg2UUOoLv1IJntpLsx7BoKjPTkw
aHHCJ7tfVv14LqDwXBzuCNNbYeOjllpZK3ADf63qlK+DvBQ83blWAP791J44YPTLJLYThTA0KOm5
NUvjXeHxnYkOmUecclJ1rt80TPQl2QmBFl++aRIxXW/X6eYOdSJyPuqQ518ugpwzYXcHv04wJeZ9
3hvg/RgCGosr5f2mZJoLTM+REaLMQY1ICsRcknYi/M8fWqhmawhfuZWQuuhnrneXKEeaEXYNhmU0
VM5oJpYhIWEaEHAepKQtQL0fbPUpiqogILbS1S9WJTftbZytNhIUdYcua7i3Qvu1V4itMArGah1R
xas98hO+pmTcsffNwTlYHEHD/90q69VmBjWF90St3u+UpzRohQwUT+/L3OpGAhZRzzWQgz02j7H3
KdoSOV5nVZEXBt6/FKg9uxdFmrwUAzRi7q6UBlg/MP9G8p9Nmj3N4VUhYOYsWpuRp1agKCt0LMWY
G+XNgS421R+aX00RLkKX3yWauFrwjHyvsqMfGk2QKZ4P/RvgqURnZw6VKwk7/oNbbvhybgKqorhn
m5NAlXbl8quSpC5vHDMA6syWXbvJiA6UPNb57+Fs+N2zMtLKtV+xu94/KNS6El8md4f6K0TVS/rz
Rb+3tRT0/mUTm0T199cYolPEa/FUzCKKh2GEart3YC8eYDuiAUz+aRV+/wECYhw4x86loqHMKkqG
cSzTt+5BdggywHlUSSUbBjipFlsmrl6NDp/7tnfENNzh6D1jtKLELtsXmDjUN7T9yvmDiAY0ppOU
a2XtTwh2VxRNxAb3mliQQDAwgrrEmRwBwUM/onugdMy7xOcvb6/h2Q+jk2lEgYDO3GzvyMjswk1F
LpQbeYn5zu6NE5xstUN/jRQEBV8zIiqwmQWFxdBzA4StqfKHL8HSnsjARXgRylx/neoPi3BfEeCy
xrg83z4iRi86BcgDZaSA53rf8yjH7VG8yZX/NZBGOrDlIQr4w9jWxtjtJ4AwS3jhn1wOVAnKtMnx
vGfXbiDVvwOhqGxFAW1MZMH7iBDL+inMrk4BCmjDnLNKYm2aXSvKYgO7Xqe3vvDFYqiofqigLaQV
SpxlVYCMd0iR1IoDUPupsv0/EGXorsFKEX4AQewt/zA+Q2oMLBmb/4/aywHdcY+zfrB992RY5C1L
ixbC8JRH/rxV/1r7WYMgeV31hMqaUXop4dRNnAgtvKDkegSdIiYptvOR8NhAspQM1X+PWebtKZ3O
v5/iUhXly1JkziUjBlsLy+KCfatcUx7Th/xG5vyCc0XWgrRIl8ofetQWlp78XFtGnqbDysj3pXd/
WeK7iyGA5EB2Lq+5bd2FH5EjL8cFnvhTJvehNRtesTJqq/gHPIuZkPJtQUvmTCAk8jBdvTjXIkUY
swQe6rlZZG9F/V1zdFlwzLdyq07AnfPyjE1ovsRkgi11sC9beIujNR6cvzK8hj0JLcL7XccISjNF
lMmpIZhmV6pMd2rRMbHF04AlSja4Eb7itteJLESTQJoV1HdWiL3ySzdJfGX018dELJ15uiKRZ2ZI
yIRDQnALzMmmi8DPhA1ZL/8EDhnAlGhay2YGHVQCHB4wPF1d7UHlum6Eqc7i3jdbQ1YMIynwd7AC
CXpAJxA/kF6DoKKBgIdhrvnRsDC8GtDErVuuUendC5ZWZanI57v6F5C6hojqpLQoTwERibMGExFE
WnnS/JMprg8SyL/VAiNnax+41mYJuo/xEREIMNDMwmhe5IjFEjc2ZJ+VyrzRuRb1MNc0bcjun4os
9j8MLaLtGmsvujrSvwKWYx12Nx+Uf3DNhYuZdKv+EJ9DLAomEfCDHDx0vqVXPqVXkFWjY1T0uNbc
us5eFU60II0PdGnWhC8QJmn/zu9+NOkB/8sxeKCbgGNDi+zyQAlc5bS/CJMnBVDM+Pe5XOwpRGwO
D182cdtMlptd3YC4MCL66dDNJHYdhePHLp+ELaHn5w9+fnbOwIKJ6KF5PFb44ZvxcKLVlawLEk0G
zyR58ksWAnYZSn0JwgR0FfDZ2HaG+YY4KOyQG6U5FwgyN1flqXphHulTjCKmUjnnW/N9fF1/AVPX
4EFS1NNdVaTzj0UioB+WrNyAkeIUXEj67k0NWD2WUazjLBxM7wy7ZovjcT3Qe/O7EMHNgogstV+Y
uX4L34IYEV/GWkRFhQ31YAL8tFKFQcE6f3LzoWwc6Aebk5OtICe4G9lgAeoxfu/vf07ZncgalE7e
E75EqXlkQzOueCOGOBdyENbWSz/GWrIyLV90w+W2Xg0oEhFJKzu1AgT3SLBEhlbpnX4HmKvhPTwy
R9GoFRXppKNQmxlZaXNEJeptppOhe5TZ5jcswM7iUe59K1JLifsDE5jVUqZU+iYlDFrUVJ0MZ1mf
/uZKK1ZzqwjiMxJM46EGjjUKGfVtIlHxgq4cXsJrf/bweqUzcAI0CkfEPpk5+j9x6pTk23EeyT7x
BN1gaG/7u0o/HLMWIZbelogIS3Pu2L2r3ZqxMrA2z5Tl23/Sj/mgIy9NMTfr45At8Plgu0aF8U2W
9rlmdKbx8zKTqTwMbpy9ZIomk8BXdXeDldUGuEir8kWjZw20Q2ix2PWzywQFpuXTOdJxLKTktWtA
k/UpHLwhgMiOayQJ63yCksiXiNTMrI4wf50CkY2zxIO8Bo15gS7EEwLhN5TKxcrl4Sr9cTcMj1Qx
hZ2oZUs7aGZzZJ/PBZbhucABIWHI1+GQLccPVm/xCmm6GPLOE+vv0kX9yrhC6qRIRYb/EeDXMqb8
2H6bIX8yoSnQtVzZzLeV34BoeR1GUw8XYRLpg6jq0VGgEfJXyoPoy17PvMKFVGbMA95xOfBPLM+j
Tox06nd6QnTTOQv0xS5yHf34Gx0Ea4UP2d2mtyDNxuGcL660GsJv1z1U13zaBAWKXTLg7IqLAMVt
jF/7KaFDiCTg3NxCppFslfvsPJ2+d04dYCCnKtpTvgf1SgPtTdnC12F5lppVhIui3brafDhfKCpj
DQ05SlN56tk/W7R+FxgeJy3HX026aEL9ynh/3my5sfUMJfN5DEcK7/QE6b7eaWmihMTXCZWysyzK
naAibuxtCp36qEQoWn2yNR/Yt1sgnneZylFsyaAkdz8IeWPYgzmW0vNa8Ry1vJMjWFYOTAag5vWR
LeHKnoHCI/Kd3/tPEXVRJudBjWtqL3g78Q8mChYO+9YsgSOHAPTcDV65iiEMRLlj+MQ9uf2rd2+R
99/Up/e8Gd9xweg/y26A2dG+UNQvkJIuYue0erkrASgTb9yR3gtntQ4V4AqsEh6BtLzM2iHSlS9K
tsEo68OVzFZ6wd3xJ13wCmDtGmYfsQI+ZrDYjbKSFLLbvgvbhpWh2HV5yKqz2GSjuiWp6v0+yu20
MII2gJIS7N9cxwDXEnfFrbbcW2AIhXK93l+sst7JXIsJzm0v/NrVABgH3qyCip/axs2/TDP4sIVc
LDXSIFLV7W7HSQLKLMDCoZtWy9Tqznv81Ez+ONB/8YbvdmwOE43/5y0dCx12xUb7FU6IQeNS7I8Z
iUEjXasyQ7JoGtq4NjT9WcrIU4VA6C+0ksCi4tNkT3ZTEn1ewOxX9fcd/QErCfTjG8fziEzfKaD8
NGl/+LceJjDGeUD8UZte/2AmBkgb1EtVxji49Sf6P8bPoZCAEkcRi1UvA84IG9ZbxxzlshVzSh9A
uLv7bQVxVnP3q3mnObxkujG1BwtZ6gpM6yIScLYpnQDU6dHnRw6JJHPDTQbKwqimhldtLt3yZjn2
dM3XMfuKAdbOXoJp6dXwn9cSYqhDLAWm+hpmKzHxqedPdrw8+QCsLooOmr8ccFGWg6xNgi435plD
oauPWH5iXJD6zT2j0b8rz9iaEQUnFeCp0zjMShKERpNQLMzHqhWIZxrj4naaT2c3C9mkpYY0mQYL
aI7ZHMNvjUm4+ppPgZFfJbBx+XYYt+IwPE2QKBMcjx+D5XDuc5bRUO5c/ZJSFaG6R9yvKnGi+R8k
O4BF3EfQGxqFR6rX8NGUQNTWRnmB+gxVzycqyUbUC7IpawAqjN+r6M3ddmXneW8iY8dAGIVjGuGE
0keWMVaNHM1oLFALTfqA+ZZDRKmiv238cSkZj/G9TIdyXnwvX87Truz787pQHkznCTEZe55sSbWa
Sm35ZBGBNSBTCfRDgk5wd3XvMHMadbQOrkGIcSQVaorEVspgHNrra99f5llcdTBg4ILBsOWSj/r8
ZqLowSLrtPR/D1Wj0nQrYQV7KrFsT/hkoXbMbvye8Ypu2zV0YXf9vRTbMmv+6cqMDSsE0urYH+aD
mfjj8FgH+lhqEgxKT7aD/uNlILBsOs0IaUsOwgjCl6YrLwZoAOk3Y9Tav0QDRWVqpe+b2QbBWR8E
nOlesTFqAPKHkVJiol6r2MDBSTZ2wtjsHNiwBtTTq2n02s0XXzTEXbs4CpM8vr5y+xrSwMV7hBa/
BLo8ReeK03PiIP3Tse1aRdT8ACcbX73VQMg07+98R59VAx7nUuMnNqOkWO7LfN4XMH5YqpjLQ9bm
3KT4RsJAooJKpEEh09KJbMKbm9rfoebVHMdO/K9zraiYleDLX3A0kK+v4p6PbaIdFG6QOkff0rDY
ghFJGpc2ZR6Zk3mlO1NpdfvGV8o1judYQbTHvCT+kX+225mTvfCErPJJDssSZkSfnam7j6Tys+Ic
DJoW810YrVzAz6EVzHlz8xWi03tnQmOBt5WaAnhqVVR5I1oB4KC8Kz5CQNrwtf1h5jAO6lMWYy+o
+HhVRGTlA5unoz1pr8QHs9BiVuNlrynUWZxC9iSLU38zilgF+6i0qDsFlgCPxQVkL6xL+5b/VAqR
Gm2jcMp6c3g1Qr+uzze9WXM4g4FWfuggin3DmaXQqh4wqst6cDkyDGVYwLN6XsXxsVYXVNhjDpNN
4TLVoOMpvUVN3s+UQ3GQJYEeP19HrszlLoBbHqWpXrDTPJnin1HNprj8IPcJmhodeCOjUPSpCTjS
e6WgX0rqvvEmBfFt9lezw4DTtag6tIncN0xRmcwPqeNGdMZ+55S8PNQyXA91w812z2wfcGRPREu3
JA/+jnqxpIG4PHxMJqh5VBQpGS7Dg7JXdpD8mhMS/oIndASYHceXkiqB/V9diq/JzxSLlqEVIqSc
tsQ4rHQn972uCyNTnobBg6hugxMUgNUdbC1XdF9vwyDpNqBJQGpCKodvIwruayCWoEBDimJZ8xAU
G8WBNlUN7j56uqRZ8T82zZCqfnQW8NZNfWM5s/IfAVadt/qWngenCSLNg2r0G3PXRc5sToTvSlLm
g8HevvTToeOh2EXzkBcIczJ2m9NY4SaEh1LwpTBS1TZIAbqelKsFAXFxkAX7xYINX8S1w3LDkFoS
ORCAAIBMAzSkqvPC5Zx1WPXB4wOb9MmKyIbix6ZmGSOAwnpDSK58n5BXHnRPPadwO/2yAN7RirBv
flXdJLh+LK2DvxEu+vxCgYS/HDhvRM25Y72INz3Fg+w+LOMg8oqFvU1He6VIOgqKe3f1ZKEpsrOf
+c85lIh6fmDnZSWTMGu2KHaHNYAOHwQE6VSxewEFxkrCZoFajAJnTXFXPzlb83h+NL7OMdEOyIvc
Bl33WhdmaFRxPoes4eTin3Z/DjjPHoEBbIMh2mofKk1RGVLUQpguL4Sxi9nILgcunoTZJeONMpuD
Na0j04H2APHdKjUNrQJfIFchuc3gV61LUf47esvZnaF6JxikkrjY8P5/Qt7rtVaNDBqzYq/0kfjl
EVHor35bUphg23leOIn0yGm+Xgv6y8OYAvqRaS1wOyH7M97yKJMelK1JTa0AEMVlprZ4zPTyuqBZ
KkhqaGkphVZRREzg9yc66z36anoPa7Qt3SZPcEfo+907utB7f/sYc9lr79JwVbQ7QNr4ReeJBt5y
7Sg+1URFRc6F2OamDFovg3DYhEvnY/aAjH3BJ1XTfENc1ktYORNYkRbFfoUNup+PcMmnKphVtgy2
wxh9k7Q2noz/ABRU6qogvkGmKJiJ3+auaw56gZ/wlM7hH2h4SNWsXv2njp0pbSOIl/8WIwPFqOBk
Uq12V284VMgU7yQZWgkCUFFpgGrOg3NCHYgT8uHIOjiTgUqgh7Sc9g/Ls8BcmXR5GFhRznxKYyzq
yolb9xfsM9tUskvcrBx/SzUy+ExQlU17UownKCHmUP5bWmSg7p+n7BnCvTnDhdI7qTnS4SV8BWZC
e15/NYwHJFrOY6k7fi3Hr2pfCoQXkoPSwJq1MnYF8M5G4a1P5hb5O/t7ZBqO0N8zV6uUrI2/jn3N
GHU0NNC5b+L8U+8lclwQTPFX9vZmp6EXg8QSu8L4zGoVuHdV7DVJBF5vB8wO2d/keyq5KLKEwDSp
SWJ/E6hnwTJmSp51E6+IKzp8jMwVGQHEqkoHtpPKYOIuBr5lv6ewCtcQIupMKEKYmPWB9ExAJl1M
Zeg29P4b4QpLL+lXx5yBnZzPpVPYVW2I1KBQF6BX8wPtjlkv5rj4lF5oSerDYTEw6UD7sIxruMvE
xqYSswGsRgDavk96QQ/jj6ptP0yL9PBtSAUCXE3L89TGEt48e9jQLRqCfj0KogSce+TR47VSStuT
DbNd2tdB72aRwcDTLJupuLxwauaPjNVbdzkVrTp4zBRdOYfDK+E1H+M22FefjEcasLc5w7UvOs83
y1OJRGews6tMswvISyJI4Dmlq7aN4PrABejYRw1qwGFDtgPt1fT2S+SCGcwPhJ9PQP3/CdXQc2Op
ZmU+ZJncsqNWIn6jMCvTZOZAenEkLYej8Ij0o3o+0hoEYWB6Y4Kd+SyJ4VilG0gTttLnBwiEr4HX
qPdTdKke9ZViw2S3d7khm0Ppl/vYTpkslEfsEEVWVxYmhU0Tc6sPZeASO/RsseyhH5N5ip97ytR7
xTiDRIxfyO1CLVv0Qw/Oh90Jg7eflbRCxMxCBYYXHsZRasq+bUJhbmEr+1/EhZRBfpH5y8WO7SI1
ZeRZFgoaHQm4Kquc0dG6rU/dW4TBJgRBDD3Cy2rKqJoMaTXaBf1Mfd44+0hHAJFWUGkuF0/EZBFM
/fHcjN7in1pZ0eO9fE3EAWZL7vjQCVdsl0LzAq255/i4ro1C/D0xbEwBvIPddWtt/VmaxY9IBRXA
lQFtYMZnPd8FAhfONgOn5VWCCS6mo9YYi1lSTAYuW/hy8EU/b+7t/BVigrDYJYWlfhkXoRckYBQS
FVKUHyqGD96AICRTslcV25LUzLCWRLqwzYgLz/auI69XCksMos35aELcOOCjjlqHHOGULBGFgEHK
IDMY2YCjPPVnOCSTGtLz9m6iYODG/fTXESA7KASI7cMYpmaYwwtLnpcErU3bbx212WJY7VAAjZx8
trrS9ZEzXAzc65kxG4tXyQzh5KTvnNRn/0VaJyrul29OhQ711KnJmIqPbk7Pdxvqf+KxL7WpuRUd
n9Uwx8fq6v7HiBfyPn/u9RytFIGYLz6NGV65hb/ngX1rj3JZgtzScpO92p83CemrP0xmWzPm8ZyI
3TNyF5mUF2y6ebH4DS73X5DolXMpzaDxKTR4Io/guzwsbkQqJu4ybDH10O65BTnqdI/C54ng7rkK
+t3zGgS/JhIfpXEAAjIDuATI2T0WqNp58tRqy7rHcRhf07CItyuUcOroDcfbqXXtRNkzGC/pQtSY
vl2p1iU6zit15gXRI4ggZkTxIqW4FtAo2yBnuKCnLKPE9+Gl7LQmj/xP5IJTe1bDJnn2LUWKXdnL
C4KOWutz1Sdqrn3ocqHsDggwKo4p33LRupYNoLj2qUgDjK2J6awCjTMsJLar9N/wAWFabr48b4JE
gy8yrCEniqrYLU6HE0C3bUzJ7e6YyZGGo+bVDRKyKSt8ANMmiZYzF+2wcJeR1cVKNSBfXPLwpO9c
iXHmclOA4HGmvJJQzrEDhZLJAkRtG3utCd8i99cc4whb6WYFRGrkKJqKlec2eLq3WDGW8Wgk3PFV
u6fdKW39dDy5y+6f3jtdxT66ngNwqHV0HU/fMspuQfya43S3YpN1MsLpK19NY7hM5ZJdsUSuHL6H
Q1Jx6gq1/6QjJr8gumLKysNZ5iVYTuawiXSbRKsFJHtyvE+D7wVyrzPWtWlrIwAGDnXRhundjozv
SnHrfVH0F2PMm7Z9epIo1MnI/VySZz+896xoM7c1EGTOYRFfoOry2MZnd3735wfMM2wB0pjIfRUJ
xqBbCpBewzG77reFKVrKPo8PB5id67XaYP2LXp68XFMkPSkI9oFFrESMC0VoTcaZXtMRtnSBrAX4
2iwiT/XLC7NXVmmlk+5I9jebFgKVeKZbzQU+liXtdAbguplUC5B44rHnDggm+uu5EESeukYrvEdl
in8xSwbOfAiT7/hbc1SfBv8oNNcSESsEYbYjuwZ387lX8AZziF7pQ+wJdsVnMI/Rd0+r90QiRJYR
/r30FDgSGTlyCJWRwl73kTKC1Rflcfwbj3K09hCEI7hsHuj37ixJblnf3KRx2vCzHy1j05AQO6I5
Dl5GNAAAe9691eeTgQx2zKRucjt8W3ZlEo7JZJSTbJhbNOg0wK9p2h6sadHizMLKf1lSUlP+k7Yk
2lgBFz2e58XxDb5qKLxbM5NTcq1WCZrGCEekUxOl8OlCbe1JKk430FmArkEi4thL1VBoVbmczSrk
LhqdV7N2iB3bdjbym4kfA5d8Rrx0NdJxW1ZT5NYDeg8tlZ0DsSS5+p8GzoG6h7Y0azLgA54Q9zbx
+lBk+PVhP4OPjBTwqyq8IN2WT2IrH8BN/Q1EU2jCHXkifxxH+qfwyg+8ymG7bQH+Hzmb963LuYFp
SOgFlJCO7uzb492Eye560xUpmkQGodX7NG/DVPNFmk778aBMoDpB/DXi8Udn8iiX6rOpiA1dll5N
4paAOOntoNUzXWLIObjpVUzSf7cZ/vgGDmjnYe5c4w/0uC9qbPxmDJu0KC8PY3wkJPFq63pMYRZt
L6GvGJ7Y4Z345QyFfCU/bjf4oPDDXf/32yhPtYqVk1OXG/NV8RskNJMrVSZ4S/H4Al4heclrDjHx
UvFiCzFQI1GkFC4IaJO6hZViZx1AfB2wDrVA0gON9sTXCVKAPI4VPRQx0behugGMb0Z6+KPiZmLf
zGca6nEgKRUfDWG6Cyp8Lc4OCfDfW4G6OfE6jjxx6oi52nD1MneOgsG40dUGpbA/lKRn3akk59df
4SEPCqCcvW2DBAyhQ/xr3D9L3BDmtJto8v71rTjGodcR+dDzdXpAjSc+MKZsoRwr2OqrAqY6YSLL
k0MvctSXkkmOPyCExwm4OoAGOEpIzxiqbkAw+0I8JPUmk1epZdcj44GlIrWl1owG0JLAaCwiXJCK
jAERrhL2U7RzYEqhYOEelXgmqrSeATw6pGgH5R5mpAvcSzMaFuR4Q+0ySb0fHXMHn7c+u7F89x1O
Y6dglmXmhW9wue2SwnNsgaMCM9Tm84YniZpIs2SXq9gOB7OLEk4h+qTkB+z5uujC33rSCVDx60hW
/tL0LaNrI4PhXXELnDcMiWSCJsJU8TE9zTFL2MQKZ7lJKgL/jchk6Y+xQURM7dSZaze8NEU26D3J
3scfNGdgTcgAF1LpSgaLCurVPlEye8xc1KqlkYuPiPmuiXjGnDzfbubJ28NqannRmvIqwZ+HjryP
WcHZzMp/g9Y2uc7vWCakLFrdNH3YdAvopMlkOHNsx4qxJ+r3D5So2CcjWBzT9U2QOhnyBPxW5ZH3
ZL1UcPursTT261mqYCGmt6MzxwaiypL2jH5uTRdpag4UBvnYFDgvBndN73QcZaCGlWOBNwISPGFM
Yhy5/Vq5QCuCqp/qz3Fn6gURpQzMLndHbSe7HHJWoMkgTRnpkfVNwxLFXCjRiyEFqUOrkt6UvWtJ
1Tz+7IugLaeMjL/+WqglbfafNk7Pp6OlrnV8uf+HSDpjltz7Y9RkpiIYoXvBT0YSkjHxQ+p9Tt/u
8l2+8NqNri9yCEkIzqkF7d6DH50NEuKDsAiUtcld/5xCwTwmL6JRG6sda74MSqc3vtd0PF/3sF5+
5zCmTCkoVA3Qf3Af7HdP1I6pStH+bifdpAMmRZOWxFtLmjeAeqUD+GJq2mUVgPY5zzgT9mCYSM54
YZZ2v7kriFXbMUquzJtz7nZij0XSO0I/LGwNfankSPuOhtC5xe0bUioF4b6ajspkoHjrQmdF+C+j
qFsS8pyFcXb86Mc/6odBtoLemQnMdwQ7w6pLKRvw6pkpP2X09KMkHLtQVgxAl7b/7GU3BK4SxpnK
WQ8b4I7DYn2ARq73Cm97rAmdRWqZhtKkmRRnCAkozXeaRExfyz+SPuOvO1AWxgDzXR0QW6a4EyVu
YkVeFwKvk+jRi534uTgz2vKjEKqXYQW7bY6EFbruGJIUtQi1muKYst6Id0/92uDYBmY/43cPpEBL
+AsOLveTQtBKheqh+4VhAoro3QyZEZTJiJHVmPm2AQtGfkvQiQguSwBxhF0aIfz91v4J4rYt4GgR
jDGLToeV3N2lXhnSktiLx2/npUPINkF7uqT+TjJLExrmhopcOcI6N4Qopy8E0ZkYrOEVSRfJ6kUx
Ouhg2DIi74Xdh5FcVsd7/azKusYzfuFmazCrNbMRboNDc90grs8nEPBqX1PXM2FFSJ+b0ditHXgG
dg/uFtCsnQMxdljlVnaMItkPZ4qcc1W35PmsKrLT3Bg9xZPStOpDirgf5zG2xhzxzJpXXe3icIz1
SSdWzEzh1ZTkK9G2bshcrJEh8sHsYHDDWVWK9xPOGUoErX71V/fY2t9tEWUAVs4jICaMJ9v+uiVY
idzacutUtfBnjUyB1YB7fpDjkoImMyndEcr8kom8I41hINmaXg5qCO1tBc0058DMJUW9vAGlRvHm
BO21ReR1QVdI35qhE/9PV0iLYMN9kQzrrHoFDvl9ubNhgUXbrGNA90VWskeyS+Cy1fOGwQHPXbyq
TbDZDDmeMx4BVUKXVbxxoMseKUBeS2E8mootPDKlUbdztr9scTmj/bVHnzCzsseT0QoRTiUljrh3
sdy3KgeMXtBHrVcDTSrcrXfFGmgFERVqs2xCA/mfEs7epnQCvISzoQYpZmH1G1wFcHk/gV2Vd6gq
ema4p4+BZNcZwPbTtmvdCntJo4moHqDZl41kbzsVggNEGY29jiwaI6wd61A5KIX04dfGsEjibQkn
woq4Qc1/GDZHyEMI7KsLa45xq3XU+g2VNzqgIWRU0M+3bBvkRowhAxvheghA4P5SWDrahwRffx3i
q61QyG45W2/mfroCsg1MoeG8/x5UBtN4dn9/sZZZS/sc9cpI9kkisL2tFZgVpwRVete8mZJ5FNxA
T3eNqGpGN/ZfFhDvOkNRi6j8JQOwiVsDDMM9KuJzsmXYdL2iSBxbwQ1LJwwSwnwo4Tbl+9UBoY5d
7hBTyNOAoV8WyUBEus/ZZRv/dTZ5GYmKmUx5borgrH6PR+4d30lthxNYvZ8SOUmlGbHf4cz2vJpk
xMxC6NGoJNpm1JHejf6LPGnXfoOrxKXVOixVIIi1T6E9GIo7tC1GkwhW7SHAlpuObEzOJXQPQdVD
PqHBpQVN4ef23TdT1M+reyt/zTS/wIgM7YZSuekshJ8DrP0+x2M8hNPyPP/RsRyXmHWLeyEBPP7K
qlsb+mB2knm8gElb+9YeBE7yTKDCPGQktrNOMZu31ariM+UIQzyetrgoGwxqE5bV9gqqklwiToP5
TLsDbwvtz6mUdKPYW23fg6yYrQxDZeNvoC05/iO7rawvcs8P8C6fHqXH3GSXl40DfHsFB8O6l31H
LOfYTlk3vlWISeMBUv1cOEXn5hoZIlrgq8A/clFAZzAP+l9EizsPppWF66gXOCz4W2UA2qWjD7q1
oGySly0djvDBxTU/F1bGUYldK82v9CV70AT6VfkV7ZLJOxzI3tZUKw+7ZLAl2+ReydQTXgeLlffA
WnZWBVop6dty9bfgl9HeoPimq3m1LFJghtzaz3GOx1m4jjR+mOI8HYwXIjRvZve2LKy8v/ByuVKW
lx+xk1ztBf9Y/UFvry590kgriFwWl7G2MrOqzuP8iFhVuWPuMsVmoCdsYqAAgo5fGXKWsXSUkxvv
6SN422tdGIZB2yvT6ME2ICmnq3R8YpRna/sKgQg0wzA2ft8q/K4fCnwZQGUfHFkQfasvhA26s3XQ
51D3RH+HMqaADY0tjI51DcQmqyxH19Hdhmb1+cEzHT98zIHvvLqeq8cT8rv2t5eZLo07WRVXBAJa
yelGymA7GXL4SRRXfUiI2grVxtXbKap6jhft02RKhibQSvyD03NQj7za0DFDBq+JoM/ZrM2H8Tgd
1jaIo+rB3QBhL0FXQmjvWE/0n8oK1WTUrzsmClqxbGeXP7PjvxWKcZdUQg4jwpQ4A65WXzJK3UkW
boXJitEChHaSnyZCeugnUY+mOvSWenSSqhDRi48Hw1LH6XlGRpOKbP79Aqh55MJyoSIVqY1mbuAh
tIp/4gPWPzjRsVCAsvKWNywIuPShJBr7iL8DBwwzIzhHhVEthUwa9iKkz2kd2u86mPjwmFSHtoAE
DZp3K1BUJLkVzmY3Vp8mfRIB0RVw9ghBw6x6G7PtxBwMOyurYI7sn3Udab683P5R9nojKBaECDjy
eQBUX0qXHklkcZNiAsDEKwoCAQzLyaNG88iOAW4iBIa14syc4rUNdDLl6NSK+NWgysIdmKROhIXF
vmuliPG1WFHiajFuGk93FptIabHWIgiZw7+1ETS/alKc/hEW6DTTAte21JfT5l/c1TyMGFKLUgl2
xPTApTTq32eh+9FKVIt958dibyiKTeBbKmJZN5h2w+XyCBfilQXM9WoEqTife2uYylQUhGgg5kw1
RAElHnawBN//4ipy7iBXBo2aGceXoV17wZpuxMVFZlnn7/fffrlIeHYpHsp8hCGiGE1EOPb3Fvx7
dUZyRxKjRNAr1LimsqAp4nZMB1YR/Y7MONj0XxPyw0zI8VpDQViFUuvs+HM8oXniOO2gHx7qPQBb
2LSdIgD6IV9VYHEtAlnELB6Gwf9SJg6XlLUfotVqXVJnLbhOLjOKnSDyau4DlJEOZ5oWG6IN0S3w
Wao1ht9pYiB/yRzpPE3Kda9eXNtgYEfEfdSH0TSMSX5VQRXjt76HXMFldD2bz3mhvd28StnR5GZi
TCH40mI8/C1wUXzjGu1j/g6gjJSQIrmU01nfn6nkFXolTNoVMt6uEkfNIovMKAh4U8Asy91+ZDln
nAhxr2kGS6PbkQhL3H6HExzRi5mLxhqp3yODGT8YkcqiYpttUj0X5tIPslE0yUDl/ce9otqi9EE8
as/hTizDn/FP61kYc9zeHq0J/0xYMC2hBpe7v8d5IkKk4+chDk+UxNby6D+jc2ZaZznklaJ4zRhm
USxfTALxjG7BROF+pBqr68JGbtBjwU4Is0OfcQkmWU9xLoA3m+8vwfE0d7YuDePXMXLOqptkw0H6
5th2QoPtieTThXdk3m2xdHT2bA9g6XmNI+h4Z/TD4GwkwrSTfSPCww85EQndY3etm6mqBSsVrzbI
MF1YRvRx4UXHG4pDwG4bG676DO4TX/Mp77SPX1fc0nl4zKum0ZO2Blj0ylc2N4l3n7HzJhOfJLxX
QbT2csLKSPFx1/SZThiH5le0UHAVBqe1NfaqRagiSlQlPBXhFlpZyl8FFZZBTFd7eHuWpl1cFC+f
iuztOB5vQzdhkUJLK96WG2+9pFO12J0FSKyO3Vx+HpkfExYlh4L99aPgQOBtSR6iExJzu0ai/Qa3
LYjjd3LR8eCMNeI3kK0WEay3mziYLW8xVnvWZ9Mf+vvEFfDQP6YtfxbvSt9OVSARD0QV3LV7iE3w
lWVelGHwBtB9NALPDLoZfabxB7LomofV5jRpKEUk90KAn/AXgFZOMJSi0FVVrU3Egf2r/pOCi6EK
1rLnFhnKwHQOmGVV5MQ0itGhhv3lgZJ8p5qZaN5C2Gm40v57ssqvmu/F0WQKHcLGR36BPKQU7eyA
ga+EaKyykTwUvEbxRrZ6IVs0IJQMgNNnuw6GJEcTTh9dUn8g4sBetvzlpQVuxzqI4WZBUeyLM4eB
qJoe/Jd6YsddLXV3ZjlumhpfOZApsI+nMerYe3T74DCnB1vf7ZhgkZBjHVaA+iX2XIc7eIGZ7Jtc
SE28H8hXi3PyiJ2isZCdVwVgibjvloJz8TPeqrzlFCx7rfLnxbOHamE2+Webje1fDLgxcj6dtECN
qzrpGQ8qYLdjW3gtyxUKuXAqBTDT5BNFqOBqxxC9CDW+QCeN1t9gltDkZHo/i/On5nb8eCF324gD
7aTSnbkSKA4PtGvYOwJKxhMtIDnVqkmj1YTrgPr4XD67YtTlasWxGcAq0UtGwqplE5+EkK0QeHdg
CuvF0FExNwgECBWSa2cb9UuwZjzMZDoTdFz8wRCPPzJ49ZIytAS4D1rBkQv71GV/98NlMd025EIU
ArfP4ZOOiL9Tb7tvScZIu40IK53cG9BSS2zc4K+KC+t8QGrvhbsDR/yfQFvC7pL9H9Oeb5d9zZam
+MTmGDo+W1iPHOqX55svXsMh6NsIarHiXcP9ZplBAv9Qf647tmiXfivcJfVunbbjBjYq0vYXFVnE
44wrc95CFDjfABRppucGOsVc+cPsOdNvg3bXZTodn09cV3+IuiN2bDBBavgOY7NuQH9+YmwkfS1z
pazxIlh3UkB1LAEgJjxNCK1PILzSNEs3QneZJmr+IYIN2zIpu5C/1Y36grAjISXxnFmNHzeBsIsS
58C5CubenOQTwLS5itLMk1IjyohEzzUzqAL00dZZW8kRKvzvedSndnhwWFT2fKWyQWjTHOF6IGs6
yeXqIf0TPvygrpgJymFdRhCst2lLZf0cPstVuEfOo3CnSG79mBX52Q/mQdoeul8khqsQkkHyaOJS
ErYgBfg1a7lggVBHjGZpF3smys+CNt3EzGNdHis+Bi7HnNWP5i63NK6Ss+ervp6K+3zqveKzaZOE
IlXMzoOqIzj4ZCKoPx2NxxO1MG/JJ5x5eMuazDUT2Ml/C1r4n7aFrNrLFXOMyTxOlDq4HOl/HTno
p9yRfHlvJ76UShl2y39A3n60Z6eTW/lMSbkwu+50xhmIVdX8FovwmZnnwRr0i8UwfBRcsB+k+p+Q
us/MjdY6He1c9x1m3funQwfLtrfgO6XGrM6gV/R/kP1WZ3pcfsSCcg+7d7NaEeA+P2QMcibdNqu/
kgPseuJNiOoc77j1LAV+dlWffl+QUmd0aK30lJrmPjKF1U6ByaTpZRsdfUWcjL27fAFUO2QRC3ox
MsXGTipoZvKxQ6cJ1IDfal8DoJiTWY4BOcMHUbCcH91HmC2FvyEa17gZr71lrhP+he43EUat8RVj
jtUJM0Dku5tkoYTf4rAbdM7oZfWcXFuRulSAzqTIs4BopyTpgOrN85qt39WWUj7lMZZJJYVZwfUH
IROD5D3SSNjODBY6bAo3oRS/3/g0xKWCJgpI7AVoYhxlq6kC63iM9zS7PoLwIDbUZ6M6CiojVJgi
RwYGMmZCXWuPlAvtnVll7xmSIvfrhEnYopghFRsaMzWgDs0cB70bMzjlwrnF/6R1gftJodpdaAcv
o3YSneZZMDFJWFyNVU6cu0nsptP/Hc9HXctm/NXOly0Yjzk5a7YtRKEeTeAye/tQyV8vvfb9DQ+R
ijVH1sdNHnntbv6tC1vdAqeFzHp2vI6f9mcphF8v73NGjEjJwPac45onRJ2EHou0bpIRG6v/5W/w
aiUDGlT0qAN0cET0N0n5BTjRcxo++nfg5fhbFN+8oKWHyw2ymtC/jV+EopLN2bqkeHbBZnNSibPE
K2Wv/1oold3tEgbv3z5wbPIojVb76PXa2lbc7aO3VsiJ40FOA2i3s93lV9bEcWN0739ci1jzz6Fn
GonFXI5Fd62YCr6LQ0Ke3wMawxC3g+1/Gn0TckVitrfqwVFIufPtGW1yd+1VjVoASSiblZwD3yAI
IBmI7CIKvs3HMHZRnAwbzhXj6dfN1qEYKdlPUnpplzxa7DWh/udoWhWoTPgWAvJtm3qqDQctd5oq
YQFqo4k7SkxwAnizVhGa3jNUc/el4kX5dFXErImyBCSsb93LAvdqGCgb0tVleB2wuRkj8npvskvy
knoAT/QWSVlryHQnUexveqOAZVdIl1KsF/MJjbDdqq/FkOaRf4GBE2sl6aeP4GvLBAyKNUMxUlAm
ZscWFOjf/ookJQ1JIJlK5EfBZ4y2jHxcOuEATBvzrBkYcfABSHY66qIRTLveqfI8JJJlgvdeGMKh
6rr37WBdxExMRAW9xFFym1pDG6OtHB+iIUsCNmQ1CD9W3gxGgiYsI27HrKgOrAT7Gur5M2PyDsaw
RqOfWZumZgjuMWIJG9moGM5vCD5LXTgaZkUGSOtd9DoQ1DJXtg90/OM7EAIfukACYXwEIRbQ5d2u
fU6YKTw08HoyIsOFns6ztmg7uP6wDaTJuRhm9EYEb58jW0dLwhWufpk+wTnW72u+I5AUvmbV5icE
D+F9E0AMMjWy3jxcnQ8sijM0o0B/DU8XaJYzfKYJRvcqh1U0DEAXG4sXVqd3KO1DBlrPkhUsNWAn
LCJa6KSpI5yCJuigjNQkCuWrJSzZw7Xi5Fr9FmaJXcVuk5D+vc46udVzpE1b0VClVCcF34Zo46Rx
sNCWnPGMK8jYh4PsrhSfr/CuF8j7yAg4CbYaY4MiXG6wNK/g/Kj4Sx90+XUnppP6DbRzPg2VKei/
PyJl3HnqLXWySONxnsm+oPaGov8qKTaI7XSIBhEJv0DzHokqnc+zGa76l0WGfD9JgflQbuXEJtLn
EaEe69YL08rYRXQL23u9SSKfsQk9oxk2CcgGE0DXrn8HN+pTTkYe7siDI0CfYNTwwqcY+RuZIeK0
2XqKY0slPYjg23wOfLl8oURJ1LO2/4yOHc8PIY9yI9/ck1YECtfvvkem2pH8VDa6KmaixgN7EWz/
e7PHnjbQpoyo1xy7bDUzM8vWEP4MsO6A4QUWVZtkXd1Xi5Y+wOjqMwojQoIafNvT5kuNaqAScB89
K9um/rysJY5+T3uZMFbYVaVd9W/EBfH4KikIsCVgqj8NFWkgdqbl9zC6J6itgayRoQeK9Zb1oqU4
DAljqWg08aY0E2OJqY0aTYwZWPAlaCkc/TWhpisQWHPhoLIfIU4YWERLSC/dVucGd2fcDdS7hda4
dKBM3IdLMbGJuEr7EphBqTQhCmXz4HfBwkOQ1gsEThufiEcFOI4wGC84pqcdlImk2qZGROC1bw5i
gX8jXtmlYjoToMG78wIkps26ZtG/2Bh5dj/9+QM08Y+CzrCxJ2/+AmfPuXm76YqpuPhPITcGPkAz
reW1Q3IjNyaBg4DeFQioricpyCGwkiSKnD+FbjpwHWj8z2leqjSYcWy0jiBqx7L5WigHFIkJWnlY
z2tUE4ra3On76UKJAuj7f77sfV0HoubCfSyVytpXNyCzbfFK9/97N/uM3WzSt1Or51k94ULfvRx1
4k8d8bVl/K6lgX9kCsSpOWN+5kcVoqm2kiPHQraxWV20OGbQzGNzSpaGjrRDiQUyZxTcNCuAShK+
sgPrf7fg2wubGOMjMZFNSmkRAgl5w80Yktbv2thD34ImElFppPbQtbD5WCeZextcdXccqgiSLSBT
Rqgb6U8RsU4jekSU7ka7cbsald5O1P2htY9B5m0QLhk7UoHYk0FdLMPXeBFAoi5c3mu99lvqu8UL
epJULa8M3xQv4IObJuw/epj5wpa+bLYRN5AvRc/tfbnkLZYy0NtEz8shr0ifVOY+6i19Fd2TadRu
IRtkwOfHFapCsJYpqzAGy1wE2KnKm297dbGX/HfEkJTDF+orfiG+kMUiKBDNn6pJBDHLOko+jDDB
+9RLaE9aDz/zDetnWJ2KCVm6tuXrnyH9uonNK9vlQC+3ygdIX/Wo3b8Jy3vbHXyl0LyJiNvIbPTr
N+Zi9/hx2fPFfhOOjPmhZ91OwZt8LRCghTCqWQvCv9skWCoeUNmELzs+oK9rsWAivMLnXd8OrM5s
u77yBII7hPdUekQJf6VBbMgBghaeRaQyPeQBuq6zzAontsEVLDdpBv5ZUNaALCPQZfmK0hFQJzoY
fejbMKNdT8S0aXH9OqHY+fucX+ikYwbUr84Il0nLhfDHjPpkKU5E5ULP21bWt1bxHCedOatuxCTU
fbC+ar7aY0lmOYzp6VQ5GC5B5ewmzAtiSzpP2RykkZ2o+2RAhPhaFyoWkvyjI8QRUUw45+wKcf3X
853YjyAsT7zvXScfaSGOgsyhYHvRU6rGkPzyzOaIk/oYpBR7mOMEPiTemhJNKNcMhRzl+aJkPhMw
yYqXhnjFegK6YEZELmHue8TW4vJD7gJsgzMRBVWaQLiKfTfxmmIPLxx5mWghX4bL2nom4RlDAHU/
DVVCb4piI9Egl5AGCSEDoK4amHI07Q7uNjpht95UwWvzzBZzRgpVVO3muMLfYThTwtEm3K1QKNjD
9RnHn8imQWTOhCwnwJ9G70cZ48toTkudZmOuDYPneNYmWYHa2xp++WRrzF7v7wg94uliDiCGSWtJ
Kao/lTbWhX8FEy71lRyxaAsB8PpPvfkbhz+GGRcCN6wwBmYqF4u7VNb5RZR6jc6vI2jkHsi4wfq2
n6gcAUWNLMFOJ4zZh3SCxEWw8YOMlt/5uD4DGzdzjPPpXNC85KxPF3vIMnioK2ZZOB+c9PzmYXdz
xqlDHBQTpa0LT0wV5OA/hfak/EvmH7ungOby+BBK+svfEe7j5JJFzVFu8maAGTbxJchVr5QG91cU
OKRpITlcNhWHBTudVNcSu1VNlMq4NNa7gtUVAzNs/Xla5SKF+CQsFwHmWpmboiZtZuoMzkHeAjfT
CkW5GoTC9lzao6tFVO8MxiU58mvc3RJcGXos2OVQQkiEhm1EiXduZ0QfLJolZqX+YuWrvbNY2R07
yoUH7zAY/JHs/lr43uZ6XpExxlxnF7H++1bJjK7swpGBY5/faCGgymO8mr83OdL8xcgWidvaJOBv
AaErKtyv2Ky3lXjvfTB7pM7F9ScwMNzdvdGs+Cj5oVSTVcomzjc6qQUV84iGamiDQJwNq+HrC5zb
0JhU0M5M8vUyWSPsSAuAERK2DsWasN0T4AqECv9yY1WAk+RVDUX0w/e9tv6qVSTTrWjUX7GraZrf
2wIGdbkD/wcGULjdPVm74B7deytq9wMJu9x8a2KP7NsH4huFFCMp0AkNwLveth4yfkYwmoNP0mub
cbAk2fxyo+sLh/VWFSo3kk4WjT+MN/6LcG0biys9WMo6h8azuPMfpHF/4J7T8xedyKp+67HOeizC
eXmpVReXSynA0KJDipqdD+WxTdRm90zUlLk45onGYvUIOa5UcjBuNgNgrFgt+Gn/abpuILiVnjX2
SvwlrqtkKAcD+YqxPyzC2oIwXP/XmA4dbMQLebH4lTuAVrVE70YkJG7jg43x7qWGS08suAmUfPZ9
lQFyEexi/JTHXhoHAoYD4EkBZNTRyOJTa7AyHGq6LB9+L6hSFo8mxfnYIkSABIItVPNynScDUvy4
vLM5P+0bCZONCLNvZEl2h6pjexWjKFw546+ERzz9xEFirccQ7jScvTjaFbBaZUedADcmzxDLEVLR
+eje4ZFkMoMM0PA7sRTDumfMLS00A/XyrEGcMKIJt0KZd5pzMrck8DmaeK3WUE1l2Tis5FGlH+/0
oICrW0XZxHW+fDipT7LJF2QRtk2VZJK+A+LIV7cO6fZLCm9aHbDQ5SN/SPHf9lVzM/5DR9dRN7ke
QRrXjkiDmeZ7lj2138NoppnDTnP/kiKwC7JTB5YMLr5nIta+kXQDT13xTyGN+aVTYChHp3Gcl1Mt
aaCTreJos9gAa+uS3Vmpqsnfouk8RSj5MWvPx2eZOVvvXY2gqSk9LRGByA7NgvESDpSZxKsw2xlY
7u+j4SBcdL7ap0ldD8MH1UnTzVxLiIk9VY9OUazaf/G9XwPM/ePHGn/3Ep/hYFLkAhI6LzGbELG4
+0zJl4P7BsixV3AUvyVts2OqfEXUR4ZHC3c/qCrcsf5RLLeZTgi3jYdrYuzKmDbNNJxcYz/aOoTn
JITwNCQCKI9WEFhh7Ze61A19rZDHzvtafHI0peBCw/hU09uuSUwF47sQNOVrQ0Uks+2e27q2M1hY
c7r19PahPucRK9Ka9+sfWjUuV+Ka1sEqjdEJGq0j1fy5VaIp95OvGXDbDWaZQPmQoPlcRN7jW7Bb
1oVmr8XCpD8ahkT4ldbJhIAAu9RdtX5fmDBtXOzbEsu4S+NMY9adRKtkxgwzsOx8tpiLFvLDqXz5
Nd2PvUlYre3MLxKVhRTCYEP2on4vIE0umyaduMqdri8dAZlkxhpInsJ32icl5tCLtxhnrcy/rx/d
Yt6kJaytx3OGwBHioyvr0Wma0sHxrHg5cHgddI79j6eGdr0AWslOYJcmfwmsEiM5K1V1g/X9yAm0
Geo4ZSWODmH8yxB9bkanEGdkqmo3+ZfwJKXYd9EBQIEnulmrdr5Po4b8wxo2ZU0Uu4yOlLAADvu3
uNxw4zU/NezvHQ4i1fV4E9uSfaBZyUZAUL40EdlGAlZDQnTAreXPgKy8ti8cFQMTjQDsvRJIVWSx
nziGUptt4VQx2PeVcGJusS0b79yzLnFBzcZsreG7Lt4WXJaKEptxJC68JEZjn+ffkXHhUnpuU9eY
KdluR8Wo8P7OV5r9dvgA18qIfisWcVhHb5ZbLMA0zj6PwBCULwY5VDE1GZXGIcqO86kjn5CqtWOt
lT+hmdHhQNM+OGGQ2O+mHSRf45MWXBEHbYozg+ctAQmaU1uMVGT6EJm3x4EOmH7j1SANyHUZFVut
CWirN7PW1twMX9ntEwmq0/liyHfINyq4jyrAXs5W8dXYgcs4mEis72y2gZwGKMrkuRhR5ce5Kj2b
ggNcr5s5Y2yYEPfD6zLQLd9MOiW+LnLJdD3rriEPeToqea9MHNsQPjYoCxveiW51xBHZQUhPiKUr
6AljwMdg3C/gnmO8dso6zbeJzOINDnm5+ndzR+oWAfM0iXsHnnYHfoPXmwUe3RzHaIjae84Lvhsr
mHwEThPMRuMYPeRSK4S5Kois64p5TJi5St5mxsfTtZCmJ/RT+EB3G2Hh0zwDzlPhoPxGUMAMn3Hr
ZabCIceECIUSLAAHiUn0iUXDdvqKLac2rsNr+ppk2m0Qk++EQZ7XjFWxzDAdd5srYS1u8fsBJlZ1
yOEKU9vnw3biBJQBOuUmT9+fY0VDKG3/KZ23mY/IaKU5E4hsHUyZVuQG2S7RnEDnuLgPHX1PPypn
TPWQ2XbaNQhmPRbw68OGxgr8yLO2pGki/alC7qfpMeJV2LTpGdl8fL3d84h2V4Rfu6jdc84/2GTv
8WDdjWUCEKAZqJG/gwQn1jHxMd7ZQNtB/N1KdFgS194x62JW3uJueGlBs6e/q6UdGeJmVR2XF5i5
AGSRND1aPxBWrogJoY3AQAh7ehwMpA5K080DXx+vc5PWHuuEhNKPNKto8VMzE5+dhIfx0W6lOSXD
Y/2cFItihHBNv33NYBBbkCppNQNRLQIrBeEwFfft414FpANJfH/qel2TW++ghVR+kFA7P5lURl3B
R6cxCC/l2oCxM1hMCP1oEJ824oTe2flOg254xk+YZryj+/Sdmbh761vGwL+H0u17Lmq0WAO5FI+A
g1tCfxyTce6LBUL3LN2DUxG6t+m/FifJvOcMyVmR+H5hD/diJbKMM3cme56gR6+FuvGY3QSx8cfx
T8B14m8wgy0WmX1wBsqYrZ7D+G0kuuQAnda2qST90kgI5KcYWTfa83DnTb424+gO1BbVYaPA594E
n2c9u4wuw6Tvwqcrkjt/mDaR2hLWJAjBvK7e9+NY2Yn58O4xn+xes7uE1MsHqK3i2o178NtKGgNb
ylqB/7J9HtlckzJyz0CGRe+XIoU9dGZXlHux9SBdD14GWieIaJ9OcSSfLHspCDnUZgkBaeZo2NJH
MualJ+5tCZj3i6P0N9uthhuFc2JCyNRgPyEiFqYIWSAyhJyszFKogm4JB6cYlwFLXqsigbRkq4J+
sm+EmthHxojTV5c6VINswXdCUbzCBCbp0VxgW7liCqsncGCubXIBSRNmyk187G5HG4U1S+N+OZqN
kNSgszCAr4hujplZkU80owiD7jqedic1TJJt0l9PN+LXUvCFwiOwTlsYHWQykgK8MPEg5fpOOR/R
nS0z80w0xv3p2VjkN1deETzrjsayaMqi+7Wql6zZpiicgrcrgU7s6AvLwyGwovKVCvHHvV7Fuhn1
jV9tohK95CXCZ/+haR6pEnAFXnP7pama3Cnc9rg3qgVMcAIRvQFD7l5q3ilpsvmvbNn8+vEILs/U
cXp3ep1xR9PIFvpLfF5pw8rKtP+d9JkkfiCplcy4mstndhV6ed8Usz+eZ495q5PrtRWb66j2UbY2
loAmt1kQbgpVyeYiirvhabmFeDnMp/Pk8Lnl8ai4yNzE4mh98nUd0NNwUN7gZLbbTfkGnhxerwy8
4MiH7ONDGsbHf2/W9VXrPNiLK/kUO024Abhn9NigzwUNALkfnqgeqn5zfU9kd/jia6iyd3zFdxA9
cB83SC2YPWAi7aYWr5oWT8wQgipOnkZVQZP7h33LnDaK1K+Kv+lC8tudeZJQ6aHHbOshcScYuvWi
QY1oYOYuPvZudKl6OeN+tY4FaAFhvpQltzc5ToocUZKuNSxMjcElpkVgfau3XybQhY6J7O3vrKIB
Y8BlUNaltngnlu+4BTZi1kLvWtBpuvF39mHde3rdBv1WN5StbeeOPI0oduG9NdOBAWaff1hA+pTa
rJhMKzslpIspsX65ZDqAIKy0AijLGrQCpqAbp0tcwggvkendBXg2NraZFKJ+tIND47sEqgqrLLtk
NLmEeyfG61g54kAvQUwjN5eKHqFOaWHz8v2z5C6yn/gbhyxjWWcc08YDpTSE8UsILEveDCqpACfM
gP3pFkMP6O7pEP0oNhdbHDkhrQjCB8jFOKA8C5O2X2DPwHs0Cr6TafiHZC1IkxlCXvUpaoFhoRS8
8q71vXdLXz294kIC8NQjw7gC+UrNgVgn1byy6evr78OqRsDwTEa/kwmj3YusQi7UdQzZqnQhwHIt
8ab0CZwC0Hvz6G+/RR4sH8WqYaFGHwMSGrUZkyUsB6GjG1stw62PcX3J/C+ajMhO7rTljnS4ox4z
9UhvnDKAMn/4QFfsTsWzx5BkzwvsP/z/QYwrGf2Ipu/Q873BSotkUjHyaLMJFtIdHu+szp7j5uLI
RvqPEAeYE1bmGq3Gd37Qrqyaut+fWt9gEvgjuFSlrN4wnCh42Xitp56zL/gYROe7NpgkdXr3Ib1X
O97h094qey0KPZOzuMqPhgeQaLNqRRsA0LDqP7X5PmlBOkf/y7HirpRtARX/IK3JSwYog+GwvMZQ
PZJ3D2H9+J22mP46B5VDw+SaXxIVunCSpgt9oBTUt/liAWlKS5wuFEOxJfkCkGYGtyGFWKbYjWqf
jAisa+LJeZ0yrJW+uNcJW3r+pKAlMuiKWPkZfs//OrFcr7Q7kqlYOXRjYEuq13WRww3myJ6d/YCh
WygAI8S9K804LD6oPJDfArg+47nxtWh7emSefnKP/fLWbBFNJmge5WORZNrAqW9YCSP9jv7ajcsB
6tSymQFLQcoP1G8B3IkzW4XVc4U0MUbenuKaMvnzhFY2Tv90MBBzix1Zge3yuC8Dv3RuTbK8o6Vn
8xya1oO4rUPN/AxVIlmoFBPWiWcyocdKP6bnH+Q69g3GS3f2Bz4SgA9Kwcs5XGUMbQdguC2YWVi/
sUi0MeSsFPZL8ZYZAp0aRwzyKbXoHh/Cpiny9XrPWBpfb7zbnYALQeOYA0iyK7TZ0NYU3SFcTjJS
TWnzPAgBhAth4xNn4fB/Jhb+WcmEFj7ULBbi7iBO7XJCLAHWT3UQRCrZsHq3vqHsPQm8ZxDK4Ah1
gbuQ4fHBDmRy9S39Gg9BRx8Xt/Y47ya3j58KD+nXK1+GpGTt9A2PQ5Jct3U+zqG+b0qdxmM0kCAE
Q++Omy9x4Pt8y4xQoROdELzSrHtWdm1EFQOR707T3YUlfdFKM2oBXV77UyyfUO19a7ztX3oXTlS6
dvxZaCCgmOJvptddVnVsjfNyObVM3lufsv2dGjaIGVRXEhuswIgoPwI6JT+/XTiztqrGPIhQx9Tk
JHv834xlhQG5hwFUFcHeM789tn/33LojCt5YsScTNQu5MLwpRD5Gp9yTcTmLbzdfHmmB3ZAzwScz
M694gIZR8SPcElX2TDsmQ6Tfb+K49oXUwsQV6x9CS47NKlJQecIATVJoOKtq0et+b5J9WeHfmLBd
jszqfCHsuY5tFhCcfJHx6qw0s9/n+zSOon91Ev+OhM3iUcPWzaqLFUeL3GdzYgGaEEGdqY+Bqqu3
/xQdjfnyrxT7IyO6sXEbiubw+I1VVV1QYRpcWm3fq4PIMU/saIP9pzvLK8wuGT4r0sXfwjeVsVZm
PmxhTGQZQLETmb715KxXm5TuH+d8YX5BAlK/qs9ufCPA6iPcZ7kBR+QyWlrR5T6hSLhqLPsGfRte
JZuMSK3p2yk8KEm53mR5cQBBJC7SwEHrFQznXQOFiLJv7Bv1vqsCzfFCBOQxEw+tehihN6EZM+6B
/et5JwcybM/E3ic7xSIdhHLxHj8BZTAsaLrlHT0F0os5fpkXfWEbzQuqTL2XxJfA2zlV5wNX9wpV
43r3q0qh9Ug/1qwvwNKl5IsTmN3pg7Wer1kTotyIYhEcCYbRHh576IeuCf1rtmCumGcl3bMF69tD
2bW8omLQjAU9KsoWEsMgryzciLXakTlUKo+wT79TggUBYIbBcwhot4rcoFHCg9Cx8iuB7zJauH/U
qZR409JvWz3XBalpGsWUX9HuoYaCFP8R71JBFyDY0jMIHOQREhm3lwCwXLoYG6XN+ypkOPlB7mcS
lceaVJEj1QiAoOyyx4NuUsPbRppZvikSzWNRGjFpg4OOExOUOTlIh2LgV+MBWgPzZ3SQ+d0i0yA7
AdYVdOoFTQ1p2rSnEQIWLZvXqbP28G9ZSr7Mnvjn7G23dTa3OYpnnK75InUB6Wg7r4yEbQiAWpFv
t82h4l+3ZcX1u6duTUU2uFvdzZDjdmvXbyVo60MVXETepsAuZj5ObVYc0wt8akGHK9+lx+7ezhks
hjhzVKwBGAX8z2wxHgobWUtQpF08ESBj72fy+ZOq5YRMhRksegPCJWDviKwHh3unc84ohJjvy3bP
3qWg2qI/gCpNTa+HUTq8QKRcBFK8JQfWqqQWaNpcHpej89nLAbwlZT434dycoAiYkmPHL44dvCrp
HfDx6nFNyGnnWgekzuyQ4U6MBcLGKM3diq3eSEhhk6DsUd/Vg6qNP8Aio2SkGE68kVo03lPpLntT
VxyuYx1uSUdHvfonAFixUDC279UahRz+2gtWBnB52cIS46bHI6buPbsKrQy7lAuGrjhmPA5q3SRP
HN7jYnx63DSBEP/oT0ZKUkVoKuVIIej/HcQ9NyBHRNs+SWmUn5epGP/pAxATBLtr7uX31UwAs1rR
7B42FT8/G7TXrmXkFQcq3fQIXmHkQ+UnBixZLWb3wwXUT998amJzdIBqyI2q7ZthMT7ahN7GJfdQ
b2g46RVHYHMtQpE7vcizedB4VtRMx9mBye2bvqfWpjt7dL7AVUGSr0Sk2CRtDmnjU9ZL0cSUG0e3
4N3lFG8deKDZP6NLTLdSqlTGwB+anl/4OJ+HnZmb4sDt0PWnA/hLGZTGjSvf9mPKKzS8S3UWqcfL
nXB+0DBnaSBWQakiWMexgDfAhCXf0Kk8EPnoJmdfDghJIWRFXdb08cFm9EE1j51WTS3EwUD1SjCe
qUgCuNTqghvEhQxg5xIZ3zpwiW3p5WPGyzZ8PYdKNWnuDRGstwrxNjP+Fd5NSNRRz7pTVqbXgGvD
HONy9vpCKe/3DmPSv0Cv/LcHxRhTwdETqeZYfbyPC/1s0Y2t2rnAyhfGRqpQlWFFpCA989OfnHVv
fz21JK5Jfa5DADgGnyGcdu7dMxtGhgSWlN7JN17d2OF8Sl6xnRferdejz7/LqrB5PhRpezt6R0bC
Aoc9qRfdMLEAfCbMH+LHWDmRCbejCzVzlnl1dLcpRobPXyOywtQj5r6va5D2+cgl6vsWh0+IScDP
pa3ij6cBc7ZSIFMklsIgzS1edNVpHbmnkz1M5BKoId5G47Mbj4tQQ5gcHeir7xTTscIWPmB8Ha1q
C232GT1yRbJJOsk2OG6tqYjbgTcCqgaUVCJo1rAwRkXfQ+hNIrKkbZliiOP7WIxL+3kG7nkBnwBF
TDGiDIFMCQwMOVQS0NCNszWLZGH+trU0mrJoaNIfzC7Lcky4fkxJhlMFbKqUuMZShhPVTmu4jcUL
nOmwNJxVXG0NdX9Yk+YXvUvKQ6ES9vLXfK64BshQVawuXplf0XFX/KFuHk/72Hnlp0S6Jf+VL7vy
63aY0K1WLJjuxOBNLQMoF2aWwofVGVbRo4u/uXWuZHi6pvxCgd+TRCKjIoxSoGC6A4Dpi/gKlWRj
TOYONEW0cfrd6eWBbzyjVCmSDkAEYdUGyoGwcdPuYtp89efAWfyXkjzXzE+Q2K/Aziwi4L6gobgf
uBts23B85yMu5tJJYgnM7jyRC5D6R33XIabYIEcqS3q4s2Hrx4BkSWZWExjeBQfAyxOc6UsRfJMZ
mw4sHcA2QHz0+/T+iBBkLiJ/Z7yu8/2udaGTV8WoQ5MaO3+GHC93v2sEjf3yYSiO33kkY96YTZak
QYS6y8SRtWIGe/DikYM74xOy4vXgrjH6xO4sHIPafyDN/DN5j6gS/6P3T5TGEesIgQFyyOf7AOlr
ea2V5BWBtgaW0FuUZ9nuXZ++tkAgY4ClZmAxwY70KtJvhPLrtBvAA6mFAChEhKC7aUsOSj00t+Li
akr6hIFhdegau556ZnRrVp0jH4UVHxjAZ6eh+FcnnSKxlt3PKQS3qaTTSj+U1nwbDVLUALkoZ7ke
S7pr1r7596UiOEoxiSRa7nn/QMOERgG28TaGVZFbNnRzVZhuNED6CKUVngkMeKRbmMRqfFgZdsj1
zuCn0PAfofLucHc1fCTHmqRcLJO6ORi8t65qcDkUqMgaCGDbwDoYQ4B2ml2EGM2l9GO55bHrAPEl
PHg2fXBlO2OWc9kmtZg+7VsimAhl+53lZQgD8dA1gKrCDNQ0Lxd3+9aNc5BebRjQTf/6SIPf1S3L
qM7mZhgUy/dkURcp/4RTKEtUpwQLHDxdlIWgtHM6b58Dh9NH7zGMuJW2xLvVqJQoIn49383VGzI0
fcLQZHeZidnKNsj6+FfZWapBKyfJJuy8e5hkPsVW6s4Yy2nfIdMeYT9xH8QAs+/ttCJ+Jr86eJPr
+QKOlwX00AxV0VRVuXAEk64RCUjIb7XV4KRerg0FA5PQoBSWwIszwkPMQ73s4DmriJDmk/gRqCGC
bj2ApaST1JxyQgvQi9DKnvryQrYHcxeISe6ukIzjgbvGbg5W7Pyz2RKLpskvGJmUZ6/eZ9JY254N
FqoEnSsaykoByoo733FfZ0MRvWK8y+OyjZimJzgGAn27n7iPnas1ZMs6+utpMHs1gO1ykU4l+GUN
o4r4Rx7822hF7m1Ngtvaup7vxre8Fd0+ut9Hz38YpV4RkWOxwt3qufIecw8rrD+os5gky1w10dw1
K/cDyyOfDBvLUJBp0Mnt8MX6wla7v+Fjn580IAzQFnRG9GKvL0vRhtNfg2NvNd5KmSlT9yrrHUoS
uVTs0gVSIKtR3HjBgw9cyMiSoA3jjpIEzvOEWhQAn2kLpfeQVzwc9LIwoEzXdll/uzKgwlO/+d/z
woNLJQk5UWPzfP7Q3A5NlmP7fy5Jt2HGYHs6F5AnnbYCJPNNC9ZYi0clBpMtl+4WxcLqZRrbv90Z
HqWKAQHqshwerryj0JddDs5ztlq5arKqKr+bbghblEHozsClMMEFVG62KWVEM09UwdWiXkR+57my
rBX5GlhOaTfVHx5hclyr+hRnQ2a/S0bKkGevvJAwTBxFtSDbbII6Yra+EDdHg/+RrNF8WgK+WjHC
gIYPYy8AYZl+VvXSkKpuKrcB3K9VpYSXH0cEXP8eGFoXKB/Brr6iuhf92D9Wvd757AvG9Q/OLwD1
qEh58f84Ne0nlNov5fHU0+m+wKi5kURCnb30VjHG7YqJKtdL2o+3zoRg0t7bW0PSrxN4GETZ/t+5
BNswPoe1aTvXbTsJTywgI6zTeIsCR8HRMdDeKfVoyKBlzm2Ls+7PzbKVWB6ZBjz3rtuUkO2+DeF0
xVUn8MFuJ8gawP/yY15NpQpoPY6Pv5OQojqVG+AcgeArD2F2GApo2vk0qbYtcvrXfD8PnQ82zb8o
vSmykC3LvcSAXGWn9u8c5BXebyPF6yekZC9KonEd1P2p47b78fF3Q1ugnywP62FYgeJF6NeIC82W
pkQc80PqHtHzbQOewJyTVDqQGqgrOAS1f06oGbdkzceBSw6B/5mCfYzCEbfaruVwnu7YZP+StvfI
6e32X06j9gPtLscI0DH5yBBkyH/7z3276RW2EpZiwaxo4zuPRdgqmnul9wY3UYteVyTq/Jw+W+hC
rHJzrVxFy3d8y7dYQRKZ76y7OMSk3htqifJrQAV4m8/v/HVaGkAciTAuRddQcDlf1OJphHrEeijm
QokG9fo7iMyWDis+LdyC75VcsuxAPpj1opiLUermkjP2EzCIaADdx1N9OIdW/1SmlxfYO3hbh+fi
X6A/tvpvQ+UzQQLxo/tNGdkOsolz3W/F/ryMPShokcJaukT2QVOJCkiLrRvuyJg7SH9B47yUF8ob
wSG0acE0MUzx8MZ3SXX9+YEk1yzWOfIP4tXb38IyCnUK60uc685VmwTz25CsMhVvUXCGc9cAsW82
qsNILP2jno33eXBzQS4xjondHiCva4Y1eAexi1r2fRPQwxTmBQYdPiaZl2U8EXlMGwiVQgIBcrQv
wzzx6wJqdwN9JYWTeqTuHaOt+w0AjRdp3xUwcqwzTT7+Q01vpMhUGcSgFXxvVRK8l0iRdPhmLTZj
v/9eWCrzUOvBotLPABFXZHhF7A2vKXX5WMQQuYry9XIgKm4/lhld3vKkK40D+gBv6q6UwC4uMha6
p73S7QMeXl9RY55GraLCbeUDn1y7+/EYnfhRQzg8KZsqRAzrSt8kRtLCcJbNcohheGhTi5cv+bTv
2S93MSUflH8BeHKBO/MQk5yfHd9c2eKSW4cBC/si2P/3ogu1r254suo3pqoN4Y2v/3E6gMtDLLFY
GUK0B3yCMzuhUMpm/08x3rtVekHas8t5na9U1DPK1ZSr6rTjtqpubIRgfnIJWJpAKjGQpzKsCPfz
Xb/6uMLwZi+D6yt5Ec4PTEkFn1MgW3sksQny3Wk70L58OfBrEA+HlPEE63c6YD62EYIPb4FOWClG
VmhRCE8tnMyXXnj79n7CMJ2lbAf4tIQ5xvgkkISh5QlfV6rWwK2LZbz7/ngyTDteXFHXcaVS/byw
Ss2Th7gpmEJGX7GTSrMlEcuN69M5gfZ8OUKzKEyKIxx2j8DHF32UkzGXCXHvlSQ+kzVMJtqKVHMp
8nW0AuUBQ4KWmrLvtQE7YHsBWrYgB9xOVFfuuqKA5PC8siju7u4yXNqqdHX/8Zp0v7e/gW1Qyhwy
0rum738K0oGLYrWFmSSnSm5ko8Pt0l4rTfRFJ7Ge3AWzdk9rQJlYxZHC1WL+sHLGhHSnRkN1vAf+
RVmzmbETdmQH6XtgT9IhcqSaWGm6COQJaNBFf8OGhHrGju0aMQH3YkoVqLHhzodQd+dp52vvA7KD
NIPq4XcID91fDHko87e94hPbIQi6R/ImNW4pyKxWWZ+Xl/ntlQzES5SwgVydgejImB9yhykicQiZ
DOop/0WpH6w9LI608VnRMjC6e7YaT/DImAlOx8+2M67m89ObhmVG94eCm+U2YthE4rM4eUtop6vX
o0y4XIXjFGDJ2qmPAbPYFCXKMZRlZkJzxnWpzfS6veHpgFVHWLnhrjZ5xgYDURlRvVLRBHnLLmAD
VlnObDc8R1LyAYbC+lp9BX9Y2E9dmOlIS9VPzVAyet5JU5l8LUHd9ArZ3HaD62FHk7eipWYbn0VU
jrybmwV9xVKpLzFUJPrR1+SZ027CboGOKqyIujhHarfihgskZgAR7SHkEw86VYKXBrF3ML+KIFD8
KwyDKPcsEObKDw2LRxjGeNK/Cy5XR5PDGd9QhOpzevvnGhhEfezq4POc1ewkc9dvINYR5kNtpWHg
sStnc981VFFOxTX26aPSMmzfmLqLiCpdQvfKmdU8sE5c0MeMImVFchDDYPjT+20kp85fBY7ceIt4
v1shePtOzR2PqhV2px/OCGXB22BPmzCjbJNTmzyP35Yl+I2iu1Nb0uNmreCdMGcFzXzKzNs4Utv+
qENUuoZkelcFH80Cm6tOmmC7w+LMy2eiMD4tUE+N3XDxmLHhDDycm1wL78ldOtLd5uDzu+sqjPiN
7yRif2UT/Ku4A4hxssCZ9RGMjQGyyHeRJb4310c4iHEJHZauvW23Z27IZfKcvV4SXnaHbGqymw3n
UWFcsurwXAow7QkEK8ruSnB9wrrEIQzFbzARrWQaYrgBkVOJNyvRcEvn459q+TuFAR0p/TRy3eV5
qGMboIw4qc7FnnqGgOON6Go9xnh7ugeN/W/Dst7C8WAnIboRvGCOHcWito54kibQWZE0xvS18vAM
z0HJNw6S9OVmo6WqYH1TEn9z5CfqBzTZ2TkY/5pXtdPW+L0wl969PAdwTwfNCUWiMgVIzi8YzRT/
bLxUvmqcVSYZZlW+d8dye2x5RrRIY2iLO+WMEyB0ukSkV6BweGotph6CQ7FopztcxGR9cwxTOyA+
UvR+9K/lzq6IY5I0jGhW+mW2rKar57OnciIGgaIRwh32jD3j2LUJaw29vDpkan9cCJ6BeLlh/ZmO
PWAlwo+O78nLa/c8pccNVIT7g2ZKlxW60wE8me2vUpngXvPeCWRGwdGlHTJInKy/QFRYdMYu5dY5
iY2UZYXjwXk0xpf8mRCx+ubdiHSfpOP31Q4g8fzO/y2xHN+KPJ0dH3ZNzHw9PRmFhrM8WF1Zw+kr
oWQ0k4y7ZmXU8u/ya6z692Ukk+widpracf0WdXfmoayDBCF5qU2W+LRkv1tRCJHsUg+wrdX3nags
vUF5fK3Hqmw2QBWI+EyPsXGXuLc2A5tcW9F5Tv1ej/V8r8gZ4XpjsTHQ1SITnDhySHV4AZ7W2PeG
3QXJkq5WJuMb24du6kgK54o5lFwlGrJlChUfN8Jm7DyxPcvme/o1eh5esVX7pkxpi+S6QQ8sre45
J+CApyNCwKdaAwtuQkx0Xo5eO8ju2VCR2sFVRY4X3BUyXiDbcng8WVx6y+E7ArAYf6bDSzIliJBm
noZVOcDMnfEghG1gcK5XcpJYqKtupuKh8qLSZ0RC7RSpk7Cj0e6eE4XtvNbLAwN2vxfbPKhz0daU
DHgxVzQFziD/MWVEvpwB13cotvjdflDiQyj+JAajjIglhLAPgznxDRsZS95oce0xJLboYnXe9EXM
E3HqJIQpBSqjZujHoNIjgyWPGYimLbTgqq+zNxilg++HoQAhV0CIG3gXOnDJSGGIfq6W58Rluftl
kxQcPF4BoLOc8LFmH/CHUGrHJHpC4YF9tSGgcPZ/9YrSugtEEi8OdWecqnkV9hh5Q7vQgLiYjsLu
9NdkqqehB/UjxVZqd/l7SlxtVj3Doa8ETiLrKbu4dTEpKlT29gE1J8ElLjR4ay0JvqT0OGTKUqN5
Or84O58HyuXV6fxFNymQez75MJCjLqXUg1651gVZGpC/Ej6++U4zk6cCWG+y+67sYj9YuGNA45ip
+EKanAF2FBQqPn+QwTKGBA4pVwvD97ENtGP4bIq65euN2VJ0advH14yTOa4p49rornRyq8Hggw3q
hVt1iAoj34eu72uKuQi9ANWOJtflKUNu8ZKQ5ojYH/Ga6+r3Ynjmex6GjKXDApA+h0aeH0K6dQeH
snurTaJZhUZaWUTF4b7rhvzmz1t/QgZOMF0k147EaGdNlL/ybi+A1KHj+lkM9zhGa1XNJo+kSXA1
Qdd09SZFjQaWuHy/UOe8oe2hKEKMqTKZ0GoL2XX4MNvGOhbCSVWlLzUleFvOjqHt6NSubBkjyCk0
scOHhhw9I1/LsvDqyN0BWHpWkYdKPHW3EHjEMMwGut49AXYwIiqlXlGiCSh7Z4NukpIrGZZgyN5T
JsTd6FPfGF8Kb/6LJcQG3uVMEk+4q5/NfsklXlyp1bOTDEd/DLfjESqRGrHIK4Z70iwBB/40Qpm5
50lZBaeWL1eu2ZnAK2qW5i4MFx+wRZJ+Ud4DVJyCA6SAzJTJVuRr5GYCWkgaMMXgB93S+wSYEe3b
QyBWWfTOWfk4XIX3lzennVXUB8AWj1eqUjHydX+GVYQJk85Yk6cJ7yIEPC/ThExCkAyWxGeIYUtw
eaOui1ybsWTSXb5dtF0ymYBwp4fAZ5tzAZG+LpBYrUyRigHLdbVaIXNW/Ze/mhZCrJ4lW+Xs/jc4
VDo8pKv5LfrruyLsgFZyWByAK56KBAC7VKT67H9zZQKhpQGpdl0I0IoguqlC5egDtaZcpMjFyoQ/
S0AiHfG4PG4t7WgKGgM91QLUklCp9Hm1Gi7c2HG/vOne8JQnsfP240X80e2wHIS3o/9HgIBMEmsm
CYrLT8iyPzlAIOHpHT7dHuNODFeEIHeZWCVHYlRDW3EjIC6dGsJ+rlJbVXxHrr5cL7Uc41+kcr1d
t1H+VmfMTeNbQvL+pfwgrrZgkbOzMYmv7wrA5QZCivYuQkukPvlchSj+AmgmYV7lu7FM2PZuB83l
bDcAbbMYlxqPt7gQTpX3jxBOYeYnY172kCxo1yi4YdlzYK3WkpypqsjfJusVW7iqMCK/eDKCfh5I
21amLCUUiDDBs6PfOlWOufRdeK2wQJz/H4G+A6vv11/SeAjZt7uk81B66Ltt4P7lciRZTVyXs0N7
a9Y00RDH7nXvBYX0q9b+eBbfTz7yw6EMJB121A4TP7xWvxsBf4hZFPXd69htqYgEObgOrNDLkOiy
PtYiq8hMnjaIC4AMvewGDMKP3z56+ofT/EQGvrFzy0Adwohq488vPIBOFJPrJho0jllZaOQCYRWR
3cGF5oqfg2RWr1c4giT0lq7cjDZOPQi2n0R/qSrncFwMBCYoaVi+34AdiZMoxLca1JaxF/mZ2EyE
pl/htZWsN5vbWaKI1rya7H0326de6aX3OtEk9n/rTKY+BxZUSrbjjQ6SLYYMB5Kw9hE1PlaTrgw7
9ZrV67ukoWPchNzohjxtlmDEFAnM2aSRcgUx10tGoYWnD8wXNe/Mx3/Tp7k6HG1OxS7ImJHV9jph
yZPe7weLTd/HuAw1PFEHQbWzs7vPjS8y2uq5mv9ve9dgbf/T51gEteDpIZZvZkhzcmC4wDj4rwAF
EoxOGOVXLB3tyhjmy/9a1RBcBSxB6E6Xul+1y1n8c9pLKyP277GLzoNOqwr7a3Cq/AvkIiptxLW5
2IU8e7dVVxpmiNox7PXOTn65UdqQt8HRq5TC4DXxfVaannRwsNMx30E+sb7psBbjjbQs9oQQEcbF
rLbMf+caysss+AiA3DEW7pLZXxprLU50Z1QhoFC3CyymUuAZBceLhk8bzdeNm+4/4TLCgkkjc68+
EOd88tdttovTTHisP/SCOqEZyvR4az0EerRz2W/NyhKi32srXfPKtXAw7p5tEfZORm/NCRR2G9U4
raCKfSXvvgZgDwO3xR5eTqzyQj9z82PKaRBfjIhhVQWL9w/x2JDYFrCiOCWXAQuFr7hyV20QCWg8
0LwF+FtsoFmyEbUPXVr120lz9KbPCY2qF/zOboGStxQqMGK6LlO7x411VTCeU2qWh7pmzG2X0bAa
sfru64AjQDaWVqcxfynTJlPVPbXUurqGt6K2r2u6jDu3P2uLSGowC9YJAmArwmaKenxSJmKP6LLu
1PLhZoySZTlSVW9KLlCcx/CJiXZQV7b91khTho6Q/+i7dzvX+bjPuDczH/1u+GJ1KtF9xbclZPwS
ElwTy7ux/jDItDQedCuAi4QTnZGZYs/NY6cH3xq7fL8Oky1HlbSG9oDpFXMXcWyUkrbIBQc7w7H7
Hcwv2toNplA+GHE4J/zjEQV/NfdZN6ftjYiL3jbKn/sHvYAo0y2sGFEKLp18CsTH66ZUkaH93JVt
BoPg9A0q8acWt+31ws2mhFdMWIzvTPiHIfVkeDWeH+eK1mTg9B8r+ZYev9bfyt/FkPWQEFP+hLIB
0POpmbuhL00fTrkF27erA9qIXb7uU3IOGMrk2L3tbrmBTZNfgxcM71dRX2QENGbhmMGliTHXhuWq
MNGH9RcKJX/zLKBAWtZ2cJPXMYBNM9jaMYnm9FElkWTKwJjAHfwbcYNqNzZwT3LK9mSQCOCdfR0M
15zvLXlQNc5PHgO3iRMxCTfk02oW3Tz73DmTeyKTzjfEOsweGhNptOdS/uCFggnFAXhUvnLqKlZs
V74LJu7kH8sqDLtsoZHJ1AhDZz9LIJgrkN6lmGkKERDeetKtqCQ2Km7D14kWHvYWZJm1M1T9cCWX
lqOBACqlCeed5l7EPNGLq5ld8qRam+h3JurERKIKKPa1f5ciRjZedz6CqNY0dMFw/TkwdWQNxLl4
uB8S65pvDdzzWPPKIZihdcZEZGppMTGMDWJq3kPQfQ2K1Uocw6xRp+XXcsB8rVVNjDS+UQx6TCUS
9rtAvxOb6WKVOpNcVKpwPb0INC7Kw5e5OfaSkiZJpX/xLVDLNz+7FQ4hHQ4ztLLuY2JQDLFeTOUo
fkY3//qjCYzt5rz6yvMSootE89utkBDm96YSW2+3n6RigqNgrC6+FbPlXNFc47Dcm9gZIXhE8Pug
HKgmB+8OOxCHRji880xp3LyEWVat81iP1iw/iaaj/VJkN6t4WQ1B2Z5Ub1neUx8kU8zGLIAp3zBs
Oxm0Iy/qeO3ZsFEG/yhN2mUu5rJE8ceWz5BWx4/+nJIUdz+gPFMHfV4H7cd/goLz+p7VpgCaA03D
A85wSVAUpoIoPrq+E+94nU083v156VajgxW3iAqMIuUNnG+gy9F/ogzQbWPt0yY9+zqyAHJWE0WJ
nxK+Qpp0vnj2owcMreOHFzDxQ0jFEE6/VuZIygVVJ7+Kh31rfalpc4fmvajXsZNmv6x6g+lZ/agw
hBAl0YuTA7xyTwhkh2/DPzQAJoY7qFHl0Z2uY1VImFBk3/mACnLJ+Dqp2CgTBGxzjL0wnsiHr14k
dyz3AH0b8acjYM2vt08XNnrRMo7RnaRsRaqCx42JtbL4grl6MxL+TqKs6oXWulx2pf78JbjdGrsU
w1yHX7+J6qwppI8/EbUuUucIPDLsxSQA/3dDxBs7cB8TKQ5vBbHtuxKQhI0KdwccD0NKHvfNCjfz
NNDSbt9wdMmB7TXNGioB/fkR5uSoTx3Uh0kVubCG9te16jSWxYSE7Lc4D2M211cQ/DOL8ZJYiHpI
CxefZKIGcU9MaNk9KUXr5Q0ckMuaFLNJPIJe93s7PnhUwXe+qCi+WQCbFtdxiVNzoUpdMCvHoew0
ekLdlvE7TTXt/2qqp/zVyAVr1YW0D5d+m3UMFg3R9tPDS/wPNwzyWvtGK8JatIHg9RawhUlLijMb
RDW2+5mB37ZzCw4lJdb90p8F60slaHNgnA4tgLNaRNnkZ4laOVEK3h1Sp/Ecbaq43bCG4o9yOPv6
cZ7anac8rX9Ah7Qm53y27Xe55P5q/ETU4iDo96Yk6auEuEoH+btrm/eT0SbhRwxJ8uTnENnGnYji
kPb9QC/8t1psjdci9H7JoZ4BQG9Mxn+iG2iu3uOuwxpwBM/lDn1xDEy9GwgdS3TtfygMCtGqmoCt
Z7jJneNBd4esLnUVFc0p/AMXQdELK0P480gsM2P8KXbOQl+d3f709hydDiSb6P6yNZ/eeoyCxA8t
9eXK6wcuzQq/HFllYXI8i8WXk5KwlkXPiKce94pGEWzMvIpgX2tjm6u9gWN6ymOhoMNvwNXVlJav
bgWociIfFXJer+i4ana/hE02LZEvFKfidfA4MnEZNmWJraTToIwqP6d1IdyqXwU9BQ0au0QI5RWC
TnitP7/xVCnlFjsmZF8+GB8uVQmxlroWdzdbku9Jwc3OlO+eoxHFUpQPGyQl8rhBS95NU6QjMPdO
X7p8GgtNcmn17lkT9GHq+/F2EPWfvA1aOtNg63O8bcKc7qJ/D66GRo1l/ezifdpZ2w4C21B7PFZY
NFNCyof1KToGCkAofQ5+HfhW6/FuHwa+JWuymqAaTS26tWZ2+bichto7oTm/34hwwJcJGAb82oo3
7sEsG/IdYM9/gRD9bFTAj/TV4QScq2YGynTIJXSLnJ/QoPe3tpIcvFmlG+su8aphbOcgPHxGHrjS
06DxQozXNHlAmw2ORx4KyqZaU3RKaiyXCve2/kO3mv+al8DGkzFi2M6h1bW9g7Xna56LodhupzJw
9MKRq7yOAsOWKSbydams30yxrO3TifZ/KTqIc+KVRL/5vHljrzNFHP2N/aMBHFBKdAlwjK+kJUbE
Qywy+JBG/Dxk+ASfPAsAWTwoYnvxvqODMqGCI3y2D0SQ1L/evRpIQzPrGYtWpDg4rOFVnPWnYbpB
4UIrYXGTgD28jSLu0HwAyrlqWJb8NKWTtqHTLxP0nnqkf8oiSA6KINaWtJtRH9wFrNyMN7KqiEUy
yw0QERgNjdCM6cc8JYp3myY8VG2lxpu3n5NQMjI4y/PPcaEQVPDAKf9J+L2vxgd/K6DzT3Y6wW4Q
ZIA/XD146BvKK3okZPsWnE2REU9PZumhdU6BkClzQq6k8ZWycQS7vj62d55NmzOO1Zj50VcZ4/KB
LbDsVhfIsSIizaVf9Pxr9Pl0ROjXmXktOH3IKMR6LvJNYQzgim5WF/ZhuBbImcBm5H7nXRKKZ94V
S+essqqGvGJ2Mb1LyWyzhjEVOxSiDC1+HYNsTDQL1q06RETfXWEJUnGt39DVQbA1ye6p/YvU+Gom
OA4Cr18Ogd3HnmO94NONPvHZCWnWo9sH2G2EBYFjICagvTkmBWmKUKSa/ZhEBiXlDC4wQV57E30Z
D3Q3h8t+B33FDRjoOZ9lRrhRaEMGMx2Jtz+soajapREA8ERxpFryaDDYLo3wvemIP1CuuzWIDQ5B
KH43++i1G2xp4lMve4jZ4RluP6HiPWus+ZTM3tz3MNE42/zx6BWDt1GL3jvcXGhW0vFJAob1zJVW
l49scGIY+l7ns7Its+4RY2An+4a1ebZFnM26jRtdnr1tDlpquoLwgNegJzkxlmChF89WYT107fut
HH6wSP7s8JrfhJiznISlPOfzk9kTC1Izbo3XOQV5hflTzeEjW8gnTl8AaCbXiGz0rLQEAuaGxYxa
sngUUeWSW2s4ObYMfcRgubYReniejgprSP73vgKPa/QG3DK/P7kSj03nNgvsp21pWhUkIf+OeReB
MeVefFPsGGh6/kM3X53y76vMimrIWx3d/vafi8HaSLVFq7XvhgnR28cJPhmJyiwpeTauN6s77cgz
upIpXNx7jQnTsYgObqBRFS9P/ggW+gvJi49cgBSo1LL6fJ+38XKMTguF3xr5FVf8YIe4V1K2qz9o
SQ+wve/5Lje/L93LwSR/ON6Yu2J36WIjiZ7KGK/qNihbtXt/TuV8Wat3jqZWGkh1v2DxtGrjQtcE
jnhl/RixYxLSw4KRAku3D9iGWUqObLa0+ChZQ3b2u+RANJHQluSu5E4FTnU9GYnCuFALEsBnSPai
4mZi6Be7SHwcB1b+GCfwo73PRETBTRFu3pB2QS8ap3aJrfmSlD9M3Er3qGcjRSJ6GqG7yNnXkroN
pVVyUaizvwLMlJLGhCobWhYIHWuoLjF6+/cblpp1FNmEQnlohdjSsgZ8rJTJ8oBmw/1hcXpi4rpt
6QhZc/gMu45TwnovtmnjIoHl5MRK9AwxQtLG52nD5eEptmOZ83DncJ9NzVw7JfTIqvAnmovYTF8Z
v9jwAMMV3Arsdo+zoLXP+Il5GwoasgeMpipbsodZQrZ2WCcPMms9Oi9diqvoy2sWdTr7ZYdkZsdT
ubwF1sOUf6ZksOVJznZFBJtlby3sgXgRy4TsbT9tx4VxdXa9eNSvxpFL8bzSnS5IgIcxNOcMGG6c
DzBetT/xHhI1V9/WGbk3Zsd1jWLI47/F6dmq3fzEmB4Ku4Vy9N8s6oBdjU49vbT4FRwg+JCY7Y/U
PKkRlTOT9GqxzhrNHtlyWEF20P8lALs+CejsuWHociLJRYVn4b0kq2QAtlfcdNeFNIyYSF0sMUHP
+XZPtTqMYw0QvGv6ahH5P3XxAIpHGTgjr/5/Go713BAwr3zbq/ni0iO5kzJBiwGGEG/mnLmr1hsV
mCfL+E1L/Lj7ph27YJ6lwstVCgXdWuHT3twsGntRcRC9qBzxQJl9OyvFi3ay33CKUgtP+kUAKPms
HknWR0ugt/tp82rx/LUKICCi4fKZo/jzP+Xw/G1IWl0ENAp5B2Qaf9KaRoGMPlhab14b0d6VMzzI
AP/AWErDAcUC9Ke5385DCE438x4OYnnnb6ZdXJBbJLubFTAIkBGEXO1hU1bMJXh1YbMk+ahHUYW+
v+YX3mrUcvuZogAw6XXKVYW8d0b1f+Hm9/qxyZkCWLADtTwr9524AArnSb51rCz4SsHEU3qVKnxX
xkI+z9pDdWxrRVRXp7vrkjxCKANtX395Na8/uCYL6KDo/dgpbmJzN7Po0+SaVAgNeiUGSSRTDUsl
I2Wj0bDl0Xf2dOX8JkdTn44dAAnQJ5wv5XTUIPa+mFerybQHDKMIyZkpUp6ltfaVNDTLsHYKtnbV
mzu4WHAVLU9DIoNh/ngGnO/DOm3qC87NKAR7314me6X73DZUP7hHrxRjFAhLgQRagkE9JD2p04dN
lZC7TNhL7j/IjVydKODJEais3D9AzfClB3k093I03xwPAF0YsAq3Ozsihyj25fNS0khySnf+Yu6l
ASAwQDgVGD5ooD9nZadu6DW56QdroQUiHW3Yiorj7GeH+etjBxP4l+4neBRxSV2DGg8z/Z1vi4zS
CgeZHN79LX4ugAS+Kgzq1YVl0cgFlNqgrfQj2Kd8USSNP6nR+qsQjVyceAgRseHR5/waq8qpjZFm
9xYO51QWc4Z2knuLY9R0rnraBTBcBDKeErAsA5yHbU/gYnhIcPhbnPCf6jpkw9RWAVkZXEmVrYKl
Pwd4y90ZXsOBZt9i5i2XDb1RShl5eV7OQoszY3nPi96aCRhWozK3JznC4MOdzR3sl/PSa8zUPm/3
1zrC74uvCi1Y/FP4eNgpYnzXxyKoBoeu/WONoEOT8TcxOXQPE3wdDiUii9GWQ9rKD0MEohPVuKGu
wajQdjIZMKAJdq7KokatZWL9JDqbYAwiToGWMKByoyh1hLfp36oMQDvdKZ7QXGF8EWD00FxY401X
R3omOr70MoOnQsUqpmicbzIQxrJ8gYarMuBP3DaTPhU/3XyR8B/xNve3bsaZQZCr4LG0zYAetY4S
Wk4mu5FzIwVZY9YWXaXHzAHjDH/QBFsL+P4JHb1B62lPr4eIf3JbxXVMQNv1GUdi3U+1qxPW5soU
6JkgCXMNdvq7aMOTCAyYP3a/L2fgLq3VrP0YyMXMYx+l74/7bVjEaYhU1f8RdoE9/GsJzJNWg/ok
TFnoJBf6Fh+256+5fGOllLKay5e4kk3Mlw+2KlA66pP5BOf5fB+3+rO4hzyBgsJ1Hgrxg+PHyukJ
1/Ii9liz9xBb7Ii7jmLvBRCV/LI4CX7wRQdeA8Ba2j2oO7rN4t6WP0Z5AGGq/8mjSbtuAyL+/NrS
BgYNTTS9ZFn9ChFhBRv8Bi9sfxaFH38LRhSNcRJequgt7ci0bjYHrwUK0OnWGiBJAWSVMFWwoflo
w7DkQsgK9NOBYmxQOobMbFba/2pvGwjIXRATtd7k2RpDSrBtTFi67tuE7h5bXsN1SFEgoWeJpyH1
UdTf8yzT7Li8H1fw+AsoZo5S8eWc15KXpaqVBDIpnM9fRcKdhpuJ5SE1V/H+nYSNCIhwYouxQ6a9
a//jduPWKWRNRIjAGdeUIIsj03v025jr32QMqV/f+Sj3Q8Bk2EPi0oOMhdOB3J+l7qYj7RtzdKNP
qA3vS07r0R/GwFFcyVimolYJSnHZazl8NEN12A+TkPup9K8UE7qW8dW6+QsY0RbKiVIDOnbk9E9j
UqQvEXxZH4ZRZdFXpKvuVDxCmRNOnKMHiJDuLprt+pyzHRHhc8JjAG8LW4R/z/Jn6qJe9DdlHa1O
Nc2sU7/6k/hG8BgnOqeIogPbOkvb42hNVgl3YaF5lDG3nnEIMISYb2VFLJeYBrr8o6ekbB1iszYA
KJGoTErSbYoQq34zQW5IRAZ1kI5xX4t6xaSmCmZR0sXjtJQEeJBV1NUW7QsY3ZntYqmyn0FYUzW8
gPHuF9E2hlKqIHlZHEr50Mo1b83O76TUmuTwSmecRsWw10XCZ2gDyUJJZS3uuyPmffzQr4SgG1j6
g2NyB/BJ8gIH3e0aXD3RSvZwLtyYUaisXR2J8YySFCCDfnniYdDza64mIo0iITFG8U5XoBFjf37F
nQQir1lCr2ko+fihHGvX+tyDgJzZbvVn98p3nJRnHoMXt6w9A8IMww6pI/yA5mrIaQfL6/W8VFO4
mZphLIkQmFoontgfueQJkWjKKZxC143mF/PZrPNj8cleEUUAxVGy/00nQ9N2SQ/qn/6wy8327686
jEGOD1NGdXxtuPMzlUWjt0zP9NP1HyE5pI4gNVmFHS+/1dQ6OUCeu91+7dHUeHaiaa1ucwBk5Y/G
8aPnXYgcbmfyj1S4Io1Yxj/zqO72kY4a9x8SOVEn+YINjiMti4nvVqnqlMMARHFCsAE2uggnW+ZK
OfrCE8Udl2Ha7luzLXjpKoUL/bPMCzKYc5WQPU/vhFwL869VHo7QFti4mTuxxPyLXdh2Cni6bcm5
AyugWaFq9OOiYODy/dtTiIqGTznEg6cZ7LtMa1zWF9QXCQeg9Ep1ryC+7FpUKQAF/pO4OFqh3Lb2
okBFqZijDQopoqYOz7TdWwe6sTn4Pk6KcRAeczBxXDrSfDshEdOlFr2wjCqnw8V8tYydefMpCPg7
YppBh4RvKf4BN/jJlOmuPmddNholdgoIbyZfn8rA6ypZSeRIIb4N7WciH7uA0r1dfna6wda4uDpr
iiJgJpg77YdXkxvau5CPS3O+PemJoIFe+zUdwFR/cFQVyAEnFQqrCgbbNbvSrD9+DxUVsMTMiU8l
hjuP0kNxmjJcDW6/7JqMNaqxognCpwSue5pkgeiFWTLP9Ub7VbijQA1FqL5RxXKznQRqKUhbfYbb
HVqfhDpKtoNj7Wu7+J0HoAVYHJ0BJE4hpXnMGkW2su+Ig0RVgISl3oDcy0aA5fcfY52SnSIY76O5
YgQSTHWkvQc+r+zrcAJUxfA5lDtaimweSZT24FUijPNoByqrAYER0i8W0LFOHA9QDZkbNiZK9jQk
80uVIHXNlHeS0lnGkvavXiPJEN/lEzhNXUmRQkqII2gBx0hS4hlqhNVjrRsSDtXkKAiURhRvdl9Q
S27zQu6vG/fDLgQvNbe5Hb3qIE2Cw/f5ABqVVTVfus9/ndazRidES3h0nP4kNzySPcARLjIKHgT5
9cS8pSBAhsKIbQ+FXwsGf2ktPsseJqAx0oxt6KbbDuNnST6s0CR1z88ssMeJF2oZ1ASF/+1OIBGa
p4jdeddqsfGCCTTCToohLWI57woXLoVlLSN7VzTvLxINO49RwdX3idh/ecIz313lDtQHMXPEx8wb
KpCUs73hyaB+xc0ep/0CghJCsImw0Jti0LjTjFGCGgk0WQz1M94KymJrkmsNmXNlgcZHk1lqrS6G
qLWqMY+/inLGdYZyEGF1vtiDtp8jq7BqBDAPz8c8Xlb9ZacgXRGKI4K2VukunDw2V1uGGeqsPu5E
xvx7vsBTZ8EDKZsR7Qn98l34fUsPjCPuBmTcQXHcjpPYoCHX6XOvqZn6Sy3nWibgMYkjoxSwPmmZ
tQsdouVW97BwRjBYyLFq8cYj+T+H8hBIQbDW1JKPLlxrD2sxCOgpBJqtzPZNzaiGXbl2gi3ruFVj
dVQbo3oUYD/GouiZcGImgO7GmPIs25+xV9LkoZoXKCukzDX4zeX8bxtdJ4BjxiF8+F3lAt5/Q9QK
7SvVAWf6yjGJLMF5KSFdO12m1sfJ0P+Qu4/tHRTJGHJSCw3u8H8kzBS4gByBu+PTtH+1y7axSVcZ
giqYT21kzSILsjErsGNCzczkiB8XRNnoWiInsAcxy893kjeIYGaA9xeJpYMjCcc7tCDBIkqNb4HS
4XBekUoflSrAsDBZSmOY+TxbKXCB0lxCZ4HH/NRLWtmx11RfFrvFSsgzBUPNbgvPyfw7+ki4yQpb
khZOVpQJwvnvQ07jRz6b6wPIGBfJ4wdaKbQzkz+spQtt4tY1SSXPCV5wkBOfaGWcclnW47ToL6Bb
f8ACa7fFJep1VpMxA8ucX18uM0cb5KqOpirncBzV2jrX3coblDay+R2PAjIt36mo1wwObStTxif8
gsUWlMOn/LZblD0HFMXy1xaQ+masUkmbr7N8ZP/zlwx4SqnDNSHQH5cgdsk1bVN1oaScpLJfjwvH
DH2WDevXOTC5lPa1zD/hMnuf7TJ7HDgEpfo6aeoHkDvrFVy0MQfOFyIlMeeGRIpexp6wTjvRxjlN
pqn+ZrHsieCucPJW8dcYtHA37RLZLEbYKC0k1Yx0dS08JdEu0FItiBnkKbV0skZKMjmHdJxKGFvB
6TYqIAlhAT6KyqY6lrRAJEBEsrkrRh4WsdZ51DuypDfyEiR0LkCIe57FiptCXwu6jXEst+QecUVT
qGBAbeOaAoHyOqLqhL4cYTqECzr9v2lZhFu/JqEmEQ1uwSGLhIWAVq7bkAZeXfS2RXAfijEsa9K4
b+3a7Ey8ppo4wN7vefoo19JuqiKtiP5iRpSYuGbCY5Xu8nn3/vAPsX4J3YMEBmE67NDZn9zbv1/G
oXChertuN02I5h1UDWX5UivZiJ2eGq1OpEUJJY9VdrFF0QNNZLVGPWi8vdnNi5BDzqOw5Wm80PlP
3K2cOnqKRAutOCXRqjZ1N+TRKwva44rjWGLrzylC4gGELb0D70+GRRHHgWc5hvfJ2l4tJIy8dfxG
gPcouPM8AdSkqoL12QJawN8u92/1PiT6rTF9wuU7C6aNcZQwHo4OkK2xl0Wo6Y+NU0VsATEj3ZVU
SW8T8JRT7z03iNlQ+w5riPLWZf9hAbiCg841xQiVwJvfX8YjsYctniLm9iEQ0He6/fh5cgjoyVpr
2VuwjlTceX2XVgpzTEQS9JsqSR7pUKAfm9E3cuGD6QG1mNBKFcJvWt2N1EcQmJUPfHcJcr9szB/q
q93E08gEcu1agSlm+fF4PvO6KP0tJkQqQxCZtKMX1OLi0GVu19VeWAowyvazBmBaonmeCDeagHG3
ywATj9pCjeQOqCBBKvPHmRNSoe+/+pTVUPwlqNSrLibL1e6P3I3wep1SIZv0YKIyxMza53WEJGTk
9w/QYXAB/hmHutls7b82nVnu/oHG3NYWw2mox0JvORiTR3WnpzIq8av665wuOgrQU51vyC4iOxPz
4RqbH39ncP+IlPNcRfSB+uObf6oYY3Lth5oI4CWT/csziPzTpppgdOBpmBrv3DJj66DX5JjsWrGP
l4RWbFwyeIGGu1iRonewkzYzmNY58Wh9EepMsAyrmpdVUfPIMoK/7cAzzcw35dqfE7BAcZVfoXuj
P8XobhwfKgu6nAulzbed4MiJt2mHeLJkwiWVl6WDOggAu88RmzGFNxKfoXPV6+c6o/hEGrIQv6HP
jTQqdZXK9VuVkL9/q/4MYfuqEPbtHX+//i/1KhEeelWUIm/FpfnMOlUDapwsL1CXXs+NcIzjPEDL
Y0WqGIVwJ6TMxyloBhuOaTQgR3EUzsJpIme4HVYsR2Zk0ua6PxsAZKu1uiXAVwaMIaSXZSmi82yc
dEHFxwAa2eyOFs0gu6hBKLgb97cS2s08wLkQH7o0rrt83zGZN4OabHJRTo7YKXowWy0liL+/cmz6
R9QOO81+reqkFPkRDdStmDVPvK3+Gidllje/65+BAHB17B/BHlmHiAbrEwV0B6agAccZgkbD6Y1s
Hiw4JYZq3je3vv3fNvwjQWiAzmx6KPqJfGKXpi9ioMiuxbUPmcGLrlxQA0teDdXDhgqbEeQCCYQU
fbaH4I7JtgaCVFZ61pRSi/5io+VZgzJ+quZIGQ88QOGqUOwhYuXXtoPcSo69xE9DWyPPDhWTUrEd
C9toX6zuvPWLp0Ush67U0YE3h9Opt/+nwOkPkbFC47hBhxByuca/9Nl9FvZIP9ZTG79Fg1/OyDua
TjvRKhXeHwqReAe1CRf4FfxiTaMn8BAjJ4jlVu/zgkFpNbK0tioJVPVRSnM/8bX0jG8Y2PtElpoT
//IGn3TGc2fNdJZtGuwYh7nY78rq5E7y5p0k3A1f/HbktNcFwqJuiKxdied47iCN395Jb+yqfcwc
R/0EeM/xWPfRmmDgD9TM6/YeJhiXt41db9j7N3CN0QqugXKNSC5i+t5JG61kjnLrg735ct4jVEVo
6J1HLCPdAT+8c8bcTy1SsJ0BSPc8ED6NeOgi0Ve3Q4dopw1SQLGGieA2TrpfBjI1LWRQFIRsH7i9
MjMXmEoNhHAb1y8EZFvOHzmWWWuNuY7Tivo7YYuHjlckNUzHr5Fz4W8Nb6u8e3+wKzPkNsy8oUkQ
6pt5qQKHNB6afMKjbaQtobp4XsCRlxpGITTiWo+z7s/vu3gw0ank0bjFhOfufN+pi0xS1dUMHmUx
846kbysXZAVcTYxRaxXm5pfbL6YsOTW5exa5oj6uow/3pLWeUEwsJhZpc1/GkQkMmuv8FoFL9TuN
Qd9gFK6yY9dJVXEA0huuodRbIWdDl3sK+rrDZ0YA6E9Ew6i37tHfWdPA7tF2k6+uZVBekKVl26Uu
HvJ+yWrBrt5whJxKOd5w9CI2FKgt9ymtz+zKB8HcHpnGoSGLgDX9LoWPNO6wyK3830vJuhgZKbOH
Xc+56GbxfaSYd4szEpOSS+xL/UJ9ve2UpZ80cANUeSFPtlFKx3ezzsiAWkDS1UnktcpBWzPL6bbR
iABXtRhcw3JSOmq65+6u2+uJjfrI1ftQRdAOsksr01eGNQhuf1klFaVOK7fhWUFDIvMAuWJfyZ2b
W+WwjpxJq7XConiSL44UK03FFCMm6Cok1EXfXgkPbKBlpL8Abz3QmlAR5yiiOKML7voTb/lceBJE
LaMsmtYbd96oJm8IrOOzPUBas1P+my1/H/Y/hcYT008vG4CbZ3i2IuwbwMka6+uH/pMQ0LiPkJgM
tAP0nhyMZY/vKw7mjA5G55lDFIaJnYIfx/XpbtdKraXygrx+vNOiFRgL8wqNQmrcZWi7M1Puv+xO
GIaxVexV7KR0rlMiqQLzjKcz8pf/wDmdICg3ZR8LPIgu84eaIClboQ7NiIHZEOpkmq5I4QG3OKyr
6UWAqjLJ9LgRPksEID5BBX030ME9aKTYMYMmKlI1FAzIHSF0ny1IZYdPPMDh56XDEOFggjUcKj9Z
jAvlP4hodqelOsPL2EmqibP3TFl64nWzHNBKTUVGPGKKL6rqHTMM3myuSQRUlcI8ctezeZGJ648n
sSpE0PG6mjat93Pw8Z/UgzSgff+yFryshgXYZ6C8brOrSFO/TDeemrrHldZdu8nJ5ViR7YnE56dn
LcXLgkkgzFTKQP3fX9+Ahp0g7T8g6KBg7/59hLlgGiTytEvaZi/XZHI+XfjpHJLfwLEoLw6RqMuy
IeDxxZeHne0G+Zf9t6o+4XGvm/qb+vECapNhNd0EoIYfcf7ljpNPUucPYBhTJTSrs9JMhlRevTDP
JSosTxhDFfiH6urQvvZA3VRJDVAZjbeHdcXMZypDHH8XEJtwkDBnxKpm60cK8egdsNOJ9j2OuIRk
7X4G1AKNnsXuAYB3Naps1UNlUZLtF+sR6gPKIyZYvOfR5DjYwU2do0GP9ttzP2p/pSTcZKZiNJjp
JsQbpFZZ14PHyAxo50o3UUs/9uUuXz5BERInPOtxXQyE/fKeaGqoQE3vmRrjpSbPirm7ME8IhVmh
5BFg7kD5IOHQeySv+5wO9WwfCy7eTEKiiqpYYSk5WnHqYs6ez9meQYX3SSEdwO/ag0WphomkFvmP
recYZgPi5jQLoak0dj0bi+kw4LkKtFcEAE8GCsbGpKerp2RQ2l0SqzLXmQJw7ZC55g5n0Jdw1/h+
CWPH9/EQJSPOWyY5uCvCdcwZJh+EV3bj9vKqrbcQoFmcWOH6kJud8ot+GjzakjBEQp/8u9HGIaiR
5a59XrTANQGFR+RLNEDy80/LGmsG5qwUeDq6kABPWXFKW2wZ/Nyu0CwJ1+YOAwrOmwxokKICgi6B
qxp0qR9s9rUZtciJnQ/I7sGaBmnMhiAsmnoyV2BRGnRmMjwJhKcwC+Xur6QobIFcV0syd86QlNNQ
U/rs7+XPQS4wZdCqly1kA3pWirfymX7YqUL8hKvFKD3GmckqktZYLqh2FBKXxz3Q6Z/4hlYkShb1
zGoC7svwEYTJFbr4czEwJqqncbqTxRxW9Fh6mup0Uo/MOCVHkPhsoZ46JNi4PCRdPbf+8Rk4G0PV
Gqr5etntVAidpI8WXl+wAJwpjNkP/0yp+VBo7tgEpHET59niDIgXWOrUB7hQy/WfKtwgvHBv999f
XojmgQbCB/UYqzzuQJCv1bRAUpJNylDeozOnI2IFCRp5qWvYp/kcel/a8eCN+w+GM3g/q3hzcBpU
qodSlEuUHOZyFuE1njwVg7ljL17+kPf9efIUJ4Y7J4+3RZnhGb+Nc5ql+NMVZs85Ype3coWWOGe8
ze8oA5+nBQNLyTQeYD2NSDv2peL3az5J9YoMgFynldO/d5Nl1Q2lislEu3DLYvwW3ptJfJP+VdRP
G2/2ND5DSdREY34NYzO07/axAEw6Vi8fiLPYHZU/qV5jdOCLakH5xUfAbLZkxC0hBSPE5PIDonOp
XKSesBheOPub+WBlOaCsLIG+F5OB9CCkh+7bD0xqBJhGaeB0L0YTlVlZoflYg5/P1nP9MVEalSmF
rHQlt15fy4PAKwIBaoeqsXXuHziUbHbGOST6RMWyllnntvpZeEK3MpgRTp+LWkF/p54h5T7ayjUd
XBRi9dyP5g0rTJa8Ly6Rji/CxZ4l8fsFgXaqh8yqx2+1NXbumSV8wEjF+2GPec9sBE3UnrBFrXYC
oUqos7bDQTzgqACxEOu0hGoJW7oMebahPBrRwjC+KNnM8hn+oPk2Rt1mYAy2piMRPfr3A78KomQU
xYr4/kLS07Y7gFZZ8GVVYvR+sBWsRkDg8M2BoiLrhcR9HnlPxQA2UvSP7oZsX/x0J4VCPuxsanZR
ij7P61MVn0Pe0txPyOMxIWf3mbU6M6WzHQJrJ/DdnUKON99whyCO1s5mku1iBZKMMHe1dwXpEbfK
Sosobkz8iru8Y5+gjbUEG/0uUvQPbEv2c/tMNYbBu/Kz7hd9/MP7QagB7dWT3XoH666BBDESASXX
/uaFyZ7oZGyxqfq20mD058kGiMzVBHs2lPYjyVl766GxV3vnVrSf45dvWi+201z88DjvXQhVJdSq
3ig3AciMHL1QkGqchoOKdQpCOIe9i9SjQ2zZsoZv9fiIbt3HljsH7D5GZ68172zAKRBbahwLlrXP
5aclXbCbpP63shpSUG9Rih+lbp9Um++dRavgfRvkWkrOmH0aqXRSXRAqCo/weurVcAoMhFy+yXya
/jCG1+/ww+YQEfI0eagbwJwm9QZ7C1NbAx9RovQwAy5kU/VqAUURGoK0J6BoS82ycErakOsz8L6v
QfdQzqfq2sBWIj3ed8cKaJE0gZ5+T7AMPPnysZUt3sdpFq91U31VW02h6b3VpZsYfnyoqAXs7MQT
ytG7am7wilRwcZVrDzkG6raIGkVoS+7BGBEwzz6bYyzscebmIUaVwk2bShPhkH6vp4CWpCnPJtii
BaPH02Gmw1Bg6DXIRlShft22wC2SzWNTmBrBaGfbppfQDMFk1I2sZEDNH7IRfuKLjOp2d9uh9Urd
L0e/+sBzl2sonUVzg5093sDOaSOFnQDrIq5aNrPHqAZv2UatYAUsDsZj0bvZPp8AnP5O9oj9NZUE
gSfK1Jwm8YAPPUrQMfkdiEmoiFG1WX+snB16zhzZI5ai0EEoIDEIMBXG4yx1vHRBciHhVX8HmJ7w
pjqNWDigmtkenAiCzj6bneFAtDnLZE2WnpcJCGDV0VDFnJFjXEIsiDexgu2HI7tc4VTKEiPZ+jg4
bNy+P7gDJKPuOk0avqswwgkMVZNhPUiqKdVIn/Wyo40dBLPJIX9Ny4Xlu7Uj7gfaR+6wRFpg0vDJ
rM9l8amAOubmXdM45qFETncMBTW2E3hYfPwIOFrIiA5C+orU/Zol+UsQt1G1ZUEH9jFdUlfhEsoF
ut+d/f9yIuUUQGq4QS+NNqQv6P89AQHVEdK9e1LhPNnbw29M884MsL2w8z20l1UGrrVqmg3HbLN1
R1tXXZ4NJSgDZcPUHzn3aUVPUzFVmBolUsP6x2dWvtnGcA/ZQIzF4SNue+Ct8uuFfHDaBr6Mj9Sy
OWgpnWRv0F3Ov/tiAhu73jT1f48GBbxz1wFBwpt79pyIW2jQckXIx984UjmU+tDKLo5R05R4++gS
Yh2wi9JclZiMK24h1OlZRisNfp3zZ81Ew94syBdw0/mY5uP+eNzJG+gb27A3X8zUK5EC45hE1dAX
RpufEUL7GdvH+76JJjArvxxndwdx8+XO7RAAa4e9EEDFp9QdjGV0mOnvRSF0ouknL5nLxTOBPBek
72xSWzKR5A2RMjSnh/dCVDbxuhjkiO1y8kYI9trEka6HHD6HZ/JPujwMJbDTJP1T1l4iIFeQf69E
0rUTJipEQa3T9v0MYbP6I2uZT847aCRkuJ8LmKnWvWc+88vTZn8SXBRaoK0+TNpXxFrPnQlvFLRz
Jgsjgl2qUKfdl16Y7Mt1bbFprzarmuh8yFheMD3PJH7Z6kXYYGHar3R8uu3hNe5yU1nfwofH/Sho
FFVFCJ91QjeuxB1d7tsRBwzzrHqRi5KXSKvJUEMOScZR2/74YHJmPdoYGxDFPbNVzV4ZhIgvzVoZ
hVCYer8PhWrD7rZxkbJAdH752TX3UGH9VwFOyipE78ljNhVIjA8BmHaDRRUiLGX39LD8JyjNemuc
FZRcIShWhmd+oAY0bNhh/g2ioiZv7ykztfv4gL9DWzQiNByvf8PMh8fvti8o3NlirI6McLg/unoW
Jsd5lyGhr71nF7XmDXd+uctBkh2hVhMg5/BId+UQbCz2KCxdodHxURPDz/Sk4JpidrUhR2kv7j6a
xbMhp7Ri5vYz8wuvpp9uCPsxo+wZkKsNUNK49FVzg76XtMKDuy8Qg2hvvlZMc1dCGBUPqI5cH31z
1l+F+NWlb8stHBq/3rCA7ofoFQ2NxAHW9Dk2iGSXCpl7I7P/AZUZ2itvVDhYivGD3liY4F25QcVJ
81zmnwshpW+rJuYWH2s7IIoP+cVW/dqVIDEk9QVZT5ku60CLI0Gx4DLgK2B2fg4dCGJV7grIOpdI
F6dV5yMsSgnq9I3ux9MksIjkf0kdvAp8JWZI89IvJ8TacNij5pudvASOZwU+RQNkIEfd7igT2vq6
/t79SGrx71WiWpj1q+25ij81SYOz6QwifoSTwJAHfiRAOMKAVxvSHZRJYo0mYEnv63G2MFT5RWK5
PrrxnkPj4SCuUfMolctTQI3NfdrMg6A+suP30zBkwXltyutb8llFtUMny7J83b2LaHou5VA43l8U
UCxICL8YXcI9LtHShW/x643x/k7IErb+Db/u2gYixjylNsbeleA1njpM0qFIvk+9NWySJrjU7szH
lPfgDAab5wwHCDzq7eONS/OmoVzuUDgVIBS8VP2nTHH9yDAXMptXlaeQL7iJWKNVeyL8GCNQ4tl3
/NbenQ+2gCcAMzTo/C+RFeXjZydoCrwECVsTOt1WMicJwbeBaDYkrqcjL7O09ucO//4sFRJZ6q/I
NM9Gd6DY7pcugFlKJk/0ZTJNJ9cu5YZvaGKEXF0lj0uFLYai7DZJCpkpSggzUNPKHNkJ2AlXKAoH
NIxZhd9YdAZPBML6HZS4Fq73ydvDhqGg9BxDo7lFP3ZScIcnyEpIrbc92M3O/5QPEMqLCVjfCUsL
7dzMVzZw4SsgHRAnjoEE9OhrlUJT5/JLfn9+Fa3U8hUyCM6z+cGMFDTIvYpIqGiyZxAhxK2s67Nf
ogOdKy2N+zZWbiVs4N4ymP6y3GTS8hoo5nEBE1oA2jIq6UC7nQ0CFvIGPfztfSSURVy5HTpDyzSq
MINUylqIZ1SnSxc4rF3qEtR1S8x/sJb3AYBYvOe7WmBrh2IVCQoJRBpq3cCEw7hkcvUUwyAagZvT
nlVadjyLmvm0Z7kV42uh8rM4upr475VtibfU9+Cov6oq9xPmNc6cfbw/vmd/ShfcA4+tputww2ET
qgvblJ7AhrV/guFQYBgGZeanNEM/oDqLtLc/khF8199ATG2Ghxqm76Bl5DzzdT3fUBE9laz+7pss
pd9VJr7raJwAXqBM1w/UmkyIBnHRFtT195GDfOOFalrE5DteorxUHj8TRdBBOZnxJtkYd3YCX5bn
LZrap6vlOTRz2tMSILAJ4ydWFtXwzPiuZfHx/9ZRM5aDNq25jLjImrS4t3L4WSB+jQjRjWHajvxi
kIPuXdKqRGonijMT/ywYAG5k3410Ftni45OQzhZhq9S6ooYIVvWy6EIDkWEXpodb28S7nNQHWOsl
q45E3B2ls9K4Ma88aZ2nq3cozD8FGXt+82hRFtZKAO8zbM6bK0ra7FQmKwA3pwI4XLbPgaZbgAhF
UxBP1v1fduMJKeyTFdSzlRVrwsc0hwzRW1vs7eskS0t2wZeIzi6TP7hY7mV6q3X2s1FLuhRSKW5W
Zii15OJo09QCQO3J91aDZazojNzz4m2MdPRPM60qdSolbqydLZB/Q4mE/M14uaIN0ghwuczk1aot
K++3/qbwCLld1MNvuKh5kmKTfK3sMYFTvzaBxtU0Oi4wkI1rF27LxVwRT/MfKDIwNb1DYd0BtM/g
u7zXr/RPxla+OAA+lKuBNt7ddiA301ypgwE6DHlbWfK8canltWGE/rO3ChU+pKoJThxhxqrdFwZQ
NMxYjWF3ymYUfWjB81QADnHFXfq02g4G7c0F5vcKvuF8LV+fkdP+Ljb5DQY1BsL3RLD+FirYCBIO
lwEGusCLLRN+rQ2u0OelFDoDESP2Iz8aetzlSstTeuVfgUWkUcwRIKpLVR5jThIOwOPKSgWGqx8p
9vGF/KCw7uENTBbz1b2/x62T/wXpA1XyBRxz89W36yU3dCbQn1hbhczFS+KteuFalrpGkAfHzIFA
FPFfck79s2M4EJ6ENyCbnbxf69lZpMyI0XEZmZs1ADL1byp5WXLdhgvtfIj6LhrYbeYVw7gmeQ13
6MWKfZpYXCFIrKNmZ+WYdW613QmR+KgiPGPoV4QZOc7O2aN+30YFF3WCBB4pGApQv+74vNBqo69p
/+4H+BgdDa9bPqyU+H9AeDyIWwhEuEpOqaoEF1JrIoXTdgNsCAtNLxMcI1TQXvi955aIEkQA1p/A
aS4pztcWjJtfhSD42AiMo0upt9B5QYT6/zKSkBeJZc6qMyB2ZdxSxd+gUIHnWYhxB0EWDw9CPoQc
frcSfFJDH94ZfsYJmPPgYh6Ft7HvPy0V18a4mdPav6M55/acuK7pvCEGu0cF3nlxEWmRahl2L/hv
wbhwuVo5T3CUtuDQc/TldeHe53edgy08zOipmzuFagRUlywZN9ZocP9rtA6CSV5VCwHTmUSOsMoN
8j/7UBaxBVhiBzujDrMiE/b+kW8KDbhz8ktULytI8BYNOtYgTEUc/dF8wwC/G40RvLpK2wrpFirf
zkQFKNJxx39C1gqewOfcEtLzK2cvqvcylVsv4F3IjZj4QcMbRoMebq58a+YmFplnpFeFUZ7DURs/
TWskV3BdM1tzXCtwwHPh/QhBopljbtXc9wUxU6Sxu8LEOwLAh6JxUZ6GgSuH3AuaSjm7i6K4hD43
IzSrwydeUHkqeGkClKdSieuxVJx46Aoe4u5RnIEDMOQu7ENyk8MC8GCZxwe/AC5z/Nww4Tn5UzCG
crAaqj0gujFtd2lanxpnmrY02e2r1Bt3IaLat3PeU9Y/XCYLmRlEo88nd9vPo6HPNL/OXhYYPc2Z
olmcI9cKsdygKeOA5YkUF1kPGMgBwK4OwBxcDjlYj8WT0Rv7DaZCdixrfGbXl37W8v5sP3wEXJ1p
35gp524/jlw08rakxC76WoXiFNAjH5hnV2HU7StkoItxUcgQ8NDqI/8eP9B2SLxZkVXYsBg1pJcU
KfvFXCNxZS5zwnNamkpgFHwPpMQL4sR4/lJmhvDPs6TUlHhx0qm4EZY7naMISAvkqbRAgbYwsrH+
0Nun8V7QPVCqWsGtDW/l09lLDVjZgeDhn/DPIqj0NblS4PdIkD7jze5w+pRQ45CDtkqQnCi+NmCZ
r0Gu04/vKyHbjU5pBx2hd9xxr82fLBawCBHz17U5+eWpF9l3FG8gWP1YaipSKYlG8pycx9tFrhbh
2swhRSloOAR50/H/bCqTciFxctBlIwPBbVTDfLISeaoE/Pf2YtJhX6EkOztY1K1VoUYltqtOqcnZ
w/wl+uVjF+WreokyVqrbrBQ9cRgk38cVTS+ySn8SonqBLOaUF96e5J9TDo3ryEg/Cpc62Obmyui+
yaz/pBsU1whxJ+XsP7CZHR1RCl3pg3rnOi7D191Aadv17IrHaliDdxpLuCbswRrBXSTtqTmzOt4X
pCO1HdPhKz4uLUZyS3wDIbQP3txCtgDDTz99UfIRKiOLu6tUSyAzIq9rhrgUBDrkO6KXIbD0ABbT
34DrSdKxpQ+SKj6/Keg0esBiUAEEWxNniIM9ueZoafOhopMoQqkDSfDgVoKWIPsB3mv186f46RNO
6JvVRdlYQKnpy95QmmPLu/FOFTGGrAKY7N+BCpn4jGJuziWHdsfOO8OHM3vmVZHiqGz2t+EDEBJ/
7Ky3SK2q4B2SU2QvgdmgOy4wFqSP4LCSS0MdDrfZ90KPdsttqApDQL7aKJWlLbSZuU1Yjoz28/+N
+ygqNQpADkgsJTxpEbzbJVV8nWMZ0Z1UvRVlFk5Co8KF/i8KGwELrHs1DPfj0cW9hb8pLmxv12AT
4CkM0Q6dE9Ub9kHio23M7gLndHwX2oR0DJqqZ86aP8T2xNCuarciTqkEOdbYpuUqJXuJmhRgASSI
ehTbTBo+pz92iNUkTFiG9ls1HVYxpnEaqlWv/GA1jH9LONQt+gfCz1y8vBu+1Y+WcDn+nXUK++Vg
/Vi27W2DueytgJ1BJwmyUUyf+7jKTXBcaotKzTGTetuUA+d2DISwuiBoDcRpepCCGuc3UXhf27c6
AulpIYXcVLqDtGBF3NpKoL2nx89YdYJY1/8L9yCj7819VcQCgLD5hSWsPX0lc79uQpsFYEss8veV
bkuPXG+gPhyjO4bn7r9POq7V7WtogfdVdVT8ilv08TGmhXIRyyz0TiTL923C6uNsRuYmaLhboZjb
gU7z5/hsQS/zdpF10fV9HSBPzYZ8RaVm7k5QycL37zx3GvNJOcXOgRY9RalyNVMOMsKPzjM2hz2m
zb8P3tBa786b3r7gfH+BL8wd5iPTA8inBI1ibEcnQLYT5zPTV9tphhlCGVrqtLDnL6WnRMTNuzmi
OSjqYBj19VUtZzrWh7sRgfVwI+eOwsZyCP7UeSYtvFkuBm/c4HEF9BaZd4oM+sNvzT0I0yCzA0Tt
9iEAlSQjo4iEFXDs23l9ldXlNrgKCKvOjoycwsLdjNbButNlfQ+0+6w7eM5sJHN9+Efb0nyV7fnw
+o8fzAjIJJSiLOiMulGSGCEMq+9OoSyG6H+Cjp2X5xCshC8Q31CtnJG+0T/SaOFPVcFbo38JLobl
Zpcb2lxSd9cz8uNRpWhI51QwTzpGqtn+M+01GbW2e1LSzJMM7zcsZH0LDUBiD8yIcSQ6g/+jNr9f
MILHdoD0aiU+XVcleoEWKzWvGynSEZfomZHxQ9z3vD+paaWyOtpAYk0iP7Hx8mgFsJH6N95hj3H9
OtS9nCWfuV3JJHUjL+dDGZw9SJxLaaUBn8/8E2wy/pRZzuBI6FK50DbvPaTgXJCX4fDRvKSo8p3Z
UBvAXVA9xNT9ZZsFKaOm+59hC0qb9ezSQ7V5rahyh28Lec0+8mBYDjJGFR7ZnHiqKftr1FzbY6Qu
WDym38Vj/QHTxOfUxk6y06hQDh4jMA1lpfy4dW9YTxv1Oyc4dGd3HwA0cgDWRtq9HLjxx0J/Jf0b
GuekwG50DMppSR3PibvdTHAil2za3KkT/5KmlUujpfTHTquIHsQ3SaF2MfHAYu7MKnQnGQYKpZ2E
gs9cmbaP11zkvDeTRB1rR1T7d7DJqi3tMs2jqaqR8HOLQ/SM2bNHNCceNYqmfXbbq0yDkQI5jO4L
rYW+YW2zDdOlN6kzJ+da+C5g1Lkps/6YZ8wfO9KGtQ5svrGJgJGaimbofBvWs5xD8qZ4l9x+wkCu
EJZ3q6rTqqGh7Cd3VnxbH+wXxOjQJ4NWanr4A+/PeqmyevjR4LVuuW8giZk95Rxg4DFPg7z15GG0
hwU4V6brU06nl0mTSwj5R3MUO9XJWe6Jjp3RtqY+ScY4mwz4Gk9La9krHVzDlcN+EkoyR1FxZIhH
BoYfSzmpkbzObMgVfZl6Zijk7sEh/f2x0GHxMhMt4s28bYr7/PHTMFDA6LROqp2Np5pLM5mAu/K+
8Ut/jATplm9uyFzQ0h/AzxgYIvFQUk7Gck6rYm28io+lrtaQLxZjcOqPwet1JZxw1E0Wl5Gr3Lg/
S/iT+Ow/STiHUYo7tfSH1izXr8DzHLXL4glVnxMtrXSv8QMhVSd7jCXXPhcR2RVEmgK8b3q+dJgc
RjLz5AuN1dLMZFPZ/NUh16I2lxBg4AR1WpVrCp4Xr/n1v7IRoe/jqFM+TcHXIxf20f2+JAgZ4JDW
tDB53ozbaaZQdVgz+7XH/J/A6FNMLA8cmmTIQpI7PyZMfTG4P6ggT/kWRTXCXhfCLZUXiGBPTOvf
fkEtbuXQLcjI8w6OFPGIK975iqOtVaKaBNAPDoH2O2yIuqUPMjgwADMqr46w1KkLBq2FbohkbUBk
0+WrOPBp9LarpEOQYRT6x3wZjPmirlOB1lp5AxCjpcN/21RywyKasqXhP/iiFAjT00tTegBaEaqU
sNtPXEBJS5/Qd9xjFri/lvX0itRH/jxv51EX52AtZ1sjtZR2vgkKryOICi/vf7FFVaodwy19kfBb
cAO0psRShPdy2VowS5ogH+Uu36lOrIqRiAeaHmF/fnbC/R6Q3eG9chUA1gJlKRNA2l4vSM5OwBcS
GWIwRy+G1jxAdpQ5Sb5/LmT4E1cvUcc1Ql1KIZrDCZ228hpKq+L90M5Sza5xG6mBmWHojez5cYi2
ZUt2cVPH70Ka4SpI2GZWOkRURJhAmie36SBeGJbelRt3BbWQ2gaVt14WHn2TDXaKBS39CNwDDs0q
EPdILE4j3QylhKrUtPbaHgIHmLuClRAm4griMum4daaW3WgIBETutdSiNoyKfbayJMcOOGhySQal
yNMtPOrdAg4ZFvBynqxQqy8hut82y81FaZV2YZE9UDZQz1Ep8LFzQwcC6oHJdgTfqx+rg+JCI1VE
wYgbwJ6/rs3UAurbDxVmirEJZ3tEfo7cbkM6gmPvJVBb0yLf3wryNq9J4SFI/jk+A/vFFBzaj4K1
4qD+zn2ppnIGGIl54SIHfUu1quy68DEiUzIui3H69Ke5Zze/ustHQFYp6EbPx2UVrLcXL4lT/c1z
ZzHJ5Tc3u169WMDtrlBf1nSi+Cn4Y6ZDRdz8kKap8+9fwVyZbLdlDzwAeymHT7Y6GSMHoUfQfm1x
8hS6gcHmoe+afSExBUHG5sdz0px5IwxcPqktyVfOdtHNyizFUdXAqsg51brkrV+hGNKMuqrSU4yM
zMxHnddk0pQlW3zSn/JKKrTKNw9MG7CNwOVx/ZNl9XY5spga+WKP7zaRIwLC57a9KLZ7enUwWhEo
o4UH0TbRigUezXnwWYiHvoU+rqLlakZYP0ED//d0NHf9nZCbcKMEPtoo12NcRWGIuRWox/grm2Rz
BAqBCo17T3bZoEe2Q+O59W0Hflh911Jgd3fL8Lpw1l8BKRAy8Y2t43yAiCfU3eDepRXQh8N6LvAd
bqruEWYZhJwhslRMy+SIjsAbXJ8/AP4c2VblkFunbZy1kwEKJiDP6EM8+CdOUqAbt2BsdAF1os+B
EJ3ES1GvqmeTSlIbR6LNeQkaqpVcqof+d8Nr4hF2N/CMcA6Zk+TWx/pqVZ8N8wUTF9Kspfvnr1EN
U+UtCMVZcz5Wconf2zR3Wzqpl5H5RtPQiZJn/nC1Fe4qHf6Sj3IFPOfZoFmUyEUvmL8r5XFidbqk
dKcUsaPae/rXNE+jSMBVDOpABlV5PBcL9NiELi82VxMVe9FBqkZ82igoe1qSWUQSD6gDtWGJeyfH
zZwtgo+by05g8TRxm16tH5kEsWMhle7wR5G0EZwjQWRx5YJgA+Gar3kvS3jO6XC9aQNW5YkGVhE6
SpOlRapa6eVaTeCdap94k3/qFClfhIUgCJPtB0l8f6Rnd43c/oC0j6BjmPlNrtRe4DjiIkh8CtIj
49hlRntMztD9VOByBfMlAx3geA9tCtxiLFQwbP6NbrZ0r57zLqLNguiddzfcHynjSZip574SQxct
XUBgZR6DUWOwOMQmtk6OCVc3ouR6w/4jYUSfWKjhxVIt8nvFftucF33cv9LueVr6wh6dZgRFxkkZ
d9BuKvaJRQbiRFqhM4aWfzR3BM94COJOLZP85nF4rlm2cJrY+SPLWFx0ROOJfFCXm7DO9NtU72M6
QClFBPlTI9UTIGavp2jDNSFBHIHGxgnSEXUjtb0fb23gHCBmUygri3fH7fxFUuGaAg2py5wVXbVf
nT2Qg/302nhz5yHONQWxDPdqHBx7JpztpaGzupvhymV5f1IN0VHOmLQ2INgVR/mN0ng9u0qy6tIN
fK378idApiUq+gRTSdqrP0iDK6mD31zIUpP+IDKzYi1FCzSJhUh9YQZ8RiMzsBqKZZbaFu1Fopvd
c72eXtcYwCOJyzC8G02ANk8vscqyiUPkup5bYHhYrXeqLh8/MPcqniuFZri9Lhv+U7UaOohGvuAM
IMKM5J7D814Rnozvdf26RX+GVXIiF7yXjQPZan8yeQ8UbP7inyDznBc6i++WdkyWcA9jjUaxk5d3
AgVE223ban1Q1ikvnTgzbFv31t/bP7By8GkQBciyc7ObcDLx8nQS65QYwzXb43Y1MKDelFQyitHh
L/MQAiKh4K3545ahQl57/mfg8MTcKwyh6iobIVICxCaCTqsB/OTmvrxr8IDwqygKqZ6bmSdaFYz2
N02HT5TFT4Ug3C/LCBOiUvRQRuD44xwHVU3igJyFVqQyIXmupqgxOgtJSyQKV8q2SFUlDjI/S9yM
msjXf4JUfyzdvMBEnBznm2eGJCqSI1W7N7SNgpFtxjY2wd7SmWvrxFzc11/rGhgewb7KqmGPIUaW
SHE0yGS0D5A3Cb9lNKs2jrslmKAjc1AmcDE6yCYb82Dc92aT0OrBNlMJyibjtQqxYc0FS+x4U3z9
TA+9OCB3p0CWtQod1kxAHKGdJn8Z+b8Y1vREyzzyaMoVaiZgrQcgfa0nqDixYON+ZrMqAiBpyZPz
I8UwOephBh1gWKUxzVGeN/8CM8KqCegmKddL0+GtoM6Gi0jiIW6BDzeXWOCDCIuUYoJ3Ye26oy0M
b7DPKzGlvIo4TNy9kN8UVs7qPRsOErQlsHJJwQMPFG9ZZ7aOPGYmjTPzm/H1E+B83z8efTNKVE8/
Fvw41WSbP6L7T5Y7JBk5Jh7sNb+3yWVeTjnnCMGZVBGcCAWnpMoA9ktIhcKdo+HlRpBykfXJCOuE
h9Qhbqph9QqEfPM1gLFUw/p0vy5uWuXh56ih8f/DApMeDtxEDiMAJD7Z1n/i0Gd6ujjPRN0iO4fu
LFvis7PSCPdDvjslq+5rsjaknAIXYVThuFP/SCBFY77eIDiMzo00GS65aHJScjbHe5H+XrJdCWn6
Vt1g5T/0QIBu1FAP1EF/QMPjl2Len4KK/bYXcEBEJ+jEKRqkPMW+Raj4xG9jkwtifptZM/LjGSYQ
DobL9b5mhRNWe2tQvFxnwsss9qaX9zsgIPt0q+/EZML94S48zCZPxiCYYU8GMVqWJOKMpV1/40oz
vHqFJqSS/ZY9WVuXcNEkkyefVM7Th1Hqe0mdD/TEBbhLKeo45PWt7eCuPxW8W4qr87p+Wnyv/Qe8
ctrjQIugelbrizjiKoOgMimhCnsQlu3Sro8jZhXAhF8mASdpvDFd34+eBC3HQm2b6aGpUu6hLHWv
S+jidXVq7/spHtYey4iMAv636pRcGh0pYM4yViPObieY8Jstv+wVFa/MI0j7I7fEeC2EbFOcslAt
zI1fhqRPTNYNWbTN/QIJLDypRK07kIWaDExmOCAsJOP+5MclmZV5ojOvAZhGd7ok9JHfIysVoaAn
XW2Z2A7gDcDW9tC2lIFJQewgnTNEgVnJgDV5daG0Ksku+2i2sQW8Sy/En7XO8zkIBV4F/cOfq9VV
NdZYuCUbpSL8kUqgYIJNc6tKUbEJD4i0DxAJ7HqRs80xNYF2XwmmFb0XahdF3mbOrQ2aDXTpDbRz
/7fnabB+ESPArYfElW+2nTSkrsBomeFhqkSCjM17FbKaTlee3YcfMmXbpC200Qonp6ri+m2dwrsQ
XUFWqyORGxz8cYJ0FGhIW73B+ob3EZfOakOxdesS96WVr4sWkJMDeuoWUym1gBoAIFjctz5Sg/Q1
pDqO7W4V2rZZDZ9z+ga0jgdgs7JNnx7tFDaJ97KXcxXLumuBq8GUa4tPyGuuXn0uIMJ3+BFdmmzO
fcVC+Ww4LJd3s6d13sWcroyrA48hjgadGurlblNEnEmnYwmSgt1D6nmJdVP+vHJB4kiqlkmy3xTb
NQhA7pwUtgU8OQMNhHkOQjvbsa2ylYQlyol2ROrRzBHupDlBZC9bxLAyfNzRm/XNIEL7QFK81VAX
H0fyUIfFEpeKLkZ/XlQXtEo1UGVXft/oaQRjpxhJih3wQrQOgVbvX+QL1APKlgj1zjNtnNRtsmLy
BWAy7PEBp+FuPDr1y4BWdRcCeBimUG0eci9GLrV+0YWl5vDsSQuYxaNAV4Za3PWv2xxJMxRA/C7F
pQPRaQ9/mbebjhYOBiRl63GB6w3OAlFPGlePKQwky6X5roJa+7aivvg8TKW7dUGGQ8drwshIjOcD
THxvmHDxJU9pjHtVI5X7sAZJVj6dcJhAr/MauTlfcDuorZ/M8pGETBzxvyW0+yoTVZTdJZr6pyvj
MPsA2UAq9p8RUiimsxXO/5f3gKvjfZ/RoqIOMEOCEjsdhRvjzZSN7qu7Nk0eThykVqMz9v/bt2WT
7Te6TQItMN0knxY5DUVt24b/IrOZQxAkW6uS/1snu/5EXVwHYHNhLLde3OWdkmwVNXtG52DpABET
M0CQAzTTOCZWx2hRUTe9SCpPHlJ1wLGCWZFnaY/B2lLQ1wp5tpbNmre+NN0oK8/isAaNRW4cTYAK
Gr2GiSqdod4AS/LoGD8EKXwxo9PPYjC+ZtRzIEXqqok0BjreXB1d8G/kvZr+ICjGrXBdGq9QKjcI
yGG/qdBC15oYAGgk20IAFhN8nNe1jvrtzsIxvAbhtHYPdHsfViuUfeRNuulCqOvHgsFnwHnuXPoQ
I9MDJY9McRpVRLiyTJIthQha/uyiS6l6AI0s0hEn09GY7Y+7M7TzBKeIoUx1rgFwOOIeL0SEWuUW
6BgM5nSIzRt0Csp3AhkqQOzZz418aIDDwk9AiOaJor9BKRpdWePkp4WFcQLW+RS/mrq5cgp6qVLv
4Q16ret7Q8HCI3kYxgss010LXSIWTA73OKK0qv4rgfO6FS9FaolZWmU+f4QPoDSabB/kX0lUYrvU
ZUXHZyFjOlxp2TLsSAvR3cLMOSzjX6jrSUIP/wqI0l7fSPFSWGejIrIUIGN4Wk+ccveZJihFK9NP
XYzVLjS4K4f5EJQgbrBfVAeFGhtGZu4OnQCzpgbmyoZ1eFu2cvKzxr6DHH3LX6j3mgOoewrA6Q9h
eqOhNXPegzJese4YeShcRuLIc4+C7PNPZDP2eJIg/GxY6+fWgDV3uutW0JuZxGLHKXQVKh/ICoNJ
ezP35MGqKLStMbwUFldzTPUObN923jypgoNTdLAL+FB7/RIJbyYxLZYtG52iJXm8zk9PVP0qXNOL
eWmlCE4vD8Zmj6MniAKnszdIfcc3n4iIxsXFXZrh7uiWFIAVkek711GtTkqi4k058yoNViV0YHuk
yotQt20v3A/vS/9d1fHzOBzvgXZvmV7z4KpGZyI6iPQ2FE8wujGM6Qy091zj89+Kwhm+LN62R0GP
dfSqdo4hlBuR7EUhlTJPGIg5kwOEthvPQAxUG1Ra8KkPJ9+DbggGRE14X7bQ0Eie1HkiULF72uxD
8yEzF2Fk0BvLM335nL3oU770rsnLyFzKjhWqAbWE4oKbTYF9TJIQco8Ec/hWB1pYS6+jGDJuSk0R
J3gHaQ3Z3ez57+yFRg7t4lAHw/opA8vdTqC6XAtPNM1Y2OgLi0fTOVkA/w72TEn+/HjvS6Ha/LWQ
H2yOIhrFnboDB7TSbFHZgISeVFkaMA/EqnAdQ/EBxXd/zRptBmVSoL7+IvQoFCnFQjD0VGmr13T9
LiwEIubQ7F39UFkk2Xkn6adwJPJCdfCGnc+GbXTdu41bVUHGdWGXrBPnt8tf+I1JiZ3kARmYV53t
zgbNe0AioUxNAKHhvloRJujarh2fMxJYp3kJmKXoLGI1NNa8Xg6MgcyDUC/FiJC6biiSLrW9yoBA
SbMdxnLjmOqgyFWLXcjskysDHSg6nFE=
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
q9GEh+JsvmQ5rAGOlizOS2Sfeis1FuriKQb0d56TUvM3IiK1MI7H3ZTCaQVJx7wDVL1cgGDScH4B
3YCaS5LgYDpEaS4YubDaLuB+4vGt+ncYjETyeTk5aPdVmZqlW7zlyBf6DSXUgTpx/UJRBQclTqeK
nmtOGslfrb6vQ+KE24UF9gPLz+CtEYv/OV5prMDVf8hGN2zyTDwYObkx+G2mVd5UjrYAjAmapTNP
ZWvgIQTd6/v+R4/xTmbjfJGtzECigo1LFEQPc5uljYm7Ru4Gx3fsdOGN65W+mZ9ISTHWa/j/Hi0H
F4T8CB0Y9BGA/TskHsTs3YtHoT4r0OcMR02Uiw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 4528)
evHA+tVn9WI2CU0qgKPkQM5sMRBEq2WONS95Ii4u5HdeWOk6qJJzfJ8yNjxT4QbvHYBGa8UPQ7Am
xcwo0ofcZKZZRrSc7/xp1+62zcKMUVCiSaKZcrlwfK67U5eyk1Xxc1ufDAY4xeKyg4KjF4o1iqsP
3dexRsyv3sVmfxZCOLf9WaBzG3hH1B4sdD82jEDH+295SHjIWslszN8SaWyVf8rS9j2qm3kfnBi3
0FIxHzqCSIL+HQFsGVRXqn48YVNIvCt+PfXr9FO5Ekhyif0B3cJD+agF2JmlymQtILSEqNnAlUkM
JAwbD1XYSylMHp5YghzkQ/oJT67IwedZqx9Xu0KVFGfVtZQKJktuwT4vyIrqYUC3X64zCB1vvZv4
CB/rtjBwI3kZKDxqJcuTbPW04z+kukBZOCpiJV0eptl0Zro0Me9gEzzWPGz8AQJ45mHg7P9xJ/og
sGoYXbfr/cC7Unfuzecni0HT6/QNvhDOb4FyxYtDedAqv89atqeCrI3JpLCsTsadWNfvcL4nuMhv
kO2wppsc06ABo3ePH/Ntx8XxKPAR/wyQTm841hsCMh2pGXgy3Ti0HoE6xBODeHcP4tF7OjUWGvLl
5Qp1PJASe0FvAUXW45LX9UDyAw2PwULpQBDrSy5qdmKgIy2rqaHeW/XgWcc6Y0EPyk1Qzjef7mgy
HtrpFEzAB7NOuLpvB4vncudchZBwUfWvkHgTPS053Q6R6aK3UOcJnf00xSohB/JKBXlcRkBPb2tC
yQhUhmIIW4Otm4/wjF50vG9UD/7StlocTHwmH8f6Ka0XOZQT8Al9GLRVKxXLFruXirKzfBJn1OBF
pGZuW3fwDdg4AflOphMAyDIvXbjnylZB5Wbl90wwGOP+A4DNrv88+iWvqJjVzO5aeeGgj/DZt6lk
HIMt9uK0PDNtgcySvduo4jEHyXkovrbGRPvGwoCexO7BzDZ5Uv9edGxwuAveJ+wepn7580os/VR4
VX5Ki8iM9Nds+47wx1xA0lY+bJeYdWdwr31f4F1pDUan3cpL2QKlyM7c7fQ/IptCaqYNgyu3cSJ/
PsOxGl48uiixE9dzTIub+5UH+CrcN763unUfqUWeaQO/T5qD41DgHcmPy1bbJl8Qo+Uzb7nEow4C
1M8mKoUZmYR+lGw1aqWFZnvjsAWeyV2/3jDlBZN2r8YeXq32Fo3sHyaDs0ickdFmPQXIw9pT+AT5
W+488Gy8NxGWW6wAUQB+dhkROdUkQ/J5WO0EnCvWI//BtovSW0ncTEetvekZz8Cjq+woTM+JezuX
fYYq31Ia3FL1r3yB3+KTN/NGV1l7PW0losiw4lFT7iDt8VdtqU8lDugiehEEaDn1EQo9re7XQJWq
TqvCq0uugKkmElAsJRWWwwWd5MS0xYZWHSto/CM2nxMZsIsTzaMBdsuYeSOCi5KSaD4K1dEMLwBj
D6ANrdh9+BKyaI67PQrtusRWMLeCRYE7OXL2IBZbl6fuZrWBnr9gCocPU4K2FeWg2RhOcZt0gG7F
yDq4uIhAaBoGPLsQVDGUQsy0NrABmVY6f9LpUro83Yox5CwxxGx5IL+Iu90O0eo3KieVGNDG48GR
K5SFtl2Rac7M49H51XUuB6ZVY549yTskVoNcS60Rc+il0ksWzVb0F9lVEm4bsOyItiPGxbxq+xuH
Bn0or2h7+XcKNDDChU81WaUaVx2zE3JoatibO71FBaQfrf/v9d/BpJhqOrKr3eJCSfDl7EDTyFC2
cPJMtBi8H3sJ7Jtfcuwstxzi+UgIlgFfJrzseFrrQNhlDet972HxWxvkhixy88zFcBb9pQm57Uud
gP62w1vxN/RkwrKORJ/OQRtKUaQn9i/a/VaIdYIEcK8C40Gxb6tja2PeZAumUZPImmQdEg7Q17R2
/hHBqd40Pyfe8caX3fI2RmkO9nxE8fcHaKjmKA9EwlDw3vtlB2nbLflB0YZMaQI2O8UCroBkayqV
mN4t89XlCN3WX+dntvZjpVJyG5byLRJM9GG5Wxh3bboU3k/dFtHBDlLvgWAeR1TDVpIX1SVnfWqI
cbPrw8emjpLR41Y1JXPDBkmrmcXgYzKV83F0jMjSPvJegE86QaT8mZSSxetSyhL6y86IPKDsT5de
Gbd/WaV/Qu/MvAU5hj0mS/HiDxfCjmtLGNnjN2C2IIoam08z5hH+kTOzJcnf4cOidF+37ssON/0k
qgsSGm5DpgnXiAjnwsgsQVUhnXmqJKe2RvUEQ7Bp3H7lFPL6BUMpLE878uxoICosKVr+1hOIVEIE
R2yuwyJWJtotHYnofHsSD6HYx8f6gG8G7KI4AE0ENCj5yS2xFD31kmQmXi6TnAcpZvjbjOcJNndq
RaauGwfs3+gk/MnbbJciA55RaXnPo/RWuMgpFm5D6ELIsK2NiZ91oEebencDb9RsxTzJCYiRVBHp
TWPucbBGcv9QxXAhJVcz3cd3o4bR5w4+7Voyrb0goYE9cm8nRtfHpjm4nyk2GWOxx+hI3+80h5nD
FQY3yhpHdOwcMzxba8keWlZmmkr83NixzxTt+Ma6FHaY3QwPhE4TGVXifRX+uPMdJhvUGWUtwCNW
nz+hqAf1EC274Lx1nk/UPBIo/RVQwQPNRkhksPCnhSR2QuAJJng4XSu8W7FP+uBPiouhDu20Uppm
NG+k6zD1d5n/n/o/nUmvLGvDX52VowTr0GA2iJRHSMqPcP5MueSzA7PbTcy4xf3HikhgxxQg/A8o
3mCj4U2rH4JEQ/7e4DX4kQUm8LOGC6uS9pUkBze43C2xWqQnZtDmkvNiBSQVMfV8cNIPolo69a0n
eGrJ8TIhOjTp14tXRqQQBSfOvId5ImpWYHfrGqrQLhVlBDzlzoatvpDtY5+/omVS3TagHYE21re2
433aqIC94U42aFtfc+vN3JhRqMOQt314Ttuqx2YvtoHEcv6sEvj8nY3GHittALOtznm1N4yCl8DO
IGRTiWYDdp3EN1ePkp0PigXAsp3LFH0ZhFFuWonDiPy4XsxFlUXPb3EfqHjuW18jbp6ub102bhbT
bGnCxM3PsRrdVS51um/aYUnagY2BvzluzKMstg9curuDE4nmsHxd9+a9ij3KN3gopPj/yUzQmgSQ
mjZscf98Kc+FTTLUNF05GTImzxI1C3DyhA+t4qC8aAV9IPEPdEbyboqyj+wb8uwcvyVMQo4hYdEp
AVn1d8R+lPWhDGugaWoPZyBvRU79ZQ1edCszTP+nitEe7HlmNIZvf18g/Df+hzrQRrKRePFoyVmP
cr8sPALe02pc7d0OOWhB6ygXMNwvZIn36vKJQEiIWobToFvTGWGmNOEocoJbo4IeKSRijnPW7tEd
IMu//NzS2Am+QpuSuW+I69ewereUGn7i7JQ6c2QLDg19/rTfnaBMoTJeP+HK9BZzlAUu2xZxxNXW
/UpH5phXM25WzXJoqZ11DQ+BxnCyi02RNG7rQ/Uqcr2FAMGPTieM2/tyDcOrMHM30FVAVZHAaeqw
qxajDbonJAxWhFVut38wVTrrPq8RVTW8uVoJ/y8bREcvP0Gv0g5pIA04zK7budEAQVDluEb0saH+
s3+qtfHusku91nfRPCzpEG/RAPCrr6KevwCvc9On7DmerVKE+uBtGtnor8bW9/6QEG2fzgTtiuup
TdSnGqAMq71FPU8k0duOu0UwBPiN7MIaRVZ03RCLcKXnNKPr+JzM9ApdVeSJeo/rR9QkmB2rTRG4
ejKMYcq4FjPR0LVq6lE3/KSHb+gXvR1GrHa8N4Nj+T8qzsuLBdb1rUFnG6OpM1hbHlMrwAIXzHs0
J/BLktKwZ4iSgqpBb1X95o2ZVVPjNErpZtCqTuSV4NRcZ7HslH6I85GgdPSzxgWsqxPSoibUOB0Y
e7DKlGYG15/b84IpyAnZmSGCpk3Jou1mprV7BLCW+mgoqHU5uEGRJAJpJ1zyS79itSCuzVUdeGw5
TPL+6uCqkiHwaBDwotv75B0X29fM1DICUNApAX2p9PnqLB1dB8qH7o3U15iO49R8PTCZkC9pghV0
dJ6iYC+Ejn9yvWLmlPAmCN/1q0mw712+WvJaS495kD71bus1cwPAF+ji1b7VtZXExWNpD/9KS1g7
HObC6NZcZxWY0et0qSkKVZ3lE3tUAw5U+ndQk0wCmH+WAKsjzbr+kZZwg2tMLy/TcC/Lyj4EBd2a
HL41t4LA49adf8ceGaM5+DDyD0KXwyH2UyJVMhbwJscbI7lDBoO4ZaxCWDhxhvxKJakhF46n8KBe
ANxdWAQaaJC2i7A0OEQqxiEPKjtIUoATxRTUfbWGZEbmBgEGkgCIRDgrxRU+Cy1KfGAa26J/zUO/
Mrgh9reBIpvvlvTJGT/Ey/nbRc7p6cvADKKsdNFD+VHOYzzuz7PaYuO4jDhVQPHsSLo7VKvA1erh
jJMqoKT3TGK9i9fgAzmWWcA1VSD74yVFl1vy+osNK0wbbWU/ELp3Q2k8eMo4fikMkYoppwuLIu9w
SKJ9OwrMukUHG9+QiGpiiAuGxPI6njBtKyw6MsNzOcDotCAqmby0wKpYq0h+iYfzHXcDiwBeYvgy
VmOp3+d1VsrBp4afHJoXjjzWKObaBovx3xrV07qMrXF02sg0EGnlISRGXRJ2l6SRCaxKObo/7nmg
qt27/YwVCpnpWf6W5X01yn2qkUxqR/KWIubUi7m04AKMvYZD50Jg8D0WJ9OAqkniVzxsa6Ah6Zsm
ktvhIFQdHnub7X+fNMOiWW9BleSLMlMjqkfqS8gUVF3wEWPDrKC/YgPNrLFwcEDTm1FxHPsRPig2
wCQgQUI287B+C5ydEh69cgeTkE+DL8D7JOhAb4XFkJk5eAP6BDAJa7yhyURB/xS7WpcSK7nTb4cf
3tHEiguleMensHLR669rHH0+d7ccuJl+Ts8bpJMdcvr4KTBQp3VuxGxw62bPjDUn2PnnU4iIW/vD
A5IXmigEGaDKNSA+A4ttQwMdjeqQ6qqBk1YLlv6Vok3qW3SU8Y+24i3vtovSqIRbDotcO0NwF+8Y
OxHT6G5qO1cmhTF6sWpVnubgfVOjxnR695PhSCsu1JS/vsrqnPF4aS8wdi/rdZ4+zLeZc4PdvZ6w
DZI37euXP2Qexky6I/0KvYbCzwLWXBL4c+SWjSWLAZGA+h04RKWtHFL14hq2qkR5ckRtheTRdghv
VsCYWScdiD0n2TwdMXuSFKrZQKp38mN8GkacGh7qrEZ/NNcQ3Ujq9gZQ4FKvULmJqMPP5irw20yX
kGMWidSPGfthrM8Vhuu/Mh7Zr6/nQlhfdU2fufia/gJHYz5bfdLrkQY/BbTC/mdIGZ7+FALaKfIj
tv+oCz2QMOjMhq4LZk1rx+FKvNW4Na/OQrWAwlfNi3xa7UX4F58A7/EPg/jz/vc1XMsXhYq5I3mR
JWOais5K3IWo52SxsjUFFkOZva5aDQrM82TsiW/C7jkjO+ig0BgogGDKsIs4hJ9IYgjijBYzOyK7
CLbBZsyV5sAp1ympPfhga2xFj4/H1jdTScWCTQIQX2YmUAvjQi5hrZ9JtJjv9Of2cnYrGm2RBpkt
/+YspbxzNnMZTrnPNzDLuagwwqJj7TQ/xGzr5zWjkZKZJSLLDjAqcFGaqZmQ+5bOKVbhI6R+ThHn
dOtlkcEojdUg+iMtXJBmzVZmbariazD9HPMDw2+4oKU1q/BgFKRlfk77lWwIRp+3phDi2iE7HDUF
0HYjKI2E2K/EOljlHJSNNF7Es6PcvsilYGYC0d5p8G5+qvqvplbki79mxSPZMfnypNAeTdlj7CUG
6dXC//4Nrf92RQvpLTT9iGGALcqdxy/KXegif62v9LGa/fMAG5NfnuOTl2MUzRnw1kSDvRlVoD4N
rwsxUcvv0hncivZpDT6gtjqT6swn+YE9kx/QyHqFCIFHYVEsLYcuQ/5orB4BohI19ar9rScep708
0+ykP1zaWnvSitqPMxkp/8PhVTYOqnyKIuFpivf5qhRUL+5RD8rrUQjyUj7su5cngAdRNveQWV6t
rwTNu8AlNqQru8jG8JbxMzQXysuim1l2dw==
`pragma protect end_protected

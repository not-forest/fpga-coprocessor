// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
iBqND8KDb8HCtgTU1kpbNyH3n4iQhq9lnekQCZck8EzASsaIDO1fAeSMx06ZbU10ngSdYdxMxF9T
/kzBIXgGKbljGNnXztuGInamtbHUgG2N7W9LI6xULJBdyYo31oTwBDyAXP+rd5Qu7DTy89cxp1wq
PBfpjA078bBAVJfBr3819+vheri8NJ/9Qtsn9Gt5m0F+jb4lhztEcSGX6Y4oZictUbcH+ppjlsXh
Tbsihp8jlHXnsb+K8cFo9PQtCXOxYuMKWZkn0TLQLQt+IU26EhyPqoAg+OPoNB6NHR1/d/O9cOmS
BW+pE/aTAWqmb2eIwwEEllVMSTgQcITCrheJmw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 14368)
mGlFgqsZ/RQwcbG1UkxgMpSqEK/y+5ynHpVb8zfy2pdWo20oHU1OZXfG4dE+BA5cqEZ3NgeRpto0
iEYjpaKn6mUFRRFdu4ev88W7AfDCxKzR8acvANV6FhINXKzMMhKydqz3PxEeL2uYJrjE/7A3RWbw
LLNjyqeDzPxaR8oCLUfdpo2pokOtlA2FHfOMRukTy2SooegX+GCLqfrDW7pWgWLPUhBDXsb6vIMJ
CQOBg6hM6TL6piQnNFHgXSA6Et7uueO1C0EhxfVT7V6RzPW9QNihOKEyQs2GnADYjYYIvlmkv/bL
yk89+5Y5gMEXehxoHF2xdMdRHtmxsH2xhqOTRoPSJATq5PpzeGYYMQrunbOSeCsjt7pgDohNnbPI
f4lPq4/dG16RA27o8yaweH09rmBkPyirNnwrwXlMTKZnCUQfLHkqEktnaOE+0JDr7aAK687KFZPM
XDJFiBtOh4xMQPicF2vpF3QX8dC/yAwYzhFQWUXDfaDfK8Ld1FWhvgcD+PmrzYZhFIvaH+IAfQEQ
rSIschLPrpXN8D0z/syizqJDBWliOiIWMsBMRsaiyk/BBHgNVZWYDvPW4aiAhADWfXo1wu1MHiei
c8nHW4QquzRM5NH90OLc0/onz/9Rb91xrK5FN72pNz9m6mOVaKnwfDcsVKdCnBDfHJYoCA0FLBm3
fT8LdVwC7EvIq5QP1DOhkgN7QHkwH8P55Y0NHnu6lMPkGcvy7PN3dMcemOMSuDc5XtuKaABlEZBp
YK6aHU1XVOChUnCLacn6mY3oTApgc6DQaXr/qjfMJ6UbtxCf4nwQ8UhsIgXG5A2UAg+kYhdZBYxB
vJIb5whufxkt5FO6Jef+a+vh03JdHetuu0QNPODBl0yuH9Gu2YjtoKa7VfYQj6cDGMXQTqjLH+/W
yXTRjhMlcth1WUPqruKfQs525+ZxoASfGBIIhUm3WsqghkQvBJpqaCt5oonpr/vq8a1k5SUXEf2v
f9dERvdhYSwLC+Ir0YrHp7SJ1TZQWmywr6PR0FGNHrHb9X+ThFjpd5t6hcnPQhyuyc5Q+pG3I8sP
yprfTZUJQDvVZgZDEX5OKcKmuZyeev+po9tbbwMd34TnuPamx8v71RSBBK0mN3RovgHoMGk12mD/
LcS3QsU4cGc61w05WG//HxEjlbozFTmnVUQvmedgT1ipIxbEcf1/+bpMy0JpXaJtP88Us4Tq1WFk
m6dLr57593BZ0jw29J4r1MJLo2R2/6uu5i4M/Er4AXDeuY4Rg7WZLBrNaIVZ9pOagTA6TejI8x4Y
ycqAc/2433ekdnakVXXh5ybZgVnW2O9wxiLhm0zL2qs7xZdEiv6VAJ0jlMWWLKb1dlUSsZ/kicld
Fxwz5/uEzu/ADAoyjowDK7rNVceuR0L4BMsZAOle4cXFWHYJwgtEK7fHMaU8OO2LLdgi6fgl3UpW
A4aZrSiWIL3a+rWVuugsXqqKiJ8lXnJNN3a5fPusciED4r4tNeOPlnBxBfpdaXs/ZGUYTbxNLuHI
DPHTvZfNJsvpoox+RYP5qzr4EyzwpZ2ymVEzo34oSs3wnRXuwI8ppz7z0Ca5S8V3gAJegDwvAZkw
RfbN7OVQ6j39TDWE2g/jiZvw7AB7z5gMEMvi4Bqzd3122PMcWRL2OUDcOQB6PC7GeUjRxypFdWEk
6PhGEU8fagff7Z2nua51UWuYKyL1AmI85X63G+IZAELDLpUdwUTjdsuVf/tvBtHMjvnEf6vab36S
6hTtYPkdg+h5PYjJqR4I9j6quYPp6A2jJTS3j08815+gjhTRlhmb8poo7Z02oUz+YajsseAVa041
6CroTuPcYSielcUqgnKAcn5WycDoKNoj6mOtbMEBjHS7NAN6duu4iLLqcFLH4zfUmoxW/0SY/ovL
hOBqv/0YGaaHBhrXf2WdDgJ+s3lMM46AD5QNsj2cXdbydIYTR4RQg+xhBA23l4upOHYrc2SJeS3a
gE5djZx+FZ4aCAMoTuH7O+qgYWSvRYO/QzyQLmaNfVN3g40XZjrH952XQv5y8rwYrNxORzXHlAsj
KHXREoaFKYDJU4ywY+rotA2ZDaRpdEl5/7HVmc+nepDYKkVBsTJvsDldKVGzLmUq4UZER/1rbvJp
nXU5osWCH0KJlpQclLAl8ZVizlY8OE8ihKX62a0JqYhqlCnogPCvZ/gRyxSFOb3IYB7O547LFswP
c13GlbXyo+J3MfZ928KKxpkldyb5yyfJfIZ1UxmProepnT8AdF8OR8Cupkeoia4GsLQmew2vsgz5
4ny27R6mgzYhW27CnBjJXDagT88ItOpaDRJSjmRwatYLivFTFcCclU+0aUD+QPS1X4Rffo1/Qnkn
ofVVsP9WL6hdQPh8IOqAl35vy9Slttas2Wgnao5PA1AFJCH6sqzhgSvVA7aSGyoQU66bdSlE5Z23
1Zlu5to+aBnc1qGdpsdI0vZ6CzxofJrPQWygpXF+wkEEZHoNjL2luZGsN9xBu+FYhUf/KRJcSRd/
P//Zro4CyYIHqcgfP+TBCPueZX+ssNFhBYMT5N1OTRPykVVRjmvHX/AqUNfCT/2s7rCPPjC0axcw
2bApRbsedOQ93AJLOlx+lFf8la6JwtJLtkdnq3myR/9f/7UgF3MtiKK5Ks6IMd4CHvlG478Rb5p/
lxFJ0Fym5vSE5SSxmG1ovJH1zHO2Kpw7+inqz5K8sVfGvqxximv1KbstNLUZmimO/C37zAdRPKOL
UO/KIjPsfr+x8runYPwlnT0AzhFLdqX2E8zrHrmzJ4PDWVHwNlrJvOeu0P8SAwXYKfC4/1UEkB9l
fXGd5QBVD3NcB/8Jdgwjq4mE0Hv1WCIgMcqXq+GDqkIFt69l6/DM8VZPHlSvP3NIzolFNp9LujZ3
Ff3dpQR2Ndi6SQHgznKorhvgzxxgA6dEEz9Yma/zPHvP9b2d5KXG348R53cY7S0egKYxMAQ+T9Hn
x5Zz/9Duwwxady2+qsHy0QQ0D8OQab6j5szqFYtiODZDh7k3XqiuFbL0OVKPb5MuWuLfKb5MGViV
+XFeHawub0uV23X8JOGUop+Q0m6dlRbgRGdohVNrXeu4uDODOAbk4CxoLbgA7XyrAs0gHX01Yqpw
he4EJZMXuDTqji4zDcwCVxXrj7EtF+jb5Fhq406fLPqkZ/aBLTCOAL0tScgDpLXr/cd7uniMasH2
JH1Fn/+nM9cd/Qmt4olODJMFlkXS4+WzM23w0bdAvsPnYt1v5s68P+r4G0OznBYvZo1nAecTJAUr
r6N8rDZWQuNlA8RCHWf8JRaXSZPwbE5i+eIt8+MoK3qzKRzNaYxy7nbQy52UXgDlfYYg9kknS48D
OI/HBkNyxc3yJvFaDyF3vTqE+hSafdo3k3SELuC0Q87YV6RI0QpHnJNg37WdB1oPL2l/jtEOG40m
TYCWPFzwfRBNdLzN2u5Xu71ZSSEs4AYPKOtzL1joogT1vg4NKUl1piuc3eYGuycxOwyHYy9QQHyI
lW4XaNTprRDG5TsmUxzuhdEMWSEhSH1ggZex45MJ08+eKc2X0jM2LgThPAZGybPc6NI+s/3BiV0S
YLzvZEvuUaZKFbWLOypop9kO6tBF8wCcZFevm0ZIvCY0FSaZL3rJy/aAhkNsa/j7smLAdMHOr291
NTEoMzDq+qwzdg/e/rP+R9naak7/KRWaOohfQLsqPqAcTdeNCOyEhVbUn51mrYQ2Ov1ycPluY5lS
gJkwnO5+mg4EQaA1RHSTzXTMdVOzIlIjuHOz1dS851KD8tcpSgXJaL58HSsG8x+n3qdcwH5umPDK
9yILIaj/06kUEbgpPRBtlDMDJZts0KInmgm/qJKPdFbZzMkR5ohXN2WGsof6jJ+0KiwGgAftyZfM
XedFvNUoc0zm9NqZdHnPNsc/wIf90NvciNmaokMPONLtNDJzhM4m5znzK2APfjLuHYMHiDevAPMq
YNULat0m7qLDlHHxcIu+ZHjCNNOa9S5SyuIMiU400e7EoQPyo/h1qK7dFpw1Al1LR2rJha8LmAsz
LY3yIHyKBOgNsihTnuAXXlYXF9I1hBirfiI9/o/Pg/P7CDrMS6AnydTey30zp0B1yuWxvw1u/gwt
+yVgv61xp9YMBhLCZLzslpQHvqHaNHuJly2FQJ36wW99RE7wcHavtH+YAhJp1ekB3PVQ7LQ0Lryx
SyA2QwMl56F+qW7IhyJJqyMrI699nOR3JJgexqNojm0mft56YmsKRRJkYM8IIuY9G6kVpDcUqgUD
mRa6LVo9tHgsDMin9LtTz7ERhqUCl1HMmcpXkYfSMdni+4Gle8X4HM04tFCLV8GIY7lkQppPdkGB
ALd+3m+tb8ns5ozD6nTocbBRx1f5GhaCKb54S4wqt/MAWEwidpvL8Jp5TYFQwrKoSnenPsK0B+sV
ELEI1GGbcITF5n6dpSDBtDm6gmKD7QxeQMxCGQBhiRhP5r8saSFXR7V/3D1ITFlxFI+7YQk3Ep+r
PoMw4k44N0aSUpFoX7pjKqIc/QDVJifE8bNdBnd4rGmU9+Gn24HMLmtjQ7SNckk85om9DoVIK8P1
mWzj3kvcTy6I/5Yzx0FOufB4FUNSU1DnQE4PzzmUaYy4qrZdf89PjCDJu0WqiryoawtkghISVc4U
LTA1AaVmIl4MhYYVEtejwc+n3tCi/qTIAIfL8PHIIKRjOlZf9VuJJqMlBTked+ehH/Y0Rr7o9Ac9
0cE3vnDXd9k1J97uycj6RZVHpgSWzGXNCKvm7lEeQY86TvAAetKibhbxoqkHHsWI9PvZhCatWaq2
fqTej5mIoIlvim2QwFAARXpI+m5wJRpXugZDh6wfZCnaMdk+tG0CWWL1gUg1KUIIJ1tJfT26nwO1
srZ+vTchN/+eTGX9Fc/TiD6fpnUecyxQH0YAoYqZaiQaf34ij4vCYk4jz/fPn+MSo3fbhPC8MiLH
ydps6FifG3D+YZGegIOZd9k6Vxzj6LYPTpxNM2hQ7JafljevT3hnuduj/wnKebwwpkcQ9Zg4uB6B
JOnYtIdNMoyhNXtU9u+/x4tOUelo5DU2HjNszVuMO2OMBLuo21jc+nmis9rBfysip2ha877lgZTn
eh/M2UmEImnp+EkgbxIF5U8armboRl9sNmCrnbYFRId2TwRrMjJUFeNsObmeW6VyRVEQRK7l7xB9
QmNBMPsdtnon9V2Bey2KYNEavnLHdUsdULcqSf0oZolEBcy5+1litBjT3PxZWzXKJyf8yRjYhUDq
AU3C9BmZ5d7nWFJDWNbmPoUjfuIEVYgn5VOA/sQdwfq2uon++tsLE9a+uFad8C1vp7/sBbrtTotX
Nfl5Qn7RE511XGKjgipcwBp8ppnoYeBGXwIOV9sx5n/Ft4kFEVVdMfrWHHjOkd0xCuK4YgUPtwew
00SiweP0HFxyWz3sEcgEA5ML7CZibh8NOaYFr66pkkhNHDfkFxjRWLPFixRWilTW4XLvTebpE3l+
IVOmnWTSQBZhFJ1zAk+g7QVm2XM93wnf5yMw4P6ItG8j25G0NHTIYQ8FQUL+q1Tt+ZClRZBpW0sJ
iFBIC3LtXJRMY861zzwfYFvGRIzPVSU/vvi/GUrk7cTSwjlEPmaX/Z2tAa2zVQs68+D3py6XiS1A
412LeFMwm2D5A9stey5nDm+ICI6BTBjOS0YsxY9N13+XZNi84L2KEOLQIR5UWNbMuP6Ix4agO9Wk
SBUJ+VYHYU1WkOWz4CtVEbURie8XcnMpQiuOAHqSOXl8gUozE5DGvSYmGObVJvKHm69Ffj/lM4qZ
waiqeD34gACBZjRRnSXxtQRXhbLv3kht/O+uJbDv4H6dOEQy9gKu/1iEUN3221eM19i4g6FYAGxR
kDg3m9qYZ/SmU5MHtLCQtDk6WlfdqaA0VUUdLiI1qzPbtr1KXMCFcuvQ0UsZIC7XS0EMAAQWBq1b
HioqDi6kXc6AkFY5ypQinfhiEMuNTcvrG3fwHtUQVCZtx9SOBF0ct9DCsiSnSkgEz7W58GpymbwN
Ztk9ZxofbqWnyGzwAz3cNhv6V4oTK7Rj+7ovu7mNOl7eRsy8hEJoHCwGVLLLbiN9b33DfIcxm8/d
zmTDS+2/S9Yug9e9+bdTf/ZYzvQDreNbx1F02OLQJliF0GqLc9LW1IFFVT3oEB8ijOpUayE4yitU
J4jf4AIeikbjy/7H/CwdLyg482rGOJBVie75MfbZ2oCqeRxm+yBBs9rthEjWkN0gaQlTSlp8+foP
91+vDn7ltg+Zq3JcHdHbey+IXlexQvS+yLIYC83O73rwP7paT7fFLi1NkjPaSgiiUuKjac4ENbvH
60zxIJTqtE02y4TZccCbIf8FcX3UC3hfhouyldZCwyy5DjWponDzQ13w0ZfSRp86mcc45jZp0dH/
An0GlXJbS1FjfwntPkrg6QypKZOnHAMsZl/BC5dLJJXxjgPBXxrphf9YuV6XA40pZ4FHwk3qn/Vr
PQ9sq2G6avlKiMBo8yLIC/z5WBxroeoZWDiY8jW2d6ozWVnAkWY+4bZqGKo8jY41iPGqhQLX0spd
E0XrDb5gVRZiSDdM379w0VI6NAlmPxKY+jNsMMb6qzezPoKK38V7soOL3nRfu5tARbzgrGCkvcYy
Fy0Nyw4PlXCUwMMKn8FOau/+/rA6jDlOLcyaNvftmGqKYRBeJfQeofvPBMPHHDP1eoLxxSY7vJCF
CEuuEo8RdYumubup+D7TOYkWms8sDGcOXC2WoWEI+q8FHSJJQXvs/O9VGkH0U1dbxVBY/l4vY92L
IQbWXTaNvrKznRNgjSHJRc9ZJh4MwVPLp0LbMIermpWIA0ebUdN87oWYSnw2ku1hPwNV0RVHovYD
/fGkp9Wd4zlDPohktZmVVsjPlmaniL7j3KGlmEfMCgbG7WJRn+Ph4AYoFYkWSAHy7/IsNmkg27g/
acfRicvOFg5Lorc3eOu1Crp9P5YEVQyf+IjmUPnLl5o94UctlX4agyng77MY4Hb7UR1AAKK4ot3N
KE1PpnMW0ZNmzawxozLZW7byaAwh046fCCUnlQIB6jcdQryTAv0ocIFCj9MhexQ3uZVsz01TwTJ9
uuWPlu3uDaDSQr5YbRyy9OokZ3KjCvJdTkD8xbqpY8cZhREhi2mNtP8e+pSXMZLdE70CZHDAfqIZ
yHdLUrE6l2N3Qln9UDjBCIkCdK5JziQX1j/lVhBVLSoDx6L95C19IS68zZ4VPJ/iXjNIIg2yRsyH
UNR+K2H301271I5N2JJKV5gZU7WnSe2y8ewF9Zr0W3H5Eir7oSiz4lJI8F7Dr3zuEnkEwkfH94QC
qSEowVJ3cJthpwTnOjDCQPj3MqViD481oKyoxWTKIosN+z5sK0/A1X1Fe83HDTaQZvrUMTdnzC0u
4vIhp4irZMAG9idX8Vrkuk514eSBQbUmGjIvyHaIEF1U6i/xHhgrhVQevuqVKqsWYJ3f0be2ZrDf
w6mxMcK4+aYzY9SmwZO1zzfW8+QXvP+p+ZzuT2CEZCxxyqyvb4iEr/vXEX8af4jRvDvTbXzlMbRH
ntO86ZIITBZlONrIQRWpwILjC1MaGNfvYwl0nS5BG63qknErXNwn/9ff6JAy5f0wz2ZAp1Jm/8kX
yo1KMMW7xNqMzwjHCEMTIjEee61ypsBCeSIy7ay1WjaRKvqyFn+NEUxvyqk4WXzEMMDZYQ8JToiM
/SfMdyVtU/xg9KLeGXQ/TujuFLPwYvs0hBOaGErrhk5nvgIv/rmDnV+w8FZjnRsCgd7p6PVG5DKa
KX2/csb7haC4xxB2n0uG9+WdYuLlAdulw0ZK4gHOUB0MDGltQYqvh4SHayZEWnQ6yKMzXct8o5wA
VnpSddYsk+OGG+AoNEdsdlLz8rdY25XX6cLMo49h8b+QEuYUgb4t3yfwfItFHlZ7VDQR7HcDnocm
cdh2EbFfvu/awT6Q1cs/u6KyJmTdQajHFZxBMkjYU8FOyhFSl2w1cNRDmYfhWlT6BpS8KYTdneFy
ZAWP5sUbttaqfYFRVJOfoo9A0SvWd8AA9Hz/h6rMyuW2/8vhNeb22fFhSPrAuidyANT4w9IDSZtQ
8NXSqIHdouSaIpXagQradNgJCKAdayjrptmEMCb0KqEQXbA23LfOALtH0twAnA2awWkkSwNtpBxM
dvINW+MO7VlrQ/PNkZ6zgEVxewwtbYrXHK5tzCejlmN7bNo+GaK5vXbVrsI7KatXfC9wUMQAl05t
5lrfhDzi5NNFDytJp7z22bfvvR9BVMGm8lGC4rz29Bg7Z+oBibXNBJ4orl498cwl2zCSm+Ga1zVh
T5AF6WCbZ1pc8YswET04ejYEZxgTHrnR+w/OH0LxxpmncMLk9sDDacLemluUIv85xtByDsCkgCNG
jMTgVqOpC3o7SVjnrbuD1+bhCNaaashZxsUOHdKjSttCw3sXBGz8W+RD1EZWUDJqH4zzvU2odHzx
791LeNMjiYh6NceVVkREnS/KLbtesUXqHfeeCqgxk8eshIAE4Gugge2G5NDNY5rS1anE7PiW5NLf
B+esh3uidlV7INa1RxUia5MCvLOW+qRYXNMUq+Xo13vaAEpNbk3AD3IEG/zGsqMkEpiIZ+MjDVfY
0rXAPyTtuVsU+puqyI0P0EuD3xx6LDC9sJTOmt+ialVitFHy7vYrQMBpAdxjt/TbwETyFPFNhd4r
kxRYFEf519YPN9BncEasRrQJS9SV0ynzkVYgxH52CJqaSg9zNbEtg3AsdDz4CCXogxvKZ684lizs
MrhMzyjV47Oa8ZuV+4W2iJV8oZBIcQixieBGFoZtmjbtvF+16cXTn7G8duCj9HCalBhIzCV1gMkV
xkRv3wkv36gffvfN2XpyAEBIa/lYzfp74U8jLh1TTUbc0emQP8oJgyVmzC3P6cYLi/y5DwcMx2gX
q9wMQdEM25vRXb8s3x3dl1kwn3lh4/DXxDcex2//1aiECvv4IjRbf6UAOmSRzJ34QT6K9RLprHgX
hqvb3W22BFnXF/UH4Cy2eCMR30xvfopT1GvVpX1B9vhrlG7sXQQ6SJVAtYh2PCEwCn3k3EgPUmCp
i/LTfxbyfZ0vxM4St+rqhYMon1AsekJ90fDNRrfWnGvsKXNwrKAHNvUIkvBAVRRkAbL+JTABURcA
V8ngK3VyueJnxM365CqW0PjWU2954vR9au/vQz2wnyjRCHT5IX0Re4QPM4yOYaArN5BVg+YZgJWY
/125fIv0gbWkGf+XddI/9GkX3e+pt0PK/gDcDhKi4nfWPJCFemoCHwpOKzT55nv4qTZ5Nnf2TuCK
npj1ZRvssTpbAFVOaq2Eg8bpJY4rdFh8s8MQLGldR1KAgcY0N8hm5s9kwkcae9IgSjEBS7P3c8Xo
io8gTDNZXE4ufMU/vP7JaaeUFCasiWWCDSk0UL4vMxD2SVrw1QBbSkSSHudPco7WEEXjtnFliRwF
PIC/zNDela/52oLGgBhVGbcMGFFOTquPoVYwYVFpnLxSzdIabF/4BkDDBGISBHcm2MbPWSmbxuuN
1tjHR7qScQJnmeFLbL5uj05M3gkJgvlzbhMB75eZo+DLcRD/cO+0CXXoxJqmfzFq6Xr2CJ5EMfwZ
w0ftxaGw88C0rQyRMkOGD3RVcXBk7quk00G23ttZMUzC8uAhtmq617onausK3NoKUA6jGakomM0H
LqIIolQYWwLqENc+Moig4zK9tmYHZLC/EKWpm9MUW/TnlhfbQwrmAHi6u76R1F8u05g0GM4gMo1+
gjVP4GoRXuV+ufegUtyUOiEyupmi8PAPj9QGIR4A7lHH3UKIJ6jd2n1TPYQC5CdXRzLgMBNCJ9gg
/sXOWS9cd8oxD5VGHvy0TjoYszaUZm/nqLMTciiKsX0m6Y2WlovlSW35k/98xwzCQPMVYO7O3rOV
3bNKB9oa/QWNcZCCTDKyqV0WfKjhl6O0gIVR9EhFzYGR0d88Nw73Wac/FC+K/EbTcxuvaJuJcwpU
YDnqdWNu9KQHGwX2CQ8lfLxqfMms0NsyR4cxBkWwsDAI/4Dg3Td8TUn9jzONSkStxAY3tVZOHnm9
2wWPE1ZfdaLN5fW98aCvDiuG9Ll6M0Ek2RM4L+q1zKIIkJod+jHaAzb4KIf5EkLsTF+NYVAJEV7A
b0+OEAcbvJh2TIH4yHipeuc7AHwzV1efhiYfND/+82qI2KOX3Vkwz2cKRwbgvRHT6uCn2Fi+9yQT
YupI5jxNJ4dXz/kLE9w1p5D5s1d/rS/8DXYzuNwnOU6GSFD9zufp34RGiUwKPRp93QZitmT+e+JK
nvD6WcK74CKLfymNE6s8/wjbCB7H3OoQaA5+VB2dT0YeGgJ0hop3G0fUooMLkIGDh02k4LZPt5mH
Nb7DI1Tltpxo4uHbomAPRrq8HIXGMLdfhufNRKKyBa/UN55w17LnbQFkj94E5dExDl7IxUgULQ8E
T1GNJrh3iph5X3bemcC92ulbKW54FXBBOcfNvHFGUf9SWmvLz21HZVfkKJ5feAA+0vy4Ucapadb7
x1rimg1RZJ28tojJMqDCzB8sW7odtS7+DGny6IENVQRDRSmhPxucC+8TGCwSDFMd7YrAH2G7Z+p6
SUvOeK9gH8XpCc6nn9PgxOzVHWfsxDEaVlMa+yOXdX2Wfko3RSnas86fVClwe/at5dhOrarDRBIz
R8ClRnCuMXBaSf5J//KdgcPjSJNaJuooWBjfWMJIKEk3HGt0k7UgfOw0Db6oAxlVjgB3q5c22NON
o5djh8XgzrH8APYglXm11ysYi4RuFxsdNOhtz904aPSxzrcACi470iS+oCEO97rVZCMWosqwDeCs
lZRX24bv5FPkhNjRGD2i4dkLQqxmGaGDwCa1pf4YEo1F9Si1lDqYVBEwRYjGy6lTyBXRFhrwT+tZ
Fw3+LgqIt2xFSCM/uc/WenP8mPOjhtQVxPSRUEdsfhi1v8+j7nxA9KR4TKtXHcq8M8Ni2F+qtDsH
NlDlYuksCwEvNWe3/xpLPb3F6vmkYa+JT1lwKU9VbOp62y5zNc8mZ8/b4UUUMquYEQJFJ0jqwFYq
4KSO3IO6gGjL9JBxjIo9cTQyjUXcF0PSv+jY6qPXstkEDVAoA+M+zDHR+8bPb3eAmeAwoBxTNMAj
wyU750LGHzLx6UsMZ8CQXq4ypdpuNd4ytgOB664U4kHGGCqbz/y5PCZG6SfMdE6R/lOzqy1FPTUu
WNj+0OZIOt9gRZml7fYAXSGEwixXjgn8fULT23bpVsUmHsPAFb3lvyXShHayUMpptOsmtHI9l9H4
3XDkaPvXZJKvGBQDWBKBxRi+SYt6aVoChAkTHVtgqBCy717qrJCKnmOkNUDv3PUScjnVdBEdM+Mt
I3ueJVWY3tErdf2bRDpGqKwfT7/T1WNzaA8jBA27QXdnLJFxRWmLeeHY8KkRDAbPnPgE3qsoD16B
tcdyHTlMSi8c7dW0GvLHDGKb0HPWsG6q6tuaOuX4kX0W/eIe29u9meNpetEkDW2UuSfRRH4/TF5i
zUpqp2XOr3RLRNSNmR71KuvqE09VgypXGjh/E17WVwaEXvkzjxRp7YaUXuiIXvaZqVy8o3D7YcqR
iU9MNfDcukmqezTE9ffTTEbzyCG/Ip0B3ShKelEzhLnaRcPwvSb0Y3L+j1+kR4yrjbvF97FQLg6N
FV60DGkdaLz7351Qcws2v0IAnRgT4wgbf4fns4X2XZRzF7/hl2eAlBHJ203rsbCu52YkcEA7jRyv
t0O8eNzo5BmusucEd8PNmZwiwOJRvpds1hU1So9Da3fhmCaV2NQVS4elpXymQDiIFqwsvfIzqsAe
Y6XxsCOB1P4Lp62FoEhme+tMxjio4Y0MbEuP3gh4ieoB0P+zhUpnyKMGH7H5SmEXSstpOIbwQ7iv
LUfXLM5hP3HOWYR5xy3fsEXPB0mm51yONfh8uqISefOtSMZlPgw7KjZCXT6vH5nJaJmee+ZtxJi1
0XzVitG6jyWgLJLLiQV8KH1veTE52Fo8jA7ljU7LazMRnf3lq62J2uaKLWzi9SCoiq64OfQc6UX/
pPQRwTtrCZVl1BKQ3Jusy0zO8LpITlW0tLqXrrFRTLMlO/OuwpxxXX+S9/iRSF41k6/qUnl9gFc7
43RGx2ymbemgAejdrYI0dz476aAlQ5S9QYlehhB1LGBzr2skz+beQz3ZIq1vgAsrvuWC8axLRYHo
QgXeQ17Oa/gBMKQmkENa7ahl/SZ8xGw+q/Z/jWoH+4EIy9f63IAXjj+WaxBrXr0aLy/11c4rKkH9
UkeFbmXEuZLmKdTj/w/f/y3J9Usm1sfCg1L258d7tDWEgONhf5pBHXcOBl/5HP0DYP9kh+8+AN8N
BLqJXkIE9T7JzqIWJJACB493G0uLxw9L9cVxXvtGzRF1VHNs6cybBfGyynolbpUraKNxVSv5RWQX
T4+7AN1OK4EG28ZX1crpS97HEg8vZyl45uFDeUatzCIoKV5zC5Nke/aN2kwNS9tECETIyaYNOefd
w8cUltHPIwnPtMekizgzU85ZJnm3NEDzBTG7rHoa+LDVTjWw7wRoAnJEFCQsjYDjHf4lAzpIegZU
P4SM1KvndC4jQ+HMK7D4cIooGuGEHaOiq/hYluiocqHT4uD8DrEV4U4e5Pj+lKEpU6AP7USTMt9c
egaF8vsmxrolUw9s+qefSBbrqQ4vdYUExlot3QWi/WtEO0xoJY5NHljez9GYzIVJbfNag9mLxHZd
jgOtyRrdAQMJ+L7VDP38epNB85aPcbHajEjBY7/az/KWohcTHh/QVG+nXWPtvG+XMwfwgrqQXHoY
ecq7ToCoWWU5mCin60hDNMg06ogEf2zwVVoz6cXN3OZA+h+zqU5GZpuiJBu8+rTkXyiBC9t3Vygq
45BbTH+LTrz2QtmZF745NfOGiuUGcSfj61mW1/KHfKcSVjvzcHuJ8yC+tvzBRBafzWctLeL474xJ
AIjGRkctSReeQe2jTQuijAniqtjT1VcTzCVwbEFa2yOL8LiTTr1wtXLvb1FVAnIMSge3dSeGSNi5
EWC5IGnWcFcyJUtqqS/DXXEZbFM9uEImb1I4IC2yX+XuL3Cj4Qo1qprg87jIdi5jrKIR32zpm1Rw
o6BIFACTL8xCYE/9zRS1xyifsb7C7nJB3V8v9NpzkCtoQHS9g1ozHwe0vPfb977kWvqJJACnxM21
OB+x11V7fy/e/TQ1uDo5TLqFuLJZaevo6i0gaiThfZ7YnhKGfeY2J8ouZIQB8Ny5LtV0iLXJdQG5
1wDRsNNi+4MHDllP6yheogHtPG5MY5v6hbZnFVSbffr5b0QD6N+OAanfwpGChLgG2ySXzQk8otg8
bucLDihbHjSznZZOH8dgviisEuoHTUF9B7RO1bQ7TskJvceV4PQRYNdsbySdnEZ/FxDKOB4Uv6I5
z19UkCQba5vk2Pd15uGKoaSkUVvJ0OufxXSHs2ZR85v9PjUXficlgV5bIM1vq7A9yyD2H9X0y36a
h4/vN+dBiOY9QUBgo0yLU+Iv3PW49a1u36hBJxEkopwfZeQ09PQhsbfd6WdcWsS2wnSHR6ufyWFO
I32tT3cHXljH7mo6gcAJyHR8FkPw+xpHXutyG4WbYy40JAKzEiKmtXX+8jbRzkyjEwiUxqtFQrQu
mp/AbZx0+KH3+JFNYMVz7OZtkny6dhOe9xg6ek3vr1ZBZUwpMvJ/iM/xV3OTaigSay9HSGp+LYLm
RLexOUIzsjwMIWQbrMCaMOS4pVnxGgRvbj5gQEV8nxk59hW/MzVLsNL30VbZC3y1CTUU7Au6908F
gUU6Q5FPDne4DFCRybghOue9nK3Fxo/RVXVUbfXBuOKb4R3SIculDZb3XXhbA3eSHfQn6+VpNPG/
rpcLebPU0h0l6wH0qzZkO8f0V28QBZTYfmTgu+oTlpIINtkX/FmM0Cjja0SEOwfTLHOmpc+QTtGF
5WWoRfOFYKpWE6H2RS5LW1AAxjNigUO0w7tf7cpRDO2Y4yOXZ1wLj9Z69kFjn/2/8V1K40yfMsNI
Iqxo5ED6HozZ30/qmoll28nsQhtgUA/yGHn6wOeNI/jQGGr51Im/wVjw9UNR8JKUHEMoKSZgnJYG
ISqFkW9bw9Y8O/tnB9emuG6nkKBHahStwJFpo3DzaGHj1BMWa9zopj6R0fN8ttFgU26tU6DzqnNJ
YRdt+3nySKPnjJbvd28pubfOFPbLPKasXbKohWStPkjGD9Klp3IHVUo7Xrxy7hjuKTiyOYDFSrHd
9kMRJB5HTN4LhxiNtW4GYrK/bdEybxxcmkA0/QVNGRxixRnEwCtlv0R81goYjXNvQiAv6Chgz8qj
LlJcO14XooHC/VJN+I3unhD7595KbGq9vfbG+JsHRuzlGloA8ligRWmHw0AW55hDwUxHXoy7sdu/
iEk2jpO116jixMrod1lkF40FIi7E2jFTfCuaGNMfYkHZMc5/BHy2NhHGShQ8UWe7Kr4Lbd7EaLOD
TTKSdRBzr6tFCw0kH09RVqgYr9Hwc2BjrPldbeHYFXiI3iFDaIJmP8HN2hFfrG9Ya44WPZeBGopY
ZO2oFV43d1lUKN2gsUd1Kf4dfwbn3bxmnp+e28tCjkNQr5FKHkWoEz1xikZid/Qm/mnTVIJq4u4T
3nHIEy/SlLG3DquHSdbucL5d0CbwaZeCvtf7kBDqLt1R6v6SWJEG0UsnoL7uMnsJ6e0VFkYWKWO9
pYuf+wbsAhI7kAdzwrXuTciizoPq4EHYrx0yRlEECH5+FFqUDdkojNRnHErpQxFCrwf17pRnSaLw
bUvjZlJEUAuO0Ro7YLCHo2ysBQCUWEZsm/ZFImfShnLJfTjffuNQE93ewkF1bMPulkWkvabgPn7U
PLt3JaFipP2F2c6Zw3ePir/jybSPhnc/lo766pwVdLJzbbwhR62cSs5ie8Hq58xmhCfaUTWMS5fZ
ZQkLJ02Glh/bZv+9Ib7gt7JSn8hL/7LsSyU0R9SU+V0rsnABysY1R25Tsm2Q/7L/KAeYJZZOv1Fq
hTbw4sD6sZZkHXqikPuJTrHwBL0WgQc75+s/avDU1n/8eKmu2LoetdUhKovxCgF+b3z4m6KFj5t2
HiX3P58CE7GEef5cS2DkIyxfSpM+vvhkgPMnBtcG05yO2SNl1L+Dg0395xOqMx/wSClrXsZzyvRq
ok3ORJM7PFR4TxRK/jef1tjeAiHsTLPqU0oRnoMIghFRgC7i4hx4hLRwDfGMIdCBA5RU/Pi+KBZm
pXAS8uoP+1bL8Zx69tpMc7Ns3u929skvC4XEfyBn80SHoFENF1+p4I3OUFvzpyYfxkOYlzLEBKGK
kAP+jZTd5kIane14Xb21VOyYmIQe9dtW1ooGrqVxn3em5KajsQy/5U4KC7INLP1AQjGiSTB3w6J3
PVuO3/fF1pn9L9TX27bAAxGsaOIs7MEXGBeyB6UMB+7azC9bhMnWgxk2fcE5np/D43JPtnGuFNhF
BcklZYhHlEd0jsuA2EWVTIX+gRs11+iR+F5iab2QvC2KHCnJGlClaw04wQyBkDiK4+QaohPyMsa3
jJwijRx0KJb8iez1xzNauwcvg2tg6QteCy1oN1DO7szuRI5+q0nGV16aMYwqkt2hfe1fjDSsQaQt
Gb6cEj3Y1YTMxPXsUPcylfpsOreUkaI43JZuIpmG/8Qjpgp6YxzAiSnxTSxFWG5eVDv9XONv2VxV
uURlxhITfbXrHYJLIKFhCUAmAiHtbC4InDS+Gq0bmdWHEi5QH2yizAUA7UrKolg/Alv4tcuJviNS
wAS7L/Cl6M/MVi9+Otz8RJ41nTY5TQ3nfUqgD/LDNiGSQgCDPUS0d1o2GxSi04CkailCDiJHiEk4
UHkbNA++Sf4HlLmiBzNYP9sFNOuxHbnD8Nco/lp4U4RFHmWAnzWDGnfErDvuVlVzTUszyeu5C+5k
AmCJgS6RPk8qnRrwPFh9Z6UZkhmUoZT+zJCj4jpXPcK+b5jaYS/WrZJvgVcVfOCwci7ZZgyxMZzL
Ss15HVB5PcKSChIweXJS+smJbEEpx/ujxy6P0tXKA9XeAjkkhYQxnIsQEdYKwnik02PgXdXCgWne
RFr7neEBjZXMs3H0KH81yRb/LugNter8ctWFMsKWlIBA95nrvGGkZktKVcQjzNqKjXFMd1N043GK
UlMg0jzmUICxIlpSeUJVhr42ZQfdeIKEntaolLjguzGQOO+pS/DdB4mFFbN/nu6/hshXkLb0rqXd
Um+50tZmNFx8mkNwuysYX90DvFevWGt9gZYgP4RbmIMeSenMpqsEudeN/dDHAD4UeaPDSTaHa4iF
bOYUOLvB1OC9OJpouKI6n9aynSgQiIWPboUnSyN2U4gNKaFQUJ1RpA91vbR/PtkY1PE2D0ZBZy6W
YWMIRe85yVeu9byCqyRuwAwc1zHVAGGo5aY+AE99kajubAXvxkJalqnOliCrfXZgtPZXjo9qLBeb
HRxc3XyQEBB8iDkc2RiAvx7B9nVrOnqABlleOO7gaSOdR5TdzZaHa631Evu6QYrmu/9eGbQFw6em
e5qG8rgzjoajNWkYG/zHJR0FDYYFMf8ikOk9SrUM3yWr/jY/a31Kw/csQIyIc0Dfjv2vMyfm9Kqa
xicy7owRfBScSw6xL1T+t9HpPxqmldNiL5QBvAsAMAHDnU07npJx0WRctE92u2NxCJhrBguV84N6
I/UnIHAj98Z1ZP1V86WKWDUXvcmsdqvm2dr2njXgJqrZdnh6nhMYI7t84v6nSnRnhuNhRYXoZJ+6
uUv7ev08g9ljALe5ewTOSeyVJNEeKBFFWfQJ1ZUI+bViJbk4bmswbjfGfyXmM26Gf9HncmMcgJvp
ROo4nJ3I3fSY3rqzuVnGTjocpyG3RwI7kyfly/4sHCQTjTUGDR+2glnp9EISHus2NL/g8UIkKftR
NKlC0gx1/HGxxPbyIzDzDPVwKmV4gc7vrGEOQGN5kL+FSHGG+RtVH5tmh67thvYlAbxamKEJjrSX
LBWE2kAIwHyhXWiDOtV3YK42Z5fbhxdxxzXsau6CvJkb3DFHOBuJ5vsqdayk7BZHeXHlf8qk9UT2
Q6NMBOKcWHqtVHM4sAK6hUyEgarOwdYbYWUf+klc34k2l4743I6vtWKyE8Ani95gVIR/AOTEg5UE
qA8qHSWp9D6F484quAxTDCbJlXwqup1hk+6ZS9cuv84MlKoRPsr7sEsQoiAW5+rZNHiCUHspJ5kZ
XI5uAQG464leuDruJGkjfU35U8DQpjieZ8etZyCCKx6ASw+Y8pNWuWqFhbTlOgbqZrLfvo/ys5jm
n1NRYVBRaAuG+uXOk3zRPgld+P6D7QmxmdjO7tq/IhZppBmhe7UggTD18Q4VVWLoSIkS3fEYNZkz
35NgP2mNLfg6jwT/iYKT4QaCL56+PETcJ0qWi8L6HiTFTQpOxfE59VA0adl5UK+Bjbr1wrKLtXHQ
T2for9/qtjTjvlDenQPWwXGeIO76LxGkX0F11FqgKQTRV3LTUwylR/N9KdTuE0vrLo85pOEFdyFw
x3U3POZP8G67ZjFn8hFdTCAaeKRmlHjBqFLLzvTGUlsZf1mITEKYMMIKfgYHVWIA54VM28NUHiWh
+dF+WOuvIYgvR5sHusNvJLsPs6IEre1vxZWQWf3WJSUMA7YLfWxhmSceHT9NiTYXIz9Jf/JaJCNA
7O7SKvDrn77EoH7gzC12wHCqI+PjJUDdQbC/sCiGu3dOh2buwsZnRfiO/VmF4G/PzP+kHhN37iZx
nUgJTEButg83ZLveJxocKUqigNx4EVYAfqHwTjd546lfAd47bpkFlZ6+DkZoD+JHMQvpPFV7hO6k
qSJw5l50sk8vV6Qk3DiCe8Qks25GPxc8ZJKaKE0/8FnOG+OXGHFzBYrkYtLSvrLBbF83I+ppgprM
pFjkf5KtyjZqdmghwH6UrmTmgIFv9KdUzMTLb7gaHkRAqmWR2NCuUoZidXHk6fCMPbHmSTZhJR4i
V5D1CXm8rUE2xezyt3RNFad5kaNfQQKvlwidraoIYKQMp6SVAvFBHKLnhK+v+q7cUFhNJiF413b4
XfPaUgSDeik/WtsJqKYRpqn8gM8LHpCCa9DuCIYCQ6N9zE5gnNEnH7HY1l15QAVeY61ZHg2OUdmI
TJOmT0XnyBiCxe9q2X7FZz+CcHCD7tv27d8oQsd0/7v4yJeF9MbAxC/JuJ3+XFlo/pmE7r4BAX0X
sUiXvvJ44WY3y/kvauDCoEIUtfdgGZQSZ7CFQtyh2giDY8iTAURDPM1MO2IXfjX5utYxtJwt00tU
EBd3NAUz5MUWSIhb6rTAPO4TM/mPSdwZQfQZV21YhjzZuYOKDceouDzGXPZlpY7sjRPPCG2oFYPy
uVyw+jHBB2CgsF5ZtmPXQg9xmAgRcSkytDBcx3iYNdWcEqFqTdXLNTY+PHZZhSlpvzUPkb3m7H5J
dnruIHuFaxmFT/s8OH0Fauyw3lC6W9YQ5y+VMCI6pGXMLLAHJVhvFOK1GqsUlmkPyh+E4Ygc1SLZ
J+2eC6VW8cJNewE+ydrefeUK7lA+S6qCqoKmk4q+KKmlFfOxV7uEQ5kgLrCj+oCQTx0R2mGP9UDB
LJ8Qsrblsmd1d6tsVQwzSkUGT+hVjTzqix4sk5j0GaEbsZqDetRpr6kDvVonCJQkliWM1KhWlg2B
J1ZitVALjFWys/671MvfjBTs6JxiHaQKsAvIHYW33fKnG696DUwXZ6whtIkkz/6mBQw17hRDnE7K
J9WP3e9RKQKBiNpFED2983bWphO3M44J+9fA1lTESroPGRc9+AMscI8RUN9Zr2ASICDUmOp9c64J
5ZWGOliGE7DEtgoqVS1oagVzwdEFUNlHvJEsrv4xu/TaFA/x2tz73Tv8Qh5Ewsp/Tev6cGmnxMVu
IgQ94tdKmJzyEogVpzhkPusy+jnGV8Xq4DnbT4+zwwe+tTWBSTHVlLMdsXNQ2htgvZoqcApBeM5m
+RciQRlxPDagDFQEsPLBlvP4YDFnHUMm98vQKAmRgTias1Kq7kHqC6HUEkM78UZTU649gpmLAj4X
EAOCn7J2CFHyPdnrWVndpYyOGtTO7pTmW9+2W/3GnqZUViPhEbKWyKVaOWmuefrzVos4oBGXYSFC
9Qk2RetetfG6+7tXtBiJIWGQ3oerVDC/ceOYYTqKL8idgGpTH3o51zyUydABLzRv4uJrPRKhLtLO
gHd2gQ==
`pragma protect end_protected

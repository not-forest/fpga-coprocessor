`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EttlWDWCVduveSOkFVBBhQ5cptVzOv9ItB4Csj/Se44buceZMu9wHQHCjlxOw1X0
GZJV5ceWoP7hcgwXmiTS+IbQdcWT7yjislsHJwymkRgJc3ZQqiRNU8NJb0wLAH2C
FDmkOiY0uH30hZHq2nYHM4W/OR7BCQaMXqRVc3jMOqY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3184)
EspkQMfUJHIg+56/x9MgwIycGZtxRI3YI5dAKe+CbnpmUYycA1+SOOXLmKMzeeMf
x81VNyE36jdDNrjirENBe8+m+zU6/iCgH7HL1qAFDpATowH7ojiH41i+QO0Im8UI
SF5t8HtIcJk1MScQx3b3Wxn+eKSeig5Ml6KOfegu0n7Efo2M6liZmsUpCydWlMYb
gnxndF/E2xfJbDoT7YEdBRrNxQiZc4yHLiV9sj04yDoctQIiQ9NMLrZPpXVmGbpw
wccQnE1iXGsu0atVeO5cJMi9jwKUPSLCJNT3WjdclHYenxZ1ZKx6y3pjPUW3mHAY
jwzj16qzNkBaT6re+mA5Y1G1riiLWzZf+qm/Aj9jl2bll0eWa8PcD59LZyjvzTFD
2i0dHEY6bHbcw8C1D3vldo3vE3Nkj8SrS53j8RnB2a9PZblPtAq4yxiIMt7nWz6u
4lbWDkXNBtk1Febuw+KgOLbUEHJeFpCaJu9lIHLK0YFBFYDU6IMbHKE9con1w9hW
62+LzT0Ksi3I7tn2uJv9mtENYyfae7Itu9/VVPervAeSLBQdO4g2qkKvkZGwrrwD
X7LH2CBneoye34caCDsRpDGERnTl2o0qbWyH4hJmTv11gYbTGMvS6QUQFJC29le/
pcwGCvr7hY0GRKw6oN+M8KLl+xndWgx+hzmVgqhVyzpefLpHKvRCRFZo1s7/Kjgb
CofhTdm1//dMNAC3NhAzmphyvxumg/kuZyMmx7vhsng+fMmw8VGkE/r2+jq8q4hA
IK0EjYVgLAEq5YRAlkwzrgWVc6HgwLZUqxVt/ZgOp4pCIm9NewZxumfOxpaHiSk/
sA25jYOE4FXZXenkf0wtvA6ZwWYBfJSrlAeKVn3stN+RV7rDRJ8mXsHouZrYEQE1
SMQkT4S9YXnGCghvH+XLeP6KE+Hsdeg0GyY9fzefDR5MIJEUSQ/4f+AAGBunZ3eW
nlqD7nuQhjKct+oY06MC2rm8WXJc/L8l8/KY/h07IB+Iq4qpJFdjir9kvyZh63ti
u1BaNr8tr9zRAqLkHdmCL2fqnAmhDO7JOIOb93/YMlxvXzE3ofoKF0abJ+5UVvDu
ZgP77qgt8yxT8iOD/OKFHchc5bk+aS3ieHmGql+6+7DDZjb2SMSns2vBX1NJlei/
d+B1W4QxdOBeuxPkcUhQ3YvG49qqEQlBQnNuzag7PJTm+kP4sfgQ3vJOPpDoy6Yb
bQQIEQLkv4L5P5HvvWpQYhM9VgTeFb9OFgJvvNFc8+CmfLvqyWxncRguGnzLdyc6
TfZyJgyx/ke9yPzXy5L8UhwrJNczN/l8rcKu362RvWlyvrDRfCXrapJlFCGJh8lH
aHSyU2JPKLAL7G8JdWK51LtuOS6wQFXE+CgxsJQVNpukIriRDu5EZESFH6ZaDLGy
0+2zYSOcssOJW9KlEMWHuqVtEMwu8zGODohRPVZlCeonInYzILc3Li0uLw2s7Djs
9ftUk2QUFU25Ctdl3zHw1l3XQHsuKChwOh+Ife4CS/nivDDIXxxDoINfRhGQtPec
AuFE8w1idwDH1eNRy84pREoAjBA+E0W1/ADJraS0XfpxRH9+9zYxDbDrMwC7y0hc
8ZhHidQaL9l6+O8kW696ofBeT7Ctdyl6GzkZHyPkEFXS+Ij2vd/0zengVbwxBzeu
nH3qZHpCVmtey8LIuolGxiB1Bob+o33rxHexTdDfyBbb9t7TyFN0WvdlfeQT77dy
qcbTi4vRjoSjdQqnyyF09e2rpyarqbgQ+lD/YwWG59axYZxF4d6AmkNT3gLvIqjI
x+FMK8H7LRtJtNyOZrz9x8RrvHzk3JudV8bNam2TT/VpjWpr0DrhpEMgLkaUoDlX
y6jQHzYzrR6kf+Y/nZy+cL3vycGSojke2zFMvzB/jwXX/ltCBTNGf24Cnie9DP5q
G+cqQ+cAVvbntJKKF7n0htBB0PXIp27dkzgpMOSFVPJG6m85AkSpXRhjSEpVzkzz
hPyLneb+P7iEify4UTyCYiw4Sd5p27/fQooxKuum89rH6hJxdE3zXVuebS+ZzZqq
L+eXVFYJgnZZi+/jCvIRFa3TY/jOb0UdxWQmW/W6u8/8m38tqG8Gye3bu2pO403P
RdRf2JVNUaAXGqhoqkWLLp9s/onmQNQUxo64O0II3LJ82EUguHFKLeFJnayPiyyz
OH93YZ9p5Mvttom/ZkqXIth+P2uuWY7IiSzSxuZYLq7LF88OIiiBB9RUa7fQp79i
TtiCDHz3it9ykAS1qqzHVFOBZsCoG4f1LKy1EMGxpkMVLUnS7g/fF2JTCKiUW3DD
68GjoClrrdcFbxwhSl98wf3r+mXzJRJionaT+j3sBvAB2iG5dFgcMjTpvyvXB3n3
OQYLJ4fCuXypjLsSCAoht/tz53FYr7F8YVbyLdajsnAebQBzGcu/Tlovh+Hw5Dma
b9akZTAY9EbitOzN4YYqJ8VeeC9hx/h/71xMcdNNY+oNzYFg+Kua/uAOPV9MltHg
ob3zgiByAwDSS2E6IM+yj5/DVkDX368beXvbnMkzREQW+3+HVwXntbQmwMF2DHG6
6sGa2OLvvsyTCQaPrrrJ4RQ5pBrXHxLLJZQj9hHLIluSycKXwoPAUBOQA8alCp8E
SjrfqQ+V1elxipGMCBVNA2PxgMz/K4UGgbTzgvgFnzlw1oMGUtCCrwwuOasc+8Ei
rCiW1s9SrEHcyPSsaI8mLHxhevDtxMdTtJZ8I95jfPoJ1wlrpgG3ZsxlPf4OUROn
CO6nq75E/caPi+6ADDMKtDkC86hq5wF+LPkil/yYmoZZFnL9ATJWiEkh00I9Rf5w
53CzLERRpzpDfxnXoz9+gpjQbL2jEyyqHN4yeldDfebc4IBbY71Bc3dgwRF8dB4v
GCLQE8IXrfHB5TN7hByWYzRFY0rRMhf79ORgvJg4VaBHvKMLN+UjVNfO0EpqXjr/
djFzXBz9GgCIgKm1iykPF7YtO4mwCgTdNGBczCJ6GNH2qwKszwfJRwOkL0qIPlA4
SAnGSkJZ2Hx8kb/VmNovQ4NSoemONMZaZAMG/HdSm7XbZGnNf79gjqJ0Q6UTITyn
UGF+6sK66fWmInbw42EJJ/olVnE3lwdEPmMhoCVLVP5o8z5pUVuFeXsykCt2s24T
mbwYhNDjlIb/NW4hdakM0lcf391byCJLscqpbT8NDWSwFwQPegCw+zQ788Xc9scm
fN0BRrR8i1iUD3kyz2N2l9xem9Fl1ZdLPetmMPG+ZXxKoX3b1rccpXqlOrwunUfV
YLG1AfSiRhLNBDE5V71AeNyCCcWqlgdxnw3e4lk7WEpi8Rj46sy0YVUfTp/Zj/Ta
4qI2ouuOxHuzxcPflYbYtJsCOLq8Cah1rHNseHRuiq0ECByJHz++tiu/kXgr6ftT
JPFHQHEUSYZiOsuI18FldOTm7VciUgKNJ6JFLzwSaZbl+tZ6bxtddHIVNMOsJRNA
t99/y6Mo6vEbLkji/8iWtVDg11EGe14YTQ5rPAuwn/c/iNuayiMaUoVaKy25PUyd
cz8G+NC4cp1q5Qe+QpJdCh6qunQ26HG6yBPCAoypZB7DF4vZILqfJzUSgrRFm0sh
gg1C54Pn0qVJkTX0yM+ocSchRy3McPtV8/WdmZjHYr6kKAXsV/aukNf19Uih1++J
DwQSt6vGVFaQLbkpd4OzqwzNdXwNAEsnQUbBFnXhS+FaNhzSo/hMVwyJpldUu3qF
Jwrn9Qx9pbYFQyHVL81j0L80SM9wAYRKP9WFvr9PlNot3Q5DsyqlauJKxl6+BrEO
bD0xx9DzVlc0ACpVAMs9gmyRFPIJsPvfC1oeDUs4/0igVSoLR4gtdZkv2yxSzQMF
p4xzYNApuRoEo0S4UimArURRKCGwbdB5tXTJFF9UPS2ip5PUJlaARozNZlPZL+wO
Gy8vSUS5qf5KvdbiYHBDS7AX9wzT8rQdYN421bGo/CIocEgp6/pVL15wsYzuk/g/
+8Xtoa2OPJ37PZYsFv2F4pIpCLB9I/U9nD+lKUyIg2QvJvMPjfLD+ZRZOJMoHcri
C/3Gq/iBHNfFQ1NcC1+lVNpNJRUdx484quOTk8ldIn9DVas/y/kF32Z3+gOWUmLr
n36VxHx5fUzl7BLXNbJcCj+XLVCKfyBlGLTjUf+oviRPPwBqxTTJxp3OaPW/VLZt
GwSLotEfoogONjhfXuQAhoAUGerzipY9m/06/j7nZC0vTQQbGSpyDGqLR5NEvv+l
qydtGlkzJMtvBv9CTF1vzA==
`pragma protect end_protected

-- coproc_soft_cpu.vhd

-- Generated using ACDS version 24.1 1077

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity coproc_soft_cpu is
	port (
		i_clk_clk                                : in  std_logic                     := '0';             --                 i_clk.clk
		i_clr_reset_n                            : in  std_logic                     := '0';             --                 i_clr.reset_n
		o_batch_data_export_conduit_i_rd_clk     : in  std_logic                     := '0';             --   o_batch_data_export.conduit_i_rd_clk
		o_batch_data_export_conduit_i_rd_row     : in  std_logic_vector(2 downto 0)  := (others => '0'); --                      .conduit_i_rd_row
		o_batch_data_export_conduit_o_data       : out std_logic_vector(63 downto 0);                    --                      .conduit_o_data
		o_batch_data_export_conduit_o_rd_ready   : out std_logic;                                        --                      .conduit_o_rd_ready
		o_batch_weight_export_conduit_i_rd_clk   : in  std_logic                     := '0';             -- o_batch_weight_export.conduit_i_rd_clk
		o_batch_weight_export_conduit_i_rd_row   : in  std_logic_vector(2 downto 0)  := (others => '0'); --                      .conduit_i_rd_row
		o_batch_weight_export_conduit_o_data     : out std_logic_vector(63 downto 0);                    --                      .conduit_o_data
		o_batch_weight_export_conduit_o_rd_ready : out std_logic;                                        --                      .conduit_o_rd_ready
		o_serializer_export_i_acc                : in  std_logic_vector(31 downto 0) := (others => '0'); --   o_serializer_export.i_acc
		o_serializer_export_o_clr                : out std_logic;                                        --                      .o_clr
		o_serializer_export_o_read               : out std_logic;                                        --                      .o_read
		o_spi_export_MISO                        : out std_logic;                                        --          o_spi_export.MISO
		o_spi_export_MOSI                        : in  std_logic                     := '0';             --                      .MOSI
		o_spi_export_SCLK                        : in  std_logic                     := '0';             --                      .SCLK
		o_spi_export_SS_n                        : in  std_logic                     := '0'              --                      .SS_n
	);
end entity coproc_soft_cpu;

architecture rtl of coproc_soft_cpu is
	component coproc_soft_cpu_CPU is
		port (
			clk                               : in  std_logic                     := 'X';             -- clk
			reset_reset                       : in  std_logic                     := 'X';             -- reset
			platform_irq_rx_irq               : in  std_logic_vector(15 downto 0) := (others => 'X'); -- irq
			ndm_reset_in_reset                : in  std_logic                     := 'X';             -- reset
			timer_sw_agent_address            : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- address
			timer_sw_agent_byteenable         : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			timer_sw_agent_read               : in  std_logic                     := 'X';             -- read
			timer_sw_agent_readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			timer_sw_agent_write              : in  std_logic                     := 'X';             -- write
			timer_sw_agent_writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			timer_sw_agent_waitrequest        : out std_logic;                                        -- waitrequest
			timer_sw_agent_readdatavalid      : out std_logic;                                        -- readdatavalid
			instruction_manager_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			instruction_manager_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			instruction_manager_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			instruction_manager_response      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			instruction_manager_address       : out std_logic_vector(31 downto 0);                    -- address
			instruction_manager_read          : out std_logic;                                        -- read
			data_manager_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			data_manager_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			data_manager_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			data_manager_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			data_manager_address              : out std_logic_vector(31 downto 0);                    -- address
			data_manager_read                 : out std_logic;                                        -- read
			data_manager_write                : out std_logic;                                        -- write
			data_manager_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			data_manager_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			data_manager_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			dm_agent_address                  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			dm_agent_read                     : in  std_logic                     := 'X';             -- read
			dm_agent_readdata                 : out std_logic_vector(31 downto 0);                    -- readdata
			dm_agent_write                    : in  std_logic                     := 'X';             -- write
			dm_agent_writedata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dm_agent_waitrequest              : out std_logic;                                        -- waitrequest
			dm_agent_readdatavalid            : out std_logic;                                        -- readdatavalid
			dbg_reset_out_reset               : out std_logic                                         -- reset
		);
	end component coproc_soft_cpu_CPU;

	component avalon_batch_block is
		generic (
			g_PORTA_ADDR_SIZE : natural := 6;
			g_PORTB_ADDR_SIZE : natural := 3;
			g_BATCH_SIZE      : natural := 8
		);
		port (
			av_address     : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- address
			av_write       : in  std_logic                     := 'X';             -- write
			av_read        : in  std_logic                     := 'X';             -- read
			av_writedata   : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			av_readdata    : out std_logic_vector(7 downto 0);                     -- readdata
			av_waitrequest : out std_logic;                                        -- waitrequest
			i_rd_clk       : in  std_logic                     := 'X';             -- conduit_i_rd_clk
			i_rd_row       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- conduit_i_rd_row
			o_data         : out std_logic_vector(63 downto 0);                    -- conduit_o_data
			o_rd_ready     : out std_logic;                                        -- conduit_o_rd_ready
			ni_clr         : in  std_logic                     := 'X';             -- reset_n
			i_clk          : in  std_logic                     := 'X'              -- clk
		);
	end component avalon_batch_block;

	component altera_avalon_jtag_uart is
		generic (
			readBufferDepth            : integer := 64;
			readIRQThreshold           : integer := 8;
			useRegistersForReadBuffer  : boolean := false;
			useRegistersForWriteBuffer : boolean := false;
			writeBufferDepth           : integer := 64;
			writeIRQThreshold          : integer := 8;
			printingMethod             : boolean := false;
			FIFO_WIDTH                 : integer := 8;
			WR_WIDTHU                  : integer := 0;
			RD_WIDTHU                  : integer := 0;
			write_le                   : string  := """ON""";
			read_le                    : string  := """ON""";
			HEX_WRITE_DEPTH_STR        : integer := 64;
			HEX_READ_DEPTH_STR         : integer := 64;
			legacySignalAllow          : boolean := true
		);
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component altera_avalon_jtag_uart;

	component avalon_serializer is
		port (
			i_acc          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- i_acc
			o_clr          : out std_logic;                                        -- o_clr
			o_read         : out std_logic;                                        -- o_read
			ni_clr         : in  std_logic                     := 'X';             -- reset_n
			i_clk          : in  std_logic                     := 'X';             -- clk
			av_address     : in  std_logic                     := 'X';             -- address
			av_write       : in  std_logic                     := 'X';             -- write
			av_read        : in  std_logic                     := 'X';             -- read
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_waitrequest : out std_logic                                         -- waitrequest
		);
	end component avalon_serializer;

	component coproc_soft_cpu_SPI_0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			data_from_cpu : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			data_to_cpu   : out std_logic_vector(15 downto 0);                    -- readdata
			mem_addr      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			read_n        : in  std_logic                     := 'X';             -- read_n
			spi_select    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			MISO          : out std_logic;                                        -- export
			MOSI          : in  std_logic                     := 'X';             -- export
			SCLK          : in  std_logic                     := 'X';             -- export
			SS_n          : in  std_logic                     := 'X'              -- export
		);
	end component coproc_soft_cpu_SPI_0;

	component coproc_soft_cpu_SRAM is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component coproc_soft_cpu_SRAM;

	component coproc_soft_cpu_mm_interconnect_0 is
		port (
			CLK_clk_clk                                      : in  std_logic                     := 'X';             -- clk
			CPU_reset_reset_bridge_in_reset_reset            : in  std_logic                     := 'X';             -- reset
			WEIGHT_BATCH_reset_n_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			CPU_data_manager_address                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			CPU_data_manager_waitrequest                     : out std_logic;                                        -- waitrequest
			CPU_data_manager_byteenable                      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			CPU_data_manager_read                            : in  std_logic                     := 'X';             -- read
			CPU_data_manager_readdata                        : out std_logic_vector(31 downto 0);                    -- readdata
			CPU_data_manager_readdatavalid                   : out std_logic;                                        -- readdatavalid
			CPU_data_manager_write                           : in  std_logic                     := 'X';             -- write
			CPU_data_manager_writedata                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			CPU_data_manager_response                        : out std_logic_vector(1 downto 0);                     -- response
			CPU_data_manager_writeresponsevalid              : out std_logic;                                        -- writeresponsevalid
			CPU_instruction_manager_address                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			CPU_instruction_manager_waitrequest              : out std_logic;                                        -- waitrequest
			CPU_instruction_manager_read                     : in  std_logic                     := 'X';             -- read
			CPU_instruction_manager_readdata                 : out std_logic_vector(31 downto 0);                    -- readdata
			CPU_instruction_manager_readdatavalid            : out std_logic;                                        -- readdatavalid
			CPU_instruction_manager_response                 : out std_logic_vector(1 downto 0);                     -- response
			CPU_dm_agent_address                             : out std_logic_vector(15 downto 0);                    -- address
			CPU_dm_agent_write                               : out std_logic;                                        -- write
			CPU_dm_agent_read                                : out std_logic;                                        -- read
			CPU_dm_agent_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			CPU_dm_agent_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			CPU_dm_agent_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			CPU_dm_agent_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			CPU_timer_sw_agent_address                       : out std_logic_vector(5 downto 0);                     -- address
			CPU_timer_sw_agent_write                         : out std_logic;                                        -- write
			CPU_timer_sw_agent_read                          : out std_logic;                                        -- read
			CPU_timer_sw_agent_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			CPU_timer_sw_agent_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			CPU_timer_sw_agent_byteenable                    : out std_logic_vector(3 downto 0);                     -- byteenable
			CPU_timer_sw_agent_readdatavalid                 : in  std_logic                     := 'X';             -- readdatavalid
			CPU_timer_sw_agent_waitrequest                   : in  std_logic                     := 'X';             -- waitrequest
			DATA_BATCH_avalon_address                        : out std_logic_vector(5 downto 0);                     -- address
			DATA_BATCH_avalon_write                          : out std_logic;                                        -- write
			DATA_BATCH_avalon_read                           : out std_logic;                                        -- read
			DATA_BATCH_avalon_readdata                       : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			DATA_BATCH_avalon_writedata                      : out std_logic_vector(7 downto 0);                     -- writedata
			DATA_BATCH_avalon_waitrequest                    : in  std_logic                     := 'X';             -- waitrequest
			DEBUG_JTAG_avalon_jtag_slave_address             : out std_logic_vector(0 downto 0);                     -- address
			DEBUG_JTAG_avalon_jtag_slave_write               : out std_logic;                                        -- write
			DEBUG_JTAG_avalon_jtag_slave_read                : out std_logic;                                        -- read
			DEBUG_JTAG_avalon_jtag_slave_readdata            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			DEBUG_JTAG_avalon_jtag_slave_writedata           : out std_logic_vector(31 downto 0);                    -- writedata
			DEBUG_JTAG_avalon_jtag_slave_waitrequest         : in  std_logic                     := 'X';             -- waitrequest
			DEBUG_JTAG_avalon_jtag_slave_chipselect          : out std_logic;                                        -- chipselect
			SERIALIZER_0_avalon_address                      : out std_logic_vector(0 downto 0);                     -- address
			SERIALIZER_0_avalon_write                        : out std_logic;                                        -- write
			SERIALIZER_0_avalon_read                         : out std_logic;                                        -- read
			SERIALIZER_0_avalon_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			SERIALIZER_0_avalon_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			SERIALIZER_0_avalon_waitrequest                  : in  std_logic                     := 'X';             -- waitrequest
			SPI_0_spi_control_port_address                   : out std_logic_vector(2 downto 0);                     -- address
			SPI_0_spi_control_port_write                     : out std_logic;                                        -- write
			SPI_0_spi_control_port_read                      : out std_logic;                                        -- read
			SPI_0_spi_control_port_readdata                  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			SPI_0_spi_control_port_writedata                 : out std_logic_vector(15 downto 0);                    -- writedata
			SPI_0_spi_control_port_chipselect                : out std_logic;                                        -- chipselect
			SRAM_s1_address                                  : out std_logic_vector(12 downto 0);                    -- address
			SRAM_s1_write                                    : out std_logic;                                        -- write
			SRAM_s1_readdata                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			SRAM_s1_writedata                                : out std_logic_vector(31 downto 0);                    -- writedata
			SRAM_s1_byteenable                               : out std_logic_vector(3 downto 0);                     -- byteenable
			SRAM_s1_chipselect                               : out std_logic;                                        -- chipselect
			SRAM_s1_clken                                    : out std_logic;                                        -- clken
			WEIGHT_BATCH_avalon_address                      : out std_logic_vector(5 downto 0);                     -- address
			WEIGHT_BATCH_avalon_write                        : out std_logic;                                        -- write
			WEIGHT_BATCH_avalon_read                         : out std_logic;                                        -- read
			WEIGHT_BATCH_avalon_readdata                     : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			WEIGHT_BATCH_avalon_writedata                    : out std_logic_vector(7 downto 0);                     -- writedata
			WEIGHT_BATCH_avalon_waitrequest                  : in  std_logic                     := 'X'              -- waitrequest
		);
	end component coproc_soft_cpu_mm_interconnect_0;

	component coproc_soft_cpu_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(15 downto 0)         -- irq
		);
	end component coproc_soft_cpu_irq_mapper;

	component coproc_soft_cpu_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in1      : in  std_logic := 'X';
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component coproc_soft_cpu_rst_controller;

	component coproc_soft_cpu_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component coproc_soft_cpu_rst_controller_001;

	signal cpu_data_manager_readdata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_data_manager_readdata -> CPU:data_manager_readdata
	signal cpu_data_manager_waitrequest                                   : std_logic;                     -- mm_interconnect_0:CPU_data_manager_waitrequest -> CPU:data_manager_waitrequest
	signal cpu_data_manager_address                                       : std_logic_vector(31 downto 0); -- CPU:data_manager_address -> mm_interconnect_0:CPU_data_manager_address
	signal cpu_data_manager_read                                          : std_logic;                     -- CPU:data_manager_read -> mm_interconnect_0:CPU_data_manager_read
	signal cpu_data_manager_byteenable                                    : std_logic_vector(3 downto 0);  -- CPU:data_manager_byteenable -> mm_interconnect_0:CPU_data_manager_byteenable
	signal cpu_data_manager_readdatavalid                                 : std_logic;                     -- mm_interconnect_0:CPU_data_manager_readdatavalid -> CPU:data_manager_readdatavalid
	signal cpu_data_manager_response                                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:CPU_data_manager_response -> CPU:data_manager_response
	signal cpu_data_manager_write                                         : std_logic;                     -- CPU:data_manager_write -> mm_interconnect_0:CPU_data_manager_write
	signal cpu_data_manager_writedata                                     : std_logic_vector(31 downto 0); -- CPU:data_manager_writedata -> mm_interconnect_0:CPU_data_manager_writedata
	signal cpu_data_manager_writeresponsevalid                            : std_logic;                     -- mm_interconnect_0:CPU_data_manager_writeresponsevalid -> CPU:data_manager_writeresponsevalid
	signal cpu_instruction_manager_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_instruction_manager_readdata -> CPU:instruction_manager_readdata
	signal cpu_instruction_manager_waitrequest                            : std_logic;                     -- mm_interconnect_0:CPU_instruction_manager_waitrequest -> CPU:instruction_manager_waitrequest
	signal cpu_instruction_manager_address                                : std_logic_vector(31 downto 0); -- CPU:instruction_manager_address -> mm_interconnect_0:CPU_instruction_manager_address
	signal cpu_instruction_manager_read                                   : std_logic;                     -- CPU:instruction_manager_read -> mm_interconnect_0:CPU_instruction_manager_read
	signal cpu_instruction_manager_readdatavalid                          : std_logic;                     -- mm_interconnect_0:CPU_instruction_manager_readdatavalid -> CPU:instruction_manager_readdatavalid
	signal cpu_instruction_manager_response                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:CPU_instruction_manager_response -> CPU:instruction_manager_response
	signal mm_interconnect_0_weight_batch_avalon_readdata                 : std_logic_vector(7 downto 0);  -- WEIGHT_BATCH:av_readdata -> mm_interconnect_0:WEIGHT_BATCH_avalon_readdata
	signal mm_interconnect_0_weight_batch_avalon_waitrequest              : std_logic;                     -- WEIGHT_BATCH:av_waitrequest -> mm_interconnect_0:WEIGHT_BATCH_avalon_waitrequest
	signal mm_interconnect_0_weight_batch_avalon_address                  : std_logic_vector(5 downto 0);  -- mm_interconnect_0:WEIGHT_BATCH_avalon_address -> WEIGHT_BATCH:av_address
	signal mm_interconnect_0_weight_batch_avalon_read                     : std_logic;                     -- mm_interconnect_0:WEIGHT_BATCH_avalon_read -> WEIGHT_BATCH:av_read
	signal mm_interconnect_0_weight_batch_avalon_write                    : std_logic;                     -- mm_interconnect_0:WEIGHT_BATCH_avalon_write -> WEIGHT_BATCH:av_write
	signal mm_interconnect_0_weight_batch_avalon_writedata                : std_logic_vector(7 downto 0);  -- mm_interconnect_0:WEIGHT_BATCH_avalon_writedata -> WEIGHT_BATCH:av_writedata
	signal mm_interconnect_0_data_batch_avalon_readdata                   : std_logic_vector(7 downto 0);  -- DATA_BATCH:av_readdata -> mm_interconnect_0:DATA_BATCH_avalon_readdata
	signal mm_interconnect_0_data_batch_avalon_waitrequest                : std_logic;                     -- DATA_BATCH:av_waitrequest -> mm_interconnect_0:DATA_BATCH_avalon_waitrequest
	signal mm_interconnect_0_data_batch_avalon_address                    : std_logic_vector(5 downto 0);  -- mm_interconnect_0:DATA_BATCH_avalon_address -> DATA_BATCH:av_address
	signal mm_interconnect_0_data_batch_avalon_read                       : std_logic;                     -- mm_interconnect_0:DATA_BATCH_avalon_read -> DATA_BATCH:av_read
	signal mm_interconnect_0_data_batch_avalon_write                      : std_logic;                     -- mm_interconnect_0:DATA_BATCH_avalon_write -> DATA_BATCH:av_write
	signal mm_interconnect_0_data_batch_avalon_writedata                  : std_logic_vector(7 downto 0);  -- mm_interconnect_0:DATA_BATCH_avalon_writedata -> DATA_BATCH:av_writedata
	signal mm_interconnect_0_serializer_0_avalon_readdata                 : std_logic_vector(31 downto 0); -- SERIALIZER_0:av_readdata -> mm_interconnect_0:SERIALIZER_0_avalon_readdata
	signal mm_interconnect_0_serializer_0_avalon_waitrequest              : std_logic;                     -- SERIALIZER_0:av_waitrequest -> mm_interconnect_0:SERIALIZER_0_avalon_waitrequest
	signal mm_interconnect_0_serializer_0_avalon_address                  : std_logic_vector(0 downto 0);  -- mm_interconnect_0:SERIALIZER_0_avalon_address -> SERIALIZER_0:av_address
	signal mm_interconnect_0_serializer_0_avalon_read                     : std_logic;                     -- mm_interconnect_0:SERIALIZER_0_avalon_read -> SERIALIZER_0:av_read
	signal mm_interconnect_0_serializer_0_avalon_write                    : std_logic;                     -- mm_interconnect_0:SERIALIZER_0_avalon_write -> SERIALIZER_0:av_write
	signal mm_interconnect_0_serializer_0_avalon_writedata                : std_logic_vector(31 downto 0); -- mm_interconnect_0:SERIALIZER_0_avalon_writedata -> SERIALIZER_0:av_writedata
	signal mm_interconnect_0_debug_jtag_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:DEBUG_JTAG_avalon_jtag_slave_chipselect -> DEBUG_JTAG:av_chipselect
	signal mm_interconnect_0_debug_jtag_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- DEBUG_JTAG:av_readdata -> mm_interconnect_0:DEBUG_JTAG_avalon_jtag_slave_readdata
	signal mm_interconnect_0_debug_jtag_avalon_jtag_slave_waitrequest     : std_logic;                     -- DEBUG_JTAG:av_waitrequest -> mm_interconnect_0:DEBUG_JTAG_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_debug_jtag_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:DEBUG_JTAG_avalon_jtag_slave_address -> DEBUG_JTAG:av_address
	signal mm_interconnect_0_debug_jtag_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:DEBUG_JTAG_avalon_jtag_slave_read -> mm_interconnect_0_debug_jtag_avalon_jtag_slave_read:in
	signal mm_interconnect_0_debug_jtag_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:DEBUG_JTAG_avalon_jtag_slave_write -> mm_interconnect_0_debug_jtag_avalon_jtag_slave_write:in
	signal mm_interconnect_0_debug_jtag_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:DEBUG_JTAG_avalon_jtag_slave_writedata -> DEBUG_JTAG:av_writedata
	signal mm_interconnect_0_cpu_dm_agent_readdata                        : std_logic_vector(31 downto 0); -- CPU:dm_agent_readdata -> mm_interconnect_0:CPU_dm_agent_readdata
	signal mm_interconnect_0_cpu_dm_agent_waitrequest                     : std_logic;                     -- CPU:dm_agent_waitrequest -> mm_interconnect_0:CPU_dm_agent_waitrequest
	signal mm_interconnect_0_cpu_dm_agent_address                         : std_logic_vector(15 downto 0); -- mm_interconnect_0:CPU_dm_agent_address -> CPU:dm_agent_address
	signal mm_interconnect_0_cpu_dm_agent_read                            : std_logic;                     -- mm_interconnect_0:CPU_dm_agent_read -> CPU:dm_agent_read
	signal mm_interconnect_0_cpu_dm_agent_readdatavalid                   : std_logic;                     -- CPU:dm_agent_readdatavalid -> mm_interconnect_0:CPU_dm_agent_readdatavalid
	signal mm_interconnect_0_cpu_dm_agent_write                           : std_logic;                     -- mm_interconnect_0:CPU_dm_agent_write -> CPU:dm_agent_write
	signal mm_interconnect_0_cpu_dm_agent_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_dm_agent_writedata -> CPU:dm_agent_writedata
	signal mm_interconnect_0_sram_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:SRAM_s1_chipselect -> SRAM:chipselect
	signal mm_interconnect_0_sram_s1_readdata                             : std_logic_vector(31 downto 0); -- SRAM:readdata -> mm_interconnect_0:SRAM_s1_readdata
	signal mm_interconnect_0_sram_s1_address                              : std_logic_vector(12 downto 0); -- mm_interconnect_0:SRAM_s1_address -> SRAM:address
	signal mm_interconnect_0_sram_s1_byteenable                           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:SRAM_s1_byteenable -> SRAM:byteenable
	signal mm_interconnect_0_sram_s1_write                                : std_logic;                     -- mm_interconnect_0:SRAM_s1_write -> SRAM:write
	signal mm_interconnect_0_sram_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:SRAM_s1_writedata -> SRAM:writedata
	signal mm_interconnect_0_sram_s1_clken                                : std_logic;                     -- mm_interconnect_0:SRAM_s1_clken -> SRAM:clken
	signal mm_interconnect_0_spi_0_spi_control_port_chipselect            : std_logic;                     -- mm_interconnect_0:SPI_0_spi_control_port_chipselect -> SPI_0:spi_select
	signal mm_interconnect_0_spi_0_spi_control_port_readdata              : std_logic_vector(15 downto 0); -- SPI_0:data_to_cpu -> mm_interconnect_0:SPI_0_spi_control_port_readdata
	signal mm_interconnect_0_spi_0_spi_control_port_address               : std_logic_vector(2 downto 0);  -- mm_interconnect_0:SPI_0_spi_control_port_address -> SPI_0:mem_addr
	signal mm_interconnect_0_spi_0_spi_control_port_read                  : std_logic;                     -- mm_interconnect_0:SPI_0_spi_control_port_read -> mm_interconnect_0_spi_0_spi_control_port_read:in
	signal mm_interconnect_0_spi_0_spi_control_port_write                 : std_logic;                     -- mm_interconnect_0:SPI_0_spi_control_port_write -> mm_interconnect_0_spi_0_spi_control_port_write:in
	signal mm_interconnect_0_spi_0_spi_control_port_writedata             : std_logic_vector(15 downto 0); -- mm_interconnect_0:SPI_0_spi_control_port_writedata -> SPI_0:data_from_cpu
	signal mm_interconnect_0_cpu_timer_sw_agent_readdata                  : std_logic_vector(31 downto 0); -- CPU:timer_sw_agent_readdata -> mm_interconnect_0:CPU_timer_sw_agent_readdata
	signal mm_interconnect_0_cpu_timer_sw_agent_waitrequest               : std_logic;                     -- CPU:timer_sw_agent_waitrequest -> mm_interconnect_0:CPU_timer_sw_agent_waitrequest
	signal mm_interconnect_0_cpu_timer_sw_agent_address                   : std_logic_vector(5 downto 0);  -- mm_interconnect_0:CPU_timer_sw_agent_address -> CPU:timer_sw_agent_address
	signal mm_interconnect_0_cpu_timer_sw_agent_read                      : std_logic;                     -- mm_interconnect_0:CPU_timer_sw_agent_read -> CPU:timer_sw_agent_read
	signal mm_interconnect_0_cpu_timer_sw_agent_byteenable                : std_logic_vector(3 downto 0);  -- mm_interconnect_0:CPU_timer_sw_agent_byteenable -> CPU:timer_sw_agent_byteenable
	signal mm_interconnect_0_cpu_timer_sw_agent_readdatavalid             : std_logic;                     -- CPU:timer_sw_agent_readdatavalid -> mm_interconnect_0:CPU_timer_sw_agent_readdatavalid
	signal mm_interconnect_0_cpu_timer_sw_agent_write                     : std_logic;                     -- mm_interconnect_0:CPU_timer_sw_agent_write -> CPU:timer_sw_agent_write
	signal mm_interconnect_0_cpu_timer_sw_agent_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_timer_sw_agent_writedata -> CPU:timer_sw_agent_writedata
	signal irq_mapper_receiver0_irq                                       : std_logic;                     -- DEBUG_JTAG:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                       : std_logic;                     -- SPI_0:irq -> irq_mapper:receiver1_irq
	signal cpu_platform_irq_rx_irq                                        : std_logic_vector(15 downto 0); -- irq_mapper:sender_irq -> CPU:platform_irq_rx_irq
	signal rst_controller_reset_out_reset                                 : std_logic;                     -- rst_controller:reset_out -> [CPU:reset_reset, irq_mapper:reset, mm_interconnect_0:CPU_reset_reset_bridge_in_reset_reset]
	signal rst_controller_001_reset_out_reset                             : std_logic;                     -- rst_controller_001:reset_out -> [CPU:ndm_reset_in_reset, SRAM:reset, mm_interconnect_0:WEIGHT_BATCH_reset_n_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_001_reset_out_reset_req                         : std_logic;                     -- rst_controller_001:reset_req -> [SRAM:reset_req, rst_translator:reset_req_in]
	signal cpu_dbg_reset_out_reset                                        : std_logic;                     -- CPU:dbg_reset_out_reset -> rst_controller_001:reset_in1
	signal i_clr_reset_n_ports_inv                                        : std_logic;                     -- i_clr_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_debug_jtag_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_debug_jtag_avalon_jtag_slave_read:inv -> DEBUG_JTAG:av_read_n
	signal mm_interconnect_0_debug_jtag_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_debug_jtag_avalon_jtag_slave_write:inv -> DEBUG_JTAG:av_write_n
	signal mm_interconnect_0_spi_0_spi_control_port_read_ports_inv        : std_logic;                     -- mm_interconnect_0_spi_0_spi_control_port_read:inv -> SPI_0:read_n
	signal mm_interconnect_0_spi_0_spi_control_port_write_ports_inv       : std_logic;                     -- mm_interconnect_0_spi_0_spi_control_port_write:inv -> SPI_0:write_n
	signal rst_controller_001_reset_out_reset_ports_inv                   : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> [DATA_BATCH:ni_clr, DEBUG_JTAG:rst_n, SERIALIZER_0:ni_clr, SPI_0:reset_n, WEIGHT_BATCH:ni_clr]

begin

	cpu : component coproc_soft_cpu_CPU
		port map (
			clk                               => i_clk_clk,                                          --                 clk.clk
			reset_reset                       => rst_controller_reset_out_reset,                     --               reset.reset
			platform_irq_rx_irq               => cpu_platform_irq_rx_irq,                            --     platform_irq_rx.irq
			ndm_reset_in_reset                => rst_controller_001_reset_out_reset,                 --        ndm_reset_in.reset
			timer_sw_agent_address            => mm_interconnect_0_cpu_timer_sw_agent_address,       --      timer_sw_agent.address
			timer_sw_agent_byteenable         => mm_interconnect_0_cpu_timer_sw_agent_byteenable,    --                    .byteenable
			timer_sw_agent_read               => mm_interconnect_0_cpu_timer_sw_agent_read,          --                    .read
			timer_sw_agent_readdata           => mm_interconnect_0_cpu_timer_sw_agent_readdata,      --                    .readdata
			timer_sw_agent_write              => mm_interconnect_0_cpu_timer_sw_agent_write,         --                    .write
			timer_sw_agent_writedata          => mm_interconnect_0_cpu_timer_sw_agent_writedata,     --                    .writedata
			timer_sw_agent_waitrequest        => mm_interconnect_0_cpu_timer_sw_agent_waitrequest,   --                    .waitrequest
			timer_sw_agent_readdatavalid      => mm_interconnect_0_cpu_timer_sw_agent_readdatavalid, --                    .readdatavalid
			instruction_manager_readdata      => cpu_instruction_manager_readdata,                   -- instruction_manager.readdata
			instruction_manager_waitrequest   => cpu_instruction_manager_waitrequest,                --                    .waitrequest
			instruction_manager_readdatavalid => cpu_instruction_manager_readdatavalid,              --                    .readdatavalid
			instruction_manager_response      => cpu_instruction_manager_response,                   --                    .response
			instruction_manager_address       => cpu_instruction_manager_address,                    --                    .address
			instruction_manager_read          => cpu_instruction_manager_read,                       --                    .read
			data_manager_readdata             => cpu_data_manager_readdata,                          --        data_manager.readdata
			data_manager_waitrequest          => cpu_data_manager_waitrequest,                       --                    .waitrequest
			data_manager_readdatavalid        => cpu_data_manager_readdatavalid,                     --                    .readdatavalid
			data_manager_response             => cpu_data_manager_response,                          --                    .response
			data_manager_address              => cpu_data_manager_address,                           --                    .address
			data_manager_read                 => cpu_data_manager_read,                              --                    .read
			data_manager_write                => cpu_data_manager_write,                             --                    .write
			data_manager_writedata            => cpu_data_manager_writedata,                         --                    .writedata
			data_manager_byteenable           => cpu_data_manager_byteenable,                        --                    .byteenable
			data_manager_writeresponsevalid   => cpu_data_manager_writeresponsevalid,                --                    .writeresponsevalid
			dm_agent_address                  => mm_interconnect_0_cpu_dm_agent_address,             --            dm_agent.address
			dm_agent_read                     => mm_interconnect_0_cpu_dm_agent_read,                --                    .read
			dm_agent_readdata                 => mm_interconnect_0_cpu_dm_agent_readdata,            --                    .readdata
			dm_agent_write                    => mm_interconnect_0_cpu_dm_agent_write,               --                    .write
			dm_agent_writedata                => mm_interconnect_0_cpu_dm_agent_writedata,           --                    .writedata
			dm_agent_waitrequest              => mm_interconnect_0_cpu_dm_agent_waitrequest,         --                    .waitrequest
			dm_agent_readdatavalid            => mm_interconnect_0_cpu_dm_agent_readdatavalid,       --                    .readdatavalid
			dbg_reset_out_reset               => cpu_dbg_reset_out_reset                             --       dbg_reset_out.reset
		);

	data_batch : component avalon_batch_block
		generic map (
			g_PORTA_ADDR_SIZE => 6,
			g_PORTB_ADDR_SIZE => 3,
			g_BATCH_SIZE      => 8
		)
		port map (
			av_address     => mm_interconnect_0_data_batch_avalon_address,     --  avalon.address
			av_write       => mm_interconnect_0_data_batch_avalon_write,       --        .write
			av_read        => mm_interconnect_0_data_batch_avalon_read,        --        .read
			av_writedata   => mm_interconnect_0_data_batch_avalon_writedata,   --        .writedata
			av_readdata    => mm_interconnect_0_data_batch_avalon_readdata,    --        .readdata
			av_waitrequest => mm_interconnect_0_data_batch_avalon_waitrequest, --        .waitrequest
			i_rd_clk       => o_batch_data_export_conduit_i_rd_clk,            -- conduit.conduit_i_rd_clk
			i_rd_row       => o_batch_data_export_conduit_i_rd_row,            --        .conduit_i_rd_row
			o_data         => o_batch_data_export_conduit_o_data,              --        .conduit_o_data
			o_rd_ready     => o_batch_data_export_conduit_o_rd_ready,          --        .conduit_o_rd_ready
			ni_clr         => rst_controller_001_reset_out_reset_ports_inv,    -- reset_n.reset_n
			i_clk          => i_clk_clk                                        --   clock.clk
		);

	debug_jtag : component altera_avalon_jtag_uart
		generic map (
			readBufferDepth            => 64,
			readIRQThreshold           => 8,
			useRegistersForReadBuffer  => false,
			useRegistersForWriteBuffer => false,
			writeBufferDepth           => 64,
			writeIRQThreshold          => 8,
			printingMethod             => true,
			FIFO_WIDTH                 => 8,
			WR_WIDTHU                  => 6,
			RD_WIDTHU                  => 6,
			write_le                   => "ON",
			read_le                    => "ON",
			HEX_WRITE_DEPTH_STR        => 64,
			HEX_READ_DEPTH_STR         => 64,
			legacySignalAllow          => false
		)
		port map (
			clk            => i_clk_clk,                                                      --               clk.clk
			rst_n          => rst_controller_001_reset_out_reset_ports_inv,                   --             reset.reset_n
			av_chipselect  => mm_interconnect_0_debug_jtag_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_debug_jtag_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_debug_jtag_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_debug_jtag_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_debug_jtag_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_debug_jtag_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_debug_jtag_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                        --               irq.irq
		);

	serializer_0 : component avalon_serializer
		port map (
			i_acc          => o_serializer_export_i_acc,                         -- conduit.i_acc
			o_clr          => o_serializer_export_o_clr,                         --        .o_clr
			o_read         => o_serializer_export_o_read,                        --        .o_read
			ni_clr         => rst_controller_001_reset_out_reset_ports_inv,      --   reset.reset_n
			i_clk          => i_clk_clk,                                         --   clock.clk
			av_address     => mm_interconnect_0_serializer_0_avalon_address(0),  --  avalon.address
			av_write       => mm_interconnect_0_serializer_0_avalon_write,       --        .write
			av_read        => mm_interconnect_0_serializer_0_avalon_read,        --        .read
			av_writedata   => mm_interconnect_0_serializer_0_avalon_writedata,   --        .writedata
			av_readdata    => mm_interconnect_0_serializer_0_avalon_readdata,    --        .readdata
			av_waitrequest => mm_interconnect_0_serializer_0_avalon_waitrequest  --        .waitrequest
		);

	spi_0 : component coproc_soft_cpu_SPI_0
		port map (
			clk           => i_clk_clk,                                                --              clk.clk
			reset_n       => rst_controller_001_reset_out_reset_ports_inv,             --            reset.reset_n
			data_from_cpu => mm_interconnect_0_spi_0_spi_control_port_writedata,       -- spi_control_port.writedata
			data_to_cpu   => mm_interconnect_0_spi_0_spi_control_port_readdata,        --                 .readdata
			mem_addr      => mm_interconnect_0_spi_0_spi_control_port_address,         --                 .address
			read_n        => mm_interconnect_0_spi_0_spi_control_port_read_ports_inv,  --                 .read_n
			spi_select    => mm_interconnect_0_spi_0_spi_control_port_chipselect,      --                 .chipselect
			write_n       => mm_interconnect_0_spi_0_spi_control_port_write_ports_inv, --                 .write_n
			irq           => irq_mapper_receiver1_irq,                                 --              irq.irq
			MISO          => o_spi_export_MISO,                                        --         external.export
			MOSI          => o_spi_export_MOSI,                                        --                 .export
			SCLK          => o_spi_export_SCLK,                                        --                 .export
			SS_n          => o_spi_export_SS_n                                         --                 .export
		);

	sram : component coproc_soft_cpu_SRAM
		port map (
			clk        => i_clk_clk,                              --   clk1.clk
			address    => mm_interconnect_0_sram_s1_address,      --     s1.address
			clken      => mm_interconnect_0_sram_s1_clken,        --       .clken
			chipselect => mm_interconnect_0_sram_s1_chipselect,   --       .chipselect
			write      => mm_interconnect_0_sram_s1_write,        --       .write
			readdata   => mm_interconnect_0_sram_s1_readdata,     --       .readdata
			writedata  => mm_interconnect_0_sram_s1_writedata,    --       .writedata
			byteenable => mm_interconnect_0_sram_s1_byteenable,   --       .byteenable
			reset      => rst_controller_001_reset_out_reset,     -- reset1.reset
			reset_req  => rst_controller_001_reset_out_reset_req, --       .reset_req
			freeze     => '0'                                     -- (terminated)
		);

	weight_batch : component avalon_batch_block
		generic map (
			g_PORTA_ADDR_SIZE => 6,
			g_PORTB_ADDR_SIZE => 3,
			g_BATCH_SIZE      => 8
		)
		port map (
			av_address     => mm_interconnect_0_weight_batch_avalon_address,     --  avalon.address
			av_write       => mm_interconnect_0_weight_batch_avalon_write,       --        .write
			av_read        => mm_interconnect_0_weight_batch_avalon_read,        --        .read
			av_writedata   => mm_interconnect_0_weight_batch_avalon_writedata,   --        .writedata
			av_readdata    => mm_interconnect_0_weight_batch_avalon_readdata,    --        .readdata
			av_waitrequest => mm_interconnect_0_weight_batch_avalon_waitrequest, --        .waitrequest
			i_rd_clk       => o_batch_weight_export_conduit_i_rd_clk,            -- conduit.conduit_i_rd_clk
			i_rd_row       => o_batch_weight_export_conduit_i_rd_row,            --        .conduit_i_rd_row
			o_data         => o_batch_weight_export_conduit_o_data,              --        .conduit_o_data
			o_rd_ready     => o_batch_weight_export_conduit_o_rd_ready,          --        .conduit_o_rd_ready
			ni_clr         => rst_controller_001_reset_out_reset_ports_inv,      -- reset_n.reset_n
			i_clk          => i_clk_clk                                          --   clock.clk
		);

	mm_interconnect_0 : component coproc_soft_cpu_mm_interconnect_0
		port map (
			CLK_clk_clk                                      => i_clk_clk,                                                  --                                    CLK_clk.clk
			CPU_reset_reset_bridge_in_reset_reset            => rst_controller_reset_out_reset,                             --            CPU_reset_reset_bridge_in_reset.reset
			WEIGHT_BATCH_reset_n_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                         -- WEIGHT_BATCH_reset_n_reset_bridge_in_reset.reset
			CPU_data_manager_address                         => cpu_data_manager_address,                                   --                           CPU_data_manager.address
			CPU_data_manager_waitrequest                     => cpu_data_manager_waitrequest,                               --                                           .waitrequest
			CPU_data_manager_byteenable                      => cpu_data_manager_byteenable,                                --                                           .byteenable
			CPU_data_manager_read                            => cpu_data_manager_read,                                      --                                           .read
			CPU_data_manager_readdata                        => cpu_data_manager_readdata,                                  --                                           .readdata
			CPU_data_manager_readdatavalid                   => cpu_data_manager_readdatavalid,                             --                                           .readdatavalid
			CPU_data_manager_write                           => cpu_data_manager_write,                                     --                                           .write
			CPU_data_manager_writedata                       => cpu_data_manager_writedata,                                 --                                           .writedata
			CPU_data_manager_response                        => cpu_data_manager_response,                                  --                                           .response
			CPU_data_manager_writeresponsevalid              => cpu_data_manager_writeresponsevalid,                        --                                           .writeresponsevalid
			CPU_instruction_manager_address                  => cpu_instruction_manager_address,                            --                    CPU_instruction_manager.address
			CPU_instruction_manager_waitrequest              => cpu_instruction_manager_waitrequest,                        --                                           .waitrequest
			CPU_instruction_manager_read                     => cpu_instruction_manager_read,                               --                                           .read
			CPU_instruction_manager_readdata                 => cpu_instruction_manager_readdata,                           --                                           .readdata
			CPU_instruction_manager_readdatavalid            => cpu_instruction_manager_readdatavalid,                      --                                           .readdatavalid
			CPU_instruction_manager_response                 => cpu_instruction_manager_response,                           --                                           .response
			CPU_dm_agent_address                             => mm_interconnect_0_cpu_dm_agent_address,                     --                               CPU_dm_agent.address
			CPU_dm_agent_write                               => mm_interconnect_0_cpu_dm_agent_write,                       --                                           .write
			CPU_dm_agent_read                                => mm_interconnect_0_cpu_dm_agent_read,                        --                                           .read
			CPU_dm_agent_readdata                            => mm_interconnect_0_cpu_dm_agent_readdata,                    --                                           .readdata
			CPU_dm_agent_writedata                           => mm_interconnect_0_cpu_dm_agent_writedata,                   --                                           .writedata
			CPU_dm_agent_readdatavalid                       => mm_interconnect_0_cpu_dm_agent_readdatavalid,               --                                           .readdatavalid
			CPU_dm_agent_waitrequest                         => mm_interconnect_0_cpu_dm_agent_waitrequest,                 --                                           .waitrequest
			CPU_timer_sw_agent_address                       => mm_interconnect_0_cpu_timer_sw_agent_address,               --                         CPU_timer_sw_agent.address
			CPU_timer_sw_agent_write                         => mm_interconnect_0_cpu_timer_sw_agent_write,                 --                                           .write
			CPU_timer_sw_agent_read                          => mm_interconnect_0_cpu_timer_sw_agent_read,                  --                                           .read
			CPU_timer_sw_agent_readdata                      => mm_interconnect_0_cpu_timer_sw_agent_readdata,              --                                           .readdata
			CPU_timer_sw_agent_writedata                     => mm_interconnect_0_cpu_timer_sw_agent_writedata,             --                                           .writedata
			CPU_timer_sw_agent_byteenable                    => mm_interconnect_0_cpu_timer_sw_agent_byteenable,            --                                           .byteenable
			CPU_timer_sw_agent_readdatavalid                 => mm_interconnect_0_cpu_timer_sw_agent_readdatavalid,         --                                           .readdatavalid
			CPU_timer_sw_agent_waitrequest                   => mm_interconnect_0_cpu_timer_sw_agent_waitrequest,           --                                           .waitrequest
			DATA_BATCH_avalon_address                        => mm_interconnect_0_data_batch_avalon_address,                --                          DATA_BATCH_avalon.address
			DATA_BATCH_avalon_write                          => mm_interconnect_0_data_batch_avalon_write,                  --                                           .write
			DATA_BATCH_avalon_read                           => mm_interconnect_0_data_batch_avalon_read,                   --                                           .read
			DATA_BATCH_avalon_readdata                       => mm_interconnect_0_data_batch_avalon_readdata,               --                                           .readdata
			DATA_BATCH_avalon_writedata                      => mm_interconnect_0_data_batch_avalon_writedata,              --                                           .writedata
			DATA_BATCH_avalon_waitrequest                    => mm_interconnect_0_data_batch_avalon_waitrequest,            --                                           .waitrequest
			DEBUG_JTAG_avalon_jtag_slave_address             => mm_interconnect_0_debug_jtag_avalon_jtag_slave_address,     --               DEBUG_JTAG_avalon_jtag_slave.address
			DEBUG_JTAG_avalon_jtag_slave_write               => mm_interconnect_0_debug_jtag_avalon_jtag_slave_write,       --                                           .write
			DEBUG_JTAG_avalon_jtag_slave_read                => mm_interconnect_0_debug_jtag_avalon_jtag_slave_read,        --                                           .read
			DEBUG_JTAG_avalon_jtag_slave_readdata            => mm_interconnect_0_debug_jtag_avalon_jtag_slave_readdata,    --                                           .readdata
			DEBUG_JTAG_avalon_jtag_slave_writedata           => mm_interconnect_0_debug_jtag_avalon_jtag_slave_writedata,   --                                           .writedata
			DEBUG_JTAG_avalon_jtag_slave_waitrequest         => mm_interconnect_0_debug_jtag_avalon_jtag_slave_waitrequest, --                                           .waitrequest
			DEBUG_JTAG_avalon_jtag_slave_chipselect          => mm_interconnect_0_debug_jtag_avalon_jtag_slave_chipselect,  --                                           .chipselect
			SERIALIZER_0_avalon_address                      => mm_interconnect_0_serializer_0_avalon_address,              --                        SERIALIZER_0_avalon.address
			SERIALIZER_0_avalon_write                        => mm_interconnect_0_serializer_0_avalon_write,                --                                           .write
			SERIALIZER_0_avalon_read                         => mm_interconnect_0_serializer_0_avalon_read,                 --                                           .read
			SERIALIZER_0_avalon_readdata                     => mm_interconnect_0_serializer_0_avalon_readdata,             --                                           .readdata
			SERIALIZER_0_avalon_writedata                    => mm_interconnect_0_serializer_0_avalon_writedata,            --                                           .writedata
			SERIALIZER_0_avalon_waitrequest                  => mm_interconnect_0_serializer_0_avalon_waitrequest,          --                                           .waitrequest
			SPI_0_spi_control_port_address                   => mm_interconnect_0_spi_0_spi_control_port_address,           --                     SPI_0_spi_control_port.address
			SPI_0_spi_control_port_write                     => mm_interconnect_0_spi_0_spi_control_port_write,             --                                           .write
			SPI_0_spi_control_port_read                      => mm_interconnect_0_spi_0_spi_control_port_read,              --                                           .read
			SPI_0_spi_control_port_readdata                  => mm_interconnect_0_spi_0_spi_control_port_readdata,          --                                           .readdata
			SPI_0_spi_control_port_writedata                 => mm_interconnect_0_spi_0_spi_control_port_writedata,         --                                           .writedata
			SPI_0_spi_control_port_chipselect                => mm_interconnect_0_spi_0_spi_control_port_chipselect,        --                                           .chipselect
			SRAM_s1_address                                  => mm_interconnect_0_sram_s1_address,                          --                                    SRAM_s1.address
			SRAM_s1_write                                    => mm_interconnect_0_sram_s1_write,                            --                                           .write
			SRAM_s1_readdata                                 => mm_interconnect_0_sram_s1_readdata,                         --                                           .readdata
			SRAM_s1_writedata                                => mm_interconnect_0_sram_s1_writedata,                        --                                           .writedata
			SRAM_s1_byteenable                               => mm_interconnect_0_sram_s1_byteenable,                       --                                           .byteenable
			SRAM_s1_chipselect                               => mm_interconnect_0_sram_s1_chipselect,                       --                                           .chipselect
			SRAM_s1_clken                                    => mm_interconnect_0_sram_s1_clken,                            --                                           .clken
			WEIGHT_BATCH_avalon_address                      => mm_interconnect_0_weight_batch_avalon_address,              --                        WEIGHT_BATCH_avalon.address
			WEIGHT_BATCH_avalon_write                        => mm_interconnect_0_weight_batch_avalon_write,                --                                           .write
			WEIGHT_BATCH_avalon_read                         => mm_interconnect_0_weight_batch_avalon_read,                 --                                           .read
			WEIGHT_BATCH_avalon_readdata                     => mm_interconnect_0_weight_batch_avalon_readdata,             --                                           .readdata
			WEIGHT_BATCH_avalon_writedata                    => mm_interconnect_0_weight_batch_avalon_writedata,            --                                           .writedata
			WEIGHT_BATCH_avalon_waitrequest                  => mm_interconnect_0_weight_batch_avalon_waitrequest           --                                           .waitrequest
		);

	irq_mapper : component coproc_soft_cpu_irq_mapper
		port map (
			clk           => i_clk_clk,                      --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			sender_irq    => cpu_platform_irq_rx_irq         --    sender.irq
		);

	rst_controller : component coproc_soft_cpu_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => i_clr_reset_n_ports_inv,        -- reset_in0.reset
			clk            => i_clk_clk,                      --       clk.clk
			reset_out      => rst_controller_reset_out_reset, -- reset_out.reset
			reset_req      => open,                           -- (terminated)
			reset_req_in0  => '0',                            -- (terminated)
			reset_in1      => '0',                            -- (terminated)
			reset_req_in1  => '0',                            -- (terminated)
			reset_in2      => '0',                            -- (terminated)
			reset_req_in2  => '0',                            -- (terminated)
			reset_in3      => '0',                            -- (terminated)
			reset_req_in3  => '0',                            -- (terminated)
			reset_in4      => '0',                            -- (terminated)
			reset_req_in4  => '0',                            -- (terminated)
			reset_in5      => '0',                            -- (terminated)
			reset_req_in5  => '0',                            -- (terminated)
			reset_in6      => '0',                            -- (terminated)
			reset_req_in6  => '0',                            -- (terminated)
			reset_in7      => '0',                            -- (terminated)
			reset_req_in7  => '0',                            -- (terminated)
			reset_in8      => '0',                            -- (terminated)
			reset_req_in8  => '0',                            -- (terminated)
			reset_in9      => '0',                            -- (terminated)
			reset_req_in9  => '0',                            -- (terminated)
			reset_in10     => '0',                            -- (terminated)
			reset_req_in10 => '0',                            -- (terminated)
			reset_in11     => '0',                            -- (terminated)
			reset_req_in11 => '0',                            -- (terminated)
			reset_in12     => '0',                            -- (terminated)
			reset_req_in12 => '0',                            -- (terminated)
			reset_in13     => '0',                            -- (terminated)
			reset_req_in13 => '0',                            -- (terminated)
			reset_in14     => '0',                            -- (terminated)
			reset_req_in14 => '0',                            -- (terminated)
			reset_in15     => '0',                            -- (terminated)
			reset_req_in15 => '0'                             -- (terminated)
		);

	rst_controller_001 : component coproc_soft_cpu_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => i_clr_reset_n_ports_inv,                -- reset_in0.reset
			reset_in1      => cpu_dbg_reset_out_reset,                -- reset_in1.reset
			clk            => i_clk_clk,                              --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	i_clr_reset_n_ports_inv <= not i_clr_reset_n;

	mm_interconnect_0_debug_jtag_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_debug_jtag_avalon_jtag_slave_read;

	mm_interconnect_0_debug_jtag_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_debug_jtag_avalon_jtag_slave_write;

	mm_interconnect_0_spi_0_spi_control_port_read_ports_inv <= not mm_interconnect_0_spi_0_spi_control_port_read;

	mm_interconnect_0_spi_0_spi_control_port_write_ports_inv <= not mm_interconnect_0_spi_0_spi_control_port_write;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of coproc_soft_cpu

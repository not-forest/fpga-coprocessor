// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
UNszGcrioCwqxJO/0r+fjPGe/QgRalb+L047+oYqCLw83X3mNx+6A+yjtQuHhvsF
Orur9/Iv25WE/B1KJrHzObwjYnSKf80zlRu0LfSZUmjcl/J5Vo4fiD82SYYDnfPt
kgueNvBexJiy6nFHt9DEKel5zhV3sxJCeHM1bapJzuk=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 9712 )
`pragma protect data_block
xijLM/j2j4pTh2803AlJulo/sjmgEt663yaJlYfxJjKmeFOhnzlGwMiiG9ZMHRGd
VyH+JoQcl8YWZvFu83QEjGGouBgPPI/ndZMa2L5PnSULArTcZnIsQnd64GsZ6HEa
+PfYEmwPhOoUjQ+y7WdK17AdOHg60ZSxCICUyYHspXFcLueuYWc/ap+DEcHW5Fyn
shvQEIbpgEbe2Bi1qJkuPzNhMykzTSKjc6/Xy2U1X22VrOB+tGoJvnw7Ep2u1uOe
ugnvNMdMVLExLb0ZbevvsKpywqhKAz9BKDoX7O5Ax056vEmXlszP6493Y0cD7Oeh
BN531+W2dlAfYM+wutlsuUIp4VK1jt+2F0M0amQjHNKSKZ72uZy/jfIhfkskqnqR
JtPtHCESSzRZTz+nZ01IozEzJWHY6UBmOzHGDfHCU+Ex8b2U76IC46x84huBgz5J
TvilDGiRttdTQR9bg9m3MNcbkyvZekerYmQWm/YSrntrMXS3ZZ87xM+kALCwz6oe
u79qO+Hi5eCyMzbsR4iaki4AyutvVvw1Lg8gaQGh6jppoQWXC2eJbgSe0IcRthYv
6gMybuE3MA4HqBDwANkMfMePyMj8Spq7xKTT/p2BalCpV6Otm2Eahy5RLyKsjWuc
X98E+olJPKMIqjOttxOEvmS2s6NoKr9fdkV1qBbECcPaXJb1nvYd/v3FECoQHbP0
DpJ9fEQ2bWOO579iZNLOf8ftCn7pM6wCxTTX93JyR+2GMMK5uuWua6opr4FVVelD
rf5gSrbmRzjy6xwQgMJM8GCkFDbNIWQtVpOEy8MyHVkwlNxqfwnB3Um8ZvDWEx80
+gW0EabZE8yFfAPrQljsuJDP4my3vKYpIJmPw92Gc8eI7OsNBdsVNqWVQABDxxR/
ICzXL4Yr7UhJtuMBjxByYdHEDaUIAsJv6jurj/vHo7lEHx2Oh8vyNJl0KBfiEW0W
9j25QsLgP7CDDf8GSXSy6PWNandabOiFFr8jlfr9ortdCNzXLm6q79BcbpY+slrA
6Q3S8tyys0JR7a+D18hdSMz6USQpyo1h2gJfo3FtjSmDlg3Yd52XIas01D/ASeya
EPmsRlP3e1dT++7XIoGYD9qlZuGf4FmRKX+louOAvd8VggLnpPA0mznuK89IJT/f
s9XsIYNIPQv/HIQ/y8TB3jF+8e2y358UnZrFUycs0ueyiEUM0uy0KRiwe/cO4hsc
0/u8eJ38ioLSPvqXojKRYmJx7skZ0ZOBpHU26j3AAwR6R9B1TARckZBUGOBAwWqq
pItZCZiOziInZqYV1UxRVJpsPEdWt0SiYrSjK7W2bTMZ2oiPiRNKV4DAXEhyZvox
OP1MWKNSx9IetRQOR0Lt9ag/vLl7Q4vvDYD+bu6eeYroCOGcktDips322PNBAikh
6AairdrqpSwRftWMDg2kTvArILKDCtuPvKzHek/m5+jgrcdv3Y16HdFfCSytkCLc
11iUbfoGFjlMHQ8OgH+1FEii0MpS8eWGqWSjSmY4C0EKj/Ubuf5sb+c95P7bPnjT
xUztc3i8FJ56IuJoDWUc5L1HsVkkMLlAs6vGc9ufbyvlPUv34T8loFkWEu1lYPoK
NPT8+Q+iyM4qTCPnrR7n4SIIhGNf44gXfgZXbjGTSymE4h/T3Jpdv6RIDRp0f4a0
R2EsiJ0F4o/Ih7y4zcM5XYaxSoCsDKj4FS88bb0KY/r+F1TA2hgeX4nwRpNDsq29
GoizzgRlXD6RQZXFx8ewUCoBLcvzoFUGjtq4ICJToA29IZ0EvPJeVsB0VNEuXrOf
RzCgTHp34n5t2ysX7mtXHmMCKrNpiePRIay8Ib7O214TzkMp2JjcrxVZjpJdYxtq
ZnZ99uWgKV7x4BuR0nNVr9seBV3E9uYyT4JsXVARTJixVVGI8+MJM+IXWJ7lrHtP
8KPFjHmE6Jd4YpMsFgs5uiOqIqxneBo64AyEf8GvQsVVIC+F1dVFPfgSL5NfsMyX
u9t/6Jgw7cWDr8NPPgm5YSgdgYLjU6O6o/QQbK/hwNLt4sSbfN0NBZ1YfO3dsDqf
91akc8b6AEX4iA2cjXdhru0knp5N1tbatUZAJVdXwUaeI4S61oDhS35KhgZoUoXx
svz/82jCfxDxE2wtVOuRj6FrRICSU9ONJJRMuvYTECTEtGnC2qd7qOHspV4Oep3l
raY21r6QpuRNwc8m35IgrHgM1Vx37+SFZWBV2n1e8PQYgPK/aKLZ3W6y1ccJdUxL
kxKNXVkhdfiEU3BuxzI/hTIKcgXokf/X86TOG05Wo1LebZ0PzSQoX34rjlNbFUvZ
2VEBUG0ntHtwB94TZ6yto9FyaGD653Uq+Mj7sxyBoLikkyZlRSwZakeNwdxISdpN
HQKFwYIycWOqCy7wSoe0ch9CUqBb2JPjdJDdcmGL21m25UJUOcqCn8uPg5UK31Wh
6KX0AMc2fnrocrpi064KzAa5D6nB4CEkFjugMOYw2QW1/ZongucY+IQvwDxVle0C
hXqkdK/yIow6eZcXhsS7yIshk6IQddDpH+KmUO+gBn6OLjyLIv/gjcXyxoMVTWta
vUHpTBFlpR67XvEZ59s5hHoxmGNDqsJoJEV4uvNtagpD/gtzHTTC1I/b6AKJ1k9G
J2HD335ay2lfPlFEURMxsxYOZydyIXILdrRmM7LgZBiYCMR0oXYgB09x+j0ykNBC
7tQLxKAgWm1ktIzHfeGqVKS1yQ6Nseq4wfrxwSM8bsgZNohKiFp+V08Kp2lanvbH
XFLHVWNNCaG+layXwPejlZvssqc0PpD9ylhlc62XT1+DCLVqVlSgL1WIkDyXxNWl
r9PsOmGU01wOQNzdQlZgrYdXtQTDsw9C+7Vh6h6k6bqu9qGkF6u/b5cP5C9tW2Ua
YEkXAyV6qjcruCvq0+/VyfwVIwMRxAffpXRnb6U73e1FaAQlAfO0f2wI6fa+JteV
rN3S5UesULTVF1RvVDXU384mxtaoRnOSF1YjnkkyLXX1xvwmMVpEDZzA7cWE/Q40
zh2bx5LmLZjQM+4HPxSsME2yDL9bLo9KsG6EBOIw8d/aQ5lzXsq7egQ6EQ6iXGVV
BGfDkD+vQ3Pz078tRaHMd5hSIbiY5d/AtKJPF4YVrTobsjF7o+IS4VxonfNx4m1W
FJTgZzdZ0ujbvTcY5msSJcl6olJrmeRM080WEOwNyaaUU+Wi/CHLNV2w6PSbW7w8
ED66xVZqjc2u3Lm4m5zeI4EdJPCGTqrS7Y98I/q50FCRSE7gax82F/lhjY67K757
Hom3K64IGHfniPZ1ir2ahzNYHskGgmVp1Ss3TKlpgTJgkYySQy8+KshfHxpoSQrA
Olhhlt+TvLHGQxEGUpCayI2e6Tl9+PLAoPkzFNoe7wGX/ddY909nl2OwfG95ji13
R8EjwGe0wVAqD+EGaDEWiCRkEOV5ytbfgSyWYOMbY1asKGcKAkQaWnqoMdVZ/P4N
x067NavsGOmvBjM0mh9I99OIyBA95UriV4GpWJP2we7RciG6YcbRdq/wfyKkl4Pe
el9SPGFsmz8reJ3BYSXSklxqW0zfQ4f+6ZylMvL217kxNYzAkIYuc2VST53vWD3/
QwaL87BY5XKQtEqU0q3kdc/g68awm/23z2fWjSSYvoJ/vZyzlSrdjDPt2D6ZJl8Z
30AI7QqghkU0EGibdRvONb4AZtpHMbn43UtHaMeHbjDRK/L6X/Lv7QsP/SJy7Mr1
GTDuZMgAnuG5F0WHygtS3NpsmmrqpAUHVP0fQeDi+hRxAlqVEOXn+eIrT3OhmxFY
/XnsAlbMJhlXaZbEtcIiPqlZIXzzRjdM287xlfvu0nGs1pFfacH/cbuTwCxNSrFO
v0Al+lNKxlxJ6ueHwFR3+AjFAIB67DIvkYCPwadA+v9E3NfIBY/3xZAqJrI3LlYz
63tFWMPNOMwCCokWI7iYE4QpvRpvcCoRhVpvshLsaymxrsk1TJKDcnsv8PB6lLTV
f2j9qtfyJJx2WxylGoNjk4HF7HHHTer3XU6X/9JcauLDtP2fxO6ErJm1U1bsSidS
IXwB0peaUAqABXTfhajtR3tXzjMHxNqPKsnpDTrfXDEzKlRwNfwDY1EIO6ln5WML
R2YMGDL4xZcOZKcqwdj3nTL2TO0BjzLnqunq8zTAfKOrytyuYiGq0V4zJ/2eFndz
uQMFzmqs1UMDrgu7l3IroZLqTP2Xqeu7uNKNY14OXvHeyZONqGCou+wum8HFVSIl
MPbe21RcJEoj1jhEDdQ5wJE+Zl7Bg49MzSxwcdSdgeLpQ/ljA3mAscIQlBz17kkE
+u3A3X+q8+/9mDllfJRBAxl/n96fHaCYgzMhsFQuxxVEn0tXLfnvyIYjfAL/1FZk
+NO388rW+S5rVIp3Gc19rvD3q/2osHxicO2TKx4deNaO/CHLLQ1knYC6FUqBXjsU
5qs/5GmviT9wOFESODnEBSzBqdEYPbfF/kFGp5hedxl3eDrQCaQw3MHh2spZjF+p
ea8VccwXnAbwHvvSkXPzH6DzD5MrC5H7/O71Z5bIBkmNGx1DNVH8G2P0sIHOaH5N
avGUdZ7m8KyxgyW3L2/GxQ/PFSAVnrD5DHoRgHfmw36nsDTtkV+6XZlBf/cmC/2p
JNDlqAYfatel+tj027W+XG0sxn0mg3wcZKG12KcgQVWjrUPoT8zRYynDIFVtWhAl
Q/72hBFqqLFNxzTGRvd27KllkoJ7o4w339gvVq3FWKwtraT1IXBD+dAyuGvipxbI
54ZqouDHV+7GBOzrX+OUykcUCtOw69s7iIsjIZrJAP37X3fpqVJ+jn/+oXs634ee
zi91/eaZPg6cn+BiJYSwo8W9TeEUL7UGm8ATJZdLe9et9Go4rLfnktvQfQeRW64T
fv7z15UleYmFYVt6OF45rVhi0z3x3Ik0JnDG9dgwxZp34DQ22lI3r22iQQaDDx6R
BQEvu262YVo55H3o5Y4dzzhY4dig1IGXE6hsEE9iIqIYFBL87H3jgaOG98Ws7MZl
BpfvGzS3yocV4oOQujDzD6VDqfBpuAhFvw1RGNSsompkOMx8WyENjYAfRtiNxePK
OfN5ishKyCtMrwpVkglXkvyrXu/K03pWO6TWYfFXHnpjBi4NgHV8SWCmZhQBz/UX
O8wqFVefjfHpHg4qzTFQVlTOY/CDuFMQtzCygDzmg8ag1Z3Lts+VS6cWyulBy2NG
cKFE+9FhIRKBZk/9SiR2p4K8LYbubfysP7uZrfZOpoaoK0ZCUr2IMWp4wejpEOnm
mwjVhbLKF3fJxPPDFUECAfGBzRRCFCSuLCfISPB8Uhu1WRkD0z2y4r8bPOdmeZ8H
CbkcevCD816pF95dYYOhf12Qq2sxIWZRbuYt6K7nTulsrAylGT8lUu3AhgLH25zj
eRipav6yp6XF3QnFzVrqUi4zhTbIkbXwP2VPBPWMPKViZGTls22u9zNEzm6DjH+i
FcT4Z/FgiHGUrmYSJhzLazzgqOolqtza2+2ylP9O6CHgZSld7NIPIRbzF1so6hmp
f/tHwcoOUyCAsoHcQWEf6TTxqQsv/U+T8783ZA925jk/Sg6EQZwCdySYVsEYfBFI
sq/4dkbQh0dzQynqZGOb+dyq7AWZV1RmvCqkcuAB/LIfntW7s8PzFFpjEUL5bUi2
Dws3VXzSEBFDSliBa5Qy9sPuzBa5kpb90PUAP2AEM3kCy4HXJXkymVD/Ae7SPKt6
+Q9jxEtKDlxvWzaYJf64SW6CcZHKuGzlR0vEmXwDvQ5oGBOig2M8Q0ce0XNGgJ/N
e7T5M1O2b/JBz7wonj7CMSp4ief0bEkwcHsEloQw4UFLC9QWHpaIBGI5u/U7mQpL
fT2R1+to5XgeoLnpLkuIwypi827pOjlzEZyGWpFS21m74y7yhQM0btVRZ8JrdMBl
iE3hDunU7ndnFpnB4zKF+ctgy93lm2NKbJ7rxS6tjeHPr7F0vSqAbMtJ9vTZ1yYQ
cgagcsXyDJ9o5g9+w4PXf/wMHVi5U3B8LPjXwLC5K/pHUZTmxAnYR35tSmDd0XCT
n84wn7kB3Tsv2wPTGzICqRC1lX/RyCLn1PBkxh0M1HokXLTbie6miOoBe7c8aqWo
LoCRSuSP7KvsFfyyY5icK6CweZZpW2ShKBHRODdM7iRSttA8asAR6vqUYciDSoyO
fCfsq+4DR/yYZRcj7CCNeKgWaaAZRII/jqm9/Mz/pFd3ncempjVdC/T+FEMl41pU
aGK68t1R+rNDK14//mrSLLyYv4Ezxtek3E6dYyhy8OkLYy73Jr9qICoRn36krgC5
QazBeaIX8ZcLHwBw0egHNzO2tZTYRDAOUyoIB5GgZnBjf8hadgMkpqJp140yQwhb
TLlVqZZOEhNwdOWY0BcdPEcxYyWRgteCo91Oi1jmRsnd5fBoZaZdfyfDEcp5Q0Iz
iVHLC7/xvkLWpNKQmg8sE0ry/C152NjNKb5Fl1qZZw6ALB0KMwSI3GF8AweO4azw
s1i1ZxsfpolybXPnuPRWkKnbZ9m3v8zyblH0dvHsyh4St0Nv+Of9km9Nn8DiW4o/
6NiluTAnJKYZdiJ27nsr6E1FHCX6RPUWTh9YxicbZvtioMi5J8fjlh4IId8TFWxG
8ZKLN5m3WtSrNjdnOJqqLCdNOFnn0YcsZHkMvQsCclUGTHVaHT7EEmwWhu2rtRcp
JMhq7TxmARw31Hm8Qq6rl1988gY1bf+kVhZv9ssqOMWzEq1dU0mxbMMvFSJJQs6g
L1ozdolKCJs8Q/bhJs1v25W/3treAGgeSYHPvzAcqEBUSGSytcy7ZCMogzWIgm+l
ZHmMa8rqdZByzQH9eU0GD62+7RWstxL3oGhTapku6JVd2RBnovzJL4D2XOHfeHYz
obQ5Qxa15Rl2Ks58SiNYXgDzbe7Lg//6IIdgviC6s/DO2I1khV8BQv57j4kDh2Vm
wRPOcJrHrGNU3N0OMxUV46LjpzSO5vJMk/hyg5KoTc+FVTGmzpYzdgB0VkLrqfR7
yW5kmIMq/wFUa6wOUuy10RX3en3HBHITFt0HvmesMPL2uyggqeanShhBwfwwOjJs
govoRzDyTdskdaVdFOmc9LX2ryRd9QaUqgmKA/JYKDuDk1Hy7iurC3CxbateuTOs
3R4awxRsKROSzPXLBFmMF46AkSssY2AyvDDaCdS3JvI3LLDNseRIMeqRQMnKIQY8
xChXF/sSiuh9BpyLkHfuuYNagMF95SIN0X9SjZky7az7yVK/eHcoZSCARu2vxL3I
CTF/14TZI1o8n4Zzb6KipfSSuRMp6u7SV3HTjQosiDAzkaJ0z0vdVtT60zDjq0Gx
xs91GHC72ZTLimfUyiQBOm3HtUS/YQ25Rr/QcL4+dWff4c5RaYYhunYGAf0MWZfM
ReiTmgrvv/fSPTr5kujd23nUsiMK9uKDTLFzJCI01sVcCVeyz3Qo8CueynNCN9CX
8e5ypIuUJV+gc5L2RulpDvvuCa50/gzNCuKXWxT1M6+jbxsb2Q6Za1+9wlG9JRV6
mtpKmfLbeGKhxlg1JP+xKsyvoWWVZgoNxJe2bYqrZkrvxrO4i3unNpI2H+eAAnwq
wLqJLvPQ8D8Ca58+79/hqT6ZVdcp0wrYCmNe4a94f0+tkpoEW0yd0kbC0HrZ8BYC
l2we0qRczCRp/4S4JgUMFzZLWnddk8qAugrsa/+eMcicJh+NHgCAcVSueQA9IHDJ
YzQOCVhXDY/ZF0R87nssbgiNJSen/yDzKwb3Y9tHZv1aE75BvuWbCDlx0UeAiVtc
GsKQ+zt8BzivuhAImVaN5K5ZiMphS2cV/g35dsbdD85/4nwjJdIDRtIvCsXaCAMn
yZCiZsxovDQOMqpRmtpU6b+nLLkZShpeWqoEjRdc6/1fP7r4rJ2t+aaWZ5iKCwkg
P7naO2mlSBOlih3ERC4D/UGiq+w9nQOiEP2XN/2VroiVnIfMmuxt+hucEAQ/Udsi
ob6c2pT0Teoc8GF3y2FbP3kfEk4OaEPO4BPE5J86pHT/sC8tuG92donQnDay47AC
X5bqHiExbV6fCoHeVq4PEuGUR17bwEAShct08d3YRMtRflnsGUuhevPASMcXB4bk
IrXmVGNuG/X3LCKbOjtuRLsJT+NIBZCwWsc3HRt/JHh97c/wqp7294ZO11nIAM/o
JdO4EzVuqgzZVbVd6gf9v+hzwICjaEz+XTjiWoV+yyYDNdSqu4r4jchbEKTupjdW
Pifmh+nT9YvmmZYkA66TBiosI1DPRI3uozCD1MvbgbX1URCVjv2dRMify6GHcxtL
E6Y0o4JmMPeDYL5gJ43O+0A28GUUD6BlLLs2TlyyY7wIO59Gs8lGDqsDQB6kyMC1
7TALxE2PrrRQuaRWonHQ6r3QTHgMAy4LjL1LFkwS2dP9RiR2XnMT8XWjZ8464Mcc
E0YfdipXnAR2TejXPWhdh6J6CKTGRpyTH6OB7s9uUevq94Axtk2ggV2qXKbBu7JB
KbF1cAuM6rS0ZdNZFWQrFhg0RBWA/trnFLNQsQcvPrdipLnANNREt/g5TrpxUown
tMTMI5v8TUDZpD/GpkNp9189x2WWCPLV8vCR4IDyI4lsZG9zwPfR+N44JZY8yIit
XNMugydnfUGV5sWNjx0UjQqrcXI1T10gcZIpoDO1cbuhaaXtlduYSBb3qvgM37Pm
Fpp6+exT6AlXl0wp6Di0eA9vNxcm+5R21Pb05uRSN7Vxlf78rU5gsGUjxq1j9qgg
9H9LqAJFDBKV1xZMmASiZXbp2CMZwDnyTdw4SKNNlZUNXD8rILh07iH1mDNdSiUM
Ml7TRYH1RInHxCqPV+BrWze4F/MpInOVYjyBmygLn6Pnq+ZPz9/ud9tcdBNFoQ5a
WBmaJUavqa4nGMPC0yizJmWZUyE2J1Yg7Tw01RhxZ3hHal33j6oIkYekpYfQ3X11
5YgMeWLfAIBdHZbKEaMDVlmHsJeMhTgse8QHfnqcbz6qh05JqME6f/hwI3kcnlZy
k8hs2WXGuDCmIcc/4vbpx39OGxxF6MGFVqPlb1iFBwCD0Jh30DBzgeMA+as09HL0
x9/j0cPUHmeYgeC/vlZBnVggDyRWUKEvoP6KdgdOqZhOFgbW1JlW3vy9HbAEK+2B
DlQg5U28YxSWmvANBCpRoTCt3UzLRIviKFbVZGgIcdA5VriA1bNzVHxKMNRPeFuX
LyhWMexOSPrb+Blvcd5gn4CZOunXz8VsYWjwcRrtMirwElPQus8JoHyq7ztFDIkS
d2Fp5GUuBt1O6GahX8Gqt5Ajs8IrdN9uX0HUG/UBD+NwOyeOKJL6qA2ZM9Ft5gz6
QZ6GD06gYOcVjCRwjUmRRy9MKlMZxRaWuMm3qX+RiLPccjhGeVuftTP1MKNFPBNP
6PaAmfLonSmhKVYfUpQyRNwoklTG3fKCGxE3VmxDe3cQajvgwrnQ5to2r6rwyG4H
eOzcDjd3k3dyVzFPQbEc7zww8vEJcKrX8BieteTy7SLAbr1jrV1JcXeoCtCFo1Qm
wHVvVlPXBH7JOnRVp36nMS3HL0/qwItQRWZNqAuthbRQLMXPUt4i9zzNkQJlQslp
4+OgQkv5zegKNzqePCuA6ZA7rC0gn+vGLE7aMjI8rzx8mhLOG0VQQN+w3MJUVPGZ
BLbq51ncSgClOFKPYyKufECuXhsQktPBepYlHUY4ISbC7INngRmqkYRoz06mM6Bk
4vNaJkKn56nw3b9GrGZeynQojzSPTnJcwvX+xYLYaehfJ6L68KUNHXK5QmYwEBb3
tzNiC9CW4RrBnsuEdzwOfr00Xfc+SBKb1F9VN9zPz9O1YLqlNIh4SPC7zIJPNpdQ
JAQZkllxyLuwDHGYVb4W8+mTakTcDDrF5XHs44oxM0CVNIUeVyAGL1ZVLwRhbgEZ
c5gjeceqqtcgc/nEe5khg8abLrSITTfw+fEt2GPg8bAhHcIImR9VdH+t/icWxdaO
vfhiKbYX1WOJ/1625cLsaMNEuyWMtlAXHvFnwgZB5PPMUVPzRvODi8WVOLeMFaZM
IIYYzcX4dDuvwaDaNGyF+iokqQ1cWxdd3aq0aVUcI4BlAQk58FsMWx6weHUUMh4J
bvd+0a43ci79XDKz+8W8yKcGKfrA/8/VsTpzhIFGDXXQYNBmI9mRAQhl9Zwp1YB4
7XeG50xsYN+dPytFYRoi8Xde29E4bUjpgQsUhjvymmy8coNtYlNnK7S1lGv7bDO0
SgbMnSD9Y8mDDF+VH+qGE+WhM2pHc0t1YStXq3kcXGAU/6sAZohGujqUwQTdsWzX
5DjObkbXw83Y4vYDpUM2bGiWFBDeo/ZMC9yf4JAKx+eVEuhxYB/XgQQB/Ex2CGOu
o1NWt0+R+6A3X5yN6ZcJRssOVrmqTbagVVb2OtllOJs12aoRR9yCEGMfu7zDdynS
R6sb8MuyxDIj2gbXJWITEnZOHaYwFM979rmoJV1KmgkKXUYf8XrJhMpXwb320XUd
2kKgb/4FrnT4+O320BFUQiJowgmWw0AeScs457FAH9G74hyCpWWs47Ag/LqQ7Ivf
gxjYzCSxetQu3656PX3w+WZEN/hE4sBTaFN/NUQbN8GqrLDFl18UIAslPCUUCTJs
kFpGhz/OiSWKfI2caXdkV+zP2u/GvxlA0hGnYFSCN/WFhY4ffz56hzDl+DrfiY/X
nQSrHJY9CnGDGEuWU5vCQLmqjG3lGPgKL14+mA7/AwZL5LVirf921CsiftLmspD2
U2TYcZM0Y8n2avmb136FiuD9AvCJtLwMTvzLXUdlE41bCoXuCUDyd0TLBxlzo3XT
47hCGeIgfPRI8yWvBUEjkgdcCSJ8AXpItt5qEZ2TCJpIIYeeBeY+K86/VTPS0rab
9OLTVlFkJKkFlF76GGTO8xBFPDTj7hibx4CW6EhvgjHvFsvUtL1xdsVujybR5AHd
x0SokmwGcea2kpNABK6OFFYPqw1kjgswsn2Z1oMdOQfiCUU4noIk5qtdrElDQelO
w6VQVjOKoocaAbEhjnG8CeCs2iTHyQYfNMlWFl3bgFCfAwJJez5Mv/NbFSXMmY68
yXOyTG1HC8PWnTeysL/+iQhP6QZ2dZVv8QAbq2BnEuq2tjfzWOJGWr7MwWPUCU5n
vxzULoLXNZ+QeDMusz/GoXsJRTBUfXtrEfAEiAHV6EdadKv8sPWt7o7Z8u6x/wsT
IOzY5Z39t+9xsDaGf84W6/wAiaPOR1dBQmLaixXjo57KK50c+wlvKrhCXRkzEq7i
vbCv0PklE88aC8JET4A0wcc3KfwV4C+YPMMLuM+tgnCcDzQLppiHtBvx2Y6z4pOU
OmXC7+7crQCcd1fc7jswfRVwV42i2NVP5+6rXn5Yux1YAvMuUJuhD1s49OLQDvTZ
aq1XWJn+1VngpoCwjf21Bg/CP+XGL+Huy/yMhTnWxsAQ5+bl7GRP6WZwqvzleydH
aolix4cQGxHVXhEiOrW4yf4Bsx4rbKJhDmydyAWQE5gxvRNXC5YWLPAw43UZD4SS
tE20GEpP8hcZK1SJ7hsrzL8zErIDnA9OZV0QZuu4fLKV1nnM5eU3YsXoZGa4UrY8
F1MFJiPm6UQ80H1Umz3Gz7lmpYWwClnpOSus3U3yafoxlKL/1o+KG4PvpWI5AY0l
v4eKGMWuUj9SwKg2Di0QQ4P9SJ1l+IcMsRTX7WocXyOeHSfeyW7JvQ9tndQt/Cwx
lXbPYdCTDH7cVpqCSNMO9ORh4RwtGQmLPkcJff0OBkffsCig/MjI4MgyFvHro8up
sTe5EaplMmxgnQj5cZwQNt8iluuBSp5N6CHtQt8qLrJC2vxBCfn6zBeCdOfhef3y
09KUjblNlf6hS61VrUspkZHS2kobPIfTBEh2vEGach55w1wfWDVhk9TYoNyAAiax
uDfV+XxN16acja6Ou2tflgeeqIi2EC2CbxXKmT8K1JHjz014N4chxUWw5Q8y/0lU
d6Qyt+KSpx10JvjrTdc+V06NXUQivjXJryi96mEhW9GCZlCbZxcDG1hxBnlj6UpQ
0jWkuTTSIX1Bl1XDsEUL7dz5AodXNuhkq4DpoP7yg7GUusehOXPmaxwwg0QrTeU3
iccI1lH4RXOBYkm7ua3XNV97nyfKDcW4fJ+zVbisUeclZeKzHo4n1BlcpyXTpr0V
Q7OqBYMi/POG5uU4OWegKiksbAnVsb7332Q4Esps377pqxrTgNIse1WxJXmL1xJw
4v1DWAEjTv4xRrC0VsCQZpyGgMHZ2eLvHzv/1FDx2gwTwCg7Q24u5zinqUajpul7
qio4Tzof39BQkuBK6WBka6DPIC9T9s9pSQjV+SAdF6efRTJVvDrPDi9GgPDJAxCG
0blHogwY4jwaHErttsBwjLRvMiSdv7NEYRZb4OmapD7urZxuIhJhf5zqpDMxZXiA
voOu/w3zINMmgzWF1GqHBExzaBXajKUsHluBufWHf9BaYSxqy2X4dI9bePbwAXWG
ofXRS0ainW7GY8BLTW5vetGxuD7eIpar4Yc4VKcJ5HeLmljNtswTmdKoB4AVZXJP
6Yt63zSfMNIl81gtlZLPeNO7VZ984PYjWfLWeITr47ggMd1/zInINUh5lILDMn5c
RANihxyT2qSAQlE8blObKWh2ngX/ZGIB1N8gy7E6wF76Fnk8rlt2TlN3AO9GIlDl
cOZU5Blqcv6XBJIF/xQRVTyrPM6DcQBSjoWBYGPPgyxdI23PNS3pFyPqohPX7zHU
1SUtHYUWpoHc1RY5wyl2Sqhq19th51O9Ok7RvuHy4hLuM84hhsW+KLCG+AGf1dMZ
AaHO9psDMnYYcboeriqMgNaew7QsmuVKRVTvFYH8GtOIpIzmhOfQ3ORE1jT1rx9T
R5Wq4FY1CmvL5hXuZEpQwsOSmT5TXK4dch80ynd4sM8NNa3S00lDwXDPjVew9nTa
z0nZyF5DpXOE+r/CD4l7VtaGHR/3Z610WcHd1t9ZJSoiK98QMusYRw1O47Rwhdh1
ruYkMDE13IPbndsGHKrC3g==

`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
X23DGGiWiJr8PsEEDQaGBO7Rh8cjyx0UFtidX61UdzJW8MRWOkNA/q/3s3j3MHHp
fauUrdomJ5Rhd+AsF4/J3U54Xo2Cjjszi7TPsoyFzEhiTPlgkEAn8loBgBZznVu2
Y16v+aiQFj8u8GgKs5A+9twaTKrmIHOKCp/rMh1jrCk=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 12048 )
`pragma protect data_block
MZG04rQT+bb/Us/eRcDQNF9oe/9J1FgJ43Sp0b6e3gFdUwt6bLpbqnZudYX234+D
3haOrlfhhoZDbRgc4P9bswS/n4pFE5Da6IN85gOKRk1NPPmlWxd2RQ7Ok1S1Vaka
v9xSTLUJtq4V4kyXLXjVDGQ7oeOXPCZPZLIm6vNJI1BVhyZ94HreKB91yjxksr3C
UhAlBtKPF6yxnbARA0trK0fz559oQMWTwWjCfdcJrREeOBiU9vbYpHwvmqiN7L3F
gLZeVmzmhejprAReKSUfsSSxwHU/WHiDpZeOQFfXwHGLD7Z+gaUVOi381dgzst4k
izzSFBKEzXWpLLvAnvpCjBEUiszChJV+o5DPYJgr2ctUipptTC/He4djMSMnbNsW
WnFsQCzuKOWidpTlXohZaMZu/kSWjpBjShTebivQJsz5KAlxBAwhRRxCORjH9RCl
sx8O7Efl1iutb/ZdmW8fQ6QXpdnUF4NaSLTuza95tL6ya9NeBNYPtPezDkWrS2n2
gHEOTSKSka8owp2Yi8qlW2L2GHBxux3L0PH5Ffz8194a0DhnnfVpBMdU48IQUjB+
1LcIt2lqAvaRaSjZAwNCDl7t0LmL4sTyfrmlD+njZ/Of/eO0NRu/nYMjjByri3XO
J8P8qZaftEnVtlYPwfPlcLyTufuL9nYNn4Y/B/Usn9cjYM5PVVTtXCoAtdmyV0oP
COc6stC/L/m0o5oVcjw6Lm9If8PKMcjMOU0SCo1B+OR4hoOP9i7dc+miWPW3/uKn
uJVJUIZyzYvcqIAz4auzkpe3rPZrZpiw4PIQkyace+9nqan876WHiSu7mumOA3Et
7Zf9RHVkrHQQVucs+Wg78U2Cxb5OfXarFgWd/oK67qvfRu2JPpgu3MOFsPnHYF7t
esb3Tq2j94/2rzD4WKI9/gkfgmRSghuyo/Fnob5UIg6FqKVU8pi+7mFRzoSMRQU2
HXaO+aGxnLjFZNRDpGG2VxXjtySfi8dKlFDc1HFkHhxusG6BQQz7gGKIC99O4qKG
mQBCcbrJIhTzesBIhHSAy4317BFhkR5s3e5j/M6zDaygcPxuzvcAwP6HGpNT8xX0
NclwojDlkQZIrv4iSRPLIFmVuqsOZSR1yyvKXgld3TqhkzqiAI9Zk++siKCtkw8G
ioArmvGKLzY1h13JymdTW+zrj4jg64k29vG0VPbykNUe3wT+je8FO/iyIHbGXFHr
YK0Yq6TJzCT1/hGuHhM2Tjd8cHh7UInlDyQ6PFK3/nLMc98GFIGO412xTL5Lw1KC
GBzhdtFS+rv98Ni5uLjF8RDSBAyJJXSI2eYruxhM97RzDC/6mfVkJFWCbTKKXGqI
IMhRx13w85EzDxZnD719DYfviNaKLU/fS32ZIRMy0c1fFtHPB0rJdMlCq1Phb65z
snmpzk3/Ge4bwnMAE96PTM3vHAKuZNoqFYYojmlXkx35Z6CF1NXqzy958MlwFPY4
8ox9lGRRbIEg7w813NYXKuQ5xTUKx91V25gft5Gi3zdZ3lJg6WHi1apStq6uP/iv
s1UDITHspnLTP3TW/ZIcrMMUtLcgrBOY0WMoLHNuCi8/t6ntFsKxLVmJdfDFTIAs
1QARJxGfb5h3Gty/W4m1ytQSt5agTlloob5NxZaKW5LlTpgqww9BWK18mUG9g0j9
jtXJJl8T0Ky9WuTMx7QC5OmOakobSWhOMRGORBmgUCQDp0fKABI/ff8HW1EmueI3
s9bEPOk/CBEBfddz0u7KFXGnUdimunB2oLyR+De0CbqSB6qjeXKOCpDgY4jvfq29
QdaNpMjKzvpdJ1HbBFOz9B2G8KfqmJuA/x58kAk5z4iY8gCJ3P7Hm17ROtoocomR
gm3MfNQwS4f1KhtCtvaqwl1u1xSggFl0oBtMUyzbKDiMzTP53hRHuRKbIZLridfQ
Z8n7RkqBmxBMckTogFmwuM2P/CSmvdk1IN0+tWDsW+IrBIcdEg+6Tq+Ss709Uyvo
AvgzviqUjZSniTBnxbf3HfC63CRkIIo/3bqVi+oaL3PzyVF1Ch7WCdKPsYRkLTDa
y9PM/jwD7SXT4wPdxQ9uWGWfDzT6keU8gMs9McvXIiFpowRT9/9qlJ4+9vMFjiXw
BWEiyb6ipGfuZLd2/Bjrbpp7Dtddw1yD4LdKWOa5Hl0K+bgL1YyaFvakpNz+3y1q
L8s0XUdKP8EheAnLm7sBYc+1XWxQPBcyZqkdsQhF/CQ9YThw+7SVKsLvU/HCu4mS
n0MVYhRi9Z76515CuHIZUnDHAIXLfw5D9O/jDA+hFTDsrN53Bwx3wjgeZpb7/kkf
tKDDAwMWcys37bKjWTNqM4x4IA/PZZpmWUAhJ6kWXHzD5g7ZxYodOHkobDTBdGhz
pjjXRVG//xGZMzwn6zZC2BfwkjR0t73EETGZ+lMFMAgjx2fI8LV11LA8uY+aHIh3
i8pSM6tcoyItagY9zTNkoTDnQTV0PoaHsdyRdl23QY1oUDFKIAggF/6qU14+hf69
lETvR3WN4l1D2YWESGignuuDyBzseMSw9SIUSTMtrETDbSH9Ho5IhSesxZ1EeVBf
GcWIIyzqY2MooHCyjV+DxGBBqql65eIhHdC7e6LYL72fv4ItGCtcWbSlFq0hO3Xt
M4OmIeVNbZBDS/v+hK93y7PVnv1/kC5vUBiWHg6k7On2HS2jMbq2aRaqFOwQdejL
EiYY7KApFduQmYmT5xaeKu1oCjvnzF15SxdzwMEGjuHNE3VFQxAhNECU1pOdoji0
QLsVNsZ/2zI7OwnMBtHSuh8ItjmrzMBw8o9v5HZvbbrla2rfCUty53A4Rerj5bkV
I30rXRnbE0UEoghGYhZb1iIrj7z9dB6hSwgSiTTUKIq3VfMPUbWwnWPzap5oXN3n
NzDFbdsGlGsXjY4icJjYNJJPvgSceTqFSpthr7JCfcEHFPArVGWmLr4wWm2HBIDI
SNoDASzbF9LJWLsWmtm5U+d3k0pqTDrrZ7Lrhojh6AJQ+MwP0f2Vg3E4LgRCNFmJ
o4Sh0c0zbozenq8SBltG3+aQfThNmZ3pIsK7L5XAC7GTiUA/gayRNbz7vxeuXqYp
xSRNYBcf7jTzexdXNrqATJtdouuncX7UnpPgcE5r50q4rsVLRCpzWj2kQ0GGHBCE
wL2OZDGJgzaUpNlfT83/TfxOX5P7yZCIHU3rB9EvCfA9JuaDbqynodcEifKqlI0C
RHKTNjVswUddAQV668Op/p4jYrKJFi/qUZaxpkyFBMKkTlIiiUePnP+P73UZULgo
8vmLE/eQk7fO8TC+gLZzyyOb4Li2KSQ9wOBuTlMzwvvWVe5lsCdend0pYQSj7Gza
IOwTO5iKQePVgNF+DJ6zmJ6TMqsIg5be0TZIOJqTXqXumVrYhPos0uQqUuQzQnD/
1cGiQBvU/hHPeg6+qtKU7TTt2lSMVqeQZ/5MhB+3aQf4jMtmZ9/a8faWAXhXcCp3
r50VeF4vAikcbVmVCb0hhseQE7qanNYpUjU61l/k+GCuFv2PPVWShKPTZsx0rFAm
B3ouZMBEVzFwof8KeUYXg10DxjuMAfglFHCmAMeO8SzDlsHI/w1sGoDVSpmIWuNd
0RSUxcUMv6F9FxKxbR6q0anfQcFf45hbem1pXAe3iqbrpwbLsvcG4fDMxrTw8/3n
XQh+SI6v1TqRnUXcHpGejMd4J1s69WiEYNFtrHy1hzaDpnSFTiSNXCavEMy1iS75
ztjzvWo+LBRu6O7nLKDJ9uqtEPf2fkHcI1JpsoEBL+C+RDJImZgdtBaOoZWGKonZ
GdXQXjMmlQwjL7WyjJj7N1AVwAZuLa+5z0eNooFTRK8+RYIJyVk9hNvKiNvcOd5a
QAPwNLzYlt8PxRfBB+r01sUhnmcZx+2p3rcyExfDk96SvoVjmzqWw+dk1J8v+CsA
PFQqjSa3hoZS8BMYgfFAXZi5NxidOaLJuoY6Cuk8XoJeMSZlUNSDIA5aISGdru+c
nKXuC+46u2dzFM5syodisWMRpfUBLWYjgJ7kvgOniR9GvxltkRxePDxIVV/XSNac
RV4ci3w9lzv9M8LIWLTxqnlFz+GRE4im9gol73f1ghbNptA5EsHyXHsGhDLIB8fA
6KoYsq+cr+WWs5O+GhKcjJPZK5LoCgK8B7zj9YzSCziVMJNEtuTFDOXT+pyDvl4N
oQioPnscye6RP8a6z3AOiBQtGKrwvN6D6k8q0MZOVTiIlOr8uN5R7NXyT9Q5fW49
GdRa3yFaQyjM4fi3qh+iD6pzw2RnmiZo2P3HdUpfQXafenA7IgqZk1EJGl5o5o87
lMNStGV0c+7BwsfpQf6881EkhZnVMWQgFbDyypmnHl7blgY41BbsNJxEtcADdEB0
DtHcfSOxutmVrzcB/b9eu7Sv3baZY/lS55YISc6B/64Toc2QL623RXc3eeNf/5IT
JHc8qnA5GfgsFlEL8R0zukUIAufqaXyaI69PYj2JNrHScyIHEQXBkhuB7wBDs0dX
/cdlostJ/4Sv6qNymX4W4avlAcbF1aWrpMTaS+StbJ0a9CaSZsfeonnKjQJ5jeKo
cyCjaWca4BLBKK1JtfcROTgVxjd2X754K78U6Qw1ekVj0lZxRRyRdd5DmMe4bhFK
1m6sliEAQuH1eZaFCKf3NngCvESDjLplzViZN+KrNkkxzXQm1tNXHLRJSKhWs8Yh
UTGgZrD+RAF90xvTtvoj7+NYWrT4MnGkzYueEJEYgU9j1/VKzcY4bdP3NzOTrtX9
uIfvcqwDEWL2dfYFBCg0owQqzBYJmYxIssvs/OwPPM2ckewMdHGVDqH4x8pRxEzH
zMtPEo3awD1UsYO70OykYS7Gs/B/ZVN28IyhADAPXscyOxiCso+K/xRXwC2szjRT
5x8qQOY7yJP9UDTPU9OsbdGwVAx38CIcr+IdwByDux+CmBBUnnEnfsm027xkX8C3
dbIFrse43ogMn0PzHynOSYfPwM9enR+YDCRxBo/dhhie7baRT+p7Kmlk5G/epH0/
wk3BoAuSWbuR96gaSUDHnl/FOCgSWUoIFWYfPFrewCvvpccnN/rLmcLRlHaw0VCb
DEQu2zOGYAOduPKGGZgz63LSpfWodnNZS19sklienJGX756Z8t/OG6qpRt4Brvg/
OF0y9TQA5T37rs2g6rCjaDHAKDW3iPz1WAM0h7PPRQLOXUj2nCLouNgHPpGuo6DQ
56rD4LTw1VqHs92QPHvw0R6I8KDKpmedTw3h+/LHBR1c7xFOl0UMSejSIHtq3btV
K1VGLeTCXz3MY0ziSOkLoiciF/dqnCG+fXRg+cOFYRWKBdOaxe9vJAVOczsLD6SQ
1CV0Vdg5EkEaa6svV/JRllIcCQuameMTbDdDaxVr1tjAPKzHhLVxsXlX/KZgXrV0
yRH8nMs+kXvYO0Kc17Su2zEqQxA9A1t72Na1Zd43QlP0Io0aNJPCmbvQqXGdUy4K
+T9u2zKw1CKxqY/h77obxTbHo+IBHv6XUOfqEJ+cMTBNdDBQ5lcH1irdKYnaGKGI
9U1PCu6+eesbB9vVyPw9YVeGk2LTOuNxjqqI6P48RHnsie6HV+LLgG5VTMzrQnTv
TymXWpYILiaKmHaInDMWaYLXKeTEu/Rk2juZ0aT5qPJ6AvjK5ZsxAcPDMliQItzB
aclBky/n8zrPeWbv+XvpFO5yacCc2ZGEEogbacBR3xKQIqC8lIe1JS4WQV3Wu9DC
wgFnpxAg2fSkkguJK9tOadDo5Hx9PzxEq3YJEtVqTu1NRFu604w7hl3tpRjXl8z4
emZU+TYuRcdrglos4Th3YjtNloVDkZPNmlaf3YUT5iHcgRn5uonk4NMNYGiFKMWG
Dcbs2UXF2qzWZ209+ME4tuZcnFrnV7UjvXHv4niAINxgwy7Ykfo5qTqfQhBJcNtR
50Dg3UX/+ShifjDrCBgWuiFR9htcTb5eTDJa4GXozDKa/X0NE7i/NT2V5iX4lUAz
dzfcN94WUm2RQzxFvwa9XPw2/NlUjDyM/L53GDMzIFmxzudB98Lw/UWEC4AubF6q
obMt6UHsSYmv4GFQWEUXcK1LDmNU0KvumRgBHr11uGUOoHpRj18wkDV93x5PEhHu
WWecFTkhP4Z1Z4tHrrQ1UgNDDVrVbjSyXn+Kh6lIAUEhYnMh2FxcCgjLBX1Bufvw
u6J1ZOxnhvcsEzl6TvcNctX23WX/rUqSMBKmXBs5QL2h35iGqVr6VcRRNrWJXuYV
lXYmp7yWE2h0fkMCv5KYl6shgSk2xF32xBHVFZlo8S1UEezHjTMt+oTdOIliO62C
Dn7TK7HaDRQImowY/aTs59sux7Q7a35d2bkYZf+YQV6FfY/jVTOHx1xvUVh+q2mf
4FiWms7qGd5b5B/qEuIflc+S7LgujrF8Df6UeLja6eqw7r8ORytn9388/ea9nE4L
3odLuDugIMYlZ/Z9meOS7DH4Hv0FnOpzZr8tqsvmVxygUF5TjX6TW5u0cDT91qUR
7vw+0bEVotyCIGY5ZQVa00ta42V3yTG9LKliok2gO/Ae9aoTGx6wnIR0+evaaH09
3tUixOrDvuMtueSaEmMifhP0+FGKVZNM1Pz2zKNK139DsTIftSDBNNrro0vzfW6b
UeVNBCLs/zLKY8m3o5W4wsDOaU8wf1qpTvJ5NzDyjs4t9DCPadFHFwONj7OtCeHY
7StjA8sRQQUv3s0HXPp8mjphVoG43Evvu+Dpi+4iL/9EhUgkH6U673e/wT+bSsGc
INaeBus3lwokOI/LiJpR+S/Xtt8FUNViydZIcdbjDOqSDEhvF5Wq4g8by8faLdU0
QYEUpjzsdj9KNiNWVipkA7MX/NaoDo4hN8/DUsfBIh3YxL01taeY7F2GOtT/jg8+
8K/WGBFDkD7CZJRRy+CFtCUQBk2QsJt1VJwI5icalso9GiZbYWz/Ke4jB7z62Jei
lTuEI83WbSDhI+9FIAp37kzWaRNn7fp3bdGDBR0rPWhNNqS1QYvXro6DdKKTuLTN
xt0JNJUiNJaR07q3ck0dPHCMxyU4kungHUAYUyrr2R0iiw2SSQyO3kjRPpCS3oGh
r64WoCiKKQf9CHrzzJ0+41zOTdByIRYa3ngi0rFA78U9DXFA9zyKr/ZEkuY+xwpV
1OUJqqhGT6TSW5htZhr0fu1G1xpR7LPWp+A+klUjZPmerXuVQSPgtmnRV2+l6pf6
gL7NV1IaEVtc/LJXgR7gHwmbKqxeaaUrz5uYmmkH989FxqzpsR+eFzV0WKn8IhnN
EHbHeFmeYcpDDRKhvxcRjAyusQzXljP9zh72vFBIpo/xfIPBpZLIC/Cob72UUSj8
F1aR5nEERsygQaSfmjIlFSZx/bobauZzoRbjjZAYNi0faqIMY0Uuzg93Vk9amPIr
B2QBqzSaLwjHO/wxeg+mJngcgo/ESVAhURv8oCFNh7oaAsuUoKyJSJYYmnnXAnVt
odR8MuET5jewcpsBCKs6XAhZ2026gf2tFQxfIr1LwUbWKEkwErbsDSyW0oonj1pR
5jUMXX55NKVX2CyfWdR/iUUWSLpjL8wk/vHZBlmU6btHGDhqNMxYw2jyN3DdOu8E
ZQvlhQzWjc8DnMx+48T+6cOF3wQuro1/2irt59bsNQTWNV1KVO5sc9lvUaB/UmHC
fYawvJp2/lDJZHAB/DqK4yyQVLyYj+UWjgAD/F9dclXWEAmSdh/ktnBG73QUR8ov
LMWpTgZyOQL6Rnh98Cm+w0mIP/mHUNPcI8L9VSJeOJDk6SIszYRJid8Q3PmmsNI4
PP+X9rRvHxwpZU3bATfMvgqgt5rR6yknvJPuYsr733SO7KOfaOULpSXWJynnxAdF
pwN1RQrwbRA/0nD/x6vuO/zRJnqAtea9EGkKj1GZ2sCbRWzhXf1sbq1rIjVJBD6S
TCIqanEp2XQ0N3yNpowPbVHadWwlDVzWOY2KpY+hwMnjF5yyD5bJypzYZi3M5FrT
yZsoluTviMByx+54QMmgNdx1oMgdQbJmQ1nf+0Qqc57NjEVjcemkdsbpoEf8YrJJ
X+fXTYZMF2hPYyMnUWwL5YU+Qklzg2AvmrGVGR0PqfIk2vCJbKtwFvzXcW/YwKT0
q72EzLNC9eELCUFPmowfP/fk8YQPvj4YefFXIIYZdCWDJ2DY4Lag1NwWfnU2xYOy
aaFqcO+HzQ380bX6gwxv1UVsHSmWrJwBysX1HJsOZP/nKq305FmVxZ/dhMu/opD8
gMj3JeYSBx7MtiZSFmp+Z2XtU6+mLFyWDat+oSJJ28O/LJyk0lAIOjFxnMxok4YR
+n68Rbjc0jkjFBJFcYIbAWdTYtx2VlprVQAK9Nv5Z/g9n2Cj4o5XS6giUAcjqYoJ
rNYgrRrilaZz8yAfwQEfI5UOaRwaKDfMObOppOvzYHjuSj+rIwO8rL/hLaQ3ArBZ
c0+ix+RUtiJ6VRZo/n8n04xEA5mKpMVR6IohPpjqlM/pQ9jWPZPBcC1FRMrwZAI1
hRaRQk1t/fBTP3hiif/pvm3V+mv5eNd48ntYanoyKnGPJeCCq0TdTk217twZDgxQ
tTjVXhzOuMHDmlnpBHQbA8R/LSPKquYQDi8rfOQVLxlSEsVfH0v04yaweZxY30rt
bs5jCX/U905yqzXxgJx4uW5wmX21IpsHyfjgeJodO32l/osVbc6XpgE9p4O2rHHH
iuaLVrAR1HLjAVRqmBdkSmeriTw/xCWb9TlYdz+NXIfpfyokCwjQI6WVhFES5dEm
FCCNkQyJ3EtyLrAw6vQv+KUx1i4JV2t2IhclHx4wi9XWfOf+bL5xhQR1n5KXvvWD
a3IN8pnhF1t2fBoC33iY2b0kW8zLSnU/Hkhiaf0Z56a99u06J6909K7r+bKYkWI3
mnAPieSMDycETfsBiCLD0iZdBh1sxYWaSJGS20U9PDPdts6KUbcMrVwUAzD7GI2k
A5gUAk3/czN2w0bXHNUcysTyC0/1dDxSsjEOGl/gGWbFJLWGnzgLm41CkcXJzqMo
TFe2d4reXpLHgRLRf+qiKx64bBEEN7waDsGELUYcXBgv5vpm39KH+cT4/R8okaUh
BsAX8tX45S5ISEt+Rslxi8zMZwjQ0avdOT3UwHbTMs0iRTJ7UhaxzUQjbWCLR7Nu
POxqIxEMt9lHnRYeArMRQDEwzh939zmsAa05SMLesdv76K9uHylA0zhF8rXk2KlS
C38DZ9PJ5LjTD4/cNKMupjYHZkJBiB1zorNw93LiP4uCTY1m41MeWuaFnhlYGMOD
V0rxXI6rf/0ECiSdzH7lR3fRBVyFsd+BgDuTApnte/sZv+dMIGBgcREORU8ub9vL
nFexeMz7lbTMzO3cImWn5oYGx2NhP8BhWrIwazDwgeSjSId+YyoExfH6CaRLLv5b
OhKIJi8b7OMSNWFOTwwdI9OMx//gzdFFAlK65/w/IkRilClTRTJc8tSmX2BjQB3Q
gbuFvxAA6zC6E+lkKhhjdQQX2dREBhZcNlcgUwy2/A2G6aQ8JJwz+GN4UE4n5B+3
cSImp6NMNjroR1rXH9H3rwhVQn5NoLu72SCEHoiSO2OygRnEKyr/XtQHK1xRV5WM
1IjydprUkCWpea6RNBetTeAVeb5ut8prmFrKFOOgeP5nUGxTzKXPFmnxZ5plRbfN
FPpJk6scysxzgTnVe5lsLXKx3Ck9Y3cqFWz0/tGIcUil3hpxjaywfSjd50VAqk5a
NXMLf2lWqYTQXxRnoDyUX6G8qRmdr30HkhLKUsOydnVuYt9bG8Fgihnn7n0H2sq6
bHmrEo8P08btMrSRyAQX2SAne7k05RvRl0yvaf2JnPyl6Wo1TrR0KIesFEt6c7Gl
94EQpQARe0aPvAVBLMUm/B34lD0d2phxHByz/EBUeU9p7YtNJ6T/v8tsKQ2vUmgV
4HK/uiNkH3UrQ6JsiZ1NXXaNW02+qYWiJHjLr18U2ZHN63zm1DUOiUEC0HYvL834
xMyzf1mwuTLNvyRIi8WcMtbO46sbfPgDYg30uGXymZa6ezvkg1Dh9HCilswDbcRT
I8AGO44HN3n7lYfl7Y2zGSW4smpSxLUlI31K4xm0c4/OlfBdDQONc6mOWOEmwhA5
NKdjJAlc8K7RM6AuI5cGALKIOUFyonb4b+zxvVe9R6xCeXgU3NzYj8j5QGQ1ssYt
HsWe+N+j6KuQ68YHtzz17PIWpY+0oZaUBfIvYk9nwcQ7TwazHIxJwWBATKsgnydy
Yo9/gQZGNhb1Ehzs/V7WM9d0G7lJChuUhCUtvjAVRBwHWzi88Q0MYNNWMrY1Vl89
FrTtj/eNUct7hMO1P+bRKO4F8XB4wJzcRLeyxXj6GsY4mCWVEsJvIJmVt2w4DRBc
5D/LKc9VaHGpAlDijV4EXIN3w02lQPCrQ2rTkDpGYHN1gQY+ZKq5dbcsU7yZNep/
IdfYrw+8kZiD5cKbjyg0el1eiPUHHfAv71t8lq7k4FbYD6nKfg6Tk9G6iP5pTy8y
7kh1lraCil17aKmeONbT9MQuGQLtmONX7HYNCk9++NgOBNT5xeakrBnJDU9Up1mw
c6lH9fSdMtV46vo+a6Y43DWl0vqsFXWE9zf1Qh+dHR0bqicdxe/ppui9/E4pmVwR
rEQY2szFo8mnWdAFalHsnPBvuQB0L8AQkpziksjSM+QN7Xa/cK8g3M2ImDAouOc6
Hp5Dd0W0bQWbk3jKKH2o2sEXHngdXbaTBe5B8HgeyBPrZPEPgkcAFWHoSozbb89k
MIfOase7uhOr2/ZhG4W0h6cf/XaXrTdYkJC24p780/W0u5hH0s82X9s98M22CxU5
QEng1ES0qKDItYlyx+F2vsYFRwg8CQND/LLhL4VpXnroGAmSWwDB7Fm21Ah1KiVB
f//WaZnzT9zUHADuU8juoYtIOFdHr5LWrocCxITzf7TM7862eeilZ+6EUuVhghAX
jwjEgeT64GS61ifU+o6yY/9fjpQrDeTlDzjTc6dyPm1Iyx+xVq/yvSxrxLXWPdU6
gf/NZWeu2r7krjtny6RbA++V+V8N5uqxOwshI2fqmeWEWs3xVYrCiAK72KJyNZ/y
aUqM6Ac63zV6WMDDOldvQDaLNdPa5H6M2CCANgARUNa/svqwV48hurbMlQ5BA94e
hLiJoIycO18s2YTbPWYwEo1XJeUbgeOH/1FDGInKp5sowkXrtjmX5ZWass8YPh+5
gYcqkRKh6BBLiCevCOFWZoLueHAbXMWaTU6IPLKnXL8L3V4KV4B3T7Nuo119jFN8
7KvDn4/urHFMGBtLmzcaTL7+XgTX+nYnQLJBpopg4MszuUmYjvQuF91wdzL6V9Nm
jyAVjS6MqizxCQ0b8WmlM5PzFAydGTDIzq+0IHK7gbktsPvJyYQEX3jIAxV3D+hx
X/0RpSzYWqygYwXVTRdn7ft+4SfsORUQLYPZPCTW9vVK3Q2MuZI1/dy9lDg0oRLo
YK26J5awqDutH56uMUzifCGWmodDHBC4rWrozfIGd7D6ofFI0HmwYtpdLF3EjUUD
BMrS4nhWqj4vuse96kNTXFR1C8c+gbKWIqSVzDUn+EW4SZFN6BCIMsw5xvSran0H
3CV9kN3g+czJpquckpiM4GKtTCLtUFYjL5xbFQH1SMP9LFEo0W/sl2iyVChzn0nL
BBddSR9P8E8ew7GjmleQoVplrdt1p4B/fnpzItsFoBb6UEz+qqy3SOgLd+jR71hj
VdOteSBqYa/ZkkLlftPXrPKCkS59ExcJnWmo/ljKdDtWVCsxNt8in01b7ZEx9L+s
EwOWYLKeWGC0r3gYHZkRhceSNBH0N0ToP0uirimDnz4VpSMgwwYeoZTLUGKv740t
2MAelrzaqbMY6OuiIn+7SJ8Ff6iNtzEXqR3fF1/lU52qRq8BeVejyvQxYZ3U7She
osrG5GD1Yh8+9X+bBhD03KXRs6h0oPd4T5ChA3HgSzWJ95Rlm/cUP2t8fye7lmdV
8kMmeuOdftZG6n0VqSlz53/mFCPWTlNOgOMvuvdOGYwiuX1G0o81CWNltt2sEooS
iQ4y5wUdAe/krVNgkDlIw9MB03p9vpXXmV7ifx50dl6tYX/AArfNPJhxMLlWGje4
BlfKVt5y2ftEl5EgWGXft5Z4Tj8q8MxFMJ1jwOOIp9VhSPYRYx1sqVGb6ofI4uq7
GiB3rdJ4xRQN0mmbEW5Pl7XKZ2wBHuVovOd5kySLV6IGeGFF/Tq2ArqYr7FQFBDI
EZL31Ua4J2OKCFgBuZk1BHlKlCzfTGMuLVe15FM7V/KslSeyaKabx8N4d0cGpJYX
wE6s0vIiSuEsRG09A5280bHab5poSpn27cTAJWvOaqfLXaB0G7gQyDbDjr/FP56E
mma3iaga524jrTjDVav6oij3CPIgkyqyHGL7X1DjALZt7ittWUnFNagCxsRIsBJ1
N+QCFllPz6kDeQO/kuVl8VT/UQfqwT4rnEuJ4mol+eG4eNSUN+3kJQF4RiYR5gPH
W5rrMTSQ5OntviLWOQmCM5tnW1ThFgvJyNtbbai/DBpkF5yg8Lh60JU5kmcyI/Tx
74Sqhr1i91bPPva/FeP6K1L0wM0ReovKrcpQgpTXhDl7mwSWcJVUd6L0P+hFOtvY
1Yw8E3jinHYPPefGEo/dhN+jsmwoK0lQGonxLnn1nMKw4zudpIqkckEJP0v7FFpZ
H4yDB0bmnkmezs4rjOnHuJwcy27bBA5t/YtxLjO6PGE4O7FvJt80kEVSoUVjVJAO
7dvJg8VzUGeeSOmDI7H5cAzYtW5DhkMeYwr0icN1zzGHGKDBFjw+AJgyzW+gA51t
YN/zSflTnuc5Ki+XIuIxPF1OdXQIrOuw0WXOlD8s4KSI102biALB0vqwf7zElp8P
WGsFLfWSkZbhVgs5KHAc3bw+bREkWkeHtK1HLXjkomKWmfXR3EYRGHBspi5RYmwT
AxBrYZHyY5SQCKOVrQsVoiBiH7BDLT+NTMJAfPXGSV1ZTX8GZjk9KjOpuTX7+rBD
SugFatbSfuH67fmjXdV0BlXcQnTY5x3WBk2fAFSpMV0KENQQMP+hVQmD1fiXuQiK
u17OIJwM9kpH/AligKqqJP4ehd4q5uAYyBlei/9h+QqyGK1VPOoaBDYPY0QvYLrQ
5Ff1WF5HKTDdahesmgSZb/isnijSHQ6/vjZBvmm/9HSX0vkwjpzdHbxbY7/MoEVy
gy+eeZyY1L+uE67wBh76ajlHL1SJFzdrSe6vBb1Gtfg0AmBkOtWm8N4dygHEJ65y
f9zCtF4KzHdBC/quRQ+WhQouM2C7gwGOETxqsrjc07BjCxOh5b3lGXnz7bQNFbXq
6POiAdna9wQoaUtC8W5ZIioVTaho0MX/+otsQz2bjxym/Btlo2dYWMC49jqcIdu2
Pg10F5+thp/gOnIzCLr0JnlXZM7P4SLJE9VWKEjZbkNTiL9Xum/L1aXPuHP9S1YJ
6Dksk4s7Hv8xn5CAz62kDU3zIf6dFnmvTckcqusnheqkvaRhI9pYHdkWSHXurJmY
Rc5tJYq5lXYUhXTiHXEjDuBYyEbIlBMc9xv77iad26Q9ptayteHghNZ6j1C4h9sm
Gtg19NW2Kj/Q9fPAC0UsAdXXEATBCdFsdZ0UQHoV/6sIl6yDQkfrb9Y4BoJaoStI
kztQ6hxbU5/K6RJ1S3kJUvOItTlRaes263K7OfIHlLpg7Bdyx8uyIoIwsnizcyNb
rcDo3J4K84/V43Gc2GMepoyHkiAf9fxAbBVu+zUPqnecpM+dYrnUfYpimgWnvgca
PGEqWK6tFneAY60Ibp3sZh9IUa7HjJNEuR+s9fGH4zTam0uoz1wzO0henGyHjJh2
iLCf5pQbQrRc2EEI87dYNeYl8ZQCbcCdqspL8l6Lr6LhFem9WZWVHs6FQCBN3DNw
sV1toXnvhSGB79vTkmFFm4ttnJFZO8WPlwKt+Npzpeu0Nv6lMhnuYST1M0xN4PJw
OsN3zSyKa6T+PQAQos6cZ4VyczCnpN0LaaOT0NFcIMKwiXyEbC/VvIhHuVzrZ4ov
Oka3XQlVeeS57st/tF3vNSU7QmxtqWMuiqRsHGntZKtts4irCycYEujZCq81XAjG
OxhH5pQmkbzFcJcoCeX3zYuv2gMTUlAGd8TtTX1hia6XSaVsaPv+RN6HOMoNtky0
m63JQ5maPILd8audg5DqagySoxTi7PEo3TgPHG68ZsAwezP+3AXQ6omr7GlNVRYD
P7tzGCk2QFcD97aCwMeA7BTtRuwKFpLz0lmKshliUecREC8MbmdPLlmpZyYRn3RA
6hntRX7EO+RouRignckswU97kSGNVGDE3fAc1gVpdUALsI3jWYg2lfPDYhbkODhe
ItKNUelUQ/jx4scgUZhRPyjT5UFwxpPU6DK6oDPWDYhQ/XJ8joawE2fyBU2pCIjl
0+VlaHriI5MXLvDWxgUddhvPm4F+8ClmrG1xCE6MocznaPpIg2m8ZtfYJRUnmK86
0pU4f9CKLJcQ/7Nw/EU07/C5f93A5ab7jaj/vMIqqcti087QSW0KVft4inidxyRP
ALp24iZlJPiAyTks8ZpV5mRfXmb8tS9ofvrxy3HTD0dSzQ1BCV1M1HJP7intlQxc
5lwenoz9EnBYa/s2travbzRW4uyAKAyFTcuf8KNy0rQ1bSzWwrYWSakgIylIsnRT
XP89+PbuaGvx1e02yRBCh37iNiT/FQcs62HsWBguAx9q3CPYwcUoeKu2mFePPzQD
ZWoWAt+b2qxPZB/A8jEXywR3OPoco+AZAElwdugTFRxlqt8jJucJyXozw8nxmRCs
P3OptJ4WPTDHCAv45K+nVvc5oyF7xZlZ3Gpghy4jA68OjHATXoXGVtsLeZs5k0eR
txtMyOb+jrjXcJD82pbrnPzJA0BejoA5Sz6odyubIKmy0lWTMpdo51BFmHg98Hh5
JOEg/387YSOtrRwAOIUQxutxjD0rbvnQ/ZGb5tXDBiG3s7kUVwmj8EdEiQHPqh/A
ftKjXEUcvGS2O+UB3SrOC8rQpGcfUIv+ESYnmku+GjiaLIR2w6XQHfCyA/XJShH8
BH+oECZs6mZPchR2mjKbU87fyszOL1JzbDTX23ij9Sjrku5R4F5bCCn+cvVMJCxl
7+E19uRM/ND1FgvxNtkFKOcF/YSeGRcC47WAzuOsrvH3P8OXUbJ2a5zUL2lS09xs
XD+Zj6bXBsr9kt8Sdss/adzlGgLw5n1fog1JsiDz85W4o36thXsT6puURUSWXLXq
+OddaQLipkaKcEEg9cleLbkP/oM/I3cQX6n08FGEDGI7bHQ9yE0wlQ5YSFj4tAQH
Fz/YhJJY4WlXGpWrOfhg4hthPJkPi+5v3cahPif5ykQ2AVLRqd896Usetm4wi+lB
EqnnPaTl84CAbymriCkTP4lQuY5tqAD/eyyd0FbF8ibP+ibT9LmXSfzHds01tloj
U+Q5FMbvfKJDvruPkKoKMVrkothFLCKn1lSTfdIlomHgb16mLVdLKBvwuBLo1IOf
H8olA7fD5v/jc2aci8HojftvXauHgImD5qY1gPj1QNFKNH61HuR5mV2TCSfm3NF5
P6huYmfn07FUhKuJNRxl9MlWuXzsp6FKGglRt8QikVQ8qKoq9cV/kq0vIk57bw0c
jYzi4oVsM3E0+E09CxdN9zWQSOhGR37RZR697iga4VHbIHairw0mRNxY+NrnzSjp
rhvc2Z7utwpnbM7Dw7b5cFhPcSWJONphPDa45q7J4rAD8m1a8aQNLnWLsnK7R4DB
DraqP59dCRr3+K8Rcnx/YXT2CnHGupkCGUO6KdRiNiESxgREPoT7N0QDLqXpA9hH
CxtAHHOeD4mq91z65UeW/2Wn8HgIkpl87QOow2clAEa4GN1IWb3HEBH8vWl/wsxf
Qr4xZJOf0fWBuCerCI+4anlD0ZWbIIMQEySqKfwBnM5EFE6Vk4a8yF6t1BZi7sBH
hRX+9jMea1eWZE+sbcb8R0hyICaCShxbhETl1W/SzcapPR2JfL24H4ZAhgynIQpW
RG+jx5QrraunykQPbCMxVeVVaRfUww1RzKRwb8XeWe0mFvj5UDrcloMUcCcMlRCQ
E2d1liHhZh6Bobw975jTgLnWQHZkSGkVHDkBiL2AO4aJVn7t6HTsVNmEd7dMXLIC

`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
4Tl6cpgOo3afU9MJrc1xJbakbZKt+88satO0iHcD/943sq5WURKPZmaILZJH1jZK
wj4WhERGA/iqvBsMJMUaBXXvRdW3RBqd45ocv6awYV24uh/d95FH8e20aOV6Cp1u
HgEXWGAwX2MEht3L/eL56fZ/Rf1YDggZNxZ3Yw0pCt8=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 31296 )
`pragma protect data_block
8zmyCb3dFVvE12Ykw7e5gH4Pg64Tt3TtKNHgAFVmMiQBElkgf7dxVw4ER2gU0zhe
JnsEXtdrNsooeJLKcwlUNFPrwKqQ36CRj8VXBVMI+DFy2bdDIhlf3/mz+34cwrJQ
vIe9GaRfjAcuFqy63MPSnPPH8ePLQed9wTOM1YVga5LWxJQIiPLfoP9pqPIWilwQ
N4y2qIN4lca3IsXas0H9ERjB5CVscamz+bzLVDiNocWbjZIwDYS7BG69ava9/cnV
bE2NCKWj5uaA72O5JgalEvAFQfR/4ba8/P+nlZ00m8mUmxsKQ564Jjwb8q9iMCA8
bQsrk1f7RMP4s0KTgbl37I9dfKjYViFtXqVeP89fy6/1NBsRfjYKaaKU3L7et4qU
5acZsYvdN8bc5+C4oM/wgX/ytsFSyD1C11Rhngmg7sx0FzdcewguAUGIqsP7Qb9f
rTYx9RTAGBK59bl1JZHPKbGBW+h0+mOkQ7oismfLMgexO8iMdfAo5UaVfr2Bnvxq
mNnBF23JfYF/62MX0khsQXxePaeQzVrnDvGpPSbx6EToWDb+Krp9wRL3LceIRjqE
JwUczumH7ETN1yFYB21pedkyOepHBLqSk9fBfWpoLopD1HbHQ+EHX5TCAo5yiyY7
b9B9cyrDvj899TPvungDxziWUmQEhRJhLj/npt79BYQrmvfTwcstjxHIMNlJUI2q
lXQwxMLNTCO5j9aiA9O/IPp5fPpCR2CrYkPkjHTe3cVYJeUYGb3HLW4bPvzsV/xo
ztRvPp1AbGdQLjma/LkjMvK9Syc4ZAdI4zy6WWp/++YICNWZgk42bVEw5K04PFfT
5sRbYgakiGIM3oWdZ8Og+26yI945tvsMQRMrqiiyagytpeYMsZmLDUp2Yd665LrQ
IoJLhsflFikdBm65fEIU4iaTo5SC3WTQ/cFAUeAQlU+2l0pF8zZUadfqK+iBcEXY
PLPRHulwB61OCSjyN2/HMjYF6R2OaK70aeMaUkZRLLtEDaRGPtdYnILqHlp51lsc
+Qo5qvfiyg/qrHuJN7EoximQwD8NljT9BTWNojUx9svFdDinbmFhufM94ecsGLre
FGtyiL/CZzFw80YqovFccRM2YcbJc3a/jGNX8M3Pfb4uti24UHWvTfkbJtj/PxCv
1BqlBFO6AQR7vCFTG2P4Alqt+qQLqbyIDrHUpbQbvOBZwi/TSUFp8gNN5/9pHGXc
qAXfhCvD7ONjtl4KSycIxezk4HhCFjVF3hhCLRCArvXFkRjPlaUUnyA0GveQ14S2
L5syj/qa0rPEk7uHSVwwKgKgUFNDJgdsviebGFQQs1vfXSDOnswzjN+jo7fpe7Zz
KUfNwgLxJvWj7MBqClFtsAJuqDYpuRajy/bZ8cG1xolutuAiwAvRZEsHIN32DpG9
dxSMHbH1/sTUFxM3dKyk8p3GqwCmzdpkJgqqF22OKiphGeb/dbprrmTtm1aoNGiZ
dhiyQSuICXhzmYRkMeWRd3g4qgDWidVsTsyMGRrRipLz/2H2UGxG3tP1QAUYhAM+
uQX2jLE9wXN+NZGqzHFT3M8Azb/0vp9lz6GWLartS9gPfp9yo+/iamkP+ZSh6T+X
flND1JsUM0/GK3MPnF4TG/zzoT3dAcXRxuEoh5Ux6HEFhpWIpEtwZOUNc9u+Qwry
I9kDBRytgLF0/zF6W2ybLg0aGccvjUz8aakWWmhWPWKLXLLJqVS7OMDQkIi/KMGK
2mZr49NHM6Tmw7lATpcgJi8OpVLqdjkGnV4cRFpJhhjjn0WPw1uE4L7QzxgGQFYz
/p9QZt06zn3ul8oHKCfX7UnynOHcCz/slR6Vos1SHp3gjdAn5xkjPewVHfnPvXnM
nZ7soFBb7f4rHUebZENixR0RAas4S5iExXJbIoXgAd4e08IF+dq/94ThpWcpOSYy
VxJ4O/th4WXC/Gfw9GzyT0BaVSmLkijsbMyOeX//q7EfannB8TE7fdBhpemkrM0a
wpLt1pehHEdyl+5IvnPG8NN3MWwwlWrNj78a5zD+/LdSgoBo+ajWWkeoqXo+2UTI
9LZqVukzt5VPrjlXe2LGv+9Or/5wPoTibAYUembT8kpW2EtlSsnz3Hqj9oGh7ZZE
LLg6LFDLGUMv637P8Gi8RGxHX3sfZPCfBpK9BP5UUpA3CflmLEyqirN9nW+eHI7G
nMYyTE8hdv59dhF7EHTTlivuzu1ufFolBKw5h4ORedrPxuYBH/OjPoeRs8XGPmLq
XUjXfqUfaPIUXnqHBeH/5mR/8RfOby53VNIK9MS2KjsEQdy859mJRWbsURT75bBu
dlFQnJ5z1KVBqaNsAMcOrFfYFwIktdeSNo+SlOM9cjqo/oIxcgh0J78VnjpYlqNo
iestxd6tHhMzx+XRsWNg5IUBp5mwJ5tBviZqvib5tHyhmtfDr6NdI49dXI6FHhtX
D5PRkicg+rFTSfsr8Hyl77Z5quJ4J93+2u1HNPzPnlzouj+nPUyoDRY3qXEACCJ2
kIvlCJ3OduH/QLmjgXmnn8TdRXfm79TwdXWgs5202DaHyW1+83+GIg0ztqLz94go
NEdEZuyzo7eHxUb2r27b5CCKHPwoGGBySPu1zKWJ1TXMtqXXohUod2+HUNbtjcOj
hohmtERQvsSPgPpQbf6XMPc90seBIj8/SXsQsZq+Qnchux9Zt46uLs8TwK+jpPhA
ybonLDI+hTrErn3m/dOYHeUQ0ByFi0QRLwAJdf7qa9u9lWDj+Hfa+9cPyCWdDKh2
CTupPBj/pYKR6/yNXM3U78hcD0YAbpeGfxmjfwnlmthDzH1LE1z5M0So1XPl7Ryh
RSkeWtAwYLiFw8VAuoGf31aFeuxPrm8aOHCM2oxGtRXmza6JZ5OdwGDHQXdtythH
vS4WsKLZBefBWobOH0Sd2VSQ+qzHXH2NHV4hpgl/dFT9kFMSDPeOU4XOF44Y71MI
WG0j8Jf8a7Hk/yBR8kG+ahdVxQrg2vhlJlSiLIfIAyP537hiDnlqah9H69/ZNLim
Ew8A6HDdQv2UE6L+dQO4NrQFw/sLjaOnc/8JwlTW5dlz/Y8+ohgNh6JSTX09UMQo
RjQ1Aga6TcDy2wtokDtv7WsVLJzfQ7igIbkrnV1H59668txNa2zOKvMjRkJ+OSgG
kNo2bBtKire2Lh03pe+Hlc1GuE1Ra2yTwyUnS6dAKrxc5Sj84rDL8u3mH06rSckQ
ESA5wCYegUeVlhzO8NYBwfLKdW835lxKq4MgCCaXxBBjEqGhFKMMflbmHfg4HYMj
qFDpojOi3elI2ZJasAC7aMB2a/pT8o+Lg7+5s4taHAJlDPBDfNJD5Jd4jSLLoYkr
SBIqS8r6D+ZW9W8ZpukdNKHec6WOjC0+JL+pYiE1XYuH00NIW8op0xRSOxHoJFWH
Apcppzd03ZLaSwtwI+mOzZ3lRvcD2KyJ+1YpTOooFdkvLcQIFRzWiD+yc7ItVPqf
l2xI0E4bBhplQrfXaHuK2pMRd9MQLI+i5vjyjLpgbymlsr25/C6lW4gPZZLKL6Ey
0f6vnDHsmbWCXqFCkUOR53FbMFpmHeF+4Zye9CTen/V4ouFmgFtvA2QeQQg9DtLn
iDBpsMeeKaZx8xgKNCE7Hbq7QKHul7v+ZZmULb+y4KUa5uMHP5tMpx9YfAAQMJm6
cPMu7Co+6RV+dqCfekqPPFvqPe9kyswWdUY/FzU/+RbT3+nKusylsKLWQaT7s7dk
GOkPuvMyz/r3fozkVRf+FcmUEmE21980bpuG23LaO7jge2qANMG+11BLJzb4VNEQ
1MYqq1tyZEUDG5qd3ZqoPCbf6etZXz0hV480tEdJq03GFCSCM6lNt4E1KfHUodLH
pgESlroScuLUyZ3P3EiatuW5kczMxcQV7TAC2TQnX6sGi4mCY6ERzC+1ZNH1hqNc
o4gOAk1wv8ObOCEtrDkCjC3wglQKKblC8co2RB2GVhJIAxmoy1x06cDde0gLGO8M
h7It2gY47VY7EM6aJqEOag5+yEfqNSAUHMmqZINbNg1EwainE0M4r+1SmQiQxaN9
yOjpAQKKln/No2X6zUV5OvAM8K+5zsker0fs5Fa+gCjuHeAQiEO3Wg/335N/Jzop
mkimsA+jA9mp1NSSe7g9hdR7pGyS0fsbEFTGm8SECDL2GYwRG+zGg12KmT+BRKml
ub07jAQpS+EfOVarcqgQuBmYXH9g7Hcg7ZjZGn8aCoW6A+fG1W3AQGlPpbGR58+w
RoVQLvx5X1Cx1g2vMs8HOvUoCkXAqvbFzDPsWIWiuxI5wgSfxB1R8OslAcRoXVvm
2aodGVbEL5Hk2mY83LtlX5f1h7XlgobkJLjARNGn+B5CAbrg/kxU6OjtfhAzpcWU
wsMxxQCwR/eli54MqFo2nUgph1TQ2kcq3PtLhjddtXbZbIJDY6rMqFeDShBDq/Gt
B4todBKspqEWouabAgX/WUAbf6RRbe2ki+pfXo9zrZlCe4cO+Jdr6/1lWdEzvkSL
LXN9LXq+/me9aVM36RYuGkVJVZesaAzb3Nxv+VWjf+TAKLC8EwyGJd2O2Xim5vpl
lzYaDVCmhfcOWLl2bYnAtRg84fB0kPndYvVvRPY0bJMTmNuF8t3qHDlehdFwYGBD
GsR8/ISbZjV+FkIdcLleW7J9HPQ9JVfaHuCKUFe7M3DT8FYZKLTDYGjM3wDeWons
6wFDK5lWzB7gHdTGpv3SHGC9Y6rD2d/SZjrMT2PWpxmOnb2HdeMsKleegIUq52vP
NLR2Hwpi8K3y49sVegBSSyh/NDQfSvixIe/hdP30iu4syZJYYVN/OVuQZhOzYNjE
/UA0hBfpdjTKiajdwICYZESo6W/zuW/ZOrHYl4DOw7DjaYxhqoufMXj123aS7GoO
UPUxwaVh6KVxCpQNh7x92LY5ZZq0UN+pmUbqDmXTsGNJIec/Dl/dS3eTWaHazz2z
t6NalhCwAo7OLwJ7XFFrQXnERJlZzAahl3DPiO9jXnb3i5Qk8DYdYjsGbv70QcgT
pt9bc9qecmb27okUVrhnhVlYWcT2IujngmgP2yqsQPF8CC1M2QjpGOeSOpZo6eSC
cPx161q1C81aWPHodtxNTjugyjJ1yIOitrEgyqKGqRrtYVi+KWfJSaueHXi5RSiJ
e7+BKuU0HAqRLLW188EefaksPyFaIJGz9G0hBKeYN4vfROEMUtoFmOHdR+cnCHZT
kO9tquHu2av5mDHI9UuLpXiaK7CfDVmyNYNXMD4U0HY4r3tl0i+1itwKNd1zoAL5
hXRwZP7gyy06qXYR8g9roQBUdEsjWQhiFardvKlPvHoH+KpsTN9lRsH1129ey4FU
JzL70J2G9Q7Di/IAmet3WLe2fW2Vy110SneKWZbjtU64Q07jx/DrxstPgVptmUl2
uP02G2EDhNZG6DMJMU1LQb3PEGlg4KEBYkznUgxkxbPmUfA/Dvwzit0vY/OdSS+5
oZQFeDCEMKmrrksMnmqWJNA9OXbbsJ2F/SFb7KBDqApcJw/qZgQ7NtjbWEukLbqV
biTO+R04si+14Wv+0451l9OaIxBvJbbOnK7LGF51MDto9BecCOIPbI5LLwDlvw5u
DGJ4qptMPGeO+U+tbJP55QHZi58E+QOx/cav7VAOh7aCyqdVVYCg11kiuF7/DxSg
5VBDMV5ZrsI4uk4NMJyRINj+MK2LXLefYcXodE5fMSijPG+XP9yGLJRoT8LhGh9u
PXOYtFgEz5R3x3gQ2Xg9BVh1zYOrD5O5WA8hKA4/k9B5MIJ/mbarWYQnPiAs3h8T
k8YjdGx/Y+zZ8/B2JBWRk+3izD+8pTFxzA1vpkJGF6OLQehmKMtXtJgZ/g4fC3a6
hPTy7HmL0Nh4SVybi8aHw8/HM2lrE1LDZd6xyvFSVeC2O6wVkhb5EX8radR1cF0P
jYRfyx+HrRtY8JEJU0fVOgUvDvjUWjSZimBezDwKwgZpc4Eou5DDUlmeSLgBcVmv
qzbkp0CBgf1atmo1SVgKS2W2MeAoqhG5izGipx6DZP7dfanvD2rYG8pjPTq1SniW
jVwNgTbudE4CpVhBQQmQ376AbmBb51WpD+tbNM8i7MsiUOjHssq0tfYcuV4E6ZmV
DTLj0t9D5M2wkXz2SycxR3bPvHDNJaxK7aLy/Cu17j7GgIeLtSrFt6RFdMjraYFv
anE7x2hv2hKVgvQWXIOZYg+AuvirQ2Uvonz/xFrqJhhzHTUzlRMasCE1/SID+nUf
XRfXyAWg1sG9oUNKhT1mMd7wVfjaYP8qsle65hChPsE00kiOB6ypf+oXePLDrl0p
WutxkmLewfsuBzqfy1wvODjyMh1kLF7/n6nH7iza2tOD693Ij5Fb0KdHjQGCd6wy
fymN7i7odb5meC5xQ1PqT4yLXoRUy8CmL4MDDkvbhtJyX4KQ9eX9pRUHutbuuYP9
mpIBZF89bi1InJ8SDBPuAo9HurF9Y+F4PxCAqE7eUTLZFiTmgNM8pdA/KxFDMvuH
pWNrFPDcuhh6Mos98dAYIlERyJIdBE6eDRpe3TSSkOWWNuRhXFpbCvl6+yM0wDT+
eJfDHS3uITwrgwR61EmUzwR2a3ExS/av9tdoytF9QvZJCsbFM7yb0cIcwNV+1sBx
4ewCNRqS3ZHZfzB/fmkNlrEUAgYCsvSvuD1gcJ+w4ypoSVUQcy/BHjEqAh/pS/8/
OozQmEZSj2w9mqMzOcmfJqnuUfhHxuVOBkFLPtsbWChbaPhdLDmdfZkwnEBxW7c2
5vbtlSIYAIHgQW8COyBeLmydaDKK3YNCs2Rm9L1Bj+vv2lYmPjLbxa684Y+717kD
AE82gYokM31wWzNu1q+KcG03o3Zwl5LWJCMMvGiOHeYqoPR2+Pl8051kR89wfUkC
iPYTVGXwp2xULgnZHdTN/V9p4GvLxlru0YaQsPqx+QDng6Xw19zhzht1gHs+fd3G
8B6uykcLTNYQ+N2+YGjdDJYn5yC037aLBRBoOvZxtTZhWdmUMZ9XD+gBeakOBY1t
Ud97H2lHXsUlQaaKdD5pgHWaXFUpjNtTHoZeC+SfZDIIcSGa+AWjhP7Z2FLIZNAs
mdh82aSnZ6n78I3xRNYsvOq2jVLx4O1SLS5A1k+VBjU9csDgXeX10Llq8AvcEm/3
W2PUU3yAoEIrmG1uTNd+QufB1s2XjNVsGnSaFnNu2UhQxo8mc8GlscK72pEwFv4x
AeKXdUh+k4Wxi4CyRVspOTPwSY6plp0tp+f3pffMZIiRX07rtnfs7tpdYGwn4tT2
fFxFt2t9Xh3zmh1ZWaFUvMp5OWKUP6hOF82lIPmrBHLlhye8NLKV3HegDWdiEpGY
r7FkRUz535JNPB68J5ey432OeOdcccsIolOhA3/MJD1rZab/57+h+8LDAI3wrbC1
eX9e/S2lrLf8jnVzRqE4yUzhlF7WId6wqrMfV4BVV+fy2ldSGl+HL0ZnrLfl7Skd
KEKsIL++MuNs+M1qmXdzjJomFQFol42dzZVwTEMU93bvb3VAAZYJ3ADoijMrxqNc
QbNsmEZXuJKUjXFLVdqePnJWpTprTwpEl4ttmFjMGW2h4hHAZpGNTHkZgW3Snq6l
56RcOlclKoT5o/d4r8unFZCJi026ogsYHi5iyvTjyek+raqTuZtFITajVO56yhra
aQLzDvbaLRswCSD3zBuBW9nV5RioejmweNWbQbTZTVa2BylDnBA3rg2zmxFT/mRt
/P+fQlJiLv5aGm3VX0155nufsb7w40TumDdxISxCAUW/SAtzz7YUU6UACX67zYL3
iyNnqYG9wDEh+Im54kWB9XohBqH3lANBNA0db5IM26joHgcUCPMTn/AdIc8K3VBO
OyOCHYGrFUC7isZ29A/6JVQIxYBQ+W9ouY2Djp+M+m63ZNn8pxGqWwk3noqbsIUm
XmXYZArO3+46QrWR5eM1P9gWnqM3vho0ItjGHz94LpszHqUfTM/mparcRfVE5qkR
35FRTBIFa9DbNq6bmEngbdJvOzCUgwdayepmbHwbe/uxT63SlgpmLL2lVsEwdPjL
/IPe5RhRHTuM0nL6ucmzuT+8VIadnMyiRGYDH7hneFcxx1u66LBB07fGecLLU4++
blXqjpwSb2s4faduxZiRcFQMmamsGn4jvZe33aJU6SWT35MfSFSJj43jkwUQaegX
e1zVIpTNCZ0sQuzfnzh5cXs14f9Jze39o1Iv+iSlzQonf8ZvCG7xewS1fpmdIAEZ
Jn4Nz0gjMfAfkfzX6lNw0DNr2h5+5UlfCP+4GXPkiWyfocMmtG9UcWwAJkhRfjbp
TfUQANlD9/qdvNKuPuLn7QIit7htDShkoUOOP5rDeg+cjoQGjtV6xSKr6vf1dex7
ZUZsrZKuHxS39W06rxxQ6dy4bbIpOQDbzDxNFtaBDNxOIrfRJldnOHy8P7hFxStt
XM2HPMcE83LXJsWVRA4wj8u0l4hOQAzhqxGHv/mQi79uXidiyPiXhe8cyEGAlku6
fn9NLKmim+QB37F2AXSOmeryEzTRcuil0gPDUp8+C/QZb6pIpNoYD2eIKR47TI8e
O9ykL4P0ISd3wCul43bJPh4V07xL3hjXIXg1jMTFXOZlMVHK0Hp1v5dQOEk5uXOv
MRnzzvHFRrq07g4Rc5L2vrp/X0Nv4OysSuxBG3eeaNE5bgfYGt2msiQYsqeAVoIl
d2XK2W7V3AhojvT9DZGrqyhJpMC9xq4D8Dc9DUOq5fhKBLFqLaXa2OTjyS9Bwboe
NEvJq/fNv90xtPU92Pe4pE6/Mh/i/6KlTsXE/03yzqt2cxQRfPxKJE0XBA8z2ZHa
B/BhXsWndab/ayIDvKb8x8QBWk14TJscVFM8qdpgtqehaDFsF/RtLVBxsgl9ga32
cg7O+oPSb0ToMc/vHln87GGT/Gp4lENp+kcf+3Cr7iO14iyFa6KbMrXcR889mIlF
uiWH8mR4UukLQJU29TYXBDGJqluorxyat54E6NVTO6Y1OCpknSYD9sht1QYeWEaS
carFov1Y5Y9rppA5lZ7jP8ruAp9+XtILhg3SthsBJ8S+E1a+QnI6csrjZBnONGUn
2VHcc+n1UkyZRbzZuW6RSyZ347oE/jMxGgPvGEzFldDXm/CJUMcpn3qEZtpxZHwH
PItMKQcGo/8QzJeBt0WWmH6oRvT17mxViHlr4Qz6hK34hddNZ8/AnM2ZNeS99LkF
jt5hsgsPRROJQiFlCiNnEYFvmVClVlHzqxBPz8X10DvvMnHEpHpl7e3dlXXoPiWd
PvzT1U+BkLrvF/KCXHEjmzQ8I03Hi0Vb9gjirJ0cPqw3uNEr8VEUd0pRghDgeWEH
eN+nfFu0O6zEXEUXlEzWxhnNY2Co5pp7+14U0qBkyuJ53oOZ74PCYTJDaSOPH9/W
rAguD9i9VgWh/7hvtMCGkiFJZKob3zHMfdzMOwGKdE/tPbJCm5QwReVHoR2kSFly
UQMkgGPO/tNLpb6BwlcpRoP+/J83MXYvfnsXCyc1T/ujRBIt/vN2J9oNaOVnuxpM
Do7UNWAxOX2le/tcspCedY49cRL2Yi3DADRqa+qt0RmPfKebgfp1NGp9QUyxJcgb
bTh+5DwW4mc1jbYP7S07eDrIvQlAxFu/dOuQaQpeNx6YGb73/QQrIEdB0vDpMWMU
YiImU2CKZYRDVHB5fD9Ii0hUY3PhutyfNn2e9YHCQYCofC98kC2PT0uFTE9VxciS
Bn/zxLsdQyYf9dQiGuFgK93v9eXUMyCK0SgzDkTpZYOCtfNUt9qKZnRLKEX4xxT3
vSqxP7Qy8dHPiGJxP0I0/sM29YQsg2xxZm4pOXfT3lQtwqIZxs7SgnBstNTWATyY
FwXsIkCZQQg5uVyX4RHK2/MCl6RKZZ2gY4QyBFI32AZSPBPeEUYIB1HNMkxEieJe
xJpVO5aAT0VrYbMswhbMYO4mw3h9YdMVDzvyllttiUBVOiy+pLCoZLez+4KOlVKi
f3eiEOaXD9G9i4p3AlqOBSZ7cT87SjDIphENFNcnWkUYNNyAIX3hGUINWOEdwVp4
3ycJN26AGZHdR+0nBRfl7YxcrGnpQlWkfaks3bvS5126Fe7BId/L36wgPmZzmiOi
4LM5z82KmPEyBQtSTdKt7saqsCo4zjLu+oR4BWDhsduMY0xC/1N8EdF8S7UzFXwm
anRMgmJsgkNab8aBYyTM322S6TYPmA9D0cWHrZk8/NwBMpJbmUDidxOSHpEUFdWs
rETfvsOLWYUCIrMlFvfBj6uCiRN/dmfGDzuvATAzpG5yzJyCPYS5LWXYZSrErEG0
H7RuOmka3JeMeAeQfFWh/uLVui7yh9ygf3cu3Zx7IiUSyMWM64Ttzgr1Uvx/QU8d
3NVWpuDTgH/r1jTCKIfzTlMx4KzIbA4HSZ43dJDAG4pNNFWk5yC/wQBvTRz+/Kbz
FnGnaCbWJfn0bDMXL/Wc037jQlEWFddWI58BJFb2tppJp2nqR/2NTxutNINQHwkP
5n+/9AnOxz6Nc1tXNN/H4rdwCiwzdPlfy9DI7QXhWmCn3NJwapgFljtbWtMO6lqB
uhx8TvC312PdEdprpo5yoUOg7vHJPrTLkP4CZKEvGY2V5PjPnFBNfsnILIzMim1o
WOjHKdaUZlRONOR08VOOphnnkE1kdFy77/KP3YiiYlSu2zhUggeOYUR80cfHlsdv
4v/vii2E9J/YYCzIgR2iPh8tpFJnqdz8nu04jiDNLi6hfU6kcT1ObklMACCUhIoV
e2Xbd/Gq5Sm0HWCauNPmQcWPminCQAajwV53aDADrUsEXDt2at7OO1XaJlvZZJs9
IkH2M6pn6DCbOMgpoYVVxt3y+4J4GJLZcg7KTYS/tON902AaqHdDEV09Hpp7pxZn
INadPSC6aVj1DrQagPx5whGAcvp5YYlBMXvsz0JkwsV3IQUn0vHSMyVUcF+Jdz/i
kqzTpM58L7DdnWfza59HdTKugX16u+Uqw+HCffkXT68CD8ul2IFn80UmQZjHW917
UR8vwIdlW5CGKermTN+1HpGXn8nKZOvJnpjzUPDpzC1J6q3waglrj+0zPok2Kox1
FyDe5FV2gyRxg7mZV9SwMkr7m7DwhMVtt8bTEo2D9Fx7GfAUUrK1vqkVmuTzW+1I
/WkyMaM2B0itrNK4o+4R8kJ8nhdT9HLbhOTW76nHnaleECn1yBBdbpc202Ldx1qs
D8d5s1pp2YM/1n5hnFxV4WbYNEwlHhWCpPM+CK96do3PGf5FO7VJg21yACpa4pKN
osvX4jQ6Y5WPPftgst6t0XMqFzdZH8ptp6hOLCD+/hxvXmUg6x109GMOgnAGfxrA
/lwBA3ENbpUfckHxNPKCe3CVQ7kZ3vQFkcyREM1gT+ujYSdb8uW/hvv/puZqPUtE
VW+TIrOf275Qg1ztiKZMj3PApAvu0fgh3UZUTk+Q6Nx+RLcaveGhg04Mt2bq/Bdd
0mN+HdYpXVLDj9xJGlw/Vtj3IbnYN2XVmkB3kxnzKNZ3oVQeDp3LpkmKdIdRmrJN
LzarLZdUzA/XBYdp5o/45vDH+peY07WpCLUl+olOUN8zF+URx/QPBMsTm+NzwTDp
4y2WTd4/e1swqcyjFYrHaqpoh6yAi4yvqEX6kYipx9kJT5pTaT+Ah2duV79K3QS6
7kFxUcwmNzXzgcSFETmbCouaM7E8gMABVGHRNhYN+7qHVDdDiGbmN2O1cISum+AD
3bDVsYSl2aNBFf2oT0tlnIJr7cdbmYT9xtFmzRR3+pd2quXRrLGzcDQKlwOlNt+F
+fc4PwvjyZEZAFBGZFwvv76tVhGfbn1EKwVD6+BhhpEwO+MdrOVUimQQYVIdt6ji
ynhbt3dyqf2kENLD1WXlW1W1L3AkvOJQIo9AmRpuYWYcGd1RWDkpFb5Wu4M/UW/g
1POV08gaQGyZXSxGZhQRUQATaRWab2IPAbn8xmMr9QNPiPXSh110xuos3zWdLOyq
TRXukT7+IEixSJ697iG7oIxenCdoVOPrSaeNGkp0OeTY/mrUrOPplqQ7YIzW52SP
UiEuhvjEENQRQM7ipHab+847qdMoWDsrLt8IzPmDV/2txKlboaaZsbrku18HySaj
KCUL1vrJmrEWMCu8xtC9YKw5uevNDF0A9DYoacrYu8H4AT2QgxXc18+4qc8ij4l1
Kkz1GIPx50NS9lYjV1Nw0PoxjpqwZuEEdihWKgK7rp4Giio+EKHbbCMySl/mdNTi
ZR66qeOHZ0VKnIK4te+MeZCI9njxchdDw6TG3FfGObhgNk5oEnwic4wY6iDy8GTC
xGRn0NAlWbRxUW/yO5RVlf8+FNi3tLyGj0GeA64bHR4PsjfD9xglarz5lNPSE3qE
vIxpCVpHMONVyItBtBX0NlaR6BASqC7bk/RsHkeBuEl2V9NGknuSFXmNCy2SHNTV
P4AnWD4NW75dEmHfYDxOkdlK94CEl50xlv6DQh7nSCpeEXu7Fe29Yr7Mf7XvUz5u
Dv4HzVcB9nunTJ6dz8WQPO9giFT5LvF/lQHyJuz+qPKJ2YX3dr+4wjVuH5HC0vUS
v+4uvvF/WSjf58Eygi1I/n/9X/Ap3+ops+jI4tTCAYbQyP4wBhCz5Unuwrm6ZzpF
QRjXt8Dcvjp8etrXbASm1bWv0Y9HHTU9sE1LdUyydblKQu1fmSdWsMKuyIapMcE4
sWxGwhIo0sPsChET8k+ridRgywPRk03JVSCbW7hzOOqaKpGflttnf96MKqTkqYI1
pzq7KzdFvYUJggsATkUBvqGzVjSMT897Iu/5mmIAhwQmge5ycQfYAXp/qxMtkFHd
aDuXdFhabOTUqo4RY9thaHnZH02FQSHU+HKKYr4qewWOxaZ2XfILx3sG85TGHGhb
yUDC5cgS2XcWhY9fKSocP99ErA0naeCZF5AWaUhymT86oMBfwyjtSZJJVNHmavy6
QaSr3MzapHGmDBn1/tafkK3vGMEIKCf3rxX34+DtKKJFnALb5pIe8i3zAwToCXs4
GsZJkugOUKoVaLVfNBAmC3UlDtJy6O0+CmDhuU/DslGLeMFdpjWv7sVe9o103rLy
5FdtGJ3kE2KVXpwdwDscNeMd2CZeZF8FGPwVSE102GGjrKnmTAYxpE8mw/ZIioCt
74SKt3WMKG6suHhSawskuY0S9EIJSQhQIqnYJgLaioFJcqsUzhXSmeVbj4WUqsmL
UyQ03suGlq1uQelGSJbu214vOQVwmz0NGYtTrpTokhTGjXoS+Cpi695yRaq5BMti
B++nOZ2W6B1RHdV5TizDpNRmKy2EUbrYmbaRAx7K+rXcti4ram31WxH4ndA9yCV3
l/yotYnswkM51pd9FsMwLJjckAQORm24+qsnmSF3m1sxiDcwbSZzt47MsRT6DUui
tFoUZSnBPZOLDYbDXbg4tcRdkT/14m1IJ/hv8Yx1OEmMfUz3IS+LooumOPmIxIkL
/OdsFmV0hLLuGpRehcef+DniWQntuv+Q+HhFKdQecqAlowLbJuaWWPhZEfVy5vIN
rJnYptCHc/XWNGlhb7f9EBHhh0O0tDs4wJiEN9Tdkb2n3c+M1rD3gAoxnZNDD0To
NIxExOloVlkyBdc37kg/HYKlnEkxmltxaACJJGTtUVBanQxQV2BA5xDap66m24IM
UM6ahmPUxQdquxRvMG8LJfpqbUyy3WX8kxU42Z90hGeSH1mPYNPjKYTS5/v0wQoH
MozdYqdCsgNiBBDMU8yNZSl/fCfMB/pwyFc+JElmewH+u3VEHSfI7mRhkAQZWaY8
Ah04Yxtu1yPLgzX9+h8CHG3/xPO4Ce406Pg8QGzhKcgeFeXi7quJ1MTZx+/2tbk1
8FDoLNKhV/PxcQTWLd7inimnr+mki28HBuriZRmjH+PC3JZbxXnckGvBcdO/NdvS
NbwZ5EF/rv6ZBTwe1gmjAyRdbQWEuD6ilEXUOqZ0n1R4HZvDgBymI18cQlwJ6df6
hZfbZVpof1kA6evqpxFallJ56jJVQpkCC32NEldpHNPJ84v6ozUK0Oysk0R7UROi
tvTwYS31a6asm1EacK5NqG9PjQSoXljbU28ZX0MvDw3soyTmJd3eV3SrKDBFKBun
qzT49fYdiItkBIubE32Prx6fFbd1DoH9g20Xow7UCYnyUpzM9+q2fsp0jWPWiISn
pN/hEjoFX1q22H6lNr9YLK3RRAP/GxDiAkhUrwbx91D8PWaxYGqwC7HsmgwHUTBo
Lys68M5AfrmMRDSDsIBHfb7oGdPwjLrb2eBivlQcxIzPp38GML9JPw3HagyIiK/x
mAb3JHMa0aAxPIF0j2gYZwOqZnR21ufrl+hHlPk/Fy5314waHcig0deFfq5l0ub9
BOq8rihcOpagdZBvSRT3jJ3sxJihM7LoBBxJQUy3s6N2lhlfOxK5/t+prOHnqvWd
VzhBjh+ec9xyO1xddLu4kAXK27DvuR2UK7wd7vR24sQS0cl+pla5OdKn6xfiZIDM
R/q7v4EyJ7dAKhyYpOFyEVcs5PkvnPno6bcqa8MEe93zmYSoM+CjDPTctt5wqdjs
ak4lWBcXkIRP6eUHiGwbASDxKYDnAxlAIPm9U2+aZZFdoGhUiJ0WDHpYi/KRppgq
dWfAOn90K/M5jZ1KOUrXMq9kJmMWO4cJFMxL+a1pU8VFmh8e55U7wuOQLfQncZJG
mxoh4uwAIMpHDcp0C2OBKFoX5QkiBSqfjV3b726Ml90hLdwojMnLcA6o5Ucmjrmy
+K9TddnnmKZXYW30MJAargLgg/N2brsOe7zDU89NFYCQgnrdYsrG8HpMwwu/Coi2
D0mOxg11zFTAaDngwKX/AKCccoh12Nf8Uc7YjQ+Qe1cZsJw4L7i5cnMet7gTlooH
DYYea+adbP+04f/pejaIgPKve+4kO4HJAIqXlSMrOKidl71bf2NslXPPz0gV+tGf
/8zEssREUPmteE3siqZ9RqgKl5jvxmLmggt9dFypAVcLWA3CIEC5PTIBYCWD9+Ze
1enkH/E0/Yrsxs1wS4jYFx0Ym4THRdtxJGNNxF5MwcV9nfuDN0zBACd0Ohjh7V0C
hZHOEVpxKG/aHoNKkSl4fkgLoJJC1CzraUF8CY1JDjAGIH78lTueG0y3M2jtVAow
6eIh74/rdrr5EiqsKgJ5ESgKVgnDBWfV5tvetbnXCGQ6M5yiUh1TCNdLegqKP/oU
yqokzmwNlAIzqh8AWqnFpvkW4JBUhAKcDFkjKG4bHrf7Edcb8GhV3dL/maJWQ1Ix
blcPydGaxfRxdaVsbpsbTAerXYX6nltaXdBJzDe9s3Qtj33zjTCEeWiiZXKGEC5A
oh9JeRecnPiMyrJ6fuZbA9oG66WhmL0Y491QZIQyPgHU25vYkS1JeeczlYbn6WQN
8Z70ctsBCSexVhvTasw9mNVua9uUwjXkk/uqDBbhh5lvw3I6KEVc3qSJHlEjdZGY
NFsEe2ChM0H+jQcWFWnbDT/BDqGq6zk20oFlNqcHlS13mwXDTSIbfMTKh1ET5eUp
KCjf0+lUrSgIhMmATwO5oLhXYrx9RSu8Tjz8637GCKU+1L7x6I9DVB71j8nXQXnp
hRhrqEj+mjO/ofW/ynvSDfY1l/oezF7B+Lq6zzImfycrnJTW3oADhhBo0QQitoPo
XVmRFvXQJGt0tvu41K5SXZd54pQ6LolM2Oa6PdtcCvC8wHChhfCwjnEvLyHrIYwF
JC1UsiIJAshPq6LJ9CCHmHz8gU6fQwo44QG/lROJLDl+kdbElUdG+26ZCKNWe64X
nuCETkorAtPrhzqt3EpPJQN4ssGg4e+m8q43XULyFocgvjUHSD9aQ8WWN1CzciDt
k26oB2MCMfskvRPb8WLPmWpyzFMCaStXStKJ5ZitRIf+9gD3s+AyYYXfEdPvs9Ok
Gri+cGRhOVcglChmtsQmMdPuNtIWWd7iKyr09ZQ/rajZZI9HGhrES0FxvozBTRxU
FG1SzT8dLmu3T95O+DuUKS1zcWRHCNOU9MfbxQP91M2Gk4sVxS/81pVWq5qKEQIv
ZzNrzZubn3ypSe42/t1H0839w/F+OM99mS5ippm/Bl13gS/WixZQtsEbfDQu9b70
uuE+sLX17vHW9tGNdJ+JbozAnW5rA23qea+cUC7Mt5S0sguUoB0rVFNNxCJZviH+
Letv5gXxDu/0Qecu9T8MS0GHIvGEUXnohSv94bREMDxaOg7SoCnuVUFlSLPSrCaz
zdISHCDsUvgNSP79OCztkzgqiNXWK12zRjF2V8sFlYUk6qEkQxYv8K7qZMHFdjCL
4oY1qSoxo1n64NxraWIO7Bj7lovPqbsEpMNgNEgDlSlELp+VLCpPLzNyt0u/waTe
F+8ksSLtL3qnCX/3aAvnuOEOv6fZDUQ+ONkLD4qkPApzxsZC02A/MMHjt50kv7r/
2qPc5A4JEmpy0zch/sZP4XZ9FyV2CRXMXpnAGTQewMgGOwcBnjVZdCoD/2uZPrcz
ZcPiZYp9tQOYgM2xXl1LUzjL6e1gTI+QJoxAcKLb5aQKgg6JT7Y6zAgmQ3spx4X2
JOj1RW0SpPVEgfn+6hs8nAgbE5dYjPoZTKN2vaDhq2alNrvAI9VyY5tKc+yKf0fh
a7M00d1Nynqt/Gk3p8IbBo56n3SXsxI/FQrib2XLEu2EzvqUbH4vGp9AALWNgvdr
xakIP4d0YgbcLakJJy/3ute8YtiUHn+5//d2tD99/0kT5YT/Eu6N3EEIivPI4DZW
/MarXuTtzSMrml6WL7wapIgn1wD/Srl4hEpF9tV8HPOcKx3074sK0ra/E5m+kKwA
+dbzf9vGsSb+Xen58WjN5ua7aF+HNGr+GpFd7db9tBRFCIT+0KX8O/ZqLDFcsTXQ
hYaibb1korv+eIR5VuUB5qfSQex4jUFkTkh82t858dWNfAPOt/G6HY5PRuExlsdw
h2jgqw6JZm8cV7/9CtYKJxDDdOstsXkhTU5kAXUmXyoQQHte5FzmMmZRMhSxg+vK
H5NfqCBXs4fdPmBOquMKPmd+9YSDqBBvK9t8yyGVOVv+nIWqG4ve9AzxqjxShpLa
SnsHlkdJYkJkq5xnqESCPMeuP0bk20OODjOc/5q3vy8P4SeUdFnlQjKht6rROjVK
95Oz/fmsbHQ7PDnzwjqXI9F496p7E7eNPtZjxF9/3Ff38pJfnsy+cwVSSmtiMYu3
0SICN92qf0zW2s1uZd2lovzOBY0skoU+9fjVWyTvK/oV9HNj7R+KB+4TW/v9/brg
Rce0WDswSwO0JCamxdpRkMCjKVHhJcHDgVITsnuasnk7m6r8bJ6crNBvMo6MFuQ5
OUMe8lhfkIL9F19Xez3NHCMkmsZduS6SWN3MPOEjSbmwBSUKbFmzECRc3nQkqYVM
WVvAwJAPs1jDivujW7Y/8tjPtXLXjL99mEtSrNNM8Ugd1ae7MjH7h0ZT2hzf0vcx
rru1LAvpNdKAiwzhM9jAgBYSMY0qIxvRmZGc/wkdmBDN/n6CZ9pTt7ODzAMuBtzy
639+FDMCeXNhMlQIrdOqtx2Il6yuN0Fc2Y6fnpjlRP2RnAwwwHT4hWUTjeKM2IIv
Q3H7vplsfSMxuqIuJZdHtS1v8Ey71xLyikiexFuE78ia/T+088Ga77bT0fOtC46e
ylMhbKZjlNcDmJUHhuo0jwxmsVuiZ8/1P3ijQ+jOCfB/Qi5vwZAuhW7Zyrv5IOFS
m+mSA1yned+XlG2LthePVmj6EewBhyJSTlJxyqHkss9csmrq7KgLvS310TIlPxLy
QmIOEG+aNd/WEVRcWarUgeZb3OwkJfYn/1qia+5mRMEDqPTdfd9xMq4Hys3SgBu9
Hr/xnkXYvz7m+dOWQ6eJkB4oUQcZ92fqWCuO62iDRYcrWNmnpRJpshU+/Mxn28r6
uWu26zSNG0WL6vxzRzYnPIf/vBKSIJ8PSXABzOK2OsVPBJdMjr+bzhH26UxUmXEg
/OB9CWfRBTbmPCLGpS/Kac8i0eGDKKdAhlupCKMeyDttt93sp12cC/2QQIyGJrN3
mBYxuFGtSrFbso0tmesZfwbfYsFhQm44btycQHoiC3luxOXuvpwsyFJxJLL0ExPj
J0e1Ql3+bihgTclBNTxzD2D5+3j8RnBl1Scc6cJS3+A7P6gjfDXxPKvVuptmaYwn
VyUb0+a+0Gdh2e+DeYmdXVibCmBUPA3HdPzZ5WozMdvn4DAssA6O9JzzoCG1vefn
tnYeDZtAgOZdenAnfJZ7Ld+D6yrnhoyUk4FvhuvuM58ZBYdqeuTUQLf6CkC9w5g6
DR4CME5zvFNMRzy7q3anLtKpBSI8Rvq3ztyaH3i2T8QazDNH5cFFAKC0Bti3pVo7
dqlOJw0ifgEP+2fIYgXTU0tHI0NISEJ3UvR3ili5lX9uMiT/1q8QcN+NWwYRbOql
yEJELyWI9QbR5ZlKv7wbD2washAGaXgp59m/S+mJM93m7JisJ2E//PPe0hn0iffJ
/hx9PafGGGc2FlLNXKlXkpANyRmIY7OpoZ1bQCi51qtttyac2HfAlReVgPPBcwkX
3jk0JuICsml8jX6KCA4W6IxXT4YOgLDwFc+NE/YIiG8eOdmu2te7bj6Dc74sgQ4O
cha1vlF+90MKnCEXM5gFKgKHtAvc+OkahnbnfpiT5+EWW5q9y07b7wdMcW7ET5u4
pEunWw7SPm6jLxBnLEDltA96Oo1s/GaeJI4upC1YXy08B8rg4Gw9Vnr0l9FFMZw+
Rvh+CKGO3dWtVzatRICTKLBgmAW8eHSbNiCqjFrsfsJo4l59rjw5A/3fsWsPOTKL
DZelEGuXcYrqwzh/1cOI9H2xLDWqg+eaB4CfKt3X9KpgvwJx9c7meElrWnx7emC7
1VxbAHjROmEFOnU/R8UH37CmB4fgz/8PJDBaKOrDKzB8WpuhuG6KHmxerYoDIE91
pmVYgOVSfTT+zZwhex5Z7sn9vDY0vaUiL8mEx8FZm74vu+yDXEb05ncMY5WVG8ep
WRfTA9rpJ+5q4mk/z5MmRlKeS6Xe5NaEhmqklheLVEbKXFsAKRia6NnlVtVI/IsE
hmkSEFjgCxy3MmX0oEhwdFocU6xb6RTb0XSMT6RQa2AlFDqg88TC5l65PUl8G/Hb
8Owtn2BLC2EdXeFiUkEVqUzG6ADqH6D01mipZN0TlpwI8eqMuRodvgdbbd2eQ6iU
48bi0QgiGRsLSU6EQ/R5WDw5TC25QuhpTiJwbCz+V1GKxpnqHDbXMnGerYKWx4So
o7lWUFgdnCq8iwUp6Rd5eb8uR7hs3oA9psNADcQIBao8KTqsEFp1A5QYCZ1ajA+t
eniKSzgorvh99HN1IcgctLSWjIIldVn7sCGFBMUSUTRC2Zz+9dtZ9weRms3NavuM
k8J5bguANywQltbQxeE8ThaaRLzakPd0ybsQDfoCt3dKVRAdMD+BKe1/t4prEhS0
j9zrbmpIaPbB67EFNzksWRWwvwhXvBgGFRP9bHJPcmQAyZoWjellbrtAnjaZBZoz
37nEjy9WqR6QBIvXDl+qSHJev6aWoGlvjzak6jitnosZRM5x4QlVTvYwCnNDHMVq
lIqyHfTGozsXWe+74sIPSSJpBNAa7vJ/8ODn/KUkOyztB4+F7EskTCX0oQLQGKfr
fa6QotAX5zXwztJ57RMBJsSBPfwyZD326Sir6WgI3isT27NlV3UBvUNvCGJMw8EK
+TOXyPCCjORgzHmSILD/QltWVP35+Y5QBaX1eZLtyLWwdKxuZZlN3PwnBAuolUL/
EIMFGegDoT9gWRV6KXLDBAyULc0SVExXXk1lDPSjuk/DQ1sHPRvuBy3UT78cpn6F
X5wj6OCnOJg8mz+aLFcYapHbtxpxVvlBJltRH4WYNh27fyVxH0J6ryLWuRc9ZzUd
xToNIgrhcLM/ujA/bNKUOuUd8e0gk4oaTpMhmfIXw25omnQ32TKSySuDnWgycaSE
JcR0LrlP0ZeLdLNn22bbJkym5du9hYXChZemMXJUWXFLyVoX3GwKAhGx7mwNViCt
L0sQkTrbILJsGyVZGmhsfqtp52e3cX13hXpnyn5i72EAGJxv94PyYiDtI9f5ZxWT
p6ygjXobuBMI8Ilw3dv7xEmhhnisfDpIZU0EZT/34Fsy/A/3NgOzOpzJZIb6E6Hr
8fcyY1bspdo9VCc10R0NeF5WHw5TlFCvB/KxpKHQwtemC+9n2bzhZR0VrKM6mgDV
xBgNUjJq9p6Kckn5WuwDhPVAIpn25Whewpxa1uR6Ohbt5L9GZdSnEh92ljBotL8x
OHRvepYVfZDfC6uVnRrR5Ej3885601GDWqfH43A4dSjZ8SKQjplTpA/1bPajxttR
UYd2HCgOeVuxFd31WFQFenpyPHTqEQtN5YbN74sQ9p+Wfzd3/Bn9TPmJn4JYdBQp
bpcaGFvUJxM4nIZXCqgiVI8LYaJvE0/UYIoQPX7D6xW6YaEaqVXuOEP6/SsTwHsZ
nGManlWZvzXmpCGlMqjDOJ9UkuYCWSc8QBkwLIExV1bNXJvnmgoW4aIcUr2AG6K/
qVDWzvkMVxypA8M4HbXiCs1biA0O0dPGJb+/x4phE/ML35od0k1s8gyve6ZvgCrh
EOERTLKu1Ack9KTXJOAANK+cp9ZyqXgtIWQ8biS94cyghP68LGWIQ9JrFM8jxU83
FnT/hRPCx5y7+bVeGTj8PnOq/9K8g6cJPySMfZTBNcmorxnbogiJB3TCK98YykBt
fGvN/L5hZjRqoXGJxDrYQ5qjEmpi7WlfAnvak25tthW23s65Zpl8aGH2FKe8RRLL
xEqYwVtPKDEn3+aWotVAqo8QL9blQIKq9G0dAYvsoVOTkSNGFLU1OrywYXYID3BT
ho0E/ujBeGODZ1zKE7uf/YYkK4YqcApHglckg4ltiTlUiMupUgDjBLn53aplWWlL
+JIRdaDdXXqHCbpQCZgOeXEQzjUTn3f7cuS6Tn35qfbPWlhajca4W7uKlEV3Iayp
LQne72BSLBJxYckWtZ4/2043f2g3NWeJW6UkKZo9Ae1ZfxwQw2MEDsr5B7rFhDXo
R2SxkGcnfKQYKbykr2io8gqGFoIXNhNgVR/gpeUp1oZIvn//HIW4Hu22mufHtBnf
Zl5JZEVPMQviN1kOxla2kiCK8Kc+PCmZZvJ564RKFhlGXQH1cXEobKDpOaeR5GVf
H3EBGjBxgQTGgTLIbaA/MWkpy7EF8/CbpHuptM09PHgZ9qlNBlMuaorVqQ6uEBuc
jw3ZncIWI7NRnRTNYokULurFaDLA+NLktLD5TbrEkA5l5mTGEhlzkhevbNnog6RT
A0mNoMiKhSFIX22MLm24JxfBij7RbGaMytUrh0Hepai2UQxmscREiBW6quF6aPjt
pxI3xWCS8I6VwNyZJVzMDC0lJ06hgOo8ARaNItOM2HSfPj2KzAOc3K05rf0qtwu7
zXmvKlsmD6kbzfWZLqCU6y/rftuD7Cfnil6bb7OZbj6DxmgDDfL/ZZEv25HxZ5EV
XeBbDcODvnasxgSaUJPMAAq8KMIYkx0yVanfqyFmxKAvCkJDnKTEyrL3KUONN7lC
UHmzBBsnt76VwDDTeBmf9Fg6ZETvccxwF0ajVBUT3kcV6El7HZlQZes2NVMuk8Ip
1O9JrP3CR3PdyO+tafuZUEzM/IecSdr/oDtL1BKG0J/HolkLOmq8O0QNP/ukDq5Y
WqSMVUc3vnbP5PZA+o4vnjXWlCD7K4aosfH8Zr0VlItvh21Ty0S0J1izgqtMNdzo
LqzlOYp5nX3IOHUKP9Ro/0Awkj7+Rlcklp8Tas/duZQTKvCElDRunJ8zKHbsKjwd
vwpyTehhzL+7FpdAMyRAhk7eGoYmUf7jZv3ZgZ9NsJwYMxdNKbt37kVQTn/ST22A
mK3MCkslHEpJEPGIYMSItOMHSAYG8IjfAyhSOREboRfhsJvqFCuxiJn4JrefYE9/
mn4TKwklaZm3a8He4C2jxqe/S9CI4O2cB3ozitA77TD2HgeDIj/IhyTUqn1Lex6w
TLThky6NptktrzB94mS3A5KdGp93ijB+WVCso5xvPOuCaVmqjMtDEAeM336tp3NQ
87sYQu2n0AOqzAau4wYPPYBcxOu4KrS8Y9cRebbrhKnsChFwqrTGx/ff7s3ARU9+
/4OrTNzLGPWs6XKCeCZUcQTZQ3u3H4tyWWhWfHwV2Y8ZVxbPbfgffKy6ODPV2xPE
npHE6BVkQLjZFMXlxAtL0Kp+Wq9bP8Q7kGZPBH/C4C6T5Xy9lQX3SBFKxd7APrtm
/+9JRFciJ8X3Pu2cYAoq52jmxUtsNbWYiJqgqfwobfJOPBdoRb24dCEXbP8SbT0/
NIdN0yn2ac5Yr5oKrswYsNEM2ngE40l00GouPeeyxkVeFiIIRhD/TOYZgf5XdZoX
3v39GbEU9SqhyR3Yqbd/CZaMQ1EGUyHXb8Exgz4eGnwDyoDQLlu9NgEhc/Qm0oIE
T0J+T08bymNze+1vflgnhrgFSQJB/YwAPu4VLtOTxo2Qq69H+IrbT6GhSdiCFzRe
CLf/jFKTknHQLUOCyASNT9ZB5/vCyojBM5A+5xgE6SzsRgt2ej7p0u0OuwVcgylP
sarYpt1v+qU0ZW2ua8jdotyrzoK+fFd70IHH3g/01lsZx5Cm8v2Jyx+9kfYU+M4w
he84BEAIHktxAWXJ3UC/vSJKptRnuhE9U0vj7hAl9tIg2r+fTrDtCSJMMIHoLr3h
nKnwRYPyujOFb7hhLVrqP7fSihQcjzhZmWO/1Vy+wg6TkmksjVitOvNQMhg1uCU0
5TeiZRdTNZfSP4lV66yqq4z171aW84tuXGfCe8kJsGuwoY2MKxo7K+GgVvV4VwWQ
o+BZJ2g/fUKekn8P8hMWT6bj2DsUX7SOZdQWRvAc82QUy3QOZ7LksxSSGelsUiZO
S54yh0T3tsd+in1v368y5mM/EDCp1zRpfGfK/Dp0xAkAQH1/aXwoW7KKfwAakODB
D/5avDSZn//NVXXDqQYnzN3mK/zo28xGXQEwLIS7ko98xLFFP/ayw+YlpHoEGQwA
6c5NLSYPQnZNY4P8ax8o4AIRPq7fiWltThdBq3UWYIeU8R8/1Nk0ELnI6BirfXn/
OFyYOqs2eT+rSwLpMSjkxGoLkN3UCfDb+CIQK9NQ3BYhIXUwhTvLqkIhc7c1ftaO
3dBnccZvnrV+1G9lQ0LNL95byQUikZGlA6onLd10I4apl8YKrEIT+Tmbuoj0uH70
VC8JHc/2YIbmbGJSpCn+sNM/i7lU6N243CQ4uqrWRdn5fgz3KvJhdtOa6SkZ9D8F
85dB/eJOm15283l59ZOB6Lncu362gH95cG6tUspRb9/htHOrAOCO8pNEsGAEbKl8
iSYs3/ZvNrZnysW0JUJJi6UKvfLdMlhxbJ2oNnBQIWjb5fvtsBDAT7WToOeiuFGD
LDGKc8CNsHlOcEtrkpPO3Gl8E/k178KR/L7xbvhfZ9WcyVvUHyOZBtZgvivzt1ZD
/skZEN7qWXN8QZdQ40B113uVtOjKW2fUBiZRNy5H5Lyg/Z+h5i03+y5VNaxk9vHb
RnertTs1wcDGQgMOMej9X6vhdAW769K4p656+M7cFs+X4ZjRliA7/pXVZQr8fgnv
Gt7V86ZY1LT3utxaSa8pDu9fLQu6vfh8NSbqcwT1BZ2yleyjWxZnfAkmAcjH3Xow
rOnd/zUY4TZIHwxupVXc+KfumYWJgKbtjmuxqbF/BjK/2OnWxlLC3yuzw7goJaUf
8hZE3bp1aoFEZntXKuJKkPYoRxew7WVna5FqUgMisX5fKo3C53oY2Qb3hG+Ph8Iq
oiOJOr05T/iUAKEXa9pqaoTtkr0Wr1tG8eW9doenf7EGc2A/+3fK8qMgyOPQ7vG/
BUqVoZsLZbh895GTegaSzb50L9VB7kMzrN6kSHxORbYyfYeoF0m9VU080xnUA96p
fRPd7ehhJe3z+U78LSAAXrS6V0/t8WZdwnHT9ooMGjzALC6DUsMuHW7BbQ44JXw6
yE81v25CGYHRD7zgvAS8MZsbY2AVMMqHDvXb4vBwyNqln5122Ba+CPx33sWEGO56
pxeOC93e33x/3OG+jKPhi6JmCbpeFC8Up23oxV+T0lPKEv80JnFVrG6gdz2VzdCy
PDYlRZ95MrQOAI1nFmK2jJU1Mi1ASvaeor1daPH/DNxQO5VZz1ZqWQV+/LYpLIf/
KGhIQFAiApkNfB/JTICdAQwjmeu5JVz30sDqNnZsR45z964Wljr1LntMaCClHD7E
p1aQHJHKzKgK8P8I4IlGI4cWwxdSgMGrnesW8jRJWeJRm0ZymH+3v1osfSVgp2f9
OUR2EEVRXsM1YVvYdRKjbQ97fGOyGigi09f5zV0nRwXC9AIj2fvo/7kqt6lqNGsX
SkSSTa2+f3oXNOMKY7bZkzirWm1n3dHuLdwajfqBBbFGLVl3OUwK0figKp78by7r
1X7jpCaw7WNomc83LWCa0YRQpQpJ5L7cD4/7s2ml5roevneOWIgmgLSiPKUlEnUe
GZQ0buMGf1vLjZdy01IHhbFaazNMwx5iffMzD1TZ98d/gSo/hTB2l6X+JjobNcfM
6fdzaGw4FgqdWAXgHf6meMEDlgi/ENe/pnGrJgVV4LqslM+rGqkqjGBtE7J09Iu6
T7n2mJWCcdhZ0wLJS8N9I0c9n7r9zP2ApHhjJ5B24QjFdP0E5KSVTqUVQfx67Dvd
hWDTtb4vZQEJfXRJGFthaF7K18RqfHLlZBWcYB9twRgEwZ8BVysYmZUqqfrYY8dL
1H91TwJkAXX3+SNWSGnLWRPAa0naXNKpeGVO8pEnqCQl0vgWsU2FPSgOeMz75uNU
Vw1z0YoHDYpzvucGu2j5SCm72XR+zjRvwrWkSo0wZY/jbY+fHvMTrdzULLZwmCRi
5pi8Crxa+9+WeYhLlClKY+LSAOjYvV1jF3FB8Qs3nyugN05S1oofguJkuZZLNgYJ
oHWJNXvBm00qPNTII4u0nziIaNHudzXAi1+gHJkqHMJk3mrWpiqxjqbzqQVh0/Gl
WOEk6wUWQuflGzwFZf3MAuBRxq4WISP4D2YUb8SNIjoqLxfVCRi3wmro0Uz9DX2w
KmdeIoAVWreMPA19GsL96R+34O6mfWHJHfxR7/FIeI3BGr93oVEKpDlGwQf9853V
+oRm50scs4JFG2k/0tJ9Ilgm6rMixh5WwVwsVVRcFM3gERUH7zQEBm8qPfY8Gn9n
r+O6o0prW2K33ESfLHat4Q9LWjmZc4mB7bTWqMDDoVPjGbHsia0M23hPgFnRoRJP
1ktL3yhYUJl7e6sJtiJOgbtswV6AtYlAJ7ikHNQ/4zAFnCpsrZFiMB4rgro/rWn6
cB8GUsGbO6V+1LFjsHNKuWkJJP3mikII2dYFSbBf4frDEVo614xPhq9jnICFzaKz
Z0cEcOHMoA9qVJ3KZogJmM0u1m2RydNx4ELFYltHdwLLW++vpTufRXWGVCch2kq8
R1c4W/rsxxG8eji2Y9LKcgtcdkqm29x2pDBeg0jWUs+QCLDQ1CqGG+b+/CzMp35+
Dmam0IeHJUph4nI6btiPtkO9rN8pg0x0lFd48Jw4BM596L7RfXSuFZBs4nCz9P1w
5MgjpWZmqNBZGzmFB36aPPVb3MvHJsz+pFgAbgKzROfTuRR5YqmJ8Ekyv4BGIBkk
3TJofaDJ2Le/OXj7dCP4iPOIS+Jp9FUb1FPgINzpVyTQ4iwvOmZIWueRAbc31DOK
nrUBtn1cFgcS4UjW3GRtNpQoilYq7CCEOqGkIhuxSprjvS6QWYpyUJRC1k9yp1UV
sslKC74qfPlgeUKCJCddkNJiuNFuDGPI1s+rKsRXd8appEskee81IZsDckeboZeK
H7Zy4MjDmNx2EnLK7T4les0B670PN9nk32hao+6RmKZT3jje5oAAg3SnmNhdukFD
SReaw/XuijKiCgelT2/FJ51M/8Y9ACL7Q6Ol/jBVnhk0wT2MhQi/bPcx4B8lv8We
B/3Yzr/G64Iutq/S+1b3lh3lUZhyw6f8ui2PCVv2baT3J/SrVSJKEyB8+OCt6q1s
0T8yIAvDxSbrAHNOgOx52rHR0x91MmxZrQOH4lqizGZ0AU3p1sMP+iCYwdpF1XYh
e7Z6/WGet3BIEugll7hAYxLO1diJ5ZcatO+IgMJMTVxPVQFxS5fo4uLREJRXrSOM
PnsYKfjowsz5FCnVgOZCvMzfS+zYYMDZLwWgwodQ7c9jRRnUOTKsTGAhhfreC+JU
zymUXcHXx1PSBmrgoCLA2AmVvui+IBguCK45FfMK6jDr463qN/s/WEG90gx5EvUg
neQK3K6dT6dPx9tvtceqWszqGH4CuItqtnJFc4xHVF6f7GGxwjyDdAgEhhLiZGQa
O/N63PZV+stbQGdB8KEIHico8K4Th9UbN93Kk4VZfOx6M3xw0A9wMJxgmSRigGTI
2Ae68CR7TtPvTgZbaDXbCvzw7L1Qvs7O1ni4cQYo8qRwJBjJyKoQT/hHEHwyh6fe
vWPSbDXMxovTlKr/VQpayq0WVqtE5xixJiK1PwEcL5FIqa9OiO7Wuwk/tIZjwuKY
HxcIbwk/vCX+1UsjXc3Fh2F0V7H0tl+uX2pm7wcCq8MuTjPGmY1FYqvLcdfPe0sz
JXxk628o+2CRHvAChCsaYBG5NmlGf8FD7arImlMksWR1KCB6V8LsBub5dQiKw9EX
MhivAyRJG4t/4JDM3bwsgbAemWM9sUSDNVj8lt5MM9jd6dK4tOBoEO7zFE9jwnQK
tLWUaJTWopFgGBAe7d8hqZ2YVe+nsxXUC4RGA75BbOp33Vc+hgcl5ya1a1knyKBP
hzR94eLXq36AgPyPMWvn8CC2qP1BJ38Gk9FBBzF2aVRDxkL95C/QvV9Sg+Q0y5PS
hPN3YbQkrgvGzXELi0jqW+RJX9R95i/VhKvHDpnFQn5S7mIk16wlRm1Q+YeuqpNh
HqXiO7rYyGD06he2MAABWTKLr/g8dJx4VEaN1bIUN8uNogysDlEzby65/LdqmDzj
IjkIq3SbiOpNI0oiyHvuxlE4DNjUxYQBWqQy/6b1nxhvQFFH410kp8HVOawQMWzw
TWmaSSnfcBaMDP2LuHRmf3q4/QieLuRKH3DT1KJ9vAorwJog4itEZnzHy/kN0rfY
EQQBVeIzyHpvlKZFVJ7AQ+HX7YCMTWdDniAN19aDSLzDYEgtUY8fu1Ke3GWKUN/q
qIgECouLwOCNtxs51ydi2wkg9TPqBTWtP7xJ/EAe8VOwh2/wR5XAIN7bz8spmcDk
Z8GV+gomRE5WP7/aq7kz+l2+dsJkuBfbvQWx5gj7AxuMNnKfQdWtA4W0CiZCnNvz
eFYIOOFQyHaRywA2JpCBuDj60fvLKT23ZeDMp0FiEkE7iyzFItt7YkbQUi7mlfBP
goT4QZHxYp2ipA3TDavpLDFqInji1erlBEu1zS27j/mdCrHvAVDigcWiwlFrytUG
TWphIhV+O4ZZQZmiLSX639klebseYPTIZQNHQZyssKky5TPRATl/H+HqssYzJ7Aq
pLI3HutQBA/NODhMGPgQKBNgktKN7be216Y/sYk3+2/p8zNmzrpxh4OF09oZdKM4
nnFlptwwCB1zfvMpyQDrkfDUYiM3tVd/Ppf9U1z6/lfeQ7qJCDkjzEWmkezDmWiA
BQnnQos1hV5XoeCS2oooWWnXoR1qnp1bYrW9o0Gf1HRdY955tj1ICUdq8lVhc0Gi
7TNzkd2lZ8D+U8GUQohV+t10Gfvbmgd0VfS1ZVRi0K1zMdmQfz/QanJqrzm2u2CV
VsA+qmk3PgovPfY5+9u/soIOkDyb2xoEfuJ88uUpFfrshZ7RiJ+MpB54Y9TTJVDo
R6jHkNBySxN1ZkG4Cl65Wsp5ITYze2wFtPlCvN++k/ZUZEMUEYDNxnKwkOwtXbAa
QTYI+ko2XqtPM8qe69QKQJ+bGDpboYb0wOMy8sW7sChTezMYGPM59cc5/wb0avC/
n3ndydEovfRrh/vmaMpvX2W+ByTrbtDoBInvHj5DYt31wQ5rV04CJYX0wqF+yxH1
W64qX++Kl3tnfgLcqQY+uAhpbChzVA1yZv+8nt4IXM/4CKjlFN3fbFcBFX308RZt
DQe1da8NqupCwzpwo9FPuSJTOhKsOOKqDn7fMDNfkt4EvXfFejMt2+7l1Y5D5rca
qDS3lupKSHXqfXqyrUpn82N38DR3bcbVvGf4yn0mA4cgDDpMYg+RFGdkrzzNdOes
HBUgxibhIRgvSIEMuDDa26VLzhH6UGIhlE9x6q70LsSkuacbu6ejMEoKARKLWb8E
5e0oo/HBW1C961kJlmu39d19Lc+NDzirO9Sa+b88lpN8z7dSNnAEX1+bQNfmVYxx
MhWA2HXmLO+C49/blaIXyNTAbAG+PBem5239UFoYdGPCv1TmonsPVA11OuCk3vGQ
0RBKWoPeWd+zk6hEB30fNB8Xhp9IQ6hRjWP+5j2OIX93iBLv2X6M601rV+n1MRK2
YgyvFmwcFY+nnoroeQg+YjxkonrDgo07QcZkovTaYQMq7g1VxMCRkqB3sXsxM4JO
BTIaGAWF6EW/RYlSnh9G3w/1yM3Mr3p00bNtL1z2n+4Pvmg5jdkIeco3Pq61Mqr+
IQW4Eef46Ec26VhPw62u4EnR9z/Q3JFGZs4GmUb8Dy/Dca+O/OQEY/dh+pzi2V3d
or4qYknAMqvSM+6rSu1S9kPW/LIGFTjbJx2NrT7jSDg54nLkbnDRe6+qh+G6aZng
GY5wa5/hJQwa8uZM7yD+18zbr04IkkxCXMIiLiuHJPD0A8EIDoxAdyBu4yJM3Os3
3BH4ZClcHuNltgjNpktkJbikl2yYrnxsP/vhpmw2fK/KZyC/T46RRiNK3+S0tv5W
6CNZ6hr7pMevyWgVM9coplzKoTn8gY9QTHZsRtCkyQM0W7Q418V2vAPHfkpfvAGb
lGS1JbS8xOhpJeXFZg4XLIIYyTikQPFDxKMRqs+72ewuvYLfiSsMd/OQALc9U29N
cJUYa+CYKcYxRtuRU05KZtwcrELG9paNbhfIiDXv9tUTuJxAiPoD2NW8/mc7HfwX
Ju4M8EtenW+UNDFGnEpMVFAaPawtCCEtv0ABXSPFb/pWrrmx6dgY7ezxMUem3Zd8
wHny+uEDOUa99ro3oAVjjST9Dl9qNo2YmeieNZC1obWQFjP4xfnqgQsz+L0FtjKu
3g+SwAqZ8YLDmYrHOw8OHamPNkuD3PgCWviPsyWYLbSLEMqEALo/bwqMKm2DL1ZA
ThdN1/Hq0DSxf+2MN2o9DcfQ5BggYZJ6tRs2EZWdj0nFEJaZ66hZ5nFsQxCUhS4A
SxMF5zhg2Yt1sGCZq8hLJDUzp9kOeaLfwxpfFNNFD2ty6tK/KdC9Y+QtnHZ1anNL
ekmh/8ypBKJo3EVQmJZbHREp+IyOTgWSwTvIHovUn04kVSj8aO26c/uOwyGrGhTo
UifeELE/M4uHK5Ks2CLd2QDSobPN1vUN5ZgACJjCBMc9UcAfPhd8/HrO8umg3rzJ
S7bbFAuN8URU11FLLL4+bJ7VP/LiaY1rJQl80U7PIdRlWyKPo7iCt98IQcfJuanb
r9iVy1HUwhCT8mIqdHBgVOWdODaVmo/pGnzxWOANtC7yyRHwvE87yJWiWRaSMYFO
DCL/QRC/l05DAgdS8ABqABVNT7w2unJraNsqnKH5MF9iNBd97i+GHQCWXLEKANq0
vNtEMBEeWZfCQ1E45TkmL4tsWr3KSoFPeS5cnXpZII4RA3VscV9bQjDq5csp+9DT
nmUPc90br4xvnqlUAoBLjoSRk/p+N//CEXIBRJpcSCNmM6UQ9Blrmp7uZSh/eJiy
5Y/dpd/Cx7hvmkboUvKlJtvpoxUtJwYTAhVTi3XwmaRXk4lPqTT49esljZSrWAPB
GKZaUoul4VPgBDTpkk8vXYOR7vvTTc57kpk2XpnrQZrBjQmwq4kpOCLzPXqRE6Tj
8wCUI1WUC1XSG/6/qDo7vdQ8oewZPbXHzVK7XOj+NMzEbjhOgdZpYrpm9uKdLAgT
vUP+fNcoNexvsrWFpG7gjDxFO9JLDQb46vFlhTjpC8ktuapLUN0q3tPtUuSsDC6N
PtU66pDE/tPecczgqMRvyWDgUAth0kxk1JGvFmfEVuRD/TvkRRqM7w0gBn1LuO93
p8lf3G9cFzCUi5kuj30CtR/HFSAGUKmQefSPfoQLfgreT7DJ5Km0t21dCQXTT43D
26j7V1CoQG0pU0xmk7HJ+dxOA9EUOLY/MvhP0QRb/1fNq5JB6Dw9wm7koA5JQkp1
8Tv4RptyppisShlJYXajSyNwJaYbBjMmxhbbcUU7P3gzxB1OpPgF69VcZzTbipIJ
1r4e9SxWR0CobQj4Af1ExtGNMPxPaOpXDFdCWMcCnbZBOpJN4HvXav62DXJBOBXN
8vN4UgjXODkxrCuAc+aKLanGVhIoNqGShS4VWswZ6mlPPcaMPxjfWFeTmXHEuiDo
pDv68xgs6Ab6nTB+OO7Ltegu/Yhq4k3ivcuq2K+8mJrk63k7vZaG9dnPNR1ZpHSD
KotU0Zl2FOoniV66yIFPaouuTKcwts9/ZradMRs1pvG/qTbGgEOqSlxlZB9lyw0f
htOJAqW/3SKMLvFrSe0lpvcgxaaiBiwz+pJXvvMbvXkQC4wDgMGqxoVumPUkV1fc
S6vuEPzOgvYA2QNk/shX/GXrVQJGAJ87hYP1dxkx64x40pOIRHWij+De2/fauydQ
DSwgIfcARLF6rlZmISdNK0GIrHPU8WltICccIALBkhF9axPAJ8B482JYhNrkbego
T2znYyxGj0X4XYQK6V2aHcqL4GDw7l6AIAeK8hd8zLcr9PYFCzySlOV2lu6foTA/
cUACc75OPLSdLLcXth6+Si9FGALWE8+4HiokK5++h5rnaIDAgH71Bh2HyFGFJRGA
kLPtuBMWw8THxuCpH2Ri0WhfRaFyTzH8i8ZxMeSwKkJVsOka2elK6vh2tkpZQ5M6
xTEGSk+01+ottCL2vktS1nz4cCf2Q6Dl+kuqJnm5saGIus7Vco0CTdu1JIlXDh3z
bVbz29h5PKDpZx1Is9K3zqFA1+kDVjCGn24DKKQdP+GxzwTwuKQYqBkA661LRTP0
7ZGMdPE84qhYJW5M+PyIHKWx50hLY3mHQg/YpoSjOpZGvi0KsHTlYnyqvcFFiaQN
IFfv/zWp9uHA4XW61JI0WXfnmxePMvlqGUyDo3pCHNELm6YXpk2tLHLht+Yp9wFO
8V0wWSXsC2l2HxbnfXCRqAhgyb4Kz6mxNxoEVcDRh49KBiYtiKufUA7//SoOzXti
tY2PMC0tdEhQQkHGKSaqJvQx5lNvjOlh0hqJ1VshWVIAyhQ5aCFcWX5ZUwRGbR5U
5ZfPL/HUcngOuEbcCH26k8UsrCeKFDW47HR1SgFsTZnqC1BeUChLxJAg8rLwFeNQ
VfC0eW6WRdtFYcC/AiKT0MHUMlUMUNgvwB30/5mQzaLSyr13P4FnKfivAXIwu48K
cmAwIlRTiup7Ps0dJFuKo1c/LPk9F/YvdWjTg0Hdh1uBE3wdG9uVc1Gknx8ROHKX
gYbpe32rTNeSx2v3CIK1/VfsHYhMDB9NmmzYs8BnuOe6mppUU0Kx6aUnjXD7jeR1
0qPimf5nCvmiQEW0u2CAwsJE1vQIU9tZ+y/gEDjWiqmo4hwCZGbbNfSotGjoj2LZ
s7sNm5FzmeK5BfzbqsWDBZqnDEPNHjsur4QzqWlcSbRe5ofjY4m1cLMvrQ6ExCJx
SahH9qM8n+eP+nRDDZwb9hsdG1z5mTDwUeAeGwBILvx0h6LCWh60fjoRi4lHo3N/
MHlAMto+UaFQmAbCTSi6m66Z9YU3kP8xvO6dxudU9TQr/ff610UZzs+EKgKWqmal
lqvpAMj7xSfsNRKcmNLit0lNdqLxFl6anILjKrMsCl0hc8MZlVyZ+u0VRoW6ZDtX
d7ulYaQ7movMxyqoa4m91V5eUiF44zXHG8F1TYGj/y/454qh2p3xnap3Q1FQRoCV
jVpEW8teXlOtOpCPNOYz6m2Y/eKGNPBJ6HA/78/91YGAcLUHE++L6CzW7nA131zZ
zrwDLjZiLrea7dPFxlHWBNHsyF1vRPipf4/Mb//6d72G6HOB+/2nMcliLq0bSWAf
tA+TVhT5LTdlyRVDX/3h0XcoXX7BmPzHBvDquT2zxuakwH3R0/g9bnX4UPlFj5vG
H+WqIliiJ658Zah/udaUo83qQe4uvnPk6siGodQFkrS48zEmwNBHqfZbFxKPT7+I
+5DxC8iuaJif4lzlUrYeZ67S29C/kRXBsbdyoHpYjd07gy+IB6o30MBbEQehsmm0
ujqxbCzhlb8ucyuFyyCAOZuqBHhAJ/HvWBEzrRhw/GVHtDuzP5YsUF8vTGvFw2wQ
3136J4aPAwVhZLhuAyGPhkOROIse+qNQGrAfLPFeWksw2HHEdLbLZmfzLSBAIhVS
CvPQimq2R7Rlpuhv0LyScSd9vrbPtCnmOFGF9lb2N7fdBsO1Mz3FWmTmwtqDlPUr
FytvhEOrNYr98oyk2q839zrTp6y6SI8FKlsBU+8StE0aloT0Ibf47oxzzXscH5kU
AAtTPRZzaAnL8t/0eK60HiEB0jpr1kJyS3OXaxXYi1MrdpDtaiI1y/px0JyFrGtV
lpC7AYo3CB35EMO5X+TuLb7uqRnnrWGyXq8WslpBUpg4w6ejrb4Q35QjpEGqg7Te
zBRlPv0ldYNuz6o0oRydmiBbji+KheribYF2L8Ohemm+DaAYH6Pkq1pdBTUjzThh
n0F8eGJfdgJ75cidL6A6Wtwbxk9LEEth1fRviC7usbVMZPRo9uyNixYQwgo5H5V4
Uz9SWdRvkwOl2AuhTzfHYXJ1ERhnrPOGfQBLSPdG3MKBfrSGGto9cSkPza/H9mtZ
S50CIYmKvbTUp9f2PaZ8WG7l48Qt+3ya699xCbAJ+XPKZobEbcvoKEANWKa11Xkf
bC7drD1HKh9GgAColUxBDb9kElysF/vMB/IrpQtRh057JfsrioDp5qHuDgSv2GTe
kQ2U1anHf4kAvsJ5cM7UX1VhK9/oOZ9o9bgkt4GUPF2xvfO3uvQaIdRPb2qEFWq5
3ar4XufZtPkA4AwY68At0SdEZ4H5I86koMArbGd+hROJK/pIU+lk0L2YRn9GRih4
Yao/EWVf3MJmHdZsmf8Q1aU6lJvBP5i5NqJ45HmaCQdHnUCHUPsiDGbT/zcGFZ/5
lj+BVFR/nLOubNnpqE4933wSOFI3llHqvkn1g/o/0qf528ZyQOsu51G0E1RSM+Ar
yMegeV5JHH5pUrInYorzBjhlG9dqI4+2+V605nOFVDsKTTqJE5KOenrdja20+usu
8ROeXh8sMAs4B0LTeZey2ZlL71qpLdrPksn2Nc62Ewg0SHCduDQ6ua8YKE4wrD1A
PUUw0zreXSGchPokvsXAuwecTZ9qC6SQN0p8gaWsH9j75ROvGG4jxj9VIW6BCrjJ
Fmp5yIAHY+FHqqJFXXLSG7mdwHGMNnI4l5GI+4x7jx65uVB+e0JYrO0WhAG9AWnj
gKO9EaNT3zcnmCj/J2IfN5LaeB23NPjB6dHOCWxTmD40iOlznyl+a64fFYfyLYlr
qjXg6xCw24L/5OLbip28W6G0FnQAi+jDCNRTq/zIIH374N5mBRZ4GPVTpoN/GqtE
2+snWAXt/gQlAoB0WYySUFFxqNSl3GN59YvM4drIeSczawMFswyNC/kYZJramrHR
gPiUWVI0U9xq7aQcYGiCex8XXkt4FzQm60BLIYK4UlSJgWrtN2k8Lvjk08FRFk2x
UHfQMbsobUDfuWwloYxRqtQS2ghduEJXZ8M9yUYMvqV4JAhsYwDe3WoIYJgHCuLh
44oCSKtGl4iUKmxuWRr9PrHogrx36wISWc16o8artXg9diys0o7V8xVwghb1kOF4
GmLkW2hhlBZX4XvApd+2B27sAuZh4Eh/22nc0mteaC4oZ/hAXSE3VvUxQeOEi/Qx
EocgxW0xPkdnBXyDYL2sLuGW1g+Ou2M22XBYRJzT7PDOPyMxQg+e02D2mQG15ZBf
LKyCk+2i6fuzsC8Vx5vErv0bZtjfjKbbaktSGJh+hO0Y1iifXQDD35qLhDzf0XPl
7zmujbWIGL2xrTS5jQexRv04doLqEFWf2+MOEQiGDqO1FrsCl+gpW9/GDAmSykEn
Hy2XVnTYoNGywND7hqmeo3cI7dRECOJO63B+xcjJCLia0plxmyFVKxniYPPxOU8N
ZTN6oWKvEZ0tmxoWmZ9+xxdFp4eZqOzI4QlyjCSWLbiEBcLeNdaZiBr7wQ3D+fuw
UsBryD0Akg0AWeE65CComW/Ksp7sn0I4g/JqT4VghQSDyyeeneRfKedXlPdxbfuD
E0Cu0UqR397fJUEEcFU62Nh5Iuq+ENxF7vB0m1QES7y/SilINX4XNzsWdLWqNUgZ
PTZmFY1t78J9kdJAI8iBHBEVLycSnQcW47v3x36gvZsVrKt8wwncigg4QLivMHKB
buxx7gqOjgwRaD2tskOw19E1eg1BGJjDN0Tjbvo3VkV+y4JIeFU4QoxJnUtU+1Yg
JmJ2wPdud9WuiNmodOZvX+XRyTyoAoYOmdGllLPyvtzl/d6fxQAchBbY/ZBA0m3N
AR7jKjhLfnHWoh0AJ2gq+6QRr+YvCTGndudkmiS27ItZssAjBoBdiuhVBFLIASFu
pbHf9KdfIhQgOGlH63XZHQhzS1FPcKPVMlrhhRRMm4DO6ZCi8Vfk5/Y+0XvVusuO
fdJMhq1fdpCie4IOKee+tW0ryKntR83dt+m4063Tcz63zRoSSJbfx9AACxDQyXI9
gj3vH14sazcdAhr/Tb8GozOphdKNVJiQjh9XiMwIrmvMYmUqKgla5VU9sRqD5s1+
aJFab7J8+FXYQEOEFcZxZC05SKQ6qpI8urjIuLyC4iK3SVuHWnfQ4qTWnsYNDgn1
c4wUP0ne4VItJcgixvwjJG61DVQVE7v8XHuTUOiDhrDI9D/v/B6MtU+Z4hZDV8lW
4kk+QHUnWL3i0oltBRAnJQVlaLAlWoFd6Rfv+MzsupsW0bOdBeufUhSc+CP+y3GB
o6JYHJ7LbU8QABX/Zuv256QX7VbNhzJyqkLRlOUSpyd4H5ZZsDmVSCH64olsasog
8Aw6+wUOnVvGLaNxCS1DIp5FPI7i5nctDx/0KANQdqVmMVM6DFu+h46TxQfPQT9i
1x2BSuf2MiF7IqgtZA1ewRS3dassDGxBjWQVm5X054SqJcpLs3TIH+7PVVChqDxu
lsNmArrSDBlEM6zo5mLkaRcOpX4oJuFEatceFW1rsgNNZoZ5nySSJ02cXv7Z2nM8
MNEK+eUgZsc6j2frSXIMO+JJ+j7YTaorodcmcO682xW+tDfc+SDfkgj9kPbmtjmO
8G7/o8Vts47niOZ+RoCxNPKlO4vebU7e1A8UkgGDhmopvYMM81pyLtyyenODVm0i
BTgResNSha4KeDlLY29fIXCyqu63p0gPKfYHut7oecLPNCYSemHbYeNvkyYvmDZE
yN473axU7V+Xp0NxyRqtSAXgHgGqK3Iuyxk8nwf81iJRepnJCrOGrYKVCUaK0aYC
7WlQ7VLBERTZB4YwO5l0vlXxxxiZvJSNejqF5hTBzrXa6z4WtHNUfQO154A29Ddg
rzJEi0YWyFZtmSlLQ4G5uGrylexXXCydD+33zq7b7JdxWB82pYMQneSclvHD0vLf
T8xeC0TBzEnvoALNM/rWfAzbxjqEFobI5jIvmAZMuQ4LKcpxAkVE1za42O1hbp3x
x9jcWL1g0BCS5qd+6i/Vab+81U8FhBnyMbBUD6dABK45rt8ZPVI9x/I2TRdznGMl
oD2/ws3Qw/fLobHzt2raLu8v0bGm4TmltBcxcrya5q5WXmbPLfYol0LpGZSFBkmm
wjySm6U6ZToHlAw5l1JFWf5ELpqf1dOffhXzdvomvaR4gYW/cT1mYcx+aZOisvkD
vtRjat6DpGxGGssjl0tUrBiKccywgtgxybBRJM5PMZYgIkkHXQCejqrSIGYlzQW2
3dqliqKBqFrwAt2IJfjyDMoAp9M9Gtmn4JkuOB6A3ZUGWwuBqmnKOx8kve+Du7fa
v32Fi27RqqynP8w3jQv8+n6EvWbueQ+4k6pgxnV2U8118y3SWjSy+RE0eL4fkXoO
WERs+Mlr1ie0vCbHoC1Q+gdAyi0o1gifOwD6RXU0a/5yXWorY/WxdkxoN+i01ZBk
HAOqULz0COGgXMSHw8zd49qj9mrjKDI7ZQB4r/0PaVUuD1uJKnJy8I1BQKfTC0Pf
F1QZmFSFkUqwK+jIQNbuSTSoBJ9y/e5PPTZGvOGosMexoEC0ia6PR72l6h5xpnlJ
hT2Kh1SXSiLopgPtOWWuxYiE4z08iize2Jk9GbGpIpp8eVBpF1Ja44SZNJ4ped5V
4vx477Ogx3XuoJoltbu1HtLUZK3Sd9ge3x7dultayT5oETAp1JY2PJ8QuU8sje0S
NMTljVpDnQ59teG7nGp/d5hDoOH7FzqhQrDn9I5G79C2Gr/89QqdIVvPYJ6czGoU
CYoYornPZUgh2CogDtdqsfQrtGHObVIM1H41jl89GgVApYgTn1IXYbQz/3x9CugG
6ZgKOcCCEfs4+OAVIIoH7DX8xQPevcSNMc7G8lpEvo1ZWYZCsmkLVX1q4Z4a/fTr
0YhXmZy53VQJ53o+UBmcI/s315IcKs0tzxobtrtQKQBFnZURJ/Aa2iEKwXPsRpo7
aLWkW4VxqH0Gm3yrLm0AbSgKLcKD8SXWklI3IxuQsSI7mFmqPz17VlyyNJpClu62
uKXWQdwetJbClSlCos7uZGKYGv45FxCqKSIQhtZqKmfSIwYYg3w4lHdw93ySvah1
ExkTGiF8M21zXDNyELqPR5dqDGHw5ysoyVoHz985zZOR4dS/vrwTxUHY/PhMrKyr
DdcBs/bRIB5J/rB9h3Ao1fDdstsrKa4Yd84xs9VTZPHEAD88bc9Uuwq2RMac4cCX
vIiGFV50A4+I32b/LL6BE1m1+TsGBbqE35riLYmvqZIWguAyGz1DtSBk6kuLLHLd
B2QqiiEWTaLQNYJ0z9Q8yc8MkQkzlv2ELiAUfKgI9ZU0VhdwxU9jhl7zmtI/+RjI
C/Crt23Jfcic3k8Y6PlyiMAewM2+x5m+nej5MxpWcALpTqK2N/SSWIIT8xfW1CwX
ZQI/vRhrqr0IQxLvTd8XqfRe0/Ji8VZQiQf7/Quxaz8y5Z3GmAY+SwmP9otTxaI9
0szUcuxtueNHpWLufBYNJbyTOOhMNnmcOqHIoZlM/oI4ci1hmPLrPvW2npkWOLaS
72vSMEkdVwuo2pYWRmd5fbxK7hqKCQy1Eaba9sxuwu63GfZL43cELKLoWclr4m1P
GKmDPtSd3j4At2pneu3Z7CgGosQhZ4P6EiBjMt7pLPSkXm+qmysRxWerWyQ7pb7V
y4khlvh36QwpojysFb5gltZ80r1Q+PaPs4viG8KtdQjHOVdGL2o2owTssrMT03FX
mIBc6UqzDlL96ILv/vag3IzWIhdxhlwCknVTlJRwRglT0PX+TOyxdqcPWQ22eaXf
bLp0X8OXp0n/jXoVo/AVBSKUYAnG8EWGBJbhWT4vcc6QbNS7bJo/bqTXEG3VLcpz
EbeBABUChNOTUwYdPthRw5b0XVtw3lkr6QhjqMv7SjRRD5/AaMiAM5f0VdpeSp5u
iWWttF7hpWRJpgKYE4Dle+9BMsBoxsnlKBZPn5H2hiDLPSBd3Kb9OiTqP2RA2eH0
Sd3jMwkMyEO+k83rapMWnVFZanIKuX3Z4Bj1+DzU30mxLgMgwBv8UQRxO52WnMXk
W3GuWFA4xKmqn0Hei8f6dg17rW8hWkzBtCVYMFmZwL25Upaf+vDjJM491b8JP70h
04jvs1a92B3cTQ4/meuKTmTpqBFl/bNjfJU3eAHwcAgzmHSiY4fXFe/CK4HRVnx4
dfe+yDBYMOm91Wa5ANNVntxTrXJzWyceJSki+vYGhned2vGEFgkhhTV45xuki4Q8
aNXaeZPUEyRtB0CtX1jkAmTfM7t/2MhuE7EhE5t5vRWnnPZPRn+kMQosnyt4ZiqK
q1PTB4y8Jdj5C2JZdUsxhuAlCKSWXfBLrPN99lNk1os5+5lmzSVGr7yeswlc9ZXt
hO8gCdHvQya9MftPo91nuzMmvaqkyEkv4ihnqLqcATUrobqkoW5bPH58mlEGNoVd
PGXoJnc89Wlqo2SAG497A/bITHDmARlS/UFoEbc176eUHUE4+pv5Jrk4tk/Lzguo
UFCDQ1umhNhHfU0ZzHtO2cbTdU+e15brDcoUlzs7lm4LEFwY+MWQrvJlktc7kDAt
pjX1d/lu5/MA4d8qX/pBC3gKyR58x9bTEYES0rzdreKGagTxwAReRkCF3cn4jp7n
iWl4Pxt6OH+jbFoNxviahU8FQzRzmEV/3826IUe/vaYhzAW1BvbLIdAgJ/CGJrpX
BQsmufglrRE5g5Ib9KK6iwrxU9thhZ29rQYwkdtYMCAY2zBZNKbvFWIwOqEVCLEr
sseHgvT7DX5pkxo9iUxI9gHa9n65W7VIxVqZZ86Z2GnQDA2VyKAmYK2ZKJl2EFEF
THJ5DIBbEr2b76kIphq2ricjv7niQZ56epck42Zm1zw9TdH4nti/vj8c2Rybnu+h
pRsm16WddnXJ1FOSI4tifJZ/TEQCHKcjHJNHqJOJmVoSNSR0uAneHKEaz5DknPOs
UbTX4zFeP+2hj7qedsdbO0Hr1KoTyYmho4vdvPjfFsmRkutiTjtI7Q0+DbqRAKYh
SUwaVvuEX3cq1SYYtgriTU48Im6Yg4QQyVMYQhp53F+s3da/OTVB/5IME6MRfrCR
xiCLyI8Ltyzx46lKqqNitjXAVlBXJ8LkQazeLV07DGkYhABvYuSBpo1yL9P8y3MW
0l9MyUp3dKONRwWwjatqg2Oz/uMXFMLDmHAuXf3jzfRhBX119hTchHdhVOq1Sm36
a0KMKhTHOGwoOQIcuoTL6TnL1lUxBHMbfqBtcuxWbpTUi9DPzyBtHdwS1+aGsMZK
ao89xGFXQzLUzypXzUphP1nAkkG8y/lsMUZmPQ8ajJ9SBuILngMkNnIK/NcsvBIR
GlcdFM+OQnJBASbbG0+hkVFK9Id092pEta8Vw/o5fKqnP9Ci4+OtZ7qL0JFXcm/F
HPkj3o7YeSxw1y6TtXIk07DqqRRZFbLv0rVvBI7HcBr3ydv6v6vKdwHgE8yXAtdS
dLxZBqHPRON8gbU9DahBkMj0KeNv2FMIflolKnJShSGvnWdltn6pJls9gkof2F2B
D5BKIfEBOj1q0MdoMZTqIMV722S9R/XfNmy3JXeZ2Ghn4f4KqO7oFL3Xzu8CQuSC
5dzCJwkTB6gMvViKtAmu4ZDFcyBDmK+3na5qAmJVqN+8XlgbigP+vgB9nCOdL0uC
kA6khwMKXxrAehBjl+Ue9MQLk5T7ak3hbTpeYxwfm5KMl5ppnCL96x0qURwT5Nik
VdVrUMtn6PFLgDBKQaE31mGQvCgqr2EDgEfwUX321k2zotlV38F2CwrkD9annwsF
4OKiMwbXu3QoFM/m/8djjDGKlANnDODHkVmbQ2qusfcfCa23bt4Tw7nF8KM/x9qf
JaeRYKm5Xwk6MBJNho8nideT8gSV06TLjRRZBZrmfwC3gaG9SqK1AjIVMXyzCGup
/JeTX7fan9dTy6WWCtH1/uuKlXbYJV7lbv9qOW6NT3133W5gtRwo6tXEw4bCZnEt
mYW0UnogoxyVvDFhO2KxkNTXS8leGy2ZRU7SGb/9OcwskqsZEyg6WFXnHzDBsqmU
wHbIVN9kcd90YmdHazIBz/eqDpc+XIO2z3rEJoSNu+pqLHms2Z5F3dYHvxlJ7r7p
xKdo/b5tSJwLj8B/Rod6DR7Qge7R7zeasN9OHD3zlQ7AYWUVT+I5s3/Ye3DzVbaV
7Llf+tuJHOOLtnqxGDXsVdUd06jqJv4me1OXGh2X/654qPVS/9y+fKw50OOPa37A
WRewtNgMYUXZkr7TU5H3WKeVCZnl8goRwcXj2ja7be/m7aC/CsNPjGqE/PyqDYnt
p5yDCbp1EbtV7G4zBs0I0rs4Tir9vFBnFjun14lPpn60Jiw6fqJS9FJW+EWZ3laP
wcvXcunIP+a/S55YxTGdnCQwVgV8E5mDawB7Hc8BLeyyROZqgqKVdfBc+6twLZhj
HqP4/hEGK2cLvyXzbfq3sRqqH0RQ4b5nVGft/+wgNd/H81MRNAp3vwT7GM34aaWM
zDK4R3l7940S6zg6EYywacXR4VSs258NdxNwDBIFZi8hP4mVYLoBRMhdny2bOFdl
+uO2LzcpZ3eokpwWU9ytElydm7AQyr3h3Y1xunzj2//q0jDmuteX6EdSVDBjUUCg
7ZqjGJNdk+NEZ3vdjVKMMIC1btQLC4U6PkVXWAzwIHHwPHT7BHND8R1f4nu9z+sV
qYS/iKqf+7S0u9y8ORhW2DN8l5AuiNKq2vmzjGzTDTi/ubeOp+jVet5+sniT7yBj
KFwsoTeohMnbtVa9Td07eaqKM7vZcGARbmkYA2p3/AeS96znJXHhJM8r7pGP/guk
Au3M6MONGe60rmd0613+WsYOl75RODweP3Xd4XBYAh3u1cTinm8lv18jLhcSrSbM
OUuVnqsG6LdxXNfsiGXzGX0JDSGwpY00eqz1utJ9l1+xENEBoJ95+oFwlIKuvGHg
ZkVYkkFVmtuUDfAdePhz5Vrj7FExubP3njm1xwDk0geInm0aNHF5wmW5Rd0Q1BQp
CBnoKliVhzMBE4TvaY/Z2FCIpGE3CtEb9zeWyr4FJpjqMMUFw/obijXNBXgMUieA
EptLyXzTWVxq3vSekZ1c3IT1elRtP2gUSVI+cYws/22y81NPkHHHF3lxrEzU/6H7
B1kMPRQG2ie7m4LfnlU75eKgWkyy5PhjFPmJkrKOC/pofcC07XeL89PIC1wdaWcL
vJtJOO8kem5JbAX9pTd6NuNMlXQ26oZR2khlB6Yhi7rwFodVh3x5xO3M01VP+seG
JZkV0POUgso0RmgPvG3D7s+6ULSBbTcM/InZt97wTvBgD+Pd/K100jhlV/+RmD2i
CkRl69cFm1t4U6JHW/Lj18orB+hNa7mbL4yDgZEPzJ/3tGj51/e3yFWs/NA2UlXI
U5PCVkckMtOYldYkw7oyxJ6W9ID7GRU6X4mPElcilOEOcSFDkVsAbfkUCKrVE3wG
fByPr1CqtETZUw2s1UhnF/2rFMj092IQodgmagZRg+Y0AWoLJPg1Bk2FxYDctrzW
a+x4ooW1UoKqQpHuRfbX2xMiAqktb4jBBXBKQTGoOxJrnb7yUf9nROJDhHaDSYCF
df0lW10dndfiJU0fsvfzUd1v7xdfnZEob2/ujGaqtw+034+bLGnjs02QaUGY2oj8
ig8F7KdskCIJDCPbDqWt7pWeM7auFbOPdSiTnCxfEhSfOViWOthk2mfT5Y8qxdoy
LyGq+uP4U72si6Jyj3i5GsBBcoh3xq6xjVX+UU1/nqlBLfzUUe68nrIfErDNlSQc
v41l1a8sBKF71hMVD8j3qtjbTwLxvcYjKkjN6pFbJk2nYkyyPx7Z6/esvfJqhAFo
D+Hfgwr8ph1cl7jiRJrDB9FcVIEN4Nwkm6iFipPrPpVxNus4g6dNHzqui3H5a0ot
9BYwd2K+0ucTySKPwUpblf/fexXRIKjfKlN+UVyNknISvqwhCcTin6sBrKpzHBwS
CINcvB7RDxzoGKYNIkOHBHA7pMp4YTH1P9WJY6e4dh1XOW0bvxTmhkNZBTaimYtg
ky649FCwxUkNBpX/K7M/pOJP+1FCtBCRPyJgIuYiFaTkN/3uQtzZek2hnT6yNGMA

`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
H251HV8uch4PqNpHl9/dSvgs4jSE5iiXrENM2uhUgcY+HOvd2w+xqWpcZ0Q++MdD
kCBja/aG33cokYgO3/zibD6cHdTt0sTT8GqFwYw1M8MbgZvtXvBFP6n6qwqTnnYq
MFsCOtaNF0s/ZP9DbY2D3V3grauUtD1aXoimy4+Bv98/n5xEwgRYY3wypr8Rs2kN
5UIwnDtBiytOTqksai9cBFjwfzOkiLQLsQ38MmkjFu5+W+gK3/5MDRWRYT9RkAk1
AXWX4/gdi82G3QPjMO2/x6lJzCGcB5NU4gVttVx3Mr0exRQf2+J9iKPpYuEMpC+w
RZhOOs7eb7x+HpvMVzANrQ==
//pragma protect end_key_block
//pragma protect digest_block
EOPvNkewwB89sToE1MWHpuge5Vs=
//pragma protect end_digest_block
//pragma protect data_block
d+4dachOH9iPxgN65l8o+TnieyQd8Q+Uw9jnjYgRemIgOPF63/fBbEPisV8dkqBm
0aT7rrKI0RqGNcx2eRIwmtnnyNuJBciSVk0/+vDZ8geJhesrmITKdVTqksQvI8UE
/J0Tduc/4NJh9OtIfBY0VsbCJ/HyCmAOjsy4nAZfU00VA2dY01AtHyhS8YyNIMzK
WeJ2/yVbwqvD4bgwtNo57Jj6q7ouStewwYROZWE+UvoVrUysWcl31l8J87JhDThg
9OzuDKYA93X4iQRKZRCOovTniq9iPWBkT2xonOcF8zqDEGDa+fHFq7ZMDEa1hdo0
RIww2jf5S45c24TWu9cSrD+4XSjj52TQo2PoNKkPk89cOypnBPt7QK10LjQQ855d
DMxuE9XZqELDL0o7WR31M9au/9AEHR6H8ZvTQq1+Gxk/9EkYH8eSSfMGnihsjGWu
UjFoisLmnQ/bR2jHmjTjSDcAkoyWJkx2Acg52ST3Xm1X/ApexevbCaNPgSnRVwxD
qPm3oxv/iUFHO39EYz0EbDIsD/KYPNofusSFKsnVmKLhrexBo+31rahDqLywbGyf
3My3W7/ZOuJdMBSpgRqkHhV7FSrHBvzqgtImrEBMFfuvufWFbPsRPebbkKq/qvOy
27UxpBa6KS177ufoy0Qbx/zwnPo/1WBBtGNQy4VZiSo74pg/CTWpR8Ontz0EzMrR
6iWyQUGM8tCv5WsLJ4EmIL7cGbx/pPnGptUPVfmMM6BXyX/1Osf3j8F+24P3xsPs
zkhzXbXtHg3U/2Di3eU4VoEjWvZyYix9EEuzqQjTHuWcLCnmnRqZQihLem8lH1WA
eSFbches727BExB7gK1lK0qwjbLGGMlqfhDyvWoS9dizD+Kc53aFwGH4CH2XuHg0
nVC0srssjS4OACqzNibqwz1a7w9sL9q6umYWM2HYS4VmDguZJz/Y7iO5XmNItNF4
yCVpyGqz3qXPI9uRAs7eKydGsMg2sv/YIDoxsaWMRgwVsDNjr0BoQgnhF9hSVCRl
Ji6K4/Z7s5W0qzQGf7Oi968KkU6+65Q6HEFLGPclghxEI2091Bwtuu+kOZ/eG9D9
8Acz8mcdNAUBLgseNOo94mfoqjj6ey+Q/EUyxiKK4BKQrKdlVtO1kWgp/yc/Vw1z
YAhvRQjF0roHFvzktivyVOx1vHD2+DYEBkIaojS33PVlzi17sCN+6nTRv24NTa1f
qFa/GDYH/DE71DVSmqX3fgDgW0HDeYDY4Rr6DUTT2oD1ms2VzeAFPPmYR38Trs7o
8x0ogP6fnOTdyNh9Za4lULKL8lYxA74nC4wevC+TMKY3VXkt//7kOqM7KTPkiMQI
ZNe4ugcLsd4vGnmy93MIS43nbUluQr1MF1J+i4+yNqzEL5RbX9kGSOywV99A9ZUX
ajUyGJGBmm5IxaHszfXemotBjmTcXHropuyjxNp1ZjrFzupxcdEn9608nvNS/bV6
BhTzfL6WzecgImyurHpZ4/HFe6CuCHBWy8HRLCevXS+OEV7FGA14CyKHkBHEi1i2
/3IGdRvIjzM3bCMvmUQSwn9K02GigJNCgFzdguXSV6PjeKpcAM+NaC2bsv39KFN5
fzNnIUXzkzfAIVOEFjG7ohRUldO3iazHqKS1Z/Di6hk6AxBsSWUWZ9hv9eaoHIEG
gms9fwQEfnpKwarVE94DyXM01fbQoqO3EC0FYgo5ncJWOc5F7iGKpSHtC1J+lZ6G
L43UWLKPanGoRB7yVxzf3fvgsPWoc3fZ3XWBWiq+7vfOWJn1NpqMB2miBIxqSqwo
vT7E/b+X21qD2OToWmHyxgqISAqJnpUI/rJglwEnIka5yAEDnYAC1u1B7SmrO5eB
J1shIMbIslSsAtAhKbZTERNS/o/w3G/1FuTVJATaitcBNz4icopgt7dfVuUfINsJ
Ci+NTh0R+XZzwxe1dHAy9DysUqc6u8fjutSTDsfURmDO+9bQLM1xGwFgq6Vo+UeR
slH6CefVHwyTw9hEpwzpxAnvhGKQaqVOUb3xWLA5/Ir0gwR5YsCJ9voI9scXBFov
c0VWvK1K00KZh8PkxltTI/pb+e6+9kQeVqn6DFA13CVzQBq4PmXbbt+nDdRsYHVO
bgVJAWbS0THV8Ft2SIL4toVNW5YF35XyryUOfQhPGsuJxHmvxRLv32/GsMNN4POi
7D8WiFemoYGdDEfVQuNh/C4fPHIbbFZrolQVud4IKW9IJQ/aC7dnaVtbdxKFYPr5
zC9IqUGrO10A74Ur4gSJElUjXnLvrBkwMQO0YCCxoJfKrxM+v3FJD2Vik5EFHwS+
BWdKLOnT0sUyELMfxl+xsryS2QACkfeFo4XSCAYhUaBc8YpxckO7t7nxiU/kXGpm
WMlgrHu8NaOe7EUboc4O3PlN0qsyyh6R7aZWqamEk+CyQmDtPOi8AV1FdX1tiOkK
q7e8P1yITvzlQ879wxNG8BZpZGldw+79xIKkhy7q2cFcXLwT4n2CgkSDiKw6PzZM
51lFqBzfK2x7MmvtCA+H0UiX+tWF2E7D3RKfhuQ6MUGodGAUKEKeLmWXs0OxOo3I
JSWptMIQr+WDs2js7YcpmNFywU/pOaPingP2dhr0nYd3bD7oA8V9/kdwQ1ctDrwM
0PJ7+HrzqCCYHcYx9vV3/YfOtMXeQlHWcex4Ky9U0BxVs6xC1WyK41/hFgAF762K
TagGeXFZ1hWOFVDEYOmwnUHszinN0l7W4zUbKhlH6KIwHr+HQmCFL+awWD3v3LIB
UYUZ5VznHAu5Embf+ShK51eIes7OZbh9gmho+ivUkfjJgY8VMUxq0saIRDZEzTd3
VZuEUChVOYgWa9FNh9udeZNbEjC0X8dvS8cvI15sTEUeIBG3gIZu3W8vHJ9HaMHa
vrV+OHLvNnuB2RDX/wlFUZm/fDzK95cmuGfXgzGyQ+BDGufHW9+o60P9a03Om9dK
ud6lrDUFWLXnc9cilQlNR5Vhqf2+1Y5z0OrbFI4UQp4X/Lp+VuaaUK6H4FGm5EuI
H5iPsVWw61YWVqnYoBEunf9IK73rPQSogHVubJgE5p4RYCBSjYvf2OMSNarpP22d
eaJMeboPL2twyZgHp3CmKtgZ6vOxHruEZ+bWkGkU9npduWSZmTMJtv7VQFwgLgWJ
tk/qdB1ikZABXuiPtNc8xzBt81SdmbHwQq9oDHlcH/C5qaCmxOwTy5mjG0S9NPGq
q9zHtrC931KfVgmw95FRoq1ThuswOFYP9BelyuXMQhlFpO4ZQy6s/lpyidrUDl3M
YQ0qg6Xr5F6eB+TvYRFEqR6vJeeoEr4LvS1lZ+52LgZPnDRLJH9ON0KsKQj/8PxL
k5RNukTrSlOgwgsshDwUNqVxLpxlGO03ihMnMjcodpD+7ihAn2M9QZ06wmHGaqxF
BR0yQ1yCMW9NrhPiQKZ0pIDnUSIC5z5RU7fEoql/vfw+XjkVcbAFaI3ET6aKD2MW
dI0X5VWY2j+iCx6oDyB+Z8UrXn58AAJlkJ4YkhiKFt2UD0th0hOgmWh2CMF8ARnR
PXZbyI/xBvm9hZkEmDUidWzt+SBKwlS/y/FP+18l1ypbtl9j3+uYK5GGSFa5IvK/
fgdReRM+rgBplSpjF2koT/0wdXzgYWm9QFtI5bxvoTxdV1jNtGh5Rp9S4JZGFn4H
C6iP4ge4+85Ap48+PDT7pKx1wJsaB1Jovj71rB0OOfp+kSH22ETNpYlZAKTAyCp2
nHCtXi8GhwoYzFwj0+KELpsv8VQ0elYjj/38eg+IVT3azfszwpQt2pk8kyEr6Ooh
hENqJGabxpdUb5hYt7i7GXyFzNUwSRQYQ3t4gtSvcOA8mrjU2KSooAvhtP7EGcYr
7pl6NMr3NToDYVJawRWRe4bsTerHqc17R3if5CV2vF9TXINMu+4SbMpOPjlfCy9V
cnQ4tKEr1eMSd14zSSwvAtoF7R11ahCnmC3FYrqFXeP/CS5bwdTLQpB5fFEfhLTg
6Po4bi/c/9x/QAue9KYnV7zS2l1/RoxAs4BlFWAYoJIQ9S6oUFDcVC17O23RK0G4
x0SM5vzMC5eIdaMpbEvdrLW1cmSV0NO4rgTNV9zpWCUZ2CdX2NQhAh5Wp5kLaAjy
3UhYbsjPuohDQiRDDtyWOTHJvFkszwRrzYVOK+ibT+ikv6Q1Uspo2tOBqxTRWpph
bs3vZdAYsbzSPfZ2teaF3yUhVgSq780h7vMipIc6lxTcOyEovEyUOfnvc6pmnGxW
gRAEcjwraY+e6aNbA0qx6o3JjQzJAW7gql2EYjUFTETZIHn6iAnFL3o1DbY1uP4w
X8ALF2pzaRDfZQeXk/VQoG689lo+0kF1cYoJCcWXfQghLVeWMo94hUtPcatBeib6
/nsNdwuIYcalHp5uzMnYKNwcz/inb4SRo2jIYujeQgbI/FqFa2CGbzcvxWNDStQF
nkwhCcLGWaOFtrJzrs8t+27SbK9frYibwnokiUHZ7H2Wh5sQsXfQHvVFeC38fZva
8sepq7dn8+bkQzz965w2R9YLK2jRbxP2HNCp/yZkD7StdwL65P/WXuRTOEfu3KZn
7Hzy9UYSVCUfSay6IT2wPb69P3vKTwAUMCkdHP9kYrTpwPdOj5SaKImTWt7ZCuOl
oK9jdbp/DYQ+IXiAmtun4hpVoc/jqMYKcKs9Aoo+AVGY3s802yO3z/Vz6xn+YX6x
beoaA82IPXW5qAwMOCr1hcscvdomQD111cALFAE6jMVKun9Qs4wcOokQ8ESGDJHK
LHKlJokwQ4oZBq9yfGIS7XH4NOcz0kQ9eo/xN/Cp3aGK8zF+9OqIxOIrmx3qRHJ9
hFjsgTm0zpzlThlYkwgze2F4bYezaULuKmTmaSrHq8vaSaaNflgnSodfLEIsYyNM
o6F2y8xQvKsUAQN3F3r0OKcxoGCf5QyZwzxl3UPyRjDxbnO5gR7UDjXKLo8jkamx
0QXT5L45YetEu6X/AEbU7X2aMpMY1CqtmnQny1MHEEQhP6bwy5Ak4ybHc6JFGqLv
VXOGQ8iGbesaJa36LAb84Z5mReup0ckK11Z5/feJhPvazTSP6GNgfZq3MGHQ64oY
plRvNrccMdiRzkginTOJ8zuTnGJ78cXMw9BMSm1B0yZtc6pdh03xSWE0A8osdjaL
s0DTrZTYzCcm9pQmrmJDkq8VO33oZjyHnHgCHAGPKxhNyhw7dqzPpN+QyJhis5Eu
s4n522hSfNenCtMeWMimvIn1CStKiWDmIsSouHvJkOHfyW8Hzk/RAsQbSlNjaQ7j
i0RhRj8k4CzcyXLxbdmA2vbaRqgZoM3SQriz9dvPU96qUt980exwZ9wu2iLUvaLx
1cfAi5D4i/Kd5og3nlzCcLWwRUx9/bFk0tyl4mZPtR1poCQ4R8xOsBwbl7X1eKZ3
TyknmfLiq8cgjN2XZewi7yxKN2Id6pUFGtspSu/+ZLQdHuYgai1E8pAt6AuUaiSy
HaTKoDg+6wJ8oL/hXDNxRBWUTbEk9XleAahGdWi7XbSojmuKlR+LRJYH92PSVkkm
S2GCl1dn8xjhxWAdMfLmJFVvxXY6Op0wfHOd9fYgRRo/YIqVFpgfyEzTySKnrpNR
2/n+vV7RYaqKWhJAlw3u6kVvAjRlaNuMemExO5b13jmK3VYqNpC+/7L1uqLveTcZ
mO4eDRZIXVQp4Woep+k2jPNSMBGoLggr6vNkZ944O23A7E1yFpltX6EY+IfMlwiB
7gT1omzqG62197NUaTgrkE7lQIR2+TOSjgcZ5ATu/b7ORpf5xti6BD7Lw2DixkJ6
ku6YC8LpUrnT3qTn0+u6g9qVg0JztmXNY8pgp0myuuWI95MMIjlb0pE4mFGE0Wnz
NOckcCTlrzNCjcOa1G8tHtEMeophD8BTRoS+njvi+wwyCen6FE/SEfAKVZVoB7Zb
Z9bncA4FYCIdwjkFFKdKiFHZgcqFzU2/6VXd6ehZi94i4k3vR1Z630Lp6/bBt/vX
YuOKQfEpkC3jMel2l7NrJxdqgGTIHWKPk9LKBhD2SPuOHpxfNIrEXSdQs6jZ/zSo
zuaDWva93iqEaDbSpZJ5MMDl5RH3ytQJbNNplxf61ZlEewoAfUzxPdY/lT6eqaKD
QPA1soohvxmTKHmiBj8xczZRz9Yb8ETJGf9WhXaf5Y/fhvm7bW3ui5avM/JKZEXS
D6TXRI9n+spLHNVvjn43J2jfVUXIbQdD4YpZpE85KT9H1KYVsJvc+x5CErwtGyui
ascfwVuMTPVhUFNap23BSuPJKNVMNiVbLnRU6FTNAwFM2ZSg2P1yGr+rsigwJOAt
bHSnQWzyscGb/ziGETdVIeW2Qciq8EfPl9nPZheWkA47QsBhFs1DtBQBiYRprkuE
J7azsR28KV0XTKO8jLvegOD1c8N2NBa5vur4SPdMdoWTVeq2g8Vi22elWXt7u49J
LmyLkZbfXyFfKgg05WJt4PCTXmIuf1OhP/DXHYAz64H7dwmzpADy9D8U0tlp0rgV
4GYJ71DT4SZi0LJzuoSMKz37APacu2bCwIwrPljeVes69gftzbOJ1VQiHjkuEhzZ
SEuMFQ+ea6lXMtqmv+BNfNv79n1GMKlw773nB0Z6Pa7jGJkAgZsNWthdJri0a3wN
6XeXTCObDHZnpk0GipaOK3m6eNZS7oGyTUmK4BRj8HdL/QCgs+CsxODHmtqwbQ1u
zvZI4Lkp5blHZHynzcX/8duK3OkbiGkhJSj7Xe2S6PyWNfmG+5ZCc8Ed9e/mB9Gy
X7PLwOOqmF6+D9U0xs2pvPieARCFCtWmpfJhwW8SEySYDZHgS72BqI3oigJdz7qH
iEyvBZojXkfD0gGtkUh9reXeEFKChZEcuIqSXOWGjydbxYkBTo/hiWjg8ESaLxQx
YOt+qvyevXWa36G1tuqIxp+/Nz40saCJWt1JNZx/wxYzgAVG5+02NvB1CaaO6TTG
TZGn5+27e/w+qc58YI1ZdvzJkoh5P0kN0CI0MO6TKuiZ+d09bgyJl9zJKznsG2Jv
IKSjmx3WJ3Ml+Oi7jc1NwLUBrVwJvXTeqo52XaVlmWQXrHNQfEc0/l1xYuRBpHxO
IHGBMiwbLFHUrKLQiH40RiqufJF0TBpoLOeEH+zBIG5cc3gdiFThQjNWRXd/tetc
h8ThRldmC6dWLwPYY2Uet2I+/w7mYS9/eJPyT0qlA8HBSOzQRoRn+bcKGsNR6hbr
UlV9IBy99AvavU+u/p7yhsecI0SxCdXsGUEuyknMhr+t+Cx0xaUteRLb+7sEx0oL
CKc+0JF7vy+ZnbJEbnKBxU+hz6FlM3gym3ldCcmOULyE6YLkOLTISFzeEvmN2AVc
FQ+mm2qoE7GKzAmQ7MJz9Sow73LM+WjnWhRNpUrdFmj4W6g1OmxtzsRsvkdRml+S
eoAG+RL5jZKB7pMxhqDtu+R+1J4gv7pJT5GgxYatvRruEFqty8kWADRFrAe1eKEa
onYTI0jll5+N2W0/PDE24t4KlOtU5BwXHIlMcvsqMpJ3deQp7XXe7nUj+RygTMUj
vbFJNJHs7gsfe41FODDdPxNGZcmS8z1oSLS+h/gvhICMLaj3/ispsjpGGw4B2wuV
BjcRlhowweCtrvcczHxptZZrsYmFE3oPhbp3ISxiPWYBBLH3qAvhp4FnqelB5qNO
DfLMft02WmZU+tXo1DMlSq87iNrsa5HsX1ykQ4Bt/JXCdwy4CF4Sqn8+MTfG6OSf
HKWbnqFbgUTNvk1JfwZcmSH6RvtBzNBAAKVsGl3F9KF9ErsVvUrjV6s77OepUF8k
FD5zlnTXUwVp9aCPbQBs1VesKedOmclQf/Tlnk5On8eUwNC8Bxfm7K9lH2wwt48A
IfpntkyJcazFMBVq9BQBkWka2oHXd6YY8QvhhZWmlWtIqRYhQg88oRHNIsjbJAE/
PfrzKwYOOGpZLqhWcF2N5dQA5IY0vERXHNEwYKGS4ioQXrXiKA68tdv6o6GHDm1T
GoOVThwFmVKGdh/MCFCeluDWfwwf/MSNIgncelKqoPT7nftb0SD32VZTQk9Ne+Vr
HEQD2ln3DG01SN/HJqnq1Nj67nZlMoHFnFN5ZP+6hc1Si7uUjKcOCjEdG2jS4zHc
nk+9MMikrX/2sEg/KsXd3seOJVXWQPgTgyRvGBFqSnCK12iMF6NFGkQ9t5VcqNLK
LfXKXUCtjuE8dE+pWtysZnAE9LqL4Qo9dOs/9Z5SB08YfHci2m3CVkoDxAuS0ISI
FkrT1wA2OxOdB6RqpiNoI1OBhs6aZZKI/jr1s3vUVu3BuE38bWDuv9ceV8onhdNR
7vWP52Kr04SpHa9edPXPfxPeK1wycOO8+KFQkzrPQgPGNzlrHPHvu9R6BCtz//DI
cPa1UolaLtkndR+4I8QYL/LVdhfne5fpr5jDYgPi9cIrT7aM6gfLeP5M8njgZ3R9
NOG4TOUlz+QxiaJFLZEtCHD/4IYjNOFbsJ3UKTQ9hi9657S0ufXqjnmRERVIZcji
xyf5xwXy05wprCERe4SDEVdDgEq0V91irKapswyvjau986PHxrssXQaE75RFaXgI
FZAhE4GxCQRjGZMwXxmJf9a8ARqM101Yo6xRb2tzgC3LOG99bD5XdiVPXjqZdAva
XnJjOveiRNbK52IcVeyPPv/zOuglzEr/EiHHaQrtWAmnCnbTdNDBb0M4oiBjcc+p
qUA9vvJ+OWUsbYQ4F32lyifTpY2l5h5JUr3KbtOyaVna56a58QA0R2IuX93NdqQ1
OdC9h6Hh9eurxFocn7/etV/17nI4sF8fVPD+0Ld7htKIg7e5PoserCX/GwSwzIOd
3DMC8Ts2/bZF3PNgvtdbMvceV+ZbZhCnmlPBAATI4qvEQdpgtDl0c49KaUfAXtwq
Ui0W2SH/GEvmQ0mDFPQSfRUk6w5FnoYGKNquECFfViZOaeHv+wgDfD2Xbm2h3+YT
iB3okFg44N2NGecOh8CCqvvAbyVpU+nOJAtY8pgDYVoDp0Hg2MVmDXrldvWu0h78
VtCkOsRtWG7iOdAxHSgenK8KZQivLIoQerfksh+ODZvI434EXE1AeLD/509/uZoM
xHUFJWZ2ILeNUizYE8nwvkJ1rVjx8O/1Q0Wqx+c3Qtu/vgG29zYnqrpmno7sEy0V
0NggEhc6uY4BtdN5ar3Mb5OW71jrUz4q+cP+op/2qXilal9nZrDTFbqJ1bOKUxqs
eV7qEDpUGNhBkORZqo9GcxYrMzgelOxF1k9t3vyVzYKWNF4xVdVIgukXUVHoY602
B91FsoUqLT/Nm0O8Yft7Bk9oYbHuE3lkxKQRjJi5kY1ZMy2z0G1tAlPFqsvYO9lc
mYgifahHnKUD+6iZnxxShntA/XSTvmBJnbV0Fl9RIbZJXR0JyxwiTvNXCemzW6fR
pJZNSFSFjqRtosEItwhsJAy40Ets3epdFg8UuSP4Cg49CGn66oahILrYQYeNG1Sg
oWWqblVN+lcOatNT7bH0Rlp05oSyF55kvtOLTtMKHDn1vd/VA14BBDJQ/WU7zmYX
9mVuvh+cB9JloL165kLwme4Sn6PJyQFnGih5ij2OKhukhn8Cp1a6bn2tPpaJZ0ci
qZuwK86+rpavW5yBNVFTw1Nye7lu58d39T2jR4fGtRvujJLJ+7IFjF+rpsxcMgYb
EU9C09WGox9te+Tb8m+h07IvZVGfqDWw9AS63JXIWDnaqg1byHXViRpr5oRZ/QmQ
VMBrIdKkd79+t/ggQPOztVQFw+cxGNLqRy90jxDcPYC6GcoPQLpf7riI/RYei7wO
uAyr6/MEBRqQGrYI4CUnvY2Vv1VGbtsvBcUFUXES2EOb5/dlOQLMn21HKDaaALqa
NHLQxu7wUobtRXZDmvVSsi3BE3wrGYijnNy6S3eLioMu72WC/iFpGdm3MOQ7CUDy
p2Tcp0nO495UicWBYZ/1asxclzakROI6Sw3MIqqGVHTGNbqSzf4t00L7BhAmpZpf
EX4z+Wc09XGHYP9AyVjLC0G8nuMGivsmU5Fe4epvIuo45y8m2iXx9vJl9L8NLvyT
9f++/v0eYVhuk0bzHTMSVPfaNuJ38OjZTdutLl2iNstSL3EsJEjWBLMLaHd39EvA
67k8cKFIong+5IqpVEDJDgrJYIun0QbJti/NlKKS4k/dcOIlswbcgLT/uL+RcU70
SgtReMWxJxDtb9HdQjvsHWRpvP8TbztekOkGWGtm6gBN/5Hh8l896ftOvn7uW9bV
x3pmAyFFGRwSldG1al6ZVLSl4uoVUR8tzlFeTRbPA6woMb+pIcHos1Pe/tnw59ta
Ftri4A/d9y4nCNZtRyg3X66fC6/9kogBnenmjjV2tKyLWYCFq/YSnIJbVt38mfH8
Xoh+XrXHH221u6DzsqPOcha8Qoi0MrFQmstyCji8p23xj3MpoYxTCoxqoOOIbt3l
noozcs5aybRckkiUzGUrt2ooAsTduwMcjrs62iUyO4EcgfnhK6/og4vbVld4ELz4
jUm8DzfUFUwjlmtIHVBMDlLIdEFP5SEeWzUuC78jEiUdb4p171trRvikmn/4NREb
oTomEq7bG6f31MDuk7kSeVpQW3iqyt+Sd8Wp8Wp+AZw8XJofbE2yHQMsn7rQ8a7R
T+eiLNOThhbOxpU1l5kuFdSLAzCU+UXR6bMUGTNqg4N1RAx4snAUeECbXN7XbxWz
H2yVbIYN7ChrgyRXb/ElYYyZsaBo0QDfXn8r3U3nuJdUihFhJ39NQusMt4EkaKwZ
zr/eFg1TaDb7vITaZNexR4jDBBOrtwH5/7YiMaiorXAEVaw5jOdo3/AsDnk/XQGx
iqEiM4OIfxQxOeMXr8uLf6ffx0ybfHwHDxc+5/mZHdPeDoBOAFJK1ucLd2ajpLJZ
zVaxw7qdHmIT/humrSgGyd9bgouhLurk0YAQbrw2pk7ML1QfNAdE72D5nGUBnO38
w0C6EQfDR8uCjMBkvK+05FMA7RYoXbNHFyUfeMFBznOWKZDa3MI4Z7Tbbob5Z5Jz
FfU3dAsSzYQ8NiKrISvr9ixz5vKZLCl4l1kKVgg4Erq+BnUXltbp152TkbYFzxO1
O/EOps7vxOLMbSuITeCLc2Aed9Dv7x6APXdGIf0A8E6F4LCHeKOx9G8bhit+A8jL
LApgiFVrUPw4BFJyvYqKayYGk+bY4WRTbY2tEZjY4+DDy3nDZUp3HvThCKDFqfZ5
S2OwHaTiXSRAPztkFJj0+OcpObHRLJ16ZpK64Xn0F1SP6SPNWWobO7DBs8RsQXih
GNNlAcqRwOEcVY1kxIAIdz+4UquvDovGTQ7GnDK679pq94UMCT6Z+2njd5viDJ6n
PAmw01oLVJlnDKTHqFS/s9Q1AKc2M+wYk6GZPiq6grEAnpwEF4G/cYyhvGFX8sVu
z/Rg8IiQwVtHyLB2l56fyDZV81I/cplHROtQkN7GZfcdX7W1B3bCgIZNDX2nwuXs
sSJZe7WciYDzatoU/uthtYJQa7P28DnSxEXb2a1T0ySnked2mxyJOs+mft3jtXRI
/Yqcm1Xb0zyMPVprlAxlGHkuaMG2Nwvbn6tDSCza6rgEHNLqCw/GUWHGfGKAqVaE
LQc1AGLX2sjc8vqaAlpui0fWw9MiX1Nl6H8Ejpcn1CKx6yfTaI5Fwx64FXCzPvPY
7Hi3BDf1N83gEvtVkBQnjGePCbZcDPl3AiTDkVpxT2tbFZ9qrr28CbpE0bTak8q+
EASLYOtc26u7y1srfxxaca9agID33ik0Ji/5qirepiD3YY+CEcj76ShDC48v+N4R
1JsjVLq+5QaXJTkfBZOcPUp94xYLeOtSECkHkaL+P8fzLTp75VjzQmzgyIqwIxJ1
l6iTrHBqJx76t8IAJ38TCn+1LJrAUwIN4r5ldoIruNEuoa3Ja11Qa83evpdnGr3R
6TPW9Z4V+xHjq1CEXgIq6zBZbkBLMdwIQgG5wvaX/ij1XmVZtqO2VMPNIByDnS8T
Qxz5O4uPMhKBIYxrpwaDdtA0Pkw/YosYLdSPL3LI6J/GjOnzpDA9w/05XOgTCAMu
KOepK8K/lr0Nibe/LchRD83uBkuSFZE+FGI+C5iNCQeXMLjxUYMLNIueJccmx7Wk
d/ItGIL8tjSv6+4BPyea6k8Oeuq60lMSqDpb61+KCBNFz7owZeTFfSh5HKroz7gC
3nYrCLY3fGm3D1zhI76yfExzTHG4Q5hZ39a8pDYKImWGyMragzTxWPidw/kJGo39
1mLKvCQQUKD6P8zAhr2IcckgfLCir/ooNfTmNl5SoDKxdVaQ4Y62qUIKckHJMqJu
z+hA/dzqsQnZ3H26Lt9mcHi8BfRniFYDgLevhYBx9o4yHOwbNiuV+2FuiqaxWqwk
IP5JOAyUiULr1Fj0qCa3BQxqoCyk7Dun4B4a+xdKMQ5wEgGF7r51M3AYFVKRiBV+
k75w67ov/0lluMeU2jlWJtkuSKv29Wrh/h/AuwrEXFb8BCrVMVWrtAzgE6GxOVEc
zFsg4zJlVb79T322qvjEDS4dqou+Gxn+4DKsPUjiKl9uF33d+qVD6ukXQohcpP75
2tL+556hvkHEC8mN1sUro5b4PxEjrGkmwrojvpEgzuazuqeDtETKU/QteQtrdcbn
Su3SCaR09z9miEOvDDOXdLqk6IqQqtPB8dwpKXbm1lc=
//pragma protect end_data_block
//pragma protect digest_block
gFYJFHP5NhKwQyBhXf13FkIz4+M=
//pragma protect end_digest_block
//pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
E541wzsHPzWLs4i2rI+cIQ5/aA7FBeYXPqy8BWCb9eobm4fnvSVlqZN+DZogYKLk
G3DGaRTbV6R/7PgT+qBQNm2phANNC6Btc3uab02xQ4Ht4L1aHr8fuDtbf+kD887g
erbBjPgi/J54FwnOSQYNdjh9mpXFRxlhGw5Thcucxbg=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 3104 )
`pragma protect data_block
vV+dyD2VxazPjVsJxpeupOucGk1vn2Vqt99xY2HrydRB4d0DXUiWvzLOETNiIhVi
k47+CIG9/S5LmXSr5r4F+Jo5kJ487JJ1EJkSMHKqiNACtLHb4VFlZITp4kkfXn4L
B25MVFLKzJdpZ2ncLAhaOIFhrSr03t4U3K6ZSXUEMdGbyAPwT92OPx+t8iJAcdMX
xSJCrGSjdwvr7Rp9x9OnsvxeT/bgXsHKYqvzLKqAi3DtKVwtIU1Lw7SCA7mX3PKm
o5vPBGyKkueKHInmcbAyS+zPYLPmAZKg+5266+12CfE1y1rNPSYbCr+883faKQib
TF6E6dA1XyblLXsm4joV+QUUEIdFRGjC0kQ9VeurZGtNQYvpfdsPfj9GL2p21jtm
RVblpz8MPKhWGq39+fzx1oqErTx3xMEb1BmX3vtEbUsthAiK45kIn7Yvmsxg9oWg
2TtgruXdH6NVQppIeBmnOWlYK8HHQOtYbASLmEZReT/Airi7trJF3O+AklfYSL9B
DQtWou1h4SjuOQyNcscKUKhgSyno3Suaim9dBDsW9IbTe38wqBUkA2VLimtmegbo
nrZzNlu3peGauq75WNfhVHNyfqGoziBisQzvPdLY2FQw+Qmr42n4/Dw3f644Y6bu
CCtKzwGubz8ycsBceo5TEg4oVASH0OWpTDIaetG9M/vGYkHXAOAshvlrzuzpP8qA
MKxOK2Cy/BIN7q3LYeU1qkgWYZhS9rPiSPWwfRzySnFkLEv7E/syU211jTgtDlK8
VHp60cueuN7QNbDF2CLFOwWPlTDBjt66xS7fagrzhEQy4b7tP+OGe8kt8aCstbTT
8fM9yE9CWbOS64QNyClTU5V+pDM3UsDGTRuezXmWtJf0Hf8QET68V4d5H6gKrFuS
DIYa0E856rrvZrvfIH7pDZUuBlGLHjhiGfL4A2q7tp85vFnH/I+u7MnY+kFlOatQ
YsADYFgyXbkRXKGkj9F1iYOoZXBqH/p+1hsHby4juweh++UiW9PDDpwpzSXhGeAS
9NWhWqknVACnav1kWM7b19L0wB55VLqNUA0V+atNsdihrbwazyKkIH0xeykCqhLd
mr93jJzwJd+qXcGV57qcxM5NZ5m2ju/ilhmN4D8kVcM1N99w4UoBzoaSwEeOYIlo
c10yLD+64HzI28RaTaGvZmJri677lRMfLb4oX1UtvDiEGIQYlBcFOKq/s9ns+X8D
8FkYE5/UUGLjyLWsPN8vTrureAUfQfXUuG3kgv8penIGt9u/DPqeIygRQ5yYk0Ao
kBnrYlr5aeZ5v+R7SIAliaT/eFtB1E/CJBtg1MWq0Fzae/D+wyL0b1IEL5gYTiAB
owysJdatUNiCOtRXQYLsKbzAIp3K/Uqh1oZahH89nfudSUz5/rzqX8bFE7yz+BZF
OyjdLDPYGAfczm+X9JOnXy5YkCNWZs7ppPS2oDkhcFND60GnA/Y8ODcdlaqLi92W
LdOG0Whj8PU5t8eSablQrcw+ZL8ENWsxMHxe7b58jKXiRcWtUSmfzRfigFplWEcJ
w4SRQTln95rGV9TUOaHUU26PwZ07L2lKwyLkC+twe8F9Ci2AJX3PqCUoOyIyXUbR
9kEjB/3qUQO42RP+5M0dXlsCO66b/64xTwkBqH6PiHROg8RvccEg1NgPNtKYC3iM
ZCaJndwXj5XY7rMxaTxHf6Lo+V3DYKZSTMgN7Gg177jihI6Dr9/Bg4ulBknbx41d
ToUt4KP0nWv3gbOvQ5hCYsmf0k7um2ZrIAzBR4Av/kJyNw/dOSEqNh5nTFILxjGq
Wg5q2DahWjwZcnsuK2GgDkOovJVXgtWeXt3ghg/TFmoEnxvQZ/iuS0nU5/jZ/4Kk
j41oc3ozBRvDBniJwkyhRPY0jd1Cmtoqir/Wy/aGoV5Ccxcb05V4Qa+7/sTxYAEx
srpIM17gMnhAD68cNG1xKtPpAajCF1l3A49JyP4x2C1EiqkXbboNoLegOJ1e+dF2
19zj/RiowZFa6mWI6To9Vqzv0nMB/pHhEnWkEpFQGmGfgbF0lHY3pLIwiRkeU9q2
wZoDeHqsLdTx08HtaubTNno5ftR4GsS9R5lDuXJvrhWQVirImslaAC7Yjq9FXsR1
ZWUn3kWoxNuFsMq+4FsOfXS0cMVXF6BdscTHnrY66aJkBFHuKJYiSUr98vcfZtJK
Q6ABW6O9mEVoTSyar5fbv4jHRubY+q1ZyrF5YnQNq5r0sR/o1286JbU+EbGoOdmd
noYCMHnwYxvTVuRisKsGfPUVOH6SowQn624ichuBuXvpg/P3g2ReUl6LtBy/9jgm
+2Vpjoj4p24X0MYIfENz/wmYGyaDcrHewb99kwXjipfLK6ABf1vNHPiU8m64Fl95
GYB4MSBs/y/FKqWwVv82YA8tGG53a7h0DWT/p6Zo6ZN0EJwmQbFD85KKZth/W8qJ
uCBZCwS/rqhaCESwo0cSPq5hn962fHDkBjZfBBveRYihrU9LseWUiyMCU1q9Rzaq
O+22vc8B6hbqB3mCNqOPVwpiq3KddfH++HIU/a9fPif+/U/1GCRmffLQUmMSdPIV
N+RpibUHKBXK+bKFZxGkrL8roaW6y0XWpdynHXcBOxnGzDhfTb1Riehh+9TBrohL
3LLd3kwDj43HKeJAS2bKyYQsmNESQpIkS4avR+E6kiZviY+eERdNIW8GcHBdxl//
0QHpiSFE0+TCOThj52uiStS+JsAObEoH13osvt4v1/NQS/QJ5e1O5TI5XuiAwifk
4zpZAVVLTigECKEz3nklc82Ast8cpN/+i5dDAJ+nj0pMsIXLC1zLbk6VoMm46tbk
EeoqPIHsSTAWtwoZ4A3lnWBMW8MDoPBSzYFbKQSXDltTnIybKYzTEV594l2nbXiB
pZyU/P/dCePKyz3JrbGZI9UV4SET/ISX/0QNapaammxRGL67HKnrKvHXEcDQcZpf
sAsFWDV1NS6UIDIGHBvEu9AALGdFzS8fM2i3hFItYvV/dfmcLvKwLKMyiYuLZYz2
U3NBIes9WFFMbQXOEw8RfwUsW/owMP23X0AIZ2eBXldFSaPigCIKMBKWUAuriP6D
zEQ6NGMlTqbKczNrc93wrTnwlJUo9gTcXiYCDb2eEUjZvbBCWXlwYUUJ/xKo2Zzs
m8yRd0AlbEmuyyIJytXg2ZHt6cEHH6+WS0xU1pXRbzQyvsRHNV8bRuPdOvTa4CFN
rggPDgkURamXM2sePJ/T3/+kgbYSGIOzVCf3yNRKvSG+vZZjyFM6i7GcYuaX196o
3BSfwdmS/eEBXR8fnBVSJ0auVqUHGTn06m13lFMI/W2MIpW3/fJjGuhvPKHS00Sj
zRrpsmUOaBMmEd17nKxRX/HfgnkeDTF9J4Q+3tM3RZS1kjbbd3/R89rG3wJ8aiDw
kyjTC/TEFwYFcMoTop5Og38AjKZhkpdqbO8lEkyumBjeXVaknlBOmuCTyr/5e4Kh
L1FHD8KdwyhuBRD2w8S5IU8TX2V5tfi2GMBcYtS6IRdEOYqYS26ZD/5oKtbnmhvk
GQitY7njqNr6F9R4LH396rLTdxIklv7dxWe0K6fvjCPebNGEBzN3Q5EJudBGwFds
5BeiUV5iBIjmYogxTWCfzv3YV+4nGNaYfaifPovt+p8g2uw2W1qIV3+goSCvk2Pc
Im0OgO/TUYxZLo9upqVUwvK6NmtWJg4cqKW40DHT5A4CY/1bUxmSFTUIHM9joo5s
WDiOHXdlx5zkFbH+L1mq+4MCmZTf6HP4DhZ+JvxPYwzIgDXif+sPjd+ks6siGLMF
EfANgJj/f9tvt0D4swoQGI8Cji7rL4vTOpYkqpPFa14DuDfPB81bp7SRZ+/YHv2c
aTWjzINV3awuPXHIiFGAuMG3kro1cEENlgaa83OGe4Dv+QuenRPP69Bl2RXpP2be
I+WS74IfnmAIKEXKF+zzaFfJMzf2yMZm0fwRZr8O2BKYdhlvKj3KfBU5tyRC1yGg
l+YBm1uaIq9Esi5W2CJE2Z4rEc8Dq8x/BCZoENT/5ZqXkrkqEl/4QqMMkoWdIkeT
Ajhnp0NkgFvakvApYg8if8PwupXQFWgtOUwvgJlabWAF0DtIi93Vk5ozVRoI88BL
shVj2iiLuFz2qkdFMWmf1X9yfneGupM5mMNInwnnbm0=

`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
uxkWU+DgZb53fq6KgPmG2pmZadEj6rT0NBb6OqYi/MoVz0sZnp6a45405gtlT334
5z20TXic6aRowPj0ng/OPNfFpPzVhD9OerTQe356D08VwBkzlOjBVcjGD1Hn+dCn
AF7rFXOZCvYBmeEY//SzMvcd6k3uTdCDTas1eErRGeo=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 22096 )
`pragma protect data_block
XyTKBl4EFsmJ/L5M4BbXXu3OGsNaZqs/TYQRMdxoVGoQJuKw/UiUMYgWtzaNlUPv
r/Mo9BkXFJe9tgVmplEgF3e24h1kbBOWZoB5nKd+6EtyHPSBG7cQxYD+9+cnaECi
O/eGgde4ielU3UziA8G62BCdAQYGigkADyOT4+oFOTpqdllr4zGsSWA/geNXU73r
KgOHTFDUMLV33y4ud2QYvJNwSXL8osKxTEJEc7SWKYI+R0YfAp/8Ytigu0TbEHIc
9mD9BepHgKvBusd+xKZdBmnE7aAh+c/3d9vRqJB2ARdxR8TAuAWybTSOSvaj4/ih
F0tQpjkI7F14utXS3REI1+O73nb68TIkkg+dJOdA0EPEa25N8TWmBDNRLCoaqYWX
GboxmhfYD6hm5n/RRMIIdFHtiOzBlPDxjH0m1ENC8ZXJRIfTW/DcXklZWs7HyT/J
sIdRaYSLckJFplxUyjXb+9azJKi0XcE37hWhhAujA70VOnUnqh5lI6/9ylVKRFPH
ckytz1Tch+1nhKjfVLJz1rxpGe+P85AP9mnxT8q6/nVIYyZbU3I7WBHLdhty+O6k
oht2B/vY73U3hI5GjA8ZvnaAH+66VgdKtcInfsOT7sSPP/GB05D0IvkNS6RmwifL
gyDW6i59cEB3G3y2qMbPWmKl8Pz003+M6oDPTfXBy0VDtfFQlxrbL6kwTfwBs/MD
ns50mZfQMn8hz6Mz07PxuBhDGemEUEc2f8oB0v0oo46EovnPhkivyGGDFrCxbxje
HV8QwXSVd8E+fibCR1PQBaRkK5WbLA9dGis9Y4xxdIrTN2wKNKeGopiy8Gz0VC7Y
MZiDEIwERwULHnoi3gM5GUw64oH8fRqgJpjSJhOS5kOR+gzyDPsfjmqBbzH+iPbp
FpbN3KpQXWvK0c8clYAc7GECgKYMzmIqQQNeIxIK87lBb6ujd/7+HDBU0X7mlab5
kcFfmBFZxDGUsLasaaN8FJiR3fZz/UrmJQ/GxDedCV1ofz6FUvihd0iSTOFYHrTz
egHIuJdAj/t1r15DqjmMa9F0IVoydW47SYWKUw1ezNmMmrMxUnNfOBm33RYUMhbb
v6f3e4DFfsRpei2U5xgrVm+jY6tSidAgIbDLk7BmI0GV4+ptzEC401Sx0zWuGtbt
JBmMcw3jNwUq1d6MestVVTOBkQcV9Vcdyo+GcCE3S/fjh0uUVBZ2/MxdDW20N5gq
A5lqvP4kK4aOmSqQv1oVHL+x7u/6ZffQzVm0cif1mzfyXpa4WXo1MRAuqpax9kpx
Ah1yWVufpc+u4yLyReDMIsEFlyxPgLWqLOkSdW5EMcA0qgSL2VVV0EbIUoguOhiD
JnVwz45K5/134MIbwyIpDTOTwiAZSOLkcckZXNqzpDjixtaUVjwjLk44SrcYF6Jb
CHSkTo4+58DMxuS2ImDcxpYfK+HOiqNKG5bH8IMUxlIrSTR4/5TPwU7KnNRhvOCV
Fq7XyHpinuyWYL4Gp02mw3zP+Q7qwlpbteFXsIc2JBP+yWZi90VlElCFm0b72oU8
s0Los6nTGZcENm7W19QfIaN6XjFc3FkNnvDmN3m0AmgtJkzjzfJQtpSDU9SgJ6tO
yuegW7Rw+907E/Sqe4oyOkMwxL48yoZCthK7a4r9P2UvEiACn3u8l7WpAICQ37bG
hTpc9HNQLjsCZOAgK++eAfud3JBTtT70R1i9BApubiMCb62bud+5sD+ut4wVdpIo
4GR2E1GXARGICrOoslnq9MlSMeb1rxfJTLUV6zeW4TRLsQ0T34fwyH6PeN6MPev4
jkLdDgeMCZvjX1+i7XOa8+Qkwkv4pB573oMfJu5o6tuFKSyEMMbmtW4n6eHoTBcF
mJ1GKTOT82xMImgXplz/7GEXNiIqk++xNEW0PtzGUUiE3+6VefNijVO+mc150uc9
yVmmUalrkkNlhdn+NajrtvHYzEOWDn3QjOR2bTHF0Z/x7Yh+iVMqb0TKNe0r6yyD
duM9Jof3u7jqTtU5pfe0rITG297zjmPayBxyamf9Bi1ElGLW8RFDlnSfYaFrY2bf
VgjVxEeoZ6XYLXNROzlIEbQFdyc7FkWh7WEQ9Fb2tJI9GxIM4Urx5SihyBlhZsgh
0WnzGx8IOiGKdxSl3MU/W7WG7+9sAbWt0odQucTtgeZZkXxJ2aoh+lrjAjlciK63
JFA4N02y6VMXKmL3MSG7kAWiyCSC762TKMTS/Dg875PNZgHjKs3dkkpi2AYLuY3F
saTiR4gBYno1qJUhz1coHq27s1Dq0XHT1qDpus9BiqbBICzb0xB+fKQZ+HKJyn26
ezIgad/IA3mB+weuQ3rc4EDAxUIn0L6qPwgVl64ZBmSYmqEvBEwwZ4yVPEifZrfe
bTw2AkBwz3WiA6UUNDl6etE6xOUXPo2Vn5bCa+SG+2ZSx9WPEnb2RNK1+fNw6iq7
Tti5U6Q/UPH6Kdf+v/aHqG+dT5OLXZIQckSaapGawJlAkC7YskY0zLYcni0pHD6V
ZpBcqMPxXG417HSIYqTvGeWm2DXbua473loucf8UK/3W7bqq/LdZ31udacyKa9YT
00jN2S4H+NAeSFiqGXXJPyYT/c/i/c5ZhW/1hzUy1O/dPUtP7SoAPxrHp2YYDWsn
qdZmV/53z8yoNY4fFQBydLBXriXjOeclKxT3hezc+WHEaJfyVofpEODQZ/Tv27Ui
ZeLIi1dSl75n/kutOkyn14NUDRkCRR7MCp2zv7Z8fp88dFkSxsUQLz9HrFaUOr+/
2LmzXzZc1u/ehdP4djzy3/+b1B3ol8FO1jJHAwXPztIxeh9PdHcDsRSGRf0xwI/B
7P1sSAqOVgdN7r57mAWpoaKWhuIErdUg8Ft+w9McuMYojx1FFKIQLt7OI8RonmJW
QzgW6JuxUcl8VSc4pgh4ThUXb9Wmv42g480KQNWM/jwmiHmK3F1zKPtDyHL7CPKG
RoRxwCqYE6XrmDHcT/mgizH6z2KwO7zaT0eKh/YlDQVAwCd6YYbYLaBtTKIP99LI
LOn8ZfI5e5EcbJDDyYl2k/xT31hUvHYhSbBZ9Dl6kapldC+zNNRLo2fBezA2qL46
P/pvSwB1fPgj/3oGt3yTbNII/DeKKHaNf6dFsAZn8ZBhnOaq0s9LMN4hqjU70y/D
38/WuTWBCmls6yKzOP+fDQuSHyLkYoPb5n7S6RXnqAOMGHS8QnVMLp2SdrPIkboE
VyQTuJKMwpGrhBxzG3XGu0fFww83CS1eRxa2teG/JCF2D26VEivgaG4Ye2GSoc4O
qFMwEdEPE5A5Cd0Fwn2+N/8sVi8efI3Dz8jkG+gJIIWtWH45EKQ072LoG19ERrY5
YZPjgC2yrVcgAObRl1Q3Kfq3PaQqoTgdy5yimw80e3J52JjXi5bzWIw6WHxaMV+L
m2IRsxPmKQk4H+36YkAh+rq9yOos0hk347PdPS03cQ0FgDts0BuTyxXB22MBIQUr
sMqsK6ZbH2KPjc7YaF+Mj701ZD5Rbt7rsxXkbPy1mYf0H3dSBH1VMBeNWGBciJPJ
Irrx1ZvH4honl3cNTPQTMvSk3hQHKV3NoftqYS8HS7PkDcVqqKEhL+IrMoQSyND1
avk5Cz7IRBODCdXPW9S9iq11mA1vqrIavcZJI0A0jzcQZAn76UPMB5RkOes713GF
d8mpmJiOdANYlIPHR9Nh7DwXPGBDJEOBGLCRHCj5NzHJoE/22BjRsiXHHxFJQVBV
VbTXmkLlRFsr+tR2936XI6GFzZabVAISpKuzP2ZahWE424zEilQPy3Jn0n1FmwJ6
9KyHkeaRppwKfAVVgqmuZ76cuTOXu/zVwySvv4sWxTvHzwFyX1T1X9iCE7sn27X6
XScV6sdfA2rT2q3x6WY6pn5Tax84259m9paVQHQK6lfcqgnpakXcSulRo429qynb
Iw1ZK4KYREOxiGHYVV7N0KH8S4s5fKyJvFopzM3EVQ4xakSXtcyqNn3043PddaaK
p9QXK+8WLS7bZgFczQ+qVZ9m/it331O10Kg6zZtJ7YbH3HIZJ1Ovp5zVIi9RTZrR
d03PX+Oe5vWth32Seps7RNdsc2A8y49gvzAvLEjRmWM9DoUTKE7OCFu6aCdORl/G
QPkCUtwFpPBy5f7UeHpeFbrMjlqAyScC+lwWmlIyi4xIEunZxAEwKGYCZq00CgxZ
2eHoF5FomXehORdHiK0HCNjGMuxnEoLZN8Ioe0fwUfdF0/G2w/8tkf+DBizlwcI4
T4e+PnR4c/rSIEYulhqbIr2uTPcCO6tNuDWxK/9WUhZHJ4FRkyOTr5ChJ14fhxch
yc//dlJxi/jnS20iRM2k1XVT2R0K80qmEVe1Tk5tyWvwDZMHx/p/0sg4tPERaDSP
lawkW1qpmLYDnU5CxrU56rQRY1MqBKrVu3ki2zQxGzgHFFZu81jbRDraTgp5sB9d
0a2ZWDPRNzAcGfl4HICSl5BySQSbwaQPGbd8DFeG3P39TkZMf6V7WYMcA0uZUT5S
HcOKuMtH1GkYqyEp9uQs4z2tePLJ33PHVIynUIGMWmCirUu+rSa020nZmowBK1lW
wnu6facOuYrrBosBHgK6fHDaa0PsodzkHLNtAJDlivk4wkux5Y0jy3ZlcLJBsdCt
BYOGgfPhVUQdlpQpon0glD9qvCIM38pLf+keDfWsnKJgBeUBcgDf5yE4s/U1SfTr
C9/64wz0zSQGC3KMUfGNx/duFJmayOoBBCac1pObGXBYrkkR6NycuLrWgwez1cmZ
6U2Toz4Qdr1c3cuOEJ58KRGRIusIG5TrCKxayuPvFOjq5xy/kdlr/v2xylso3jAQ
t+pzGqKm2lBkwfoYppx1XaPclaPE+DC+wcfTqPbq9vnB9YquEsHeOR64UXNsYo4B
YisP0yZ+d2McEd5aTIvONcqCMrQyyc58w/aemDzds8TIscQP7mTkYsAB7Ukt9Dgx
3rcuFIDGxB4XYX7C3xdDIcXdiHNxPza/58oNYf0jotdRm/aLBLklR2fxX8rm3WdE
MsldsyL26JeobvIBbX51YcjT0ih/8sVmxFN7V8ifrvoTfIiVKNiJQ8Bd/NzOeJON
0tUOT9l/wkwHCDTIMw+o+d+/cU+m7pWW5cs34Qumacq2t82iDcGMEOOE5vBeVKpj
AhXwnsMELzrN4RExkmpUyaNQFBwgPoVXWT8XqpZgLoi6RG5eK/8O7+z5yPl9ZnTC
BrelWzGn5dRuhAS1+F3u0L7f5C0SqFuI32PgBqbwR70WDXKFSdQ5w8Jo4kvsRdWH
A9mAQVbldn28brig/MzUvG+tn1/UMEa4pipLuFKniamJv5+TlTYlYHJZfg6e2Zvj
ZxGCCrVvFXCjNMhTS/qlzzKFplBvhG5rLPcZXtYBJDgYnqKql4PaCdJDwg+5f3rL
EFpLVbxwCFD9C5zRnsDlFigrneCYI85mq2AJYKkjilsA5myTkAFP2PfsVIxe7mUD
srmHK7KKRMJDhW8LecGlHgSLiqDTHosnIvB4QWbChwJilgVBB8IHw1sm9zKxQxCG
C44hC3EokvW4hFcSPsM+cMkZBtMzh+fFWExBYtiIeC8iYhnMV6iPtjxgYARh5kvO
0wiN0DFRnLehtyP5mZbGEW7Jl+qbqMlTudVT3gyoO5VHvDVv/hLztRQo7WKXLGNT
MqTSz+xIDHcQ9SHF49bZF49NQmCVrhqvDeXZ1LLFjFP1PI5yH+rIHjqpJuQpFfRB
an3qbLHOqLBbeH/qjrhh6lwnB9ihrgP+c/0L1q0/eojsMtIr7e1+xpcOtvkz1Th2
fe0Mtr4eOxkIVdn7a0kJOfoUcIEHY8S6HFLAbmxYzGIQjmTP/UiD3zXLNvsdEy6m
DF6xxXYOlNb/l1gMsvFX0nsUkX1NVsqCwRXW/2Th9v81CH5AC34MmWM1eNPd1NZc
c1YNK1efE46mNxWiAc5G4T80BIJW+WFUVOmox7ZtcvH46WiP4f70fRtLn+Z86IY1
6Dxg2HWQ44R1MLG8D8Xw2Ui/zxaIM3VRCBE45r5YRL3X0dOFyoCvNEoIViU0LyCK
b2w/TCtfp6GklIICK/fXzCRIuO1BYoEZhSuKuUp5ov/ue0vCJUFTKvEMKLUDFEnB
NA9H1nXG5R4CTBppXSV1BPjAvzp4qk0Va6JXSABjQCeQywqblKzGJA3ClohmDzGa
tqaDjj/arPHPH+fqP5i/gzicrK4BslCHrNOeYvhg3LaJQ19VV15pv+YJE1oe9cf+
MMXn4BUyrw+8G29z19z71OiwldlGlv9yYkbB/HzhId05C5xAx/xSKrEoT6P/nKsf
eQ+iHQiYFtYyfE0ONZQj14HNuHYt5tRDhpstndb97AiROIvSQFo9NGFS6CPSsHoq
w1EaJiPwwJNlngu5OXipFMOBlQ7sgvup5oQFeoQMNwSTgSBLa9doCokMyHo3Dv8Y
OFKuxSCk9SszorbBui+d2zuCFeIqJsQBmqkXpYg1m+Rl8IXj/ZFUTvQg/6siP+nG
IoFePfdeqyXg7LN4JVWjKm6/C5SekySo8qhFd8eI0UK5MLRQqcAI8HuXq6lmfSXD
C78mFXX8XA5JXzGOSTwyGz+MkWdDi/mvWc55SGKWAO2D0yU0f+pAtfadcOLha5vR
dJVZMNaA9U0UMR1t2v7Ns1LDI6mGQyUNcs/7RzDf4pXUFp3nyTD+ygmb3wXIxtW7
0EHyCV16U42WjA44z6vECqU39qZjg79ldkvtWlDsqfpF/FAlZxbjB6Cm4QclPFoJ
yp6SgK8+DJPvVPCvfYPVxVf+HueUgMQZ6VCjRl9iEFyJX+wTA/Tq64P/PwMpY7dn
/uGWkx2JPyBzwqtyUA0nT2Q2EF3XS6VNlGdlIf+mojATecQoek9y1eFoxnAQgAVT
O5i7lz9/6rjdM++kC71sIVzobxJJ3hgkH7hWTVcHtaePPEVaH7bncGv8+tpsxTVd
FVEV9G3SrZFK49EoD4VW2F3JnIej/K3v7v8NjL8vxLiN/djBtigLx/l9FA5kUata
M1PtCgIcHAY8ThtRuLQ8x9ySBDAvH9/b6a4c3PV1ytt8wMrVxnk1LSdZ1CMAu4Ey
3YRVeRNQE07bOwGVtXpw634L32I98YHCbT9NMGBK9ug5VdpoCeu61aVIRL/zJY2f
DmCXCCR3Sssd5cCirtklF6vzNLgc381jboijExjjW+Q25pyWpTjktHqhC+gig5o+
7Enq/nqcwFhhqNByTnjYBwZPuYkNaW1jygXAAdrd7KNYTxX2KgjCbyzMJVYa61vj
fTBocKzXjEGfq0UCquiFfkcHd1JKfnP4nk4X9XfvlBp0W0Uds0r3t0A7zmehhWNj
f7IU4sYot2dlFpe1rWVt1OwKqCSjXk+2uZeDfiLC+bTBozOhctMYsf++MKQPgi0o
A1tFgpIxewmiWOV2llw3cyGFX7wN5ITSjhbR+iIvFQhv92DeSm6BH/7KZO26jMG+
HnOJeMISuBqH3Wa/uNJeFykf/eI1dMxWrIgRlCcM6ZO0DcF/gn1fOyjsxHHoJJ5b
u/GNvxN8VmEIdcCRa36vrEEzViQ4MCPL5tmbYk0HHa9dwcEFQqnyczgkE8N7ajQJ
aACaLHU2qX7o2DnLTK73B6SHw6yiyMpeDOlhBtii0ITl1hinaHbENxcjjNjUogKq
S1HbgVUZqtaprWSTJcdBb2fOJsEhDam+/iV0mjmwTpq8Qv+YmhV17k4P6ZCQkD8W
ZI2mCCTG1saz8rVB7WGyiBguIAHU9FrVP4aAdv5CTG1iqasg9l5tjtq8fPit3ZKT
ceMiMt17E4lbILB65Cg4NeTaCNyxSTkkzueirj4Di3dm5IxQ07MuolBfQiHowXbI
ClOL2bSSrxMeWjUyHcUa5xuUx7L7mtjfIR1TcMb3zVfEDecp9AedXJk3HGVXIPsk
j8TqEsh9puKNGdWp5Jl6h+Qe30Muf412kHeIsRhL0x0ifxCqixM1GH8+lXll0cCX
nFjDGu2yya40psyUofXeEWjrdxBOZdth59PWSCHczbQEdbSKOwsMl7UfMzTmNWXG
3bkVL25IbpTiJ299VOFoFCvHpLTSj2FMnl0WB4Bpfc10BJRQMUrMZiSV9xGE/fVg
vl26ndY44+LxvoHWCBEWpw3bALMGFGG9ghhWq1+8+0IGwyLiVYCPRXK5IS+bidkb
InNq9Io4GvH+FGD0ueH1ZIotsQ7Q6z0AzVK608aU3xbByijyz4kE1VvbxdmMhBvg
IkaqQvUoZ3kucgcaD/seWGJEH6HALazQ3ueLYmbONdoqFBoqi0zvK/pIVtUd3/wd
ZoxPSXODdHY+FPZkqZ0Gfh9NR+d82PuCuVI3Y+Xzry/JkvCVwtx2OkdrxFnGzc/n
yiRi25+OoQbHNIslPFuYa8RC3kBnR8ri19Cmz2lNZR9Xe7k7AZZLkixA3MaZOcon
CvKf719F02DJ1DhMtbY4LDqbx08OEBNOB+qppvCalppbjA7poXeUAubDTBHtZ2vd
PgGPSPuIbL2OqXicCCKX8h/IumZbtrswnQvWvigzsQrp9M1pNq3n21XoOTaUMzgq
/m2UIx11Zvuhnlu7VWmn8LtY5geqR/wAMzpd2deCWg8qUtfMWVETMfT7SWY1m3IR
awZFn6b32lTsgix71cY3efzArbvpDKAEiZ8smCFFNq0fvFvgw5Fp065YSjG7q8gr
1sAbaf48hC7vsuWoKh7H97D4ZQUearb3pBCbwAKYytrSHqhtx+4vWCzEoa9UzuVw
yeCCrlc/Joj4grDxnqINmDQ5EzceVXyvubUzEHY1wwSCrYgKrvcWM3wPZsT9DVCU
l1Kn7l2L/tDC8v2YvWYZDIR5+q2PrQ2HSdRBect6WT6qTX66IRWK/awJ1qiI2aeZ
Q1HPCc7IUVuBunFGoW2jtRTqdf8m26c5A2q/gRcMvdvnw/7UkpsHGxvISJQf5S7s
iPHNEAP/GlMwnqYTlLDDDoOWh5ya9HM2lCwclNlOp9240HAEhH5SnCUqlkgZ//oj
tR2eTAhO/z8amzpEcPKJ+W47n8B0BhnUBMD959iTokano/8akBCMSKjVEliBhaD4
p9SwprY7PI604LgtDiL54bTEL9defhl0COHSQg8gWt2wAAvCIfOk3nF6JSZFfcw7
ulgOEPpOrXCF/AG5cEUYRbPvOQv3Eyy/2rjhL7gxM9sG9Quz59qhpGw+hIUtDO/O
tjQIEIru5Yfu8EzhKb93Aj1P1BnTyQCRQerHo1PnMTnK73w/LL3EmbmPmdlWZM5G
CGXUMvwdR0/AJFQH93J6WZ+mCD/tuLAWLCt2Bvi/12/xYDmfKzpUR7nV1L/gSqjt
ZSmdz0HIGLw/YHlKG87Tan0PcNMI7M4ETXNHJPumYdPb3UTQme82mce83V+OmZs9
91HwPkAQRL79iEfNxJ/1b05CiWm9RjycFduMw6lbaCcIDpDyuQOfXacHSjxnV/cg
hZE5cFT1284pQbHm5Itdub6P9EGkPvwPaPEEPJZGIhlODmcCb9WGTXyPaywLhxA0
sQ5D64SR2JiRMRugOCLCGNsAiBlKRsdvBFm92RT/frdAWQxq9HuGVpo3IhAhIrK+
+Xuma3W6d1uAEDBTS+0zgmhykwFYTbuisS3nQZRZouv1X/JEYQLB+/PP7frP8V0f
QeYKjto3A40tjO3KEietdJXZr1r/DGZ8nuV9NmjX7CB+fbv0r6KBCoQZAh5ZGcLf
+6AqBRYPjpxOk/KGcDVdKFgNaiaIlGVd3dDTPrh7HvhjaQ1v4iKeO9UnkDoVR7Y9
+bj8eCplzv+rxNmZYykNW99SiQJ3gWI7PFXFw8xlDlO8KoPB4J/Wv+zqSzqPxBg6
SjrzFxt1gYS8Zpc1D6TSf+3oVOll3zXUOqIRSmfAz0+T9UTopTiP++qMpesndApW
1ro3UqzHqSatnsSH1BY5Ttm1T+VfNt/Lm5C0nQulboFC7ak7GZm9f+aK81KpqXhI
mctbtK2TUFJeFiBOY1IW0mtGppxGxB9LF66Gh1vsHG32tjV0VHUhRJpR9snERaaU
udAKFvvB7jnLEOnw5/eIyflGj/ougrPh2l9oMq4X69obc096wI1ejgiKA87b8qVE
xHphIzVkfBKxdZ6KDUpGB7ZwVxxt2J7AGwdDcarmePdNdJZIHrBiTDE3OBvoDS+J
z0pduuoMnSAjrER3KrOS8w2msAqs53wM7VUCjDya4HcgMsDnl7kWl4+XISNMSRtF
qvq1EuOCV+DdKpSBHgTg1jeVSy4CNXBVSDDHlopj6EHXyekS3CIE2/j3aV0pfRy9
p/XuvcDY6VFUW5F+DW2M1pJxNaSTduUylOwcWUXOQmAlGtQXJPyUQ0FzyXSwq2Gs
rpk+PO2MLAVNFSkL3QM+T52787GrqCxukKjvAuSCpV2Mhn6oWcB4+Wfs+m5S2qTf
lK700WDaatxgsqA7USDVv6IC8yT8eCcsH0AssRxGlx4/+nUmcrJj/oXVcgSAbqhO
GV5Oe2nuQ5UrcZESogBn64jKypQf6dJUUCnHxi8r+LkjyEtNSfL+ujLXQzqE1K1P
aLxLm2dJmnedbzT5KCq4ld9K2udxeoq+UH59aWhSXWcLZV6JXklJVl4qajZ+smQF
kYsvkDImjcTYcYn1LKVOuudXBHjI+IsKaKighCZfgXCek8kD19Fb1FG9/Og720mT
WQQfybiih/cP3kx1rSyFx2fPUSeLNLR9gNFk86bodnF4FNUvlXJAJg81f/8sX6Xn
W2uoW6rIbBjdE6U/irQP9s/8Olsxcu7IVP3yG78paUo6R9hnNGxTlEg5s7MmFqVd
3vn98LhcAUq2g/fP6cA4VcecmyjKHls7CvtfoU8ojLQEt+wvvFyK4PKQELbiEGNn
iLgi+f07YUvdsaR2dM/efXiCI7NmMPnbX7Nq1yJUyvli82HtaTH0M+zS/DddauhR
Aiu+v4WaRmEaLgR7TlWeu+s97Cw3MZ9GWZkqvyJ9Lol62RaT5sZDDwo6g0WObcbt
/wy7yo/HP+3IG3aK3ZOdwYPuxwvZYLwb0KpPNaMZ5raLm3D5qUQQ+uTpE9p4CH1f
8I0/jNCyiEe+s1MqEuVSxuM81UBp8oHd2wQfIjAs4x8D0iIZvYphQdUarN1AJnVw
n1HK7dgPldonbmDJNR4mn0D9wFe9j5FVTRbJxV6YYGqBZdXr57oGLMgFKsIu6GcL
393X+/YsczUbHB2ShZHFbPgydBiqzmvEh6TGEYZhDjw+ouh3vqdmJWlA/sRayZuQ
LcoAP7JMf+nZ2MMGguxkCkPIo2r0VASpKr5w9hG8Oi3gaTN54OuBFBmbUyr2wnBb
wLrbc5rVEoLp5B8jOaoknNY1zSGMZIN/JsFfSMlAC5TsFS5hjhgjDrwpzAv4zNfj
1Nlm7RgtMsH6hAOuVkkS7Ycuv3kFzXDMuZCP/jrYOBvBHR/DJq8G5d899+i0zUug
UE+PoEq2BVuTvkf4Kjgf0HMN1p6JoaSCzN7Vd8iI6ERUe3Ew4kPns3wP0CDt2Dl1
qgeljBxJwMh2nZGy/jNzhhiy6pJxMHrheQfgQ4xnjgsxHxyiW2vrFkPfm8r+79YU
SWZajYXsfXu+svDaRxVkJI5h7eQYK8XltTlnxSGAi7BO0nuQKHm3B3iVPI8IUiak
qN7PnTKvMlbtmFckkD3zpwQiaxDaDncoZJdiBixuBO2O7MxZkNjtWq1DQRl1xoS3
ZhJfX3rBSA+MilqJAfxtTucZ78VVh7BlwslOSdlNjDw6vp7T5dQIo5OZDRyjI5e+
4WVgQt2BkP4KB/UXYvn+WvjkuGZte5rxSWNn69nBY5+UZpegl1DKGA2LxpCRq5pX
ZopmR5WXQD2i2cJoROeooJnJyAUcwCQF5XXeuKTQ48lF7zpyS0fmqbEaM5kwLV1k
UOeiLUO0W6jMmggSq3VGBYsvq2CEAxGHQqT/BFLscJ1aMPNBGC4nXhuutczS9p0M
96aRt8NWiWaMzqPT3o9n3/h39IBkYrjgf/aOrx4w9/N1FZ35ryrfHle7zTtoiGKA
GwcMakczjjwPvf+ipVWWRxeXo4MYlWZHBSNcPnLJ0pE2fCelr2QqoigHSuGDLx0A
bL8EP7c4MqkfgUfa1PECJcjrjhWp+1RZeewjMjetffqdziAnVRbdMIGCUTTk0nIW
C0pj7+MxWiVi1G4R6VrNDwwOE1w/Z+5dz+wzQypXP1OMX5JBGy7TW7sN2CLCQA3P
JqJsOripqYKfzMuLJP7Tx8f7l75hqke97LpbJG0R8HDqPM3shj1QC8WxyVUbXXMS
1aKVZfbw1D6skF2O2BFXvb6Aydvt/sDi1p3PND8mWkfrwc1YEmFltWONXoBFjSyZ
hvl6X/HP2WXVJBAtoxuZix5w7PElbMfOKzZBzY3EQNJGeq8IqPAOnYdcqdg+8Qro
COwNI/oa3Kx/oT+bBGbhxo//vnaDaVjiZTgX4qDWTCy5+YkcaBlepEGLC3G8gKYc
C6iK144GQNDK0MlFhttTm6LVIC5cY3dYrz6moqKTrm0/Nc3Vdc73AdQM/44x3qpV
ypXwV0rOkESfN7boQmCReYrnRZSxW2GivHSfLxxrI/ulir7yhzttqJn+/kmg/HtR
RWbF1LnfruNJZ0MYyqoqJ+yJ8P+9jTADYS2UsrTUS/9BX9thnQtdWDkqxrtBAcyc
f6lRKwbGywXsAcQ+00RMeE2miSVarS6a4+0M4L4EdXDM7Yb9UmrzZqUTGRMH0aJx
L075Pp3wBQ/KkFntaBBgenfJZeXYalkL75Dn05An7n/LR5Nu79+WfWgP5pwgjV7R
YebQy31YR8qbTiHsHEp9ZKjRsr/bcr2OB3dPGASJUJXiqCQC/NVn3Os/Y00TJQbW
bdDlveD24PGDxhLkcoNN0j5SdccdjUj1rL/FhKGi/IOwDtESmtHr0EXRBEsdl6Ve
f52aihWIBIUUAxQ4hdVKEugpunYf4t55pmsqvMeGqgt7dWlMdyC4sRIv+jrro/P4
7AZwyh05CdzrM1fi/YcryEzoMT4eFfDlJEEJSlFd6W6LAGvGYlJOUpJEef0gEMgz
3W9js6/IC1P+Oct6UQr0MQa6YRTU5FhS9DUMcf0VPVkMqe9C84EGEw5S+hPyyt1y
cn/BjG6UR9Ae622BfnuSE0VdBEJlxjAy4mSz4vmblI74+/MUR9lBIypqsCTHn64q
X0NfHkW7c/X+ZnUQE8VW0kNcrmDOmyI9x7IpIIh6VWArxOVbQoLDcJELLl/QlPIT
7FvNm0Ls9CIqHN76RSFNFYsFfLpNV/xKwCk0/mWfX1biycERvzuhA85WdWAtIKez
ceUvL+aS6L7iBImhDZZe5cQ4S75XOPWJIZi2JjqEH+KeF74aKBtNGO5LChzHjc2M
5SIQqmncf8S12cugKkn4APRWMxuMX9bHWgBGN3n9/4D3AvpRp3D4j1nq8vfPrIgv
Su7IGGr6E++YucEsER8rH+CHEBVNbQGXQ9t/sYXoRuFkbysoaV2am3sAhJAXj6xo
9p+sNsIXc6UFgjh32/hTsVgBLRsHtqow5bzhgmH59adgfeKcGQRjEHlfBw3QXQNG
Z1wwvRDl5PE+PISa6IGnYOakz88dwLvrErsqfD7bnBnPhHx4SewBAzuW0rNCJQgO
4NeVhFfx2swpdHLg8kD2l1k8LAn9hopolKN680BwkDxBgLJhxTSZ76nm24cXpd28
HxWuScwS1Z5FY9BGviJZh9Y9/Of4M9x7+ZnxzVHH3GQzVHG1FkDnpr17VkWB3evx
ws/me2ES3v4ObOLXzliNAwg02H2aztAEGOUXUPzIzd7tTlZUvQ/9YtkM2PxCyq01
1ixj8+2dJeBDDYvRjUIJdJU+G6fIYO+khbXBM1b/osAbV7mt6zFwbBIP1ICxlY2i
ZwMP/XDjV+aeTwQjrmaMjF2KG15keJwkkT2pOS80mn8Mpp+BFmXiGe+lc78Kf1wX
D4H0fln3X9Zp9Nwubz4RXns63Ib2Em/9kEocVTO28KX0Ff6VyjYOu61SK75Talx7
IWeB/yFPMfi5hu0F2oCmn1WEcBWgaJxADty/K6Ubx6M+oYSgeR5vOKdI1XezmrmX
DDrxn7S/20tESZsyyFXYcifINNWROBoyYP8cdztCLY/ihA2XXB0Govxo8EcCVisQ
/QdLY0fBrCngBvd6nIxMfpZRVGWUQf4WpiqfSODcxNkMi515jgGIxr9ihx3dGZf7
Rh48Izd1k01P2dVhE97eu6rYkU6rcQieBbq12EALuUA91yXIjTopGY2TopC8oK9A
mnM/dVUlFMvRDpJf8GCVITzAkfNdqWxBEYnqdZtrCpbVKMUMU/l+v2Q2B9PCk36p
wTU6KLUlIhAkImX5NrrIrENj2lhK2omLQWnLYqpmqiE596N7A3tGPkKECD/klz0e
wJQAJ/WKV6A9BY+ORkTMSCSx95C+HrzGcxvc+hCttE2OqZVnRILJad/I24Ozq13j
5JFGkC1H86emLv+nEtL0CCbJCqMDQTnYYkHtmy497BA3kDp+Li4PJa16YWTrkKP6
aK7q3ddSunLukmJI2WD95qS1vx5WfjZA4tPSQDQxag2f7OpveAh7NFy3Ix6Smvp8
ZRtmHU7NTJlWpQ16GBK4d8nLj/PtDqTN6QOUWHCsJFRR8l9O0KyB+5MfpTA4Jr/a
6pT3FryTqclk+UWl+lkShH5BaZ4T/OVCmRaoLzFq26fsOYB6hO+w+hwVoGCtUHZF
WaxdYi9BlPgKjmnLMBA0pDH2/MWRANptB9EBsUcR1ANRs0ZQl0iz7ydvXiu74bX6
xvzmWWAUNb+OXN5SwfaF9zkMN6yONG4pIPsXfRzcDSjeBjhZym9C/to2wg9zgB0L
YSTWv2Fm/eNQB8u3umRfJaXXiw2QEiqFjYH2yhjBH11XPTwlqHQT5u41aeVWj7xS
7DGVVeeWwn9R9nWhyHvEwPvaDuWd4Fq08mBL3RDY3w+lOFVVwKG6QDRcvNwlbpKc
MTNiYcA5H45LPl0jTWuJ/FYLVtpvQQ+mRTwm34kkPRwNb3b3l9mQktqe8N0+a+mz
DSlXzZ/COKKWAnJchoHw/vYNkqsIIPpTjvdOdLXLNNAxez/oGN+QIsPLLCIo3K58
MxBIHE+DuRaBvn7IMaa0a2R9mj5ILb4Tnf+waPwWA7hoeNvlTBNcgyh1E5Thmfgi
SzuzOyYBGTcyl4dQSZVbKHzXu1mkXnbZLT7lNFuI1qgMW4oqu1OESXsIOC2LZZ0k
Dg5sMdzRN8GFv2g9u9/C5JS3I8xPifw8OF55B/c04q8gPNM4omS1F5ixPBw9WdHr
rplqVbcHC+M5xhLrLcL79OV10a1sTTyIYsAYDNZxJwxNBAGPfdqwAbgSPDDQK0Oz
rvYp7GWlUR6GaITR2peTVrCP50usE5Vtjtv75Y3YxQkpcreTRKSWT+3hOfyjWaYW
GpStPK+8bT/+Y8G1/VZ7pcWUupJU2iXLN1NnDj37fOm62Q5ay3SvVKQTrOjyS6zB
7RYp0TIa7A2HG2R6nMJC8y1TJSMZUroYduoZYZwNTqZzhcUtgJB6LYj+o8dNqnND
XF49LJBxl2ZuzTDycNiEClUW4Cv6tXW99fFnzDcygf6FbvSM9W2QcdiNIdQ01e5Z
SgBanCA+WeBXitwp/Bm/8pEcLWHutVw/k3JYYmmvuWpqzzPz8H1k1c0Hpp2iDAlx
ihwdjcS2/+LZNqXbakgqnZ+1y0PwKLEQNb3xcZaYrZAwYCgC4DEPDRXDSLzUIiwy
EzDDgni56KcATOgQr2ipEGfPyY1fcoqNLJ+BKYzh9S5WqcTNGDGMX4FCwxC8eC8b
H+wHaWi3cDpuVdMdBeqvAT6s9tI2pbFigYgcLLPM48uxUnRGYZ837OooxfJiVMm5
8WC1aGADn5wIlEct80dc0oaZtQ6RbUIR+MTFuWK5XAPgEVqnT36veaySZ7yjBlzI
fevPuWek4NHL1317qNghiM7AkKzAw3VktJadqdv8HI4wTZcAF5pQpe/Wlb0smKif
MDBJGtX15ia94YMYdRkNA4SKTJTozkCJKpKmrY5HDF/stRHiD7Paj3G7KJAH9MCu
rDgnv8kxXGAdKnGYwadk9X6VWaXvE13rtzbdnMzAlCsBc2EDgQyvIS6Ye61PdMew
WuTHQ9EJCOK2tsbs1lAdFZpRHvd4bh9raMG8wz2eKEiLRukWemEAEbUC5awM3cn5
kAGoB76hBrLjBEGakKwNnZXC0W1k970TnjdJ6lbM9YUbbQT/Oi34P7z0xq7RyG3m
SWA6XDWvGHFwx/4byhRWoqtlHUm5JE1tteV/3ANu4vA1WQkLBZfg2Au3gP8dZtRS
be9vcobYNkTIg1IQ7VAtL4FRSOIEnVbXwLtaD44adA8FDQmAfzg6UdVEWZCYy2O4
Zw6EFTwJ9ubXHEyFEL3T+f99dIJy/NjaObLxFSnAonCILhU1v3stINnOYfmGmbBn
1wL9IENEpvXlMJPxDGkwTeEZ/ReSuM7O0n+MKxNPyijpqLIpUJRCExP5TLweVTV+
6xnLX1hte78OUs6VOFdTXsdZcuu3bjt6X1t7Bs/jr4kRd5kUXhmhX0DXyYE8Qfh/
tIxFoyZwAM0p1EBvSltiFpLsBZ3RGFnxp7Pf1qRVIvdXLc40iQpf39mrRxDWeXv3
Ort+dgC5jewd/KljhBhBqEiflmpSROCEjwf0/drThwhOcCb9lPPn7/o9a1J3l9nd
G7hnwsi416kCaPfWIaYuVjQAAQl7O0aiitXkDQ9SS3jaEI006ZAh5OIf76vZ6yPN
U1wMbNf9N23bm1UFvcxD6DnEAXTBamuMxWwSLFi713CIw0zeyzI3bPTir8hVPPRc
qhlWPKKW0XwfqvrmjD/zK3bNwLSQnLDbO4pHfnRnRkV977aRoEeOdBAGkeZmtbYJ
WF7w5YwnXTGOpPTaehV4d3nZgjlGtbQXL5aUe6XEp8w01oCTcdBrGEN5E/Y/4EkM
GaNmvsiBY3dkvA2HdDgvIFEbv0KN4iSHfgr09nfreOabLg9fWqFbo7vJNEmlIgwl
jSecXxio9spz/5MY3nsslYW1LTNt3ECH222fPp7MJG7QGYHHYQbDCwHibBPWV7rG
9aVFuw4ENY/nzwI6qYXso7eHfzcuSZWeEMNvX2xHHFCSMk3XNp733kfKmAQBtsZC
P/kIOclwH005PXqBMevvtKBu66RZEoVX//i5rRgBHoU40Gy/oPhmzE7Fi6ZhO6R8
5d2ZULFeyFS0NxuMaMTjEagg/fMAI2vR/vTo5ySOH2fSuLpvuy3fhQbe4TF+QVAt
4yXRA2jIMIuqm8DE1MsjP87bCaSxivxNUW939f1yEO/gkEYYlO7zjEELr++O+FlG
hhFIQyDDuBe/U96n4F5XBfEGNbuicim4+Fj8It/4JjISK4PXmxEwdqAqVaXQBn5s
UoOzRr/oN9DVuqSwjmFXmsK0M1qkkLNYZ2d8knYJjdVRpfKY44SPgAijiMuPqJmU
d1bpd68TnO/Jx7194I3HiMu8rVunytgX55gpmsrk1OWbVyefeUgdgPRhNSrBA/Rd
94lKwoTNxBzeOLEcpjcUKkd4nP06uMCOa9fRjqvzeAYwre7QUtRiyXUW8G/GKnw8
WD9R4gc46F/hnMOihvFn87tIlqmTVllJpS2YvcNq64CNTdhqQ1piZahqh6RcxMMq
K1eHwwknFbQk9keLAoSMfVVQJBHcVFbiRrZUQCxOde3qy7fNQPA8bE3iU9SpW/Gh
bDwkl+RZbv8HlzGJ13Q0eeWtzIQHkF/10hjgjzJrXe3ppon40BqA/GUMJhlwvvV7
p6ED63weB1FfT58k2kIcM9TlWP5RmY8PNSJZPME58/C8HbF2nnnjVwjjw2bJUWXE
ALo3huMrIrz5zMbGRhd1eSy6xQnYrX5vCXse2QRFjZ7GE63/YRAzgfYz2GWVWGVr
DGQln4hcYH6aFta6+HGG1W2bHcnvLTgiK6IMHytdCrJTIdHf8LBMmNYpQNwZ7UlT
ER6cst8Ij/M3lAofH8WSC/+HrnM01rZBKgpo+MvSOiGjgfgHQfT/yd1Y+Gp7RsrZ
A1G4fIguD9RoOg01/a8QxljcxKyGCV2LpLfwESem0WY/TM8IFLaNKMKSg6gx25J2
YnF/LQT3HtY7vLRxuH+FE7g6L7UsVLryxlmiWQ6SihEu+IxnKQ8sLupULtBXiqM8
ruv+tw9g5lW6CUfxZEqRR8GyYazKHYU2nmjxbUEvpw2cwICKovZ5k4qNsd7rJ72O
phFDkgrPF7KF/KelLI51j0PO897q4tsJLWm12RMMYUjudFGYIBf+sl2TyNZPwDTP
e8z5Pyp4gwzNvdWfh8wFj2xQXO/nCW01BvEiGMUN0xZ9cQcVyQ90uiQRQcd6PY3f
UQIQ3lnAsqG7nkPgTHhv42wakGqZkOcQ2aCbKooe8NCE4EOoNVQTiCnr9RpirGAg
t35ut7Z9PFim7VykfL6piCIqm/cK4dfVelkij2tnNCweszrQnTP1mEHY3aAiGyZB
eKEwPHqUD9Sv+UFMAJVQNpVGhV+XPOon2CLHsJ6lRo69EtKFulFkJTVM6Sq+s+tB
YRJSRbtptTRCWZc0NuBAuG0amdLMzehnwu+RzAY5+43C0zFTHCbydqZsmmsmceCu
58jFPQzwgHtdjFT0+AE9ef6lSQqrw26G6vXTNwVU4NhBVNKTcHpmkRBLVIa/q4hK
UEC2JV0CeRh1bT9rRe2hDh8UAQHnxPsksdVT8lZf5XjwrjdKEkm3A4rwVtrxAGyj
WfBuBuVPleCf9U4x3vYiHq/+9CQMdMjVcSH6/iLBnEJ8u7Xvb7r+INYasXhOB0Ta
bQS5fcavNScXNSCTMppcfPFB/NcOR3nVFu8ELVnucjbYiHmucYdrsaCVNwiwWTXm
UM8CnLVoFZWd/gp2a2E1L3rp094wFHiKfJ+93YYhwuGPdSOe+ccIRFRpwQexNq77
eb6h4Bt7YaM1HGE5kyZlBdAfAbKEyiZ75U7pbPe6PtxkT//C6dfK3JDl1A5aPOX1
g5d6PvNJ+16guLGlEUx1vMENz4v2ZSzLTc8S0nTeQsU0kZPiv8o3iBkZDJzjLvgg
09VZHbJZXkmkBno+8aYM9yo0z+epagdQuB3F14D2ipyPONu1RXlUZ9oMR4fl9E91
U78fEpzCG0ALOlYV2dJlTdznFNmhDErU1KqTyamPbVqqknkZXMMYZsTKSGxUTHIO
TON20H8tMLh1Mb35TRXsbUCQrp5zgN29L2+SMKtyqjFeY9nIc60I4LCbyTKyrG+l
XaHzT3vwZkcOo2/5TTHcrFHZXWk43zek0Bu5kaUZiSaoc4/UuD55SEkEOf1MuebW
KA6V6gXCH/JNxqbLr+7zzR9bEaapAns9v8w7PiV/KNPDILFqcbRIXQlBGIw9GIMv
gpXkHHykCd1LiTH+xkLyllKZTYnb02mi8N+PXHk5oxKH5Wi0Vpz49Fpk17h6dmoC
i4dZqD4yAHaoVTvtGEHShYFVFtFFrRuiy9r2UZDtP7dpJl4/MsXMLhH2+fSK/h6+
APDJ2f+z23CUbnuGNd2z2Zs3qIQD/zHvfD+TMyaWYv8rgA5+o+k5wusmkedDRhhw
jPoNIrhBwXjPhwU2K7hDoynxyut5o5PFgWM7J7miPSE09bhJjb3omxs7b6T6Rlop
3+93kdtusGX3ib45znB06WNpserrQLxKMJ9mi9i4i0PXm3qx1u83CM5NBxOg9HvV
RinqTfYUiz4bL9aa5gHhzo2FHxxRJfwKcwVRq16/VWBC1HtxaLS6jyN+Lsn70Kvd
im+XJ1vAlYZ1BPtJJJCqZXAsB45X2Q2nVa1jX//0crE8oW4172mcL4fjM0pdvl4n
Vsz9C3psW6oVNNHYD9zWBkUYwKv2GxfjGdtsfRhl9m001v2nUMl0Ee4sN4u6cw/S
5nvKYdwUzmfPXEjUnXYWl98NbCNTxUXYRkdRLIGgrzN2BXNkywMdD3pUqeuc0u+e
CDwzarBvw6VLmn2UXdvlCJqZ043L/hS7oxGrN3G4+iPt2m2JNI6C2lVu7lRZ85pO
YWn7mL9QVc26CAumIe8kUz3iV9Gatuu3vGinPBf/6I0XdNBf5LXkWKByYdPjveMl
+E6HRmR+YZ+ZZQK29gg61r2Yc0VH5ij1QN/OCoLpyfaZkULnZ6LOwoD3H0s5Dqdt
8qXMPo4HNkMhbvJmNDTeWzpAd7ZQ/AEv8pGNynlkX4SQu68ILcohFwWKXb7W4YXA
CNhx0AksMlkLZLxapg/cbxNMzzUyW7ixPSkSJl99mY7vSqnnfZDE1CVPtupi/0e0
vfy6ukc7juLzhWJ+3xYxxkZrADIJ2FLVUBy8jzE8ngzFutxxxaqFrKr91J3/30f0
wouV9ijSS2iaSSmqPpeY9mGzZsE+aCeltC37pXXnlA2tl/ZVxnevDI3TTv+8H/3Y
EDxeN/60XXKH5ZzdmRK5GRjp8Xo3C5WG+yDKhNVouxflDkhc4kZoQQGfISLa28Xf
plSw0cA62+iehGHC0TcBSvFFbzxDdUmeyxc3t5CHmNffjkoQsfia9rTX8EVBrgXp
1HpXR4K/JSL+WcYXlVd+zDe+45CHmBb5lnlE8yeXjfASu7gZTpnUfBj9wKxhzwPo
78/0N3ZtvLJDaJs2wIe/rlfzPpM2fRYzqyJRTN2y1YcrQMpPe1aBRq2ZzOruN/3J
yVji8RF+rAcAm0zbtybY5sQjyx0BHOZitpryiZHuZJFa0UIhfZdii/69DQDZDlob
G8pQG3Nis3eFygO+LUPK4d57rrAx2iqKInjrdHhoxQBClCbMp/0SWZOCvL5czOoV
JCT0dYwTFgO4cZJ4lUixiGTD3PBR35repJyzWy1Q89TllNreIUF3PAD5ieX2GRm4
y4AAQBLhKYeodmqt7fZcW8ZNTHwnUQ05D0Lu9m0gyUgYmO1bBmKTTuROg+3RU5+Y
ZFUF+Kv13SQYtSJXtEGV2hGBqqaWZVB7xU+IXXIoCM8OeMOHFUYjD6IdIPXPHDiZ
74uY8g/Ykvn58Qd+x6vJQ3UuJmXIPPYSjS1AxNTXypSZChocgBG+hnMpwXrKGVug
jlgp5KtNC+q6KA6AuY3LAVpKHfc87SxWRCCit7VViuZ2xWPt9xP72v/BlZURImyT
7o5CV+t+SNHtpvRGUDPrdXGduwl953l2BJfD3mAWHXdFr++8f+KqPoFV3BDfw/5y
ttMZ1Sby278s9OTActs2KVkeZJAAmgvRveTIArSVlDL2mjuIO3gZKxxUJgrXLu8L
YCc2CmXF8Un/EYk4WuSkROAS93qIdDE8TapGivdiTr+qDfhjfTZ8g/1NRbihgvhC
ZsUG+kZgQeTbKKPwM1bJLX75NiixfzFdP48vPHzkrFl8Wvb2wiOr1CMzCYFkV5nE
FjNw9IqVD5h5o3wq3LBW2gSmvKPUFMiamdwg08aVozwoXUOhcARgNaIdwTs7Z2f4
UeX52JwiIcyDg8R3WtxILw8CpszdZID9TNN96D8Hmm+Yewnk+kA9sdjWwnUd5OY2
HqzoRlTiJlrhTJheXxDUlqGKUHkN6OzqpiV3/+4uRM9RFFCz7l/VAZ+ccMt8O3LL
cMYdzcHogKiRj/DBdIjMqqrVPbDTNRW5yTOW1uSKZfTs2HfvqhQKvUrJIDntTWlB
yAyVexaPQ+gjDckYHZEKDVgtkh5A2/MC8ZWVT6noviBNpxOThA/GtGnamqR8WV9n
FJZiCrJfzsi9qyY5LiwRwUKbFXPWqYQCeqKvmbdYwlhjE+Ze71Xqt0HfNBhsGuVY
BL70wuFp4kFeNFnh+1AewNzaUVnNVaSi7JVRmXdbOHeHRm9uqslz3Gv6quu25hSY
CScYHgf+w9YaWDtATB1l0keIAjqnuasABG5L1uW7e/4bSz+KEIZEPRuAgUlxSBnO
3jG4AHAm8z2jyc3uYQcKKl0JdkfVDthGzWMTDMEHzsXbhtXdWKC/PCo2OxSwbw+U
5RtK1aGcMpdIo3U0LRu0s2YjeOlQ4HDeDmeDmvESkXPgotvngbGw5Z8yehhkCTEs
RrcG2wy+Y0PPPLxocvO7M5POw62B8MRHz15TI64tVWMrYP4pGcGXyoiiDv7KmqsP
IeCYvPaM40+NwYrph2MTc0aL5j2trcLIP0wPKnI9UNCz645uohxp+RBp/UMMFwZE
VvpJuRJVWLl6IDIlZx2H0pXqx8itLLY6lbeEhNqsGKGxw4wpZAkvPLZcZsnYW7Ql
oj8+1PnFK7qiG74Ap4fTwd92jIK2o6tcHKl/ALN5+TZsz/Bhstg5LWeMT6BWXY5C
8fzrZaG/yJRJacgsFZcdqxrMfAJcAF3cLdTO4OKK1WtZyHyRThw7aHO1bXpMeTiP
0InfQoFO36JisNs9yhPUqd4TnupCSQFhuiYDQBwkS56YXzwhBs0iXNzVH1r1rilH
xqMoHGr2VRjkdP6C0ZzbsYodOVgZFwc2xsr7Ks6+MF7+JE9V3oZKl8Ki5zkNFISz
9YSc8kKzmvz7oC/6e+9wPWiBky7zjXr7fyrCJzF5FpK4wem08aROOJbgufoK0gfc
GCz/jzAN1X6vDP7MAIwwg/y4rBGhNL9G5vhl0QQ7eyvc7/zYjR1GK3aUevGYSPue
fz56gLGWE95xtKwI19a7TJYBLtAzST3JxGyROlXElfkuPxrrrbOxqHAz7BDSXIwl
CP4dbknI2HwjakfY3dnJyaG5kP7GRZwqgfOx39gttOvr/uz5xRT5FVJwonRXEyMp
We7gmaaztOJ89Q2ihTts9Ib4KrWuBos3j1ssyJKofhlYRsUBuug7f+RAgf77X1+b
XFdmphS4fKw1jRGUHqLaTPRegDi2boOHMDa0vPY1OY54Z4HvyzIUx3bQuUtqRJ04
XtOjnKdwOQ6cnr72u5VK7CCvp4W/eO5q/FcdYLKeBVzglwrw/tPDL8Z+vrNGD0ST
Xz3glBCijvkz8tEnhBU55VgzlPucnSxbrBR2l8nWsJcczjzdBLQUbse+myVNWTJj
E0IElKzujZewYR4WJuoiOIuoPZO1/vnycMU4Sanurh8xhqkb+q9pwEfeiEmqV/Ih
5m9cGjG5/3Z8TRnEL8Cq0mw8RkTLX5RYCbl/muDm7iRD2ybnkWULTYpaP7iF9ddZ
jzMzx7Bg/VOo2ysTjn49ZbBY6J9nOVLOGC9ujXkoN/dKugWHAIMR3Fe2QzGyv9EP
6/ZI5okLIJe3eUShzNJKwQ5M5PsOMAw/Qeyf4f4jyMEZRnC3EOvL7KDbuqF+cmNz
wA83I5yOkl+V51NXGUMLNFj3FrR/Tgm9LH4L/zxvzMeEwfeT9VFwPr8tdTrK0iXF
MU6HFgQDLwLCz9rhJkmQTPOb7todUgfGAJZTX8loqoktYNaveZF4Ww13HkIfJHs8
2WVEmmOSKXZlxpd3ti+MkwloWRj+1XDNISNftwNWOhqzcF+P0kBjf4X7N40CHCv2
5rLeJoV48kQIq6OkSDkP30pugy5kJNSATQZEfo8tBnzOsPMQoaywMvoPzT/A93py
ivXQcbApxAjM8Lu05HVj9b/ttRl11luYpJc1CkNSSJkD8sviYnASAVFD3RAoQwXX
UHmb14zee1+FE+Ive5CEo/JXTgdrVlLgNvZYctzIM0ftNfEyj+7dYaDdaj10oh0L
YwzdCkQOchf5SKBC49P3SjPmMflaLbE8aoBI3OotpsjXgQ+KjTfMhWVHBUQe3ZaZ
iSYkq+vW7HPLljEIZGBoKfyWhjEWs5oCpNHNObrXXgSkAOmFyGD8tHFz0UpA9Kdj
i619vM4r7NAw1XC93MarvpbE8D4P0JwbZxXAYx6QmGpiCt55cajPanY5JxYOznR7
d1NQ47fyxYgWcNBw4G99eXYOl/Gt6TAmWSZQT0NQphcZF6zsREiU2ywyt/A4OgH4
PdL6rdPAFuJmAAJ3JvuY9/syia+Qqi0MvCgkGKH11Vte5/0hGlgE41WIjYcUnW+F
KJd19m0YSv5a2wbXDA/ixuYPGZYryBVKstqV2zthx9dsvF72M00YnRKN0tjWq/vK
x42kWCZeJdA+2j4uDVXnUkO9YC9BAc9h1Pw7AIjUx17av7mt1Sl2SoRLPAazrAzW
pfYxznqA3IZEa/R/qmiielCvzvE6yNZrPwNfcoFyR8lUMpIY45yyhvNRTPLG9wlU
O5Hp18kRXNXDNq5MlrNBBrMvMHccd0n5xyB7tGaq4gQdHvJwnDeM/E+fcDTr4IGt
XaX8eRhA6jo3zVug0NhTXKswePCLJ31XVi5w0+HJzD6eOFVjl5scpvBWWEZp2N11
0hHNg2JXwAe1ByCfZBj1/8XkRdIFDFLlnYZ8pVq2+L8rX5xX+HUGxv/Aua1XpTXo
+jhcTLtMKSqEVghBp6SGsEcqWp6cVlbQbDU0KkjEatrTGMd/Rk/IJyr9FecL3iU9
uUKnIpV9C6GS1uHm7fyPAsKz/xY34z9SMkY1fq1EE1IhN3csnwc0JAAGSrnjS5dL
7uRa3Co9O4Vr81frLzSIObq/MVKwvXCeC0if7pNx9IRBmvxSNzTVH/miGZcVNbo+
cJUSd92uxd4C6rBJFvS9hr/zksq60p9WBbfkju6IrgWpU1PhU8ytB0XFpHor2mvJ
dq4BU058BdH3O4us9/BA3df1HHrbfZaxl5q3EQIZYM0Z2pAh1QWeyEiCieiTs5gI
pWuAZ5X/e4dCZx8k5Enmj73G25PbpQ4RvyLP1fdd4QyFmaIEIbiDeH9cT4k3kjWL
awFMhQsHDH0MQwk9+jUS+xYvDGmGMjsvEua53TRQ+CcBtG8qMlRQ0PYPr/GXegc5
aTQJg6d3/9OP7J43XMA4kYyzAfag/z7LmvhanibkuRc0FY+UITbfWBKlenBsZA0q
b8PLwxWz/qsoDoiH/Up3XSAb0pu+hx1dwLsfdwtqgSHHsQU5d8s7w/LAG9vAX0kf
zGlWKRe4YdqHy7YcuFz2VvksljHr2nzyhoiK/gbJ/ljpGlRnStOtMSGZnB98W5G2
MvE9c/XkeOzMLOe3Ihnm+vwpXNpAXh1uJr+dIqaTJb5qOTEHozVxLSkxJmRqIx1l
KlHSyWJiuVwAL0ms4A0s+RtknKiVqbNGQbNGmN67qZdxdsfaMSGP1AshfPAytEjp
S+se74Ah5zx/X6R0tiN9LhpxWFA+l8ugOFg07sLm7W7fHF3zCocY7tTuXeTfBA1o
b1yjs9q2trZDHxDtlEAAS7W/KmsEZqoiTYa5TsJuUZbvPb/PXUdgh9smYH3BgCpA
qjFGbM0MsMtb8oH5hdy/UyXBzA7L7QnsIhtRdGWTOkno002z81p2apzdYhI6MKRg
EILHrt2aiU9vzz/E4nqCS+6FaWAuHvJD7spAhFPAYGhKmxYedabyMVXXrnd9g/VH
iEV04o5F8SWOuMQnoSoT9H42Z3bI97d4WcclIq90Lwz5H/6ZMB7ECVdTNov5oQ7d
KKpAOAfyEJLa8XUqP9By5QO5mh73CGhXXZT0xiiNyl9YzwqsltDtgz8GqFdKCtmT
vCcheHwoB7oo3Hv78WPVZ3prIaZQrbnQioHeEqwsqWNOBQSzr+fmbFZsai17sYzK
LuDyKhUol+5yWi1d1qP2FIzbTGXHirbp22AIzTTPB7w/+IrVVOeS4P64JReIDRps
0eqUmUZbulphom/NtPmgKvhjyzC9sP0OQxM9a1dA55yHPVSTRKXqmPlnW5n3Mo6P
cxgo3V1ZsoyzzD2y0s1Qy6n9zuLtMVzSNnS0Rvy1+xCblnDs3vdWisYtpJvhJvqP
CGkbVyuv19kYRR+TrMIlbsVyLmGIzfgcIoVwebH+kygYSnBseR6s2NjJIydZmc6/
1gQkEL6MJFb1D58+8I6/kQya2gTvRTKesL6MflHaz3RfEbv42DNkmI89prCOU+yr
ZoQW/k8HG3yfflHgH39FmhqlFKFQIrARmxxD8bJ1t8/KXcxeJiW1EK6GyC0kkrP3
y76O8QZvTCLVsROTmzXyCZUtQ9kQApo7EGHUZm7OhpX6OZDlAIZU/16DbR3izZj5
HBP7wMbewktAKgNUf+JPARS1eH4hgL0alw5gT+iUzOTqgqRm2q+doDENexk3TFbv
7kDgjynyuI4193ml9lVZZx82x8sLzFIqklWFfKl3xxM5M4LKdTQKx8ogOJXPtkBK
0YCj2maFG0Uqd0utNK/Axnjrcf+SadkmKoJwCmkWBuy5FraSIG4ZbiQa+FbmkKyy
YHUZlOTUM78HUeI05NjeposAk2/2jntxuHTDOTOtLs2eO7RShmdJTxf+9Y1/lYhY
xcwZZK6lsbP8CYajFv3FCgZepqI6Ifrr79fSkVtt7oX7LHViJ7U8UwJZgNWq5/76
8otq7h8mxx5ICCIDgZ54mChx6/dbhPU0EKd6VHHIqka1JeVmZgl2VZAXaDUHRudJ
XqxUxFo2BVWIzsQNpOXHSJWq1Mgi/9LKgJFfeDlC0DcCUNOQpjfJ2/EMPhD0gcGk
IxZGytw4Lpgw756ky1e2bssJWLg6r7u9zayTQptXzv+PQ6p1LPvkIDL6cM65+D61
7u3s6ciYvQkc6Xb/pwf6E0oj2U8Qz63mk+PiPa8ULTs/cVpyDOht768+s7PBMZQM
jWP2+4ROI1BEa/HmVfud7RjDYRyYZLQynZWZT04XfQEFqqkTPp1DGF0D1XPHddX9
SiiY2zXkZl6QX22KVN1+3oamMeT06eUn/bWz1clW8qEgppGhPnMJRWgSvaJHE8yf
hPHgmutekZekdcDl6Z0GR6HN0MamI2Jy7tJXH69+3xRoHbM8xi/+d6t2xG/m2jEf
sE0r6I0umN0wRN4TuubVqCwc1j4kzMk3IETOxuX89misJaKGBnexahLAYUBdNacm
RTqfMXK/xfW2OgM5xOd053kFMyLjTaQfN7l8JOAd6oKDpXIAS1JQrUI16CQ20zGi
CcqE/2ykJonl/cx9M5EMFrGvIQjzJ00xe+kvTiuJyRqkgwGuFumWHE/2sNSsi/AM
pR80PsSvoMZkFj5vzE/Zx/RubupxmcRav2w3iRfoLPYsXPCAlwMPlW0/fI98PU2q
9qCap9OJ5ZaSjZtTqU/zjEWv8NMSa20QjMf21zj2B/Oo4zx0KKA5DEtEvHmqrL84
iPybx0BBCsJm6C/k5Xrj+EOBU4hfbaYrbUuL2uG2+U0B1J08gWfibj+AosCIGPKB
u1ogWYLEuxRVbMlJ67kFyQroPJO4D/164gMvmg7dAzWBrE1VDZorU0YQr1tbx1jx
mlQ+Y9/+RZCwIQYFkiRj+xkU1bmjRfOYzlZVEK+8wyh+uOYq8eCp6cJc79NWmyu+
YzXhqlLIBoBz4gJBIFMO6qN5IhEwEwUAcQKAPZNL74DnVCymoXs+74149i/+r2m/
2zvrSR5dDQ3p8iJlAwlBojovT0LDWO322vllG+OIUR41er9M2xmvTw3AVTW7fWVF
3yJPiyQFaSZuM+4qRMwOP4YNqaCWFDPAP7Ap1I0txDa3Yj8ZZ1c8XeRNKZMQQ/VA
1dOyrPC7IBHP3PnLokrnIN0XJWyhjyIx9Gp84grs/m1ZQQg5s/P1Smvaa/HHzqBk
ok+wjuByIWZO7cpuY9IQw1BUEpHRmCivNJVqTGJGYOp3g4GihzHMrAklqiiJuWuw
P2h9f/lAfB44IP/3aefkQOzSJ0SDUJ//NBmGe4DNPynLttTA1Uz/HKC2D+pfPDpf
TBYX6PSTLJIs+ZBEF+1u9sk+PjR2tW46G5pMAGFI9wbz1Yyb8wGzQOqBKzJFb9MX
4aA7S2sHqnRzgePJ9q+aH3L5GDnAoqMkhzEpKiY+66lXu7ER9HVQerI4Rwfd9OMr
12Bwjb5LJ8Zndv63a/CKT20/W91VHhaAlQ1XtqtM+I1/b5yi/5ddyyZ9ySkjnNpO
r035n49pGEbBuR6pDvVaUs/2qr8uXq4NYjfUeVdEXdQvxAA+Y7vKLHOve587MQci
g197ly7DchXeKAXt9FALvo0/nUQUdW5+xr7+CEmCm0GoV+utbHQ7sUqi1NA2MCSa
UvNl9csO+Px88C1ZJuq6vk9W1VXU5+c1s2QvU1qbzmrCqgErDdaBCHARvTJi3/6H
Z+wGBHGtBHYniJXJGjWkeLiqeXLlMiZFsAzrIGONK0jeitkccn9iv6nWG7JFe/hC
w2bH16PIKINDaCyENTIY1wfRZdT+GxwTK0HiwNPmkTuJI9Lms58aU4MgwCwVGDW4
D6aoXmSr90cS88EpO9r6Dt+Ia/4AGIRMGM/ui3Sn6Xa90fep/LLf9HvZAikfjR+x
iHiQC/BWGhSbOL+KdHgwQIwtpDtQdWZXAgP3yMkQL1fGJ7xiJhrxHagJB8KnoMYX
9ZGDr8YUfM9CUnlH8F67AmX/0j4GL/+XGZI0TALbZJLFzXZOUdRqN4DwHUBgXcVA
jbDani6dSgwKaZETz1Jr7WUmFM8ShyVz7Na6E1VvRKC8/OqLAhEtHC5KkNTuTZKC
3j3M+zvksfC2zOu6VHTJqIULDtaZAPOMcnuWJzZBYb9cg7Fzl6b8KK+eExV1cE9q
NP5+tZbnK6ieUD51tM1BLDBO8GnJu54zGoV2w/Rnwnt799BNuX3lEdqY/T5wXGEo
RAIYg6uhnajemjNOjBKEzS/7VwyaUUb98HD4/ZqOkaEegGN0duBTMzRpf9Bjh08Z
BQSZ9aJM6uJY+fbg6xs4rMGsq9W0XtNvC9CPGVwhBD6ymYr7TND782sSnEVI+tcz
FWsjE2pXbgI06lFGleEa+CPJ/YzYErTYeOCR5EdSzWg3Ven1VJkGPcay/+I9YE3Z
nqpaI1JtyI7gxrwANJYYTARDEegS6IiePw4zPQ1Cpi86nBS2MtE63YdxrwuwwAOU
SSBB2mMJlPfu7y1CcmYyxqH2iy1Cln4L05UPXE4fY5/Wrt9LZK8YiFK676rpiQp8
6xU7tOUYzUkxFB4z2EsfB6gdgiXqmVQZQBjARniurNN0M6I/dnolga0WXSNOGtT/
8+AK2KSSncFjmn78CfiM32VDemJjStOeWU2bdt9iutk1rxzOpTfkED6401Wee7LJ
3Yv4Y9NVuZbqPqlNKOtrB6f1rFUGhVgAKsbguSHQ+m/r29ZCFh7MTquc1EC/lpxA
+u5gXMhZ4inXMJlnDUJwDOTZv0vr6PRIEo4yoI0Wks86OB8KKY33PaRWY9Udi+fD
PWJUduBbjr/ktaAFE0L/bABW2fDJVMv7XIXNG1viHVQpa3Xi9+Df7HzTDtkp3IGV
iEnzE9+JSWRDJno8mw3Y+XB5Vf8Ir82hdQLe5ljGRcTr/LNWZC+iBviuarhsQaR8
xDnetqds+KErZEj1v9IDNBVEwGY9N2fSOV3D08vnfknU9A6TFKYtDu7rBsTr0aPA
IClVBYcaKWjqAuu/LjEAwR6X7lwbk3VpCDvwmLvtYpeuOFsm4gzZ+TE+/eM7VojA
55NAcUktuMwTqXZS/HDuqv0gOnCFJoOKwT0ZVWsaAeCorPh3rRVU8a+e5DAmSrBP
3N/JZQWqRLfr+quBaQKjGmp30F7kkMnd+gjVWTANqc+1jW8fkk9ZUD12H+Vn1nyU
JsW33RPMks11NLmp2917ow==

`pragma protect end_protected

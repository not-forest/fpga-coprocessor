`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Wz7Uq/BOal1o0c5Ut/prlrBl26VgIpNjyHUfRDALtbBVShj7ATNssjlfGXEP4DvP
2VuR8jCsqjszdbPL/bWVbtfWdQTm8tQJs41oSonPRXPVZdNB9kdUuJF4wct6LE/A
HfAyF+jwPoKkPOg8BqhpgOHfO8PobH2TcR5nsg1BUPA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8816)
MSXEd9HJogUL0TySJ8Kxc+Y1R2coTn7cbqRyrJ4ZTqqZNqW1M8HNnVg60Rp4gUMO
fBObKBxcH8CsQtUQhRWPhOZxSRhWsWb4xbSOrwVbqEb1YeFrb5qE6CoFtP/vh/vX
TckR9E0TyLZEJwiTNv0/rZaKSx5K7jfru6C68oRahn3InWFJuC/IxWdY4UzjnOlI
7xpnrRfI+hAtytx0ptwr01CQMDB+IMj+/pHIFRMIh4D0Xd4tsI22uBTGrY2ZZkt1
4MrlRfNeHriP2roUAt16lVcw8ERmltQ63i5dbAYOssQF/jwEfXUrfWAsx3w0QXQM
etYxIi6UCW5QRipjPHgorjJ45UKgQGHjiRyFxy1AsmeNnIyAmZJJbEbuD8x70MGk
NWjNBL5KKdG4BRpJJnNNdb19zSHG5shcCDrVQ1stdVJ8iA6/ccdCkggmYYhSPCDf
J3xsVr1PIWPOjKxbwDpI6lkJHInSEVTcmumMoTkhYsGTtauvqiVb15VDb3hBL/Sn
vqcRSbvLoCYmq+aSr0s3BHa/X+FSddqyUxEMnwurgDopxrdL7ZVMlg49IELJxrb9
mRC2fVe5eNrkcnDB8nWD8VtWn3N5m2uMrwdOI1hfshtcYlXfzTZduqwhwi876wHf
ENXIR213CeUzlH6V6VWLlaBrP1mFdwOEKKr3hP73u0DrZq5zwbuDHp5r0Wc3s4rF
5ZrI7/3fFIFjqgubAkz9+cW3KykbMrwXdZrOp5KaxbU4qBkHdhbI8EJ0abJhOiii
jHm/Xv8W1WINw89jNPRrJGQaGUIGBK96MiEVB4UzMzHwgQxMZn72oDW9bycihNTK
wRm/MQ0n6gJzSG36H5cH/Twd/L8CI5K5wOZKiJi51lUsASkCHL1yK0CfyydmzA+H
mFCxQ8++SaWRzADMPSqc1SnSCKhUMpqErUgP7kYBQgmhWKJUBumeIDvw22ooe70l
2jak1dF/3S78jAvnkVb9akOF8JSgLjrVar5ZSXP4iYhYTIeCwZ+3mytmTF+5yZu3
CnNyqwpkorYFbqMoIq8KoMp78RNr7cb645lN4IF8M0/V4V3C2QFfmang/3weX7pI
AL7tfGb73bnferM5ZfJbLfXflaLzfTFrjTSGVvxOzyFygtbGy1E7YBLnxTGMzEYg
P4N2ZSfu8JvN/6UqfYkJy40s1LyjZJvZoTfi3kKhiCpfSlqcxatvadV1tumagWAf
X/YgRbT5aey7/HzPHBPcEaUCybSDf0VKNP+rKaGo6oP0gh5CQsjoRekFEdPJ1Pp7
/skjl+L02PD2iQy+uz9XafdIyr2AaP3Fklq8gOog4jOD938YPoJzQNB7GxjcIi7n
JSXNY33ubwZG1raJJaNc5KYVkxlHmMEZcsqnSZqSWmgLx8fW+c73y39KM/ERgrcl
5BlFkfWCtC13Qp3LSsjmB+36agIYsy8O4eqcvy100iBJB2A2GvqL+eNI+0Ij5X9g
bPq/d7i7ttUd+AujVbJ7Nm09A/au4j86lMQxLb6KmavZopHUvhXZB2xFAoSSG2C4
Qzp+iFx0aqjKlHf0mXr1DuDhiRPXN6LvOs7LAfFfpRzxfNMs2cUQ2ftBT+mTNxtC
Lrsny1jbxbV4gA42sZSKchgYsZiK5s1h5jOGBN6Yyg3kWjV7nvq3DDE7hXi4gyuO
g/LjOpALgR7qPA5FRyAPmGsKCSWWqt77l3UDJbSZ6871fWGJbJxel7rwOqKayac+
+y5LNSb0Y5KoAAONZbSkP7P9mYehlOl7W/Kj8ZLd4JzYZnuQ4xLjwsJfyfTGvRYq
id2HdWE/kekxy2wXppG40D612PuOmn5GWGd0TK+Hl8QEihjsP8j+Q1c+XGtA7rrA
Jii2UKdeu5gso09u5/KTiF6lNEuA0Z+o7hc2pHgh9A8Jdf+px4EcHbYhNLg88VQb
9UvwNz5s/f+lWcLLlipX5bLJpBwlPAkJWPlB6a02aqHGjvF6HCteqiJoZktgK1ss
Xzj+0W/CgY9cFdXuRzGP5HMiY6T4C8JOT8dGH/rSZQJOVZmHPkez6djP6Csq/usx
daCwLHhzjkpTUzOgY4wPJTKFPG3/Rt63bnfpfz5K8g8DsQHsrN87czdvNX6Dbb/z
onMJmbsL47xmVbT/R6FQ7bRP7EMvylvkdoKWd0qUXiBC25nLTmSTI9c0rEN6K11H
mI8Ql5oa4ihyyD9ZmpRsZ7pK7HnAQf+tjjSdOCoIVm4CyuL9AnhzXMWd7vFoxfAt
lsAQ5wYwfm65q57n8bVbZ04sVn5MyHGqMWe1wcyHT2kRlO54GYxxa/dOqCle1teM
BB1E4coJ7W+8EaX1r5SNgRUF9TzNdnRcj2SaFldNCrr9kg5lxCei5KPT7fwVk5Zm
idlmVg4wMAwEwm1WCCNAJ2PSAAIzQA0ssCn6cGRMamQUrv/bujKDLNIedYaCISEJ
q6uOhYCERetc3pEcFj67T4PDun9JUP9aH5BSc+KQaKEV7B3uryTPHRK1FLh/DE6g
wUnCtmQSM726XUmNYgLwhKnRCpoy5ckPeDDv5OeXGQkl0haAgQQPHyElSRdNuRXn
qRMkzpMIf6n014URwkbnRUvsbxPRuW2auwf5bEaL3hw15fsKjOZe02TSGa7NydJ4
gwfaxzmAhRlvx8ri10RjkOyOBEg2AwCvN64IRJaKv9a7meVb2ShHKb2bOd4ZO07/
N8BOu2xoR4D724k1K3uWG/hhiDMzWOM5EfmtyqnQDPkgUTvkSLJyxEFlVxf6fmuC
Nz6msQ43aHSVyqJrTohPHAxMJ+OB9V+FyexMBKzsPgxunIgZJ35Q8LaRS8N4UpAh
MEuf2tJGAqJCHP1ptIDpqI5Pzg4rPk382Ilu79qeaN2cxmx2CzZ5WNgVzyzlJsAd
d39MrxY+PlgjDMtgW6OVZRQhnGY3WC7cxaPIikGU1Gxz8uYLQUh9tCHP5VgEGbNm
tsVfvTPT7K13aufCPWo7ptUsj6QmErmoIUk/3PGAplsCMPWc3rTKf47KBPpS/wIs
2E2Q/vv1l/50n/zjb2fbUYYmVD6A+lxjfL3hKdqPYBuakzwJ2DdETtnmbEeleG81
ED2AZG30ne5MPWo7e9RbQuj72+JMMwhMIfnypwEwUe78xDXs2pcO9b+QElXYB7r3
ciurzefIQ1aPiQIy575P9EdYRQIqqsZWZdTHh5lBi8qUUumGSQbby4CUBCCE/7U+
xdfud5zkuRBCI4Ah7VeNjdLpTxpq3I/rqEMjn0gSGWJKJdsmE3KzCwT94axmgrrI
VPeuYXeCJQpsb2sUoUc9jUOLFN4ohziWiklNceqJJdPbmARLNmy2rlGt+BkOxbHW
m+yi+rsCW4AsM2bLHmBSIjgZowD0rzDhsuFehEoxnvb626GlEYQN46iNNFFYCu99
u3LJGZteaBSgGKU7qrYZRxbo6PaY7jngqR9zBRirvDu6hbAqCjRNww9J/1JyLCHy
y4AJ5BGZseR0QgtJvnkbEeEvagvXYzQQ0tAsL1jdV5QPLB4GaEZdSzOcbRVa5k0+
eg8mqIJ7ZxaJf1EG1hDLuWewz/EtDBp85t79gB3lKMWmKafGX49MsFJ4eOQZYV2W
0VH/cf2N9Jq09kHegyey0aNv5hqfBn9wehQbutiTuhCrnorm9dnS7QKGQKift0mN
IxxMeSM55N8cmY5h+2bpEsRWAgmYVcJKJmqCTthKhI97cZpOeMfu6f1f6bMCmCyc
bcnHfgQV8vCriwYhr2jPpFaVgbgGctDteRD0KU99uM78UqOlE7Rj8c78//An3Rks
YL7l15pObNYYkXikcqDRIjougiXka/0H62EIVXdltQo2ccGdrNSS5uWYHfbVd/aL
xZ3TwP7xzYuv0DJ5IY0Ia2gmcIQUvEsm2Nz7ufE0MH/Ut6RWQS6Rs/MkUnWHu0vz
6mFXlMfg9SlQY2OqPPN+HeUa+NDISPUIUfAqrXa8eXNPzRhDd9Cuid72J0z2NsYH
B87o1rMPSI5WsxpK5W96zTG0qHCm9OWvFWTPPk2hCLzc/oBWLpcATbqCxb024wAt
/KsdF1J08M3O7XkzAxsEATgEDU2RRIj9jp2uoI6eDjHgiLfPyPPMJDNhLOHbne+T
M4Y3Ps4npaSDaFZ8Q7PDmPKSFHme8qFN2reIaWUNDBys7Ui5B3RKmPPDBBLW5Ocp
8TDm61jRu7hVCcIqnjEOzC7d02TdNfbgBLmxNesV+uhJ+qvF++xcBpnp6XYFIAGI
/7idF4sp0GbnLeaQsQiHvg7PTIKpCCB743IktWMZ0XZKjRNzh8JGVG887QVfK/Rg
BDJ5FnKBNlac5gkHr1VYwdNS8SO1J830PC37V4NvSJ2MMtMWXcp8IHA9ivNQjfrh
hbhudvNm7tBfBs8jlfXtIWklIuVylGknb32FsleOrsGvc5YOoDgudyGY2MLZ29hj
t/AX6lUYj3Wpsco/OhBwEUS7ik3olZjAqPKq0SzVQN03H8wMyyMljCK5ZBIAcJaa
qoV9bFGe1a4tTP0NASFevNAkJmhLVJul5YbO3GTAnWJD42BIhaDYTI5GGUWyXABh
AG8sO2H60/cFrRnflTYyCE8oegUxspv4mUvhBz9Peo2B9rR9FSP4sdRCEW4b3gc2
RMZBJ9Lx4yJJCN8UjWfnP9ReSaDs7RynCM81s0wvan8m0s0wIlNioRetSFVlKvaa
7NF2kQhr9O799aQHtz535Ur6292DFO6CU+Y7yGMlNMbV5sjBIyhWdDSXYLaaOJVy
uM9j3Og2UVcDAjpWJUFuIcFvtMcBoCycv2VpXcLm7cgcPpNigUpkjQ03gP1vWkL/
jg0Q+uwyfF5f8J+crZTmFbPqOFdFPoPHMSw5b6O3eD+eI6d/vt2IcJbo5QXjEr7b
gA3psxS2K/clBBateZ+tu7V7qWAqNag8SMrYmGJUZyyZA2zZ+zuPfxVakAQR7TZ2
5AgD6vSagQFu1PkTHO9QZSlPcEu9cgwVFWPfu9/r/+HcZwanv75QSXlnzBGT0HLB
3qHer+J4C4ESsL2ANlie6LWKRUc+K1Qe90ddLZ1QKWpEewxBEXiRJ0LrHU7tvRPI
WxMw7MwkzHGZeBBHUMih9GzqNMpNqzm39ZiFnR3TD/Ul44qch/57i1jFu6tQdNxo
+1xJIgv/CGHvjFIZJgiZGWW1mNuQ0B5TAQCHnFj3ZBbGdMVGsQ+J6ThycWYjG+2k
5j8QbpiI6PuQdWfzg7rBP7nJxrZ83G9TNh0vU3FNPOwWWF1z+4R/nrijlUtkW94r
xKtidKnTvruv5JFVT2yy5I4tbViaPrbuybCgE7EvLl1s0pJ2xPauO3Tf+BsZKQJ8
6wpvSqVEqqaVVv63RCZgnQEDLrdPcxf+R3vMf1rbBz3TtUofVhxIZCEFwMyPwhjL
Gqh05UhaxPiEgJHQGdncTQvGAp7j4mBYbAuJR7tuQ8KLUw45Likp9AUNC1/N78v9
ZQhmd+v2Xz/jCuJ+oKyGUhHpFM9zGBvp2bkfEFS7B7p8xvOizWptM/IWgixEnw4P
fsvAKi1vyn8jE3pA9p0jQXRjewRZ0Z4aZSh7KaW0dDTCcCJ64TTotZibdy4wHB0f
BgqoqoLiJerp1Vx/HVuEU0aLyyoN14lJ/rT7NyV06/Qh42XtLpo8VZOdw02o/kib
qV8H1D9gqZ75ODXnYyF75dMRoJyu+DbKPdy1HNU8iCmo4d25RauvFzhNidGC+g/U
iSDJ+T57+F6DOzfwY6aR8rPXk4Nfi6nkKaoq9xuB7l9sL6KbSK6RsNNs1IqjgpW0
wWFKhledXlH9C8sMxsy+nTopQITYgL135fDilJN8eBY83JNkntP33SzwCbj1cJWV
plrr3Kvj6EB4ElO5hPTDW3OZ1HNJ4Ud4G0K/c6kZk4ir/t7pag9/SsM1OBLn97j3
nKLXrtt1AcCWrhC69R6XqSFq7ODPyu6WBrUa5iNXfYCuFQk4lRq6rJHS0jq6mvKv
4gtq2nucyWOfxx7LuMAnd6aZPSk9JvmzYHv1WAytuuap65h+FV3Y7qbPD8kzkixJ
6dRfiXNG7NazBG+eOvqtM7x0fyfKXP2SWPLGNE6s92O5tH4rLtdkLA1y6FMhorLG
AYf947NV4SSAIPC3Z3pONRGSxAI6rE/1lrCKyMRHvgNlHWR/JzTrIS56o012Skfi
h09vuQu4gdg3yF48AZrZepvYUtW6tARgqC5o4EuNZW8YzTkSG7DtHuGyO9AfOcQs
mI/WacV/cHPqCetYfEqIDIi2An1JAda1BF9Cc23ed4xfHPpce3xY52OmXBtmV65v
zQ9M3F7PYRwOxC4v07AP7UPrNG0YoHTNk1szZfyCdeA9xfbdePdogbJ9TfUrv34r
GS02Tg7jdspVxbZR+PeiXQLAnH0C+oFvI2K17AqMhys/SD1vJxNrSkDAh9DZOFcs
EPXKtYPrdXyJLv4UzJtT9DRBNvDnNHspJJ3maFzkOY+eGiRbMkjJk26y+2cJZSoh
y2waWRzoenVr/oU/LStmcN1OLVPoya2LZH14sPrkpNvFz0pPTVMJTHF89uEmelXQ
zOlKgnv2xA3zlQorjT9HZFRRW9dP1YzClm1RkTqvkS1somnvyP6VEwYNyoHWGwAF
f3kDWLk/7LxksUfczB1u1qQxdLsB4u7lN1d3oHnhgzc705XgEEqnwkejVUzd65ho
e6PvM3PKAHVREzcPBoeg5uqaxExbDLUrWOuevBD2RDpBXW9s6goLlM+hgY9Evxdh
0OtAvhw8jgsORMHkpP1pvo6FrPXiDx9bv7katvVA0kAqHCRxgo21BiJQx5ybFky2
irS+pLOXEHxBirJN11J5jtQ4arZWI7n48bdxLlGNiyNSPdIR2RjSLCXO3jXAMdHz
ovBJS6Oo2e85eKc5nFzUzP+ly9RP7Kl16oOA7bmVmtV8ZeJxvJ9dS8aIqGVwGtdT
wyHzLsYPZyWNGikq3FeK763Gn9qUeEkdB8HEqvY8il/S/xE/nAyvM/Ac0NAe8nHd
GDZ4mbliQTBmLitPbkL0uo3sT2/slOpPBm8CE6jSy80xBjH9bcB0maHLanttK/71
T7Bg/V7NJ6NT2Wwsdk1kpRBr/iNrXc5H44stPPlRwpMxb2LAFu1Jun/MdITgPiQm
gWAAiwbHmWwN7GtaQae6fSHMqwX8GO2Bu6Ydu38zYUwcG6JdLNrtX17hDyIcEN/6
u3am5V1brfq8nOC7ZeB9XXx7BA4H0fUOQyxTf+yypKZhCZsem9IbmQ2VjyJoBZmS
jF9vVVu8gEQRII/rzfWbaVrg2970j1ZiV7TpRcPjRkQyGmKmo/LkzQ03LsWaYb+H
UDeDH1eRFELoi87+z7IwdDx/MjCgCxWt7iygYWvG6w1BTLrcBGDAwPK3p0ZH6nMa
ggnKsxVqUWPm+Q7K+xCxtPT/SJYb2FJoZBhMCqvikMTw5+zgVOENJv+AszwYXgyn
eD2CYHgZbncKllne1TymYLZHFy3bwdYzccSU/LwOouLDRIllq1d2Ao/dD5TMa9/Y
s1lanPox+PE+HJL0rJfciOnKySeSiBh2aEaPkMMlsgkrYrzCjNphpGi7qOftxcWk
WgksMRWMtS2bC/QOmtNkQXZqHCnPWMYvCsoCQQJNtM34TEp2TWQL3RPOAawBtzSx
XVAgDgJcdbBgAa6ksp9qNGDJbPJtqZE6WXIFSH/nRVUairUhsvu1PkvB7/Y1WeQD
c+MVuMvXzSQHNB5go6u/6CF+DZRbQV7IMffBaU69ZGKAyawEqc3D6SNwz+BMziX5
N0srWJtOq9T8zsMEhzcbCktSFQA+hm4fYl7KBJnk1phBiBzrB9w5LhoKlqv/nH5h
634z+7YewEyid1Zz8OubH22zr09b7B9NL8F0P7kxo1TqkDl7QjlEZ5Kh4Z/M5ZdQ
ZpsGgESuFlV0muWYrpwFC60d6uAd165wrr3YAYV/HZoFSqvoE1pOk+702ezgNpS5
ZFI8hlNE/3kaUN2brWxq56aw1T5V1oMTOgL32tUC408SYlirmiczLq9qTQk3f+9Z
pwR2cJZP+3FBZC0HqiC8V0P2QJzM6x0AhnzbFQGHMz05+6MttBNQLd4c1JyNaDPV
2lSniAyrGplJyyhUThN6evqdDbiE4heZ2kGK7Bs2vCXiovc7aTi4+8YUnFC8Olvb
4oFmxUFPotsvzrdPD42IOejg9JR3nlT746Bo6gsSD+eGEgoSYHcX+W2MympsXZ9v
6ctihlZoOa/QhyNOr3VVNJtznhoKYiM9FtSXcvqPqeFJclIDN8TNmOCz3VVr6QON
5ZSbR9vg2pwOUzlt3Q9n+tbeLXtrpZ3c0Tv/ScugGwxLbxdMvWlxPd2MX56cc8om
GZWXgc+B2pJey+g3na6CZ5faQly0WZvi4d6kLWLqOC+2mZ1uz524iPugqIvNV80a
kzsxPahXIEFhkz1xsqsRE5LwJ4+0ohWkiysYfJCUuXNDgiP1CPLz67Ha7cT6AFjd
kXzDTHe4x58LCBuDG0RQGmmUNXuzo8bGFK8iX5ZcwUx1E/J7/aD7QiAJ1XNBAPZU
fwOVFKdXfPpdZueYqjdSPTCBarHg5b0wf5eRr6ngQJGI9eJgdQupx9zf+4wHDE6p
X/xwdCz9pcFBqLjT8lTrIPcjfsWmu7Eu+gzDEOaZ+HdTc2Yoh10gVEWTdhRYscIG
mlneQkbLTEC4ZVUalv2D+sjI/yywNXKcEctIylOfmMyy1mAPOYolmqLpupBlDHrp
ib9NtV+WsZeuIThHM25Eks8Oc6QNnPh32TqFMDui6M5l75R6ur+DAy89+/6M/Ls/
VtyKxFSxqTZb4dk9NOrX4WuigDhBLCUH2CCscj3y/SrbrHhQy8HSJnw3Catai2OI
ZCxBG1cfrQfwFLs/lMiGD07knpyCERGXC2lC27sz7eUrmzXwKFfqGOZLXIU13h8Q
BwrYZaIMObGuhDcTLtFsss+QcloeKxPa+LmDLNs6sbYxvmvLv4V6B+x6QWawAgAB
AZf7bq2A3/cB0niPq8RZq6jLZEfRiDjtJKGvHgvU+a8AHzQ167XEHDyqEHSZpydn
puTkmdVgZVN0k2ngsYaOsdPA6/kIlNtjumKHM1uhph3QE/0CHNXPt9AZ50to9AQ6
Vs0E0HF0a6LSvp8hiVCzSFOgYX92O3yyI0ADPCGD7jouuQWdnvmZgzcLy5EDRhBy
NIUEKAWIRRBevKRnRBjTIGV4yJHpL5UOeeqBFUUGm7/Yp6fPatx+8TOthbkI05yI
zZObDiR5lAeEi7bKtNsFJLJ8beyGV+dW0DUpoHq9o4bxL6YA1KOBLfZDwzyyBNZ+
XzMpsZnFPXKQQXvorwOIu/vgZlz2MgJScpmaRmrHHMHVQ92hLioV+7WLhX+EhQKj
0SO6n2jt29iGA2OWcb3yqvGTxNEorGAOi37VV6Svaf1Cy2RqSBVzzBWlW1lOPnQ8
Jm7cG/XCYWWUtAmjmseZzCpgJCZgnrkWaVaR3DOsF/ovZpNMb+y1n7s+0OWvSLbj
5LegWX9cqJxMRI4NS54p0IM5CkA5iJz1rYB8H5+XMw6LQOREs4vseiVNOhXRFHeR
MHxcP0qXXnvRfxvUU+YbZK5ikptORS9T88niaAgNf3uOmGM7BHIVYaWwoI/ZQ6Lu
SE0iE8bY3sA3aF6ARROTLHIv18wjYh1BaSyM4Q0i+bpzEt0uHaBmQvpKW1X7gd0r
vA6AGfHSyrLnHDSKfN9hYwMIf9MPhEaOB4f1GaKZ4jnrf6dQx8JwpeGcMUb+7nsG
2VXq6+dS+AySb4xJeJ/KkPTOE9QyiDiuoKnbv7fwERcamkvjR6p2+NY5xe1h5zZu
0sPr/b0MgjexkQRl10gM23l4xlsOTMk0ysOL5VTMBtWnPFOBqTlyKzx6iowy+rpa
/oEZWQUE8qMpv8AOKHQV+nrioEZBapg1AA9VpfQjBEzJ5fWBofPfOJB8CtzzyNoT
pB9bwgMojq+i8UkkPv/7ay5zTyCSNCPkYyVSmeDzwhpkWA/Ka0DSCba06Qi2xIsy
xRJrs1FxMprnHtIETAJ6LcLE3uxL7yhkEKng5paDJXXONbARpngfPAHe11cKS/w5
cR5FrbfstjpJhClcqeWHPGGyXq6q9RaHtoO59t8wRrZXnJ2TOXmOtn1ndoAEboee
yZ72BrpBtfXwF0PiEoMOLQuZEVj0HOf9vql+pUgiBP/hxERBKDiDBxVEudu0LBMV
D1JGa4MYiYcg+55AOdY9RgLirXO+D74f62KCtHfkfe885NC+RsW8S4+P3MAoHr0y
2bwwAOkDnawx/yhf4uoX1zqlJraZHTbohHHNF8v6msAnlrT4+T1CcI4GkYlBSbON
fxBNDurNdxdDZRjNYg+vx7sJnmjuuikblhvNvUfc22SWvGWzFk21+HlZky9izdis
Vj5t2fvJhpmXmtbbtmIGVXoACGzQSmU2LtAhXn+p7wv9/t9mHcAApOsxS4kHGI4b
Slk0HGuMIRwkGHUYqIvwOlyXdFjrY8acjy+UL3ruWf5K7RMUPmVoaocTfomV4yZR
CJXDhuaqeTpJQ278ccsoUFry/pGYg1KVpXk74Ix/ogCRj1XybWDMt2o0IblUoAYz
QOOkwmPLoJexDRB/0bZc/GYKCHbwzFz00pG3RNBh5cSc3qc8GRZ/IA7qy/YCHvvJ
T3nrk8AqgomIqEA6F1uerxt98aOllFgw7Sf0Qx4YsivVwQ166JHxUIeUsCDsITmT
fmmOnRsug9Z9Ave8g3w2NXxKPfUTgDSKiK0l/qg/gS1WwvHLryJ+0YNxZ9pKImcm
W3WafKSX9ycTA4kmXJ8z3aen29OjW7tpV8MtaY5UR6M/pVD/5o4xN32wAHFV5ATj
Mn3pbS5TDlZ14HDie+IOFPratIcyw9/dmv+b+oMn5WVkCIvf6RxFq+num51dAPun
jruCQ3qSM01D4X6TTxtkdSjkHYMDK2MrTk8jBW1DERAFoCLgo7LLX6CxbZ0hUhDE
Z/pOjQ4MLIEOqdr9YMJf2NNO2FO9nfb5WOA5JIbQtMmPTicKJ0DQ1MqjldITy/yS
XEAwTsWs8kyLFXacN7mEcMd3tknkfF9BmMnTXObLLLIw9EAlZCbgJJ5k7SA1jz7o
Bw6Sa+xroj3gH1oO9xmtzOzNw4vFF0bjW6Mzi2qfExy9ImL8yuZkkjj+if6nepR8
qbWisAi7pJEPDc1JiAxOSc0AbbEQ6fyjRRHNhDkr9SKTKv9nOXVZoNDKUbp/6Sfq
v1CnOd+O46GfekbH5iACKj5ENZEF8kNYtYJ3NDXSc6Fg8v8jONEdMJeA0zJbtwIH
4GecXcB/D9MppqxvhvjAJYgLM1/45dzkXljcshbg4xKXI8ZDDW+Rp4pzyDB8JqTr
MDG9DxQM1i4EntmvXzLOEC5WGY8m5BBHsNV/Vvr0lckYCvEMElnPn0oxofhez0Cv
Snn5/MeO5JhRNq7H7kov/UQDqPzqb7LST8yiMklsXmNJLc3hZO90zXmneATzqvTl
x1BOwCf/GtTBzECVF/XVgEYO37+qkergg9aHcq5twhQzlm7BY7ZqQCUIIPSQEiEp
K+2HZTkyY+GnKkLVjOADVK32H6EfE1WGSU7JcznZT6kb2IbGOQUXctijZmO++04v
7qSA0i31zUMirp/h+z6gsJBFGLVX9LZjIhG6NHHYf8yWaQbsZmjyQCzgc2WoOlfS
5zNZRKtBjzmA2V2iVLC4isJpLHnRZXuNs1i8EGeQLNp28FcZlZBLMgEU+bECU1Lg
qgqEqE1mZR3UGCX+GtaZJXqi/TyUmRn5xfHTvFlWPGM=
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
LdEUDgdh2EhVBhSn0dUllOVTMo/Xg1YYsuCKzHp96N9luW/SkmyyuAHSg/Etlbc/
Q8IPta0qx5PKrRlS278Z0hbpI4WVrGllo3ykKbBCutnPuhxtKg66lq+5+d7zt+OP
1uzSJjnewkqVYpqtlLCk/zZlTpSOOGo88PYUuAHptXI=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 7568 )
`pragma protect data_block
FUSgE7gjWmThM/FxT6zBrJxS69I44jDB5PQlDSB/BX7WJT4n8VRVV5uGkrhHIiBi
W5SIAmIr1BWFOp8FsRR53WL1vXCzN/IL8DGrFSUtQStq7y/VRjg7eA99bTtZ10ye
IEd0gLh4qw9hR2erHSZllgrsOU/dQH5GvcUPNKaDosAfkhqw0lo6PTzVKne6xkC2
mCyxtRikG9/ZM1wQ3B7c5lPqAPtjzhbhAH933cc5X2tP+yOR+AnOJqiTB+cMs+Sn
mXymTpSbcBdYS+VAXT9AUwCxoo3UFW6IHuwJFoMZWYEula5QuTZ1RtB7NBohQUPn
ChKoj5YA+u9x265PDPPfuKw+u5qfjq8UcQE1aN94E9Nq8+H7gmgnqVthZxUxK5NB
68NMXJlYdbev3SZhULhh5jTVek9s5GQI4+X4n6a5qs/P3G8rI3sHKqiQ0gdn5ZyY
hdozcZX3KqJV8DG4gm7EefXzl0H2IppeF1FgWvjXqlj2WWforvDRcEeiP1Zrt+DP
2vBe7Qsmt8ve+MJb58D8fP1buucbSN9lB5zMuX1ckHlX6s05Iy1tLU2KuvfZaAhh
yY+OYHkYep6ySt032YO8z2kNw+AxYVIqc0dphkvQnL1rRw3wHNwNP6ZNMcNTKIHe
U37JjRyds2dgr6Vx5qp43TrvvleZjZ3xDxi9vhGgk4VDXOQSQy2sB+Crhcy4Zyck
HgGjxQrdGEt+EPiUJRp3rEbJ98Epe7euFkw28a9bFo6I//+RLXUjgbIbElnUGPUj
aje8QduwVOhAnr5G3IDklJI/1vNu2i65cj3TJ1oDEbmFY7VP6MTtCqXyzItQyKdg
PHDzG+o47s2rhkvrxPqlVlx+Au7YKz+HcOHFdObyIslj3/E9EtA0A+2o66wJe50I
BWIp36nbtxEP1vWkNbA4KTh9WStiK7kzUe2Xxf8anCHRuhntxdyvpQHrw//K68vX
o2KFZYjYZThnWI20jOlcN4GsMK0dsd/SMs0Nux809l2uXbJr0lJhvDEjsoPHrNqp
ehrCAI54WMoTbzgJOgyxEMJfBKZ/0ZysoCXtf/ElyaXpYvUnl61ZOGmPiCH0Q0R/
y7IoeovXu+Si1LDftEcjBNS6a9S7LWNeVDJZ18sVRGFXvngxzabf8MKG6GjmDF2u
ldh67OLnERfmaoIwZvdrDrK96CFpCf2HgTGoUrYEgO8Z6qTSzQL9d9lIinNi9fSx
G/+NH+j5ezzFkvkYVxlH0qsdYkKItFTcyI6M5FZwjJ5YAKq0SMG1YwHWbakkhZ+x
ID2VU0d4rXR6hMHjtTm+tT7uSlLFdKdrQ67K1FaOW4YcboHNdaSin1WTDRrQYxW2
BnWSCPwQKFSfA7C49rKTXMiQzLj6vrZFFdJzbIgDBHWp4ud5awGYTpKm+EGWYuCM
YN5m8dBrY7+2U20ecJzfkFRJDSrFotmumfaIfxNct2AUATSxo0HWIzDICpClLi2d
Ju7amwRlOQ5mrwKWFBxs3eaDKRLQ841eHIHF5qQjswl+wWke3qNDP2gsNYqplsrH
IDXMSBMRQBD1fH/AmEPIpU9eSq4JuLt/bdMWTvKLthJ0IJodbnAcW6n46R/E6B68
EW4PJ2/3FZmul1KbABzMkvRe9gbrgdqFuBpuLwRT+YAYT2kVdLvfqLcd8juXf7rM
OWRrndMy9Lj8tSRRmwMMpUhHmbcMfp8UYadVMJSCqBzFQAZoOxOlNRKL1vXkAGPH
Awaizw4RhhGpLQ/opcSAdnLvUiNZF+CTp372DxI9ferpEWGe4U8Cs4vJQ45W+xAo
tUuIea+2CnjR/CiIICm7QiWQf252FM4pRbppjU4SYEL3uRCfRwIbSy/HTRIcYLXL
w5cGL6xIfX4RW1CrvcNthCu/hQQKF/Iembejmmz1ty7hT79AiNWpAK4XMcD9XJ+x
yLwagJz2a+iz1H96u83SbknhKd7HG+x28WS+oi1IwQEeIZVG0jnAllgHKQlaGlTL
zmL1C9OqnsK1awMWiTzfBJ5W/PjveWp7RxISPr2bk0ZhEuKlB3P1uVdoDE1+42AV
faLK5XA51b5cBh6NIzggjAO4FLLUWQX2dvpNqmCEX5Sfphh4ExgWXUbdB8nFbbDr
hyLf5fLkUZDECE0jlEXlZt5xNLSeY7rgE4dvuNEN7RvFzxTxgP6a0RrQIMpq7w5q
tJ6rh4ZlH84LLdYvc4GH7Pd87P+3YwLfO5CRcnAL4xQDLqbgiatdxBqJ0zbo4SGx
i16Jw2RFLqTdJknrs3wLCAN21vnznqdS0BGp7yY++utJrhqJAgKdKS9w5MT3Hivp
QqHdLwt0loJagd6vaIhHB7EmpjxDLpbZOG+iz08amgq81eTnKhmU54i8pcThq8fV
68eFjInT+CZLp37PeRrHBOszNvu37vAH26VcmxJjpZ5fS7N1uZQWk6BgtBxtudcU
Qnrnd8rOP4UDsHuReke8p6RCZYR7z5posTSM7S8zOA+NXsMGdSfU7Ex1HewivVtu
WHqkC/TmWd7BRxSz2ROHuHXDY736hB43y4uqNj1eibGzga4YkNSdkXtfKaZiKG7p
NdgxCkzaqfLnNO0xNbqyEs5/NuaRg4/g809S4yw9kj0a2ipoM229v1Jfv0Wixw33
EixC0jlaH/8qqBlb5Vv12130hjCWL68PUbMrX952GaW92RY8vgVudWXfsHy75RD0
pqN6iBcbGnxMUgljtgJYRrPyOX4ZHKHaSIOEa15uhFbUgV2mnhlefI81eg28+iIZ
pQoZXISYoaLYeIQGk7aDmwonB9zFo0Ew/ZCZpo/F0vlqcNgFDKZkvcs8hU3W0Ije
DhVj7d7Rbsk1oN4oJOKoA9LYWOmNNUr3gctmLRRzw8gTNTdZv74r9t3vkFG4XnO/
KbtIk3MEhmSDGDDjR8gMII3BclFuiPJd1D9MOWprqqPfIHrtsne4yTCNo/2ATNia
WkK4HfVu3jUTIe2cWOLG4a5w6hjLOkpjrHCsJ47hk4iljzVk8dE+syaJyHdz69Hi
BdCtd6I+DBB3BlDX6sOQcd65XuWi80pOaL071K6ZBbZ5dTtQ3RyFX1q8sDBdxDhT
lA9Q4oS11WkqMKxgsDsv0TWpM4j9xIgdRAv/ztx3qFZUHtUoI/7zkNBckKzOPcse
X3KgAONdE62u8iwUPhwmpXfJKQ7wGJv4C5jMsPrOrZ1VorE2c0rpVhZ1vBNFxg5B
NwJzdZ9limBGee8kNqqsHv4Jj1wR0yCL+A2mCUbdu9WdTL1TgOLq2l+jYp0qmhaj
36vT/sQKygYpqe82dfcWcPF786KdUcdFzB1ibKRMpC8AZPxvrpojZp4kn9rHztmv
FujDrc4OjSXSlj8nltG1XP4V9DcbhCcL/uwuPV+lDykYHgEhgIDxOJRYFxvV1cl2
byXnS4o0jOEhwM5qJb8sR1WUQTGlHUuGePgnpvPTuQaUnP6IJYy2uSpk9zhINVCd
UpzckIaNjSQ88Vnhupl13vn1fPNkBWKpCKob0yl2dyVxE9CHWgMvIRlFjCsfXEmV
wzprrBabZzWZ0DGWJ55f3NE9o0YAYMuDdXTSejhBb+9Gb5qqKJDqz9fNkaDJl4h8
+qk0OPbQLcAb5g6kdKr07/SXC13lG6zQK3vE2z61DgglBCMC4IWwuK469OMzhQWJ
/3AaXcq1bdTEZPKO2pVN4Wi+fh2Q58KbQeU7DBx+79+n7snEZaPzkvSm9vTr/HKE
4dKwz/sA/JipdXkOgr0WDjbnRX+NnZAaXkwqZfGIdax4t+14j4f95NJ3ykVu0R+J
yUzeI7OtUOjPY44LxerFaERHnMQK9JT906a6cNL6iF+M79PCAiYaCl+Wsy/hEOvx
NndCI/crHpWt9sCrLIyNcLY/r99OGtvJ5A3/YXqCOd3Idf/T/exYr1ijwpkrk40B
sKQU27nN8UwX7Kr6AyvURqZ9Si6UuP228feqmuIcvn1cr3p6XzlgQPdk323RLYgS
DuZzKpOhfHUzkmCPSlZX1lgu0fFqSAUaDw15FBFSy0OMQT2GJT0JibGzwr3KlEHS
HGTP7qGjd/X2fcc6otFMpYLqiAOliPxfmX2vetuVviIldd2jmlST15U0iySR4Ytr
/TkKzk+8opsVZpC2c+knTZuB1Ty6eM9xe+xjCinS3SvsD05GhFKf7Hh+qR5RwmLG
LAvuIQqu3DthTdZOdxZ2B2bG4HQ3Cg4DzlL+TYc9L5K1/fD7xi5uchyVd2LQt6cB
9k9KG4Ym7P1SzE4Nw7uK5vf7lPlunFtdR9YR8XapRt80b9Lxf0dy0xaL+rLV2pnV
wqffqpTDaaXUC1j8qamxC6wJs7FK2QJU8RfQgC+uuSxEf6AOFyyrY2cPUH0TCLS/
mffOMJdwHC5Yad2ODSsfTbV3pRX1fwMRKbUtcd82lRO4BGxPEz/aksYjMR4uRs3b
JYyUlxKAJxEn+PqgDSCwlIaKPEbXxfVijbLhIffuqt0JLqVG6xclyD6IYc4Hou18
XkB35GXWuPH5JYc6hqDxuaHchxvCSElUFYsIhAUw6wSp0dTh+FuQrYl/MyvXLrCJ
of1mb+nnvSO2fbvwKDNf9UU7wO6fyBJ1vStn0x4QuWpVI4YVDmVLjHH4ykWBptj7
NwvWRnjD9QtyY4e86yriTHUn6S9rDWljcwSkxIzDqiW5Q+lDw7ROSLPdGZK86meL
hTNXw00HwHYdIOVNt9T3K3ZKj6sTHANOSTQLiENFQ50rsx1zCMSQC5C1r0ZK1ETF
zIrBe+qOfqGjqSyYy7+1/cdlbs9A29Kk2l1QR+z6O5n17MbcaRa03Nk3yIAr5X3W
3efk+VszG51+518mPD/w9jpNtY8O0VrKiVYOIBXgbpbG+b3sY0qzAsWo2Xang60R
iukMsfj3/IMyPVYxSaVqPCB9AQIspXT1JkdQaScVoMkpZqK4w8U1XwH9qrgDIg0S
xBIV+LqEjkyzz72UrPOoOOMNqw9Zck+VcgtcSEdzVi5PrF/LJbY9fRrUZDMaV2M8
n0aXQ1DHToIRrmyHoZIykm94BHtMvJlzmf+1nz9sBq4kYLrY73U5U0HzwivnqVy8
7y/2qJYycwl0jI3XqGbs7n3lQXqgi3uiXEU2k3K/1nONfsSDzOWmRjRgdJbeT6cQ
D1quUJ1Qiq5QsoLHnjXp69utslmI1KNa0abFsZNf1ZqPpUjg1Rvw/ZFQVm0G6r1G
KoiWi4uVNFxUyP59lN7O3oRn2EoS0ACaaRGbcwvBJC7UZs2fEMRIDRlBtMzT5E7H
YF3EdDSh+1pKlhQFFuNznEWX6UaDAhwAR35hRzd0YRg5vtEcs91IoFPMwZjooaSM
XFSx22F252clAGXRd0sPiic4Kn9iI/a92epBk45hUXH6S38C0LtYHozgFgbw4vOb
Upklt+83wr9BzEzZTO8bTpHRfNh9zhGl895qTad1Snj9DtWba8qbu/NkcljsSqaA
SxSfOlZHoasyZ4mNP7mFOF86B9M5kMhi6pq47FyvH2RrIdHqeGFU73Sexh3eOhp/
UVIC49ZeCgOYzQRYQZfrEuKI/wWMzHeWZSZiHy4fG7m+GHosZdhZuG/bJEibQSNp
p/6RdACM5+v+vhuUJmPexCC+bda2dLjlQm2w8HJc9vMpeJWR1xS9NfzKohSZiqgd
D9Nu9zzKXoREj/vMvcoPEaTAijcp25jrficsdFotbOiCgLjn7iY5y7GrO2NRG5QF
xbGoTl+1/fKF+qj2EgsGiDA0oAMrxfV2NuNEY/K3ExWgM3WpzueTtebrJ+u+/aKl
2CEYuvvoYbxGKc4u2x7mOnB/nOJ3Wy4l6JTtjbseFaEVL35iajYVuz+o+S0IhkXr
qSwEXcxDURQyp2NuoLbQu6B3yl7uhm2GrE+a7HtYeR9VKrFqPFCkF3ZgA/3mvfz8
4o3KxChPVzdB0LkkmSKvEUT2M1ry0LVSH17pNiz9m4diG1GFUxdCLCsZ7gwqvArI
DFA3VVd2O29bKIg3aHbKxTahXChzON0nAM0V3lW0Y+ZvZdZkR7vP+tmWfy0Pkv3Y
6ebs+hP+aGEaMNvLOsbKRxI1B1Z+BVqvHBeqighxUJxegXX0P9P/nmlC3kh/uIM5
OtNpnztyZ0G+Sj/GVc6liEIJz+70uNGesRUa6YPvuaAYnKpjjVmsZ2C0Cs1m41YQ
F98uE4U4P88ho/J6n5TR9N4NpDoteRacR2MhslQJQR0eYX0hVH2AybOhpGnJ2xEQ
m9h8JmckD5aFdJRIv3TWemtoNoyZoFOB+N6Eq7GSKtBfHXx//kimun9xJWoB4g/6
gIvMhOsa1ZbTn/OYVEJiSxXuWh18uUM5AnZsv9vssstGc3t8fGtUT4N1Eucm291H
lBLfWNri2X4gi/SkPH/ZkeDBDjqY2jwGmzjECXBvFPgQJDUdHV45EeO+vH3P9fz5
435Eht0/fkZ3vwqlGTm7qmbaew5SIyh8PQKLjRYrjOQ4vPtzIsfFE48FiY5aJ5Fp
SJYd+7rLYTgmzQUiKaZaWa6FPVDNJZD90YqQJnhudyrUQRHF8Snwl3JNoclNRHUv
Vm0d8DPSfZxprFwG5uk+BDmEx7aHZAKcrulGIQPWFWalR2olKuNxjq5QrbZ+/uuE
krKufPle1BtNG5V5ZeFsVHdOJ4QR48upxzFgZ9J6Gu8Vgnww7hBEb0nMB30YhBPV
FQLYLD4t47kQN46klrHZSWfeDvNrfV07Wzse4Xeqd305iaka2TN/6C7sfk61Fds3
Zj28R7ozFzRlXdHDtq3PZfdtOER1uuyfaJ00AIEdAQDs3QzYK9K54wdBR97NlZqm
FcVBBeBDDW7y3nfWo9e8aEDlxMtul560XwmqKGCwMSZJbLCV4ANhTOiXrCxAjIUL
41GO65gYI3dPLhSxv+MGJVGLg8REiQ/NQiM3QTMUyWPAHlog5Fc3c9y0QOmgPU7I
Y8lov4aQimfCovpLES7Xt3laQ+tGJBJOseYzhx1yAkV8cxnJWexYlMd/ToWReFc/
qSBX+hCJTRPBhVQOzjTd6ITvmwuh5Wv8Hbqg1e9SK/lH7MGbDZ8YsuWb59mupj2M
+aH5nLLyPVZJWXfaaoii0ov9gwVyHZ8yb+XC7Hr00an6SwUkGGZ1/GSc3CMjcGwy
qxZ4KxKGecB4l8nhtWZEBZnpUoAFzLjGsTpAZRGJxQBJo+n5wWCU23Gu5wc1N74i
mVCUNfChSwoFILJHNjBgDRahiVNPnEnVU1L/dPUKLi66UZDjolymBtsjMFj1bWQM
K2ZXKlkRcQ3FOTDQHSOvPtHwCjTHcpNPqp98xPcRJS7QcUwc1kUjJMfvo4Rgrdgs
I2/3xXA92YhaNjwsL+rH+UojMTBTUSMhvm2JnqsNyyE7vT1otgtwKchee5lYGnky
oDI1WlJi/wop7D27IfnD6eAUuUMogdASCpY1lMuVohpphEc/KtaoEY28jzPnJ640
3xh5/1dzkuSP54ExQnx1xMkxzPRXfbKOJ5nc9ThWi2Ic2cRgjNQrsrzcwR9lHFhk
Ua28/dI6LeEMqcWX6x7xYLuOEY3rnySGYFPiLPfdutgbP437eqVM/PzL0HgLDfAB
7qdfo//11bUfwxAtBOyiMOSc26nm+UFEnK/Qswhc8wNU7ikvXFluYsJNlCQP7/hZ
hsNithWFlU71mRBONQRFOKqOmJ6SWtuyakyUhUB4B3lgf+t5DKLE7L2A+F2Bl7OO
P4XTisyV03+eZvlLwxqPGE5iswndIHQH3W9tpgD9oY30UAToczrLbwchjZPit+XU
Viw3LE6/00sD6xwGR4GDeN+ZbsnpzBD8igfnnI7i5RLY8Hc3xD3FdLUiAm6A5iOL
OaSF6uD8QZXeDKz3bAxnqEh5EEFf4fZoIWw2sapqr0ekOUD808Yxu0L1eOJVN7Vo
CDAeo5ugtjMUwjDbEPKgdpRiMjVOSkFksmMKIet9f9Sh1OaLxkWvVtCw4VOjyb/s
1mMuurY2VxYZqiQHQ8SJHxaxw/vJ990CK8WL/A2KZ2GNWet46ziJxFUAaYIaXwPo
6wbWw0Opfc0JXraAH9920mums03MxGJTnun1SikQl162H7VvQ9zhUCZ3CFh24uQT
j47rX7upLIXIxePbNBvi0YzpFWihyqtJF4kV239kCux2fYjecHrxoEU1JSJ/xBvO
mDIZpJqvawaLwxhGHavChTwyzkLbqFRoQN5IGckyUvz6sbxyuSfwFArYDEEBrWk3
DBZgoTyCFNCJ5nJWSRFD0X113M2WKzJ3dZVsGOdLH8Ivm3FMVv9cXEkJgX4B39kq
zcXBxy6e9/t2A03AUDGRl6QJg9k0sxji/JF1t1OqcFEPB7r21q49ZthjxNGco3aw
1kxuElsAZzfKO7cu+l22xXf2z7iMO84VDQhckTQB7o8yD52C/xdjKTA0Wm1B87et
VrCQSJYEx9sXqkHJOSKSxxXI6OB8G8IQGVMOV96sPVdKf3PX+HMjwCjo35m3aEOe
/a1PTzBQXyGGoDcI5QT4yv1oTIT5czq/+wSMjyKIdQL9Nm+g29ZEXQVKvyr+NgK4
zVEZ0H0VztYshmUFtNPA9bsc9qnTzwbSztwdkEwGGClAbrhn2JbdE0JMcxKw4yUu
bLvF2+5yEG2xgjkTUh8Suii8GxFCUQ3+qg24xkRUxIrNU5F0FH/NfBCQrBwskG+P
0jkknT8715i4AWpxUqc0MQ2Fgry9//Q1+zrBzJhOcN45KZvLEQEsaB9Vn3buwbbP
tfNzcOBWZhkjCQuVU8L34kb7UBIjXMl6tzfNvaz0ly1vHsxqoGwfanWNr7XyFJCa
wGZFHFp3/ItOw7IFFMbdGdzs1PLHK/eDlzo58pBnliK8BAr1tF/ntABBfKPlSfUk
xFXivFkQWNFTiCqD+Ly4YdUXdFZwikfc7aGJfsPqm8YNPqVr9+dBP99avjcGAg9P
VNAtmEbfqBv6kkwYBPXlPLPRAqO9tvYbhW8aiaw6IdSZO/mPfG0RlpcIEl3DoDWE
CguUwthveyw53lxHydRo1F0W1xjZYougaz9Y7MvNUqhBdqHqCI2MYYfx6EJs/dat
m6klhrtSsef0ExnYY2rDz2iJxxpAU+x3HEQPOhR9suNP9a12OLbRQkbhWQ4K7GyA
hpMEYgEnG11BZUKnQlMF2mD050Z8/vn3LZBAP5UN/ULT4WIbZXeDSV/r23qrlFEj
iPI1eXvTGxkbv0U9GmEdXxMcQ7+HMSSNULapQPXLZnlPwWmYGh6Aa+PziLgh0/YZ
O5cogS5VtchVrJxXh/3ZxYdX6tgJnvyGUuejl+yXPYloO09r8gWObJJ+CWpi3uBI
3WIwzDONtgSx3o+RMcLpjEjNC58ZlfZ4/NRB+8sf/b+W3HH8tMkd5pKl0ydbBAem
nVxz0MKxgwJ+lIbIVrK1VbnrEbykW0wF99bNdWkoijhtrcyw5MK84AAquC0DSFXi
DXZ3lpU2p2gKQn5enK+3CtQBzjd19fAmIEDnEubCeitWx+xmIMAXymhlGcsJa4fH
cjM3WEjjbynLHlAklvHfD6yHY+HjG5gUGEh8836Nt91h3G/UbegPLB2efRJnsMi5
CCan3l66ZiQiAFP+H3nSyFOanwsEaLZtL8Rj3EG3SVabkMyKf9LtIf4wxv1ULqEI
wAHIqLAG94sz9b2/hM/ohacUsN4qT/ieQ3CYDMi1z77ahyEPkzX7vEg2FvsEjXZj
COBjbrTfE4hn80GGqJ44yKgqeaSwil6pPQSP8Y/6F1+dO/QOBs+Lw9Mmed+55DWu
VZU7FCJleVqx5duiNJIzMuNkqfik0FS7Ov74OuroGYjrwwPxEehLjh9H8qGNLrBo
6B8UbVc79WwDaNwDcai2E2KVNqKDikg6sInncFR4Om/Wwl/DtqkIwL2LfkxRBvTY
8jVX1FWyKK4aG6o+3gX/JGU07qjU08+C1mC3qwk6LdCXWPmjBp6CyVLNiHa6cTMv
5j5ucqf/lN4OndakOrTcTFAApebtPWKGntCR1+rlJ2zgJ0pEnIfF4gcTrnqz0fzt
v3+o8GQAc1/RJQJiuDoyeU+FoxdSmZ6FDk9AT62oN7dsaoONgDV+S3F4cYU4/Cy+
ECzwMXtCDKgTLJfszUr2sLeR3rLwXoaQC4JgtGcsBk8=

`pragma protect end_protected

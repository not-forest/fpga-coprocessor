`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FM9Lq5pTwa16vWtIn5rRz3+kfsIiIF5UL3HnZ9F8z8iPf1QnJf3Di9AiP/RHFO7H
Q6m2+YrRijS2IoX24Pvcu1NSDAZl8i9hoZgUcb0gn0mG8PqXJCrE53xm22p0dgzL
tDcNzykIVpi9EBs4JVOesVIpFy0wZvdzPNZuC4GKJ+o=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12128)
ch4hXm617RS+HvUH6HuXCTKoEhUPbfJRU/CKc9tjNjFvOf7BCokNvFeJ3fQvnUhv
Jk5sxx3+K7/6okiC3xe0xuaH3VK+sm1YWfIhUH4M+bqdCYpwYeM/FsPmQfkRtqvJ
+lPnp95Dmfx73EGNJ5l1llmpn9R33uFaDTApa6S7acECIO5HaAsuieUEc+bOKI8U
42ox4l5Y/tToXJIylidgGWvnV3PGQ+4VFDe0q2ma0D4gamosIliI2h4pReD+gWAq
u/6oIg9/Dn/ZnyChwLZMA17J0GRAvvskPkB10rYucbdLVkQ0LFMm+53LkdgR9twN
0pNm7/nbC/YWdLoRmBqEfnFjfFWbKOPKZhm6FQkXZ2An1Bh5Elaft7x2CwH07AzA
xP8nbZ8q6Ln6qdLU59c0dv9dVsn1tjSlmKwMB2PWUE8jK62LYYDmXk8tC1/JFX9p
8QInqnh6NQmE9dusMscuFSsCiNl/psqFpWHW2GMnNw3OuWFuqnZke4GgaNI1pp8w
b4ZtE5aI8LcQgYgppHRmwEUTjiRGTVvgw92NkIaTslo78ktnkdEfZnXVs1Oxw+P1
y9rILqGPa0CKwSg6z5DdwUZtCD1NUURRFZvxW0b8L2I8I20xG0JhD9UphCb4FO/S
028illi5lZ/vnhhtyANo99m52+hyh6SnNA636rnZW8G9o0XJ8Miz6Se48ysZAznt
K4O3NITTHxGKsBfxx28iih5bSneUI3bkkn9klIO+0HL9BVnguhz0kIeZb5vY9GhH
Qi704P5azAOoHXaNOdY9c+jWwwc4IhkDJHbn/Nw31LxNOtzDKLfP27fdsk53pDbg
p5L/RV7Jr8LnrdZ+dgDyy6+WjI8ww3+IFDKzAfLODKkxqSCxLUtwj2hcVyiUf8lR
ztWRCuSFP3CILBkdDwbkzx0AQOIPGUOWXo7Hg1rL+lrSorttAizbMkHfQLNhODl+
tdCRCi8AesHMGSqzS5KTWjejZV344oLUYBIcgbNuiZtuyAGivkzFI4jhsxxYFNzh
F8QX3yUVKEhfsCaPZLuERnfyt480tZwyKZ8JQo2BpjUk4iCZZMTRUAe5ncxJpALp
cK3xRNfpyyXntcgYiGuUmZOmmGIkgQvEDFE0T2L673DX8qW2NB6uHyhJfrlvEXur
jrwU3iEc6GeFo1HjdCfksDBd7eEocJ8EJ6Cj3sKGi9n6PIxPYnFR9XUQuNDdCZXO
/n3zrfvTwoB5DkK6yzoVSY2W/hoEQOdbBu3Aocp9uMhnU9iH2qdvht3opFQhSb5J
PDklsLbCILNOU4PA92/yvfITaCwEWFARQ3WZ58/QBo8R9QwZokK4PBHpSYBepkwB
dwigl/EJDa2S7eZk2+zXoxfH5l8462o6HuGo0SKKQDOev5gIYiUrBazdQISS74gR
3YCuPwbXlAHKnA5GkFW6l63oGZW48OQpcuJK5xOk+S3bdrfmICsbDTzBvOB3GqbF
Iv1k8B9i/XrrnD0b2m1QbInSVn8tQY9Bh2cuEZ2TRqmoD9I79Z0Zw7H6nIvA8xU/
tEuW19sVDYRUnXd0sUr5dNQdLis18eVUHF+n+qru2Obu+7j2aX0OHOeiYKnOMN75
nNh6FYRcJdzub11o/c2HpW1MK2dN1DKs/43kefsam5mbOFw2MT57HmB1RBIwfeI1
pA/QtjCb2WZI1+DI3/62syZhbDf2DTfxDlV7wZ8sX9PN4o3vhvD7RLkqxLSsOOPj
qNotcX3JtiKUCnoNQvMkAJx57/7dzxr1uUt3oKE5KJ/EfhA360TU7I0ywo6DEuIa
0T88SG50Xz3krFAkOVbYH5VcvWAjweRdXbpQjHsOqbQyh/ZqwDb5eoDwxwVQ6/pC
OkBpQRsUr8R4JnqIp7keKyv8b4oHo8TO1yBKMg7uyCFhNqS5zXy3H4O01ZRb/v1U
3lcO4CUbdaip2/Kc5tN6/2H07KyxUamUufzyBkgOhKi4UNGDBrljjqWjGxETWw1t
BwrdZUag1dCcORX/489pnK8Tbm6XvpnKq4Ya2eP/n+UvHSfGFVPjl4YT8KS+jumQ
6uA+JvxRODunIalmXrdh2ehzP9Wy11cbs9VIlUiWreTm5SFs4qSLLXI1ptlHdSpi
zcOAt/EoO+kpUuK2jI/qK+cdRjJ3dTOMsP1RPNI6Cy3RVaxAM61fE3b0NUqqY+jp
EqVA9Kp6wiZCVgqeG7S8Uflj+CpPSTEFQQ/7esGw2tp2778eCLKDM+QyNzz7OLd+
X4zjnSNsw8982R4Cvx0N791Jfhe3kAAzAM9ld6QaPJzldMQsJlI0SIyNr4c7L+C3
p42hvoi0zDlGCh3sAJ7ugzkzZcjMKPXlnYhNLamJ0srjWglGUu6A91PxJ+tCmy3f
ACSQFWm7fpSEGiXe4tk37+iZy0BQPtWoXmlxHmiAuLUb1F6PGs6jvqyJ95ceohtO
pI/PxeorDRNMQeXPQ/KuiZSMacRgljtREBHGWkAvgLWNznnNAqefozGkhGYzIcUx
PYlyW/63J8GeFqsiWFuURiJG691W5oYAi8oiVGW5kEUatoXb1yXsnauBv/VQ1EcU
IAcsRYvj4QIp/XjlPDVf2PnyHM6OR4JbEbIH88bgqa/GKW44ACMflB1/kqhEIj03
HVrlGklwEslL5MILfg5Y7nLwes18xUmFqkSnx08ip5aUEwBR72gAC3ClRS8PyQl5
aYMjtmFge+2AsTsEH+Zf5FLeugWeoDLU5msV6+0VoBqV0WFXp1sDTjVy/s6M9Nqk
+rmV+e4qxDiXjhxLx6EPhjZQWx6CHd7d1QYXlZ/R1Wv0rkDnmGLRKUQwWUGvJ4jZ
VuygjxSrNtR8ip8/1Hg/gRKbeqtj5NHcvogIWxAHsi+45+UKYqS8Fz1H8g4aVjQL
65cJxhCmwpbsfy9WheoLnhD+p1n2A/iXSVX9dLnoLjDlbuSo7/tpUpmaTMfVHAch
OAKlaOR/5X3KZQRvTlj/3CrulXRASdwNT2LypUc6Fs4XEMsYQepuP0vOQzmh/Nf2
9iAzTmkNPQyMe3MV7NbNHgUevpYeDr7ZLmSmOiblX1P22sVskfcwdZVyefw3KC2w
lT37krDUBHLUg3OssxCwgaAJ9zsx0nNflaWS0l5WNECyyPiyVIQO+nRpzV8uMZCh
9gkXLuuYeTrSvlJu8ZpoU7rpSNobWwNK+nmPJUItvhkMDhFVzZLcep3XQMyGL6uq
a9bWm5cn8r7nBOMFOssWkfDCcjAARxh7ucLkXdlgJPqQYpmSeBtnu0TZNXCk9Cow
reEm1kF2EVYGEjwuZQMtTvguQn5dGofgArpU8vMwqQW2LJNZta/OKG8UAViCv3LT
3CCW1+WM8d6n1JxKfCXTvj0Z3WFRLh4GpzZgtgCXHLlLxtJspskxH6NlM107wm5b
4Yz86grbEN7v0vIvrBY/GkG2GxqGpox8HvF6E5u/BrHj73P8QUwbFgd31XP69VGE
wH/0+CPN0+cp3R1M+ynWdnBHa3hlwTL99oTe1SvZYVnqwXLdlSfw7/V6VBGN863T
hWY2VXYUEcstV7rPV7kkfCZeVCvikwRLwR2zJIseEs5nKmaD5/dwkjEO7zUQ3Od/
8DJXIaGpwfu10IvLeIOpXmNzQHYTXSN/e1AthMnEvdrXKacwUHFUwo5VJFzl/L5/
u4aFmpe/p6Mx/O0/gnx2ZiDR6EnU51+wLmOXZlkmQ2804LPKANjJP94/P8FGt1R0
oJgVkeBQmlSw2X3rEt7cYEceSMMJ8EcD/wYcfXm9QQ81SrW5JFjsl94ppOBWa6qQ
SKUiRcA6745iQGqS4afWadqG/Xs+R0uyxAJZrKu4MHXxezmr5PnG95dRjygqO9MY
Bw6ka0H+Lo2YYIpSG1PrpZXLq+9Z0hqgbF/esoSMN7MOeHIvSPFodkNV0wufcGmA
WB7Reo08JavCZMcSfBrNrSvGfwmgS7Soz9ZKY86OsJFMTTw+HSJmERkzhuC52HPr
H6xmuFmwFdF/GEQmRKU9Cek7rXwwz473tgy4KtU2Me7tc4hVvY6t/BK4gnQGsJDm
I5w+dY/BKxZ2rnn963/oZGnKpVlmSlafPwMYn7W7cfYr8tn6BmycFn2tR6lC1QtS
NqBcp6zzQ0At20eI4pDtxZN+dFySWbgf6yC/LTvgzFimGi4vrIELwLtjMzBo6/5n
zOg5WgFklURi0GM0K/8lNdLyL0yws36iz8PP9IFDoq772DHXRo+tWgTCqJgNAMLW
12G4saYZZXiOE+vsAgCe9cMqtzL1N+BHSwdzUlKtm5BfDshqgVqa0itR10fJDuYD
Ulv8NPXj9CSe/bX7gY3BeKa91SYoV1cbkrP+nbQi7l5IeDMHVsFLwVF3A1+guMK/
o7S3Yt6h8nWyLKDnNFZPFnh43MVdZpLFKBh4Y0QMJRen2bf3KweK/kqi1MZBOXrs
J341RhI1ZdhVNC0y2cKQeK1NKM4k3lr7QxCN0nDXFqfEisYOcFCsYEqVRtwoKefL
H74qECemzSR73bljzZK+FNXM5v3ZnfgN90zktwa6YWb5NpuhrgUQc9dRzO7cUxtm
P+hpe1kbUNeGwA/gSnTQfaw6QKeIil9WM5h3wt8joUotEhUJY64xYhdrTNCAz648
GHm0oszZ3Ip82JWUetuSJB9PwUQXONzuqzZ3MvxsGkfqz20Sjyd5V7/BTugavt9N
Vl0H0dkcNxF4bXn2pSARPZQXRCU+X1yQIgylT15YbWvbIZZXCnNb329AnWUrSg/J
B0jnR3oFuAovuaUX8VeJuzk+GiXWcOvbJNj7cV8avDXjDqpB7X5ruKVZ/ov32kQE
uUqJziwDNaPXhJfx3Om4Bmx9CB2XhuUkvWkjtu9l6B89+XUBjbGtIXprMbfBHKVe
i7lvkROU/ASGw1T1SjIFz16aZSZ+SBl3m0nETQvgDjQaAd+NVi823FNNVl2DtSY0
m7SwJFw720ofBvFFuLGoxZxFGAQwdwd2rJFY2BlonWT1Fh4pDfJTXpkVaKPywwhE
kICPmBQejBbuHOZz2csU75She1RYcaJmOFhesaFNdg8M8DkG4XyCsIrgNjzzxyA8
e1dExdZwKZnsbVWEnM99vqqcJ9zeEs8mNSqNHsSnxlHShFNCPx39aHG6MrE+PI3z
RCoIQ9eGIMs6sq7gBUw1KpKA52Zn9/AVznx0GOp7F334h5TbBcNr3FwZx0whD/4D
+t6AqxE72d+dcK+u0/HOTBqbqAqj0dYgkGILTjPkZZdOlIAZdfI+Z7IbZSvOZmmR
rYBhZWaT9865XagrJE2BOEq1Cj/YKSItSkeKgaMTKkeT+kXkFH3BKFLhm6hVbtJf
Se4Lrp2rOKXAbDFxx+9FgoE+wJla3c3YfYxDPDOXXjR30X8U4Dt+FiZNbkH5iuTO
1DlYzFYgnhDBIVI6s19rikTKyh/aGXXuUKTm0jzGW3DLQ5O26P7HMlTI7MvDN+Gw
WBbyL60Omv2Lqi68fLrUmNsLVSV3wSmv8eM00H1izT1PSTyrWCRFG6B9TUzZMM7q
TTcv4yD+8pR2Xcr9WO94m9Jm4XREEKZIaCepesEMEnqauv9PLvim1bQ2F2LUj+JM
6swWwtKclc0QHJw6czuVY0nyBYN66K1kyJD1yEFU7uMhXkjW7QY10YmgleF6QX6W
TeLz6fTxs2MqkfFZcFoI4Pv6lpxM+fIAnraD+kAYA0VwJFqBwik1vD8etKHWW4Yk
bXMMrch8KfpbWIkDAORohyn6OAwNyY4DSRk90iPP5sn/dSRoChn2trE4gKreZTk6
m9jF7iJJH8akD7ELzbJGlPBdbp+Ub5oXS/norShbrkGNvssVcYyhkLnjsz3U/fke
tKE30ltVHLcIbrLF1mmNsLRWQd4xr4lAVo3HHykX3v5aiFWMFYSSWC3xB6XbV2OC
+uN5FHT+YgziirMRGqtRSxUHjvf0jijjvtua93GW6RobetqMxvFVlZS92QhenG4F
LQr3rjq+7rjEjiJZRCyo4qHfBprFzOQq/crEE7Ii6248eH5Fg4+sp6VF2B2A0gss
PZKWLW+RyLhDiYcG6NXMAxmuvaIRsHR9z2BUrg6xG4llLpnm89M0Fdwa3GOy4EI0
CbND9SpeG3/iiJNF57tGbHUFQRUY/Pt6GGhcoATbidcF6GtVXtdzYhNzdwIqAwXu
rRpHfYloYjVfzt8D+wQW7J/cfoMXjYq9BQRkJ/ItvPsbBr5dhhs6+joau/rw/Sgt
5JjuEQ66WBm1RHg9naxCvJ0O4HF2GuaN7kiLskFMSuez10xeTqHow+VMR4Egtdv/
qk+LTvmhxQAvwFpjpyqk2krKhIuNXFeL1RhmsSnBWyKtsoPNKwCeLiRgUZdqUm2L
FIYHcrUzpNaGIshV/G9b1MrcqOzF7mECuinuOeV7m8Xmo8+G8QtcYzT+qTU+tJoP
XPAdl2ps4Nj0SVhG9SiJ+QFZfUavvPDtr05qPz/ICa5dXDe1t9ckbNRTukiws8Td
2Xch8Hum8vypYlGsZ6l6jm6+tm8SMYaTuZRVFqus9O+YSUM7BVL+ObXWqoKXYDWB
jV3kr+D0U+KWLkEJcofb5C6QQL1vsIAZt7Ij6QpHExWYZHcf0N1Z7YB1MFicdgo5
6rkaS7FV62Jq8KFMwI+t22DLsIaLhfEqtNguufh2qBFyHufL69pSrCDxcKkJ8Mwz
IAjTuQIRbRSov3IyhnVrpQq3qJ0hRur9V9ke0BHeOFNpsasFwq7djCOQN9tHWeek
3JgqJTRjKIt7T1+zqiDLBWv25eb6bET9K4L/mK53n8aH3tR6svi828pudunA96ic
hX1y3ypDvocW1A9rVrgAknqfslin165RV3Gi7oYYnn8iNa5xjmVRlLQUHOgeTSFK
6GRw++bQDMms0NKcG9tmZnqF4J5ZSFEkHkPlxNaGP7YuDx+/B6SkLP5bNbWiI+BF
sGz/LCXNNGZ48iIczVKNRFH70TCP8jVnvL2K3mEfEyKnS1rkZQVxnxBshwss0W38
eGIzhPImFSbylKWVCueTvahAiuxgc/MtbxOeE+p4W+7iq1tQMXpDKtGQGaAhTCBm
52HLIAQCEcAzHBZTCkbgBpM2iijLy+d0F5pjBkgWGjjcc4M+CNYEs6ek74XFvxj9
353Z4vtQW/tqmISjJkG3dPnGILCb7rOduKxuEijwlIxSvrN2Rh4pLH2ybbds9Sjk
3ItLV+CWgVNHGWRhC3IpUmqMk+bA110nIDgHfwgc/Qtdo1zTofHzABhRs/ddVWtp
ISQ4vp8Op88qfhyeaXRSF7YJ4+iMi2XhaOdy3d7zzCB4PoJwxJ+xItiUTnRuFMjw
dgDm9CGksnBSCNsDtUqb/mmOBaJrnwxI4Oc4Pbd5iAelS/dBAEKH38ZhEaP7PnC7
vm6kY49dv3FIJC51VFgrdu4RiwbkVYRQUc2rRxtVNzqCwfpVxeu75ZYBgP0D9rCL
943iQY63s7YEuRYhM8Jatc0TSIaWN32F4nIh7nSTVok3irxWHPT+jGKtkoBFH54e
ZV3BeiR9DN3vu45KgbSoOjeNExs7isXzdxsM56MQ8LsO9kwU904wSupnRNKMtsxk
7QRjklO7fCu3TmbpTWBcd4i/jb8gYf08heZUfBvDjEb+iqb2Ir/zGQzbEQN5UuUG
GM5MVl9pzi+lzknUKI4YOSwKFyFtkbOBBY4iF9CnR9+KBsYaFhCGq7oGM3pautPq
WILrSdSlhNkk7+kGhpPd9ZUww+duY7Tvx77HaslV9RkFpLN5TWBEURKOciNWO910
8vS3UO2HK6coeU/ukNLInLc8V+30zLh0vSbFjKOErmQ8vnU0FFAVCcEEHgS5VdGr
iEMGlkj3X1q4kgzH79k8wLurVSuYcNj6cdoMBL6P/rUIIU3rsGdIGK5HPy9Lol8F
WTIN98RoqCTkfaoAbIfKH0QvZo389Zgv3SLIukomRlqX6n7nVLITKg85eANTQ+KD
L8h5gXETGD5jFlekrHbAvCes50gjwdlp0jR6P4HCqZ4crcvXFAtvta0EIrJPnwhD
m/DkDZUvA1qXTMaHCb23XHvrkQJ7NcFn/WBP0XZbj12ZHD0Ux6Jo7KZVbwa/fKCt
14R5zRDnYpBHTkeIRwS90DNmLovRtypdEz4yVC0fL9TGiyNzv79aRsWSnwkMGN1R
JnH5MVQNIXcOgXrCXADeJTGR5e5Z3vYAqHPbe41Gbu+WMTEdS4z/hQQuWu0ftxJx
QcWV6Sovv+gMvU9Xm0Hd4SUG8dWqLFg0rCTBX2LGXrjh7kAqt8FReWuF1z9YAEeC
CqRYiS5opOAJ3jt7B3kieYOiGc2AEyEX/Vt+hRGCHIfZMe79TCUr0fwXuArqEylz
KiL5vtyhaaJn1BExkiq6L7Oxm9SPYb5IsZHHLKRxzdkhdvaXEFIi+AQUZd1CJSYi
eQR0WoTp/mgdZqOPhvprzoQtsycYG67Kau+iJGQsWuI+zi5BdktIztITkXfCC4+4
qfVyz5EeKWYi73CbGk1B0sFrMxtMC++QewcHRrbvmSCStUSFO27LB51db3ZRqYnj
QPFEA7DZxC5jTs2UX5m4C+zwNhRVRYaZiiT7ITO7uhirDeDP4K4eyB8gBBE7PwEX
F64JMQiQ7/Uq4bdFbJ85cuilCYY6Floz8EOcGyH2p+n3LRNQEMbjM0DzUhadUgdF
CWsHn/OtNGJ3VaMhgLMGU34CB0zECqsPmL7Sx8cV7JRWdTEMhzIqj+6pdVOZAjlJ
bNTAyyCUXLDpv99omRA5uw/RO7k0GKf0/GKNUrWWhrS3jL24AG/mSpIXeImM/yiG
/aPCwqqcQozEQxuvV25F1/s3DR1fAKFe18W7SCb5k4Elvjcb6x8bMJ4RxOwDEHiM
8RemxOO2GfvNPLIZkU6s/7qAJvn1Ve3L7zLUAxjnw9rCwRJPgNr9PjOxG3RhY8sJ
GXAu8qHr3MMbDcMcST9mQIrI0Ov0jnqrGDH/NKetDW7ZnnmDnkB7t7uYy9YkMCP3
R5vIRZ63ManTrT1ca/H+s2oe7JUvRWvuQdb+4POl5l6wwHFDCfIRxdVFDyQmz4nb
MGo1q1/17ndEwjdu+q+KHLMuyJj7mgYpcWy0loTXRHr9bX0aVV9rsZG7UxNQz8g4
sUn832aCcWpJeBdj74kv2wa/WPULGkIVAC8ERgk1vGacprVo5AmDtfNas4KoKoZZ
fZNAebGGVxrSXeJ7ahEqIzJ0ZnPTqLoLf7PnTlZtjMORWlA656ZCTX9odCZ+RUCo
5vLiMrXf4al/XQswuVQsMcryq7OQW3r9iLHpgWj56Wn/udbjSWFWU3Y5D5BCW3DL
oO6jOVzaSXMTzSSDfPi9p25rkdGEZI6BaI2B/eYxlTOkpvqYb8JW2lPSKchd/R6I
jj8ExYBPFoJgQhwpppVofALkheOFAsAN5ZCbhnchM3lDwjk0ctGAxLD4ZraCVKz9
7+UdwiksUbcMgcbdINCQ6TKv+o7kKeL6rOEn+PKOqNRCWhDSGZarBTAR7nTxjqcg
A80emmbAxN9fPxvKPbNy0H6ytVXV4ILpLk0rlO236h42TzHsRx6KyLxoZMPbED41
lOS+XbijrZeisTYYDiZzhEVTI3CHQBhgLUlqSIJFUmNr2WEXqQAI+XseA4jHP5Tb
vI1Pu+4ChmGOEC2yOM/1/b1ONCwd7dk7it3CRN7bKczvp8ZbWq3n+toiyixnowha
i0AU6r+5M5cuq647aLDkC1vnzdRQmwUCFESFBDtcncVOr++dR/ZBrwWm4aRMgXxZ
S2d3/nTWDz2x4/h7Zh4a6s1TWkOAOX2DzwMQ6ahyS0lT6vkIbqafhVjCeukIYvE3
Q+YA52ovom3AVS1tiK7rdqhtVE86vEv0zv+l7lWv54s6vWSlYyqaOtMeZnX608nO
Wz3tE4xRVdCM7zMUtGCYag+rX/K4oprG6dn0d9+/d3tE0WjB9t0NjRL7uTE9+azJ
11fW0jcmDHa4ZckXoD25SjECP/Qx06fWhDHQPffTzpzktRdoMfhTwhaI5LFvc7rN
PqFY+ei2qp0rqZi9/EirB+ON58lAw3SCmXSQuvLF/MDNQqFyoD+Ylh1dkdIPbZED
mVIboHoC5kekk0Jie7iMafV2CvTXeaG1EoRIiNbxZx5sMCfzaJaAZgN9e/24eC6n
PKoRk+YRw4B4dv7MIi6Dqpj19vkHk542Z7kafMwVKVMCzzHzLrkL2OiGWikwFz30
SA391OZP7YVpocOOn+F9bPfxUx2+cFaHPZd2MPPqnYE7v+vtH2+kJERjcoLqEq8K
wPGAp46xQAT9tN0UBsIRDljdRiX1MiuOD9DCnkqttf0Z7NJeNXiNQAls50wYUFm9
yLDFEXWi1oF6vLKbh8UgVoCDAW7nUKEop0NCf/lO8Tx56U6HB2OyBALZDyjhBPRm
vpHEdsiC5jHZq52i7vuvVgzvkElWQqaskoItjhEzFUWoAjWhw/asNp3ojUfErO0U
Aq4oUefLFhdVKwIVq/R4vJxw40X/YUPdBM1+/MoVN3P+f6QwVOcmQN7OFs2a4Qr2
oiMUw7rg+Y5soGdqYuNYl7AyV0A0NVvRGQu3Vgo5k1izslZUaAYS+83tavsN9oKY
sHC/nd9+nLQuGjeNvY+qyqS39wQsHWDlGIcK1SraIFD2WvdhYAPHj0LO0oDyygHW
WzG6v7xo/ucrpt0faKmCr5uWDGe3ShMYJEfiH+pwkiJ+VcIPJYRQ+ut0iuA38Iau
u4qxFqGsyCz56DyrT0E6nvBc7XZkrUeH8QMM5ARIO17QCfjZi+iDaVcEbyTVddmq
bwMMb5vEOSohv+ErotRbJZvVsBODFNW+jpGzXFpmvVEVJ+teKXEV4ydSZHM7IF3g
OQkQwbCSIgnLrkwgmLifrjQ/bwhbh04cItZGhZIEx0ySVwdS0t3hG5VLMki5t2Ye
VMh/iHPA7M+mf56GnuChDFvTtu0kX0Kh7NtIB92Ge0ABj8w38aYwfRgNEwEbWWcv
KvhV5V1QMchV283EgSJhX9UZwY1qYZhbJLl+rN0HlAHtZgElqyLB4hVBJUREVIkc
glNmkmHn6R79LFszz9CMBLiUdByIqmlEcUPTaaq0l4gnect3LK/1UhJ9KKzlbxFu
uon+V6UwKdiwoSAlH1F21wiOIeWddOM1cfQhMRMGr0xkaSo7YRhsT52WytWKLHJv
OrOt5t5jULHAkMI6ru4efW9iael7KK/k6vlxj0vIitDW5Mij3MiJZb7ChlSp2U7o
tyyU2/Gpx7BBWXKk3kJtIwxRXkzrbkfRFBg5uCKHWvmUzzz9DUsi6zSJcPW3erZa
w8IOtxxvyXNqdp8nNNr+IzQ9Eu35MjaD9XW6diBA0phsOtzteewrm7V+XvuAp2Cw
5XkXnFITGvpQTNVTX75mGHbhPgurTf3NBFaPvZAOP2royAvcsx+OQVDST6cveelC
PA7aOmBCpVkahVH2YiMXOWWbLq7FVIYk7CF2E64uG0p5uCoBZrtuALUeSdO/2lcL
6Vsb5R5tegxNhZncmK9CT04Sp1RaDhsxMNFZq9tsVA1Tw9ULTBJ4Vcvh5eqLRiz1
MK9DNRjBxDsmLMJx9yvmFm02Zx56aSfyAg3w5aK1B6u4RBkrPXJvy/IHLvKw1eoA
/qQkHduSz5HhZkWaX5jopVR9+PbC/MVlUb63q96mP+OnfFGxyc5h6/7DTs/TWskD
owoHZJLvXJgXv2eHYS/aSYESEQWEbFBbh0YPuRISQK26Omugj/cWOafGwWwF1u7o
RDZ81vSU+yFOUSk5wjrtSBrTbsOfw7wcPwAgy8R0N+uRpOE5Kx3y1+tnw0XIBdK+
HBZXxlkT4r43QdOWZOI+PcZ1I0ZykoLu+mqoNuo1QzWx3GQ2hOMHTAKM+4FDopm/
WZRLlQFL0v6isF+0cyLrzlt8Dletii6p/6UKYUvmwQqdDRo99TOPpO3saaALfWWG
5O15IuMBMTblUXCLzWrWRSl08Oh6UDTl9xj4qYqyU4AmCt1iz/AvhHtF+dM3XUzN
GhEo+/tNwMNYkDNv3dpoCIx2oLtOS5imtQu49omHlETnCVyVJagmLlUNAQsyl4Cz
/ARhePvdTkXcmhLXAOoWtnEAnWVTh1FrljONCwAW2njmGOYbKVqO0rnGp8GNeDO6
yBQzPvfLf6foTfoq0gHQghPMyW+6MVIeB97ywnRrLBYhkXGFwlU2wgFBgWtSI4n7
4EKdsiYOBkMDs8C5iIABLZ4HCMx2gvKDkzvBoIK7Ux3Nwxicl/cC8ZMkEtt1PY3S
7hnO9DjcUa/MVpUnSVoZOqCVPC6G9cgL3PJfLeRRI1nnRLzHXff30UJcFFUNxdKu
SBgIpNo+i4DfAt2923OTXi1nkxHTxDTDdo77QBr3I0TN65d3NbhKHu0QWcZew09E
pokHLizw/l1AIuy5BVOAEuxkjfwbbAZv9QNPbMcxMexQGUUzOcKW5oEAoDenuNsL
k0eEs0b5WQKLaOSiEPrjhVv/bwi4J7dDhfmCcYTXPdy4DLjQjdbMs72NTE39Nmb+
lV9PsLHX2Eqwq6ZHwq6kJ2gXC1HK3/+gnDSYA4QsUHKdH78rTCMSJuTbXZhh6Khp
x0zcvpp8BplAQ8U02jt5gynLV0kSfTDLV3717lDWLvnbfWVMrFJv0lpwia+frWdX
8Knff691BIeZ6/eP4Z9Jh7aEfcUm57PrPWJh9Nya8xP1pSrMVaZOOrbAQFL8IUNC
JDnYjs96uvbjhSBZVg/e+79I4IhP5yz3MNqCmcwl6o/uoo14FF0ejWKzqqfTm8eQ
z5Rr38Cb0tvGVpiLVymcnDH24lHMTsjqiqHvbKQ1OnQ/3ebAGFOAj0p4lEVXpLZF
F2cwVDQwNSiHRUess7yL2/RmUdrC0mwqeGr1xY6Pd2dlknKY0nJmG8DKathP3W3O
bOia2QzU4k71aapMB7Uwftz+kTTYlb5xwQ7UqTrM8N/W2thJ7T3dCSAGyKdqyK1x
lFQv+quVCcXJbScBY6ilVJYG5FPU0M9iq+R/YISn9L4J/tR0jQ/hAtmgnQelqF2h
16tHJeRLnicS5CdSMGUBCHM/QGPmojLE4Fy/h/8p2z14yPEEhaXPNCk+RHXrogv9
oMl3qzKPv3DhlXEktbkGhgijfF3JlrubGJufwmzHsDlL7+RAYVh7ADzpv969c4IL
+y0fj8MHeLINaDomfxtDYrh7uggDxG8lNDuotfzMrZtiUJIKS4CHt8GQFFJ1n6Ma
lD5NvIBOfGV+bTDJ3AhZz7uZIwHJon0NLIAWUa2fpfJ20nQS4W6/PZREEB/e+XAU
E9VWGx4Rb+ZY88G1g/NTiDWe1qjwe9cKN8aEXEfr7IHKOPEo5pP3qt05Zw0Ryx23
Y8gqs5skPjz1qhxhbNtbvgwgtesC6tQjVkEqRDCIQZE8+U/PHHGJyTBJN9ILxoax
L4+dBB/q8qQMYCL9w+1ihXMwc/jtlyamvO6g13NiHczS+2uSYbquh0fqHuXuTGMG
lBJXllzPi5CoqQfaQPcR4ehgG07/gWdaH0zNVcUwWPAAgq87hlhY9XR5VZYAI5n9
1Ae+MGROYcgH4Jvbyx5sT+kOWrsg8+b1WOHC4G5XN8ZQHY5BbvKL5lsEZjybVx4r
glCSZli9FLs6Oh9WAwVV6+q89on7l1bl59YhjwRWOFge1BtD0rk0agSphxJ2puER
4YaCXT8Alfpx6H18HbghEem6PohCjD0N053FIza52sZIBqAiXgqgypwWMxhmtYvu
QL+Y2hX+15Ypc1vm2vAS3cYYfw+9ooJOktvtcsyDamfijFiINxtwbaZDlrnUSR4F
FjNa/G8oUOwIjIcxZR2Fk5i+ZWpamMz8XIyTXdjEP+1YdvPbTGvMC9ZOXUyaGw/H
uL3DQWqLZOpLb7dmrHPDnDfTuKZqHLkV1EjMq+l+XWTGtilFDxgsR+WPjFCfs/xh
eM+d3KyoC7L+4kaopgzECjJ2+Ew+LzTvklq8z0FAE1OLQBG4diHixwvoWjPkPOxZ
10H8DJtUoi6gpmuiRUT5Hyhmznv/PC5wb9S2ZP+1gd0GjOYdoBWNK81DW6RJc+XN
yxiyUL/EEwn+AFUMZzr3wpmBzNafOkl7PLsDeg3XYAcQ66SnJpQHzvyEgZjQwzx8
8WSToH1GJn2aS/as6WLJHUlH8Fy9XG3YtfgTPNzf9E8Zy2DJ9eAgihWXksstmzho
O9LGPPDZegivtobmvRC/rXDSvQFtojj44FKKC2dwQDbHAabuPOq087kxpT690EKC
sMqENZFQlYUA3GeEKMk53Ds9wUtRBjczd+tqAnNRaUt7uYHYwGPqA9I7Cf8b/XHi
RfnyeOmcS5J3A6bMW+l/M2eXQF88Y1e+zsGLQyUZ7mIKAvmn6fCoNtx+L/MWeFDX
qN74wGQW8FE10ZhEjPJASic2G5YrpPTSiIlKykSKIC5rujkUNknXJrYEZhFhQkeU
WT1go0o6ipmUemgeqLUhIIVIP8ycV4bLfwGY+ET3kwJCSVfWqEfnfxrrklz/EKgZ
c8fMSBn1yyALyP0TYDpOR/20lCZ3ZrfILagDGd8A4uRiaPDXB2E6dfs5IUZ5Ug67
4LLGauNWydKCjKBL+V2KZoMFwNs3dN+FeSQ41EtA54lr2yntzMs/76FoQ8wldM5V
6NGCECC3GiydJGgJwJkdKU6BcEvBONW2nzUzeb2TS6qAo6inXiEx7UcBlwbbOozw
KH7sXaK29nF0aBLfsGrGbeNYWCxs4eUa8BTX5EtYlXkxsTohzLnuFok9pOWt2kTI
ggY2bAicRHkPfqHuOqS2MHp2HdiJiH7B0Ha3cxDc4CcOKvBCEiuGfaGoX5K4fwk1
jnbRsf0+14V7heG2EE0LSL2UCMxn16R1z20ed42ism0QMCpMJKRnZ9nVaaNqlXyT
w+1fNwDcXBqzQJHTw3+MZL9TCw7oDcZYB+P1JStR40fhGgUxvXBh2SpYfwhlByuj
DZMgPa+xFBTFfkUh/EN2p03pcKoqNPJq4vd7m7pV076KLVi9QzRSDoJLEjedNbUB
hsq4NL3QzdxwuxALkBGZ+4YuNUqgjCsFn3S510Sd5/znpBrf6Jn59N/gGESoTXUL
Nk486xGFWyOMbb205H6mG3sxkROZaGtdYzq1HKX75cZkYB3eULLJLS5Ujod9braN
Uiphsr31wt5Me0Z1WVNDaIOW/H1eWAnJ0w89uJVABTeUaZ9Fc5NFW5TJnZ77yoH9
lrUapNY9uJU2bfEbJdRAHq4AlR/godkg5CXHnRikX5ckrfRs55xovdGYHsVPgwPM
Ml30HwD1uIOFk4SpZx61knNXV/NRvUSc9IUBur1VeaFeACtVW1L0N2IdqRBG+vHM
Oev6mIhbFjaInOZwoth8xMpMhpPlY/xQ9t7ibtJOLmgQB17YjEJKZi7fqpn/S967
bHuRa17XiBUGBkRaTKw4oS3PyakhhMIOEOtzWXUTr2FPFVeeMZtZf3OzZhzA5BbN
WWzT4fF+or/WZILRIOnZ9FVoqrb8CCUcwcK+lxVTYiH34OzuIdyN6mHCxGJtiYyl
Z0IBvH9NFkTDW1tPAPHGM+VNtIUdVflNQseoO1VDkbAE5tTWjJGXPLW2DPMTD/yf
a60WdnIOLYQJ4377vkzdfKPN7jZ28u07EBmS52lsxnX87cMku2t5HIhNBJBpyag3
fwPEB8mWPn5a8VR1J+Nquk8FZJ9yhA3RFumgHwjKJ6j/LGuKKN1bIngKqrjTQSbu
ifAeVTIU9EeRlWQgMhxWanvN5U+z25k2gBergv+MkiPDabqYrfelmvdXNS14H3EQ
Xk/EwFRacDAMQvb0fzgk9rf48RbZFL0r1hQ//bb8T9oo+sFppuSyLJgJF5G8eQtK
2E8DYAIMG/bIVAr7Y+nMCydoelaxfqhMMJDBR+aHG7gAQYzXBwARYOLiOObaRnD9
qLhRE7Q+eKI/bUfFzmTGmngtM1DjFEShgTsLA49UW4p5CM7B6UKBAbFs3xLfSzVX
7bAF0TmQIYNlOkZHpUnybxCI0LH/jKp54iajLygUubpekscOy769SLpEb+BoxFMp
pcDH3vKpTIuDc0PIc4AGeI5Uzjwi0LkemouNE7UVx9/7KNnhfGtSJ4Nt8+GMytv7
HVKm9wPA+Ca+QtHhZ7W5+vTytzSo6r57EuRlhOpwkWj7llUr315X3PwxcHnf3Nc3
4YzFrigejCSb2P0S/LjVYRQQix9pmub6Ths5Mhsx174=
`pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Cb54eceGaWVDjvAnMn4TgonBLqf5hQ+uXg3ZhN8JNWhvKCEuQ2OD/s8dFQOowMJx
6AB9Jhq27RcNqdLxN7J4p6BquVc91G3BUm86k9hMUej3AzYfy6Rli/FVl029OiGE
WI1ar28qs6AX6q6MzI9MJLL+XR7hliXvATQiSM+JjV8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5072)
mZKZ8W4/s8gowpZMZ+T6HRiKYJVKVjgqyVuh3DXRNLUiyvWVbqRl4Wlry21i+7UY
WwYHF6EBcadoQq3OZRcHSHLP6x055OogZHz5LCZ3F3Q/rbT0BfyXCnjuFBzsKYQu
X5vgYlQI3R6PRkQYc4lOdVrqcjYibCjnYXZTbjIVbXo2VFqakNvN1bmZQVg0AYkl
fwxUmHq6RdhYtVpH0aIcWHOzkU6Dmp02Bu2Hnwb2r6sz2xw/ou6JeoMveldE7YoZ
FGO14FpcvjgNqoKnQN70zTNivvZrSKa2LkWPvNcmevSUW/5hxee2jlYs5swKEfVz
IIrdukJXDHbL1jDUnvgTwqSN/e4GeQ6hqXzKIGi2mXbtOi7SL1XaEfKQbRncWuSq
2cPs4rbK/4RAddxDxKYH91rqptlx5OpHJWkLcm9w7Xhu+UJICrAb3j1kcAYen5ME
EA2qDyN8ze8Qep0BHrF2AtxUWIhCk/K+1Lc/u6hpv8f6+MAIXt7c1KA79iE/5GnX
UOU83rM25moCAxFWUUgoeb2bNYPimmfwHP/rdqYAnsonkApqi9pOKuy/hp7u2AUD
OTCnmE4mEDZeIqzG8GvKFeabQJvAPGWheBxjzr72f/Ud6bQDHrUzYew33E44DyjW
7wRo6aNavvE7uasML9yNHxbGv/3I1L/h6/1RT8y+qyoVAjgEXPMy02k3a4NgN2Hd
XSDNON02na+CFx5frgDHhcnEYqeX/KEby1p+XPsVuglBUq+uOGFMtwfmbmRk1+Po
2T8MAyve2HNu829koCqPOZW2lsdKuZ+Sg59wym5jBJPaWWMKTcbQMn/+KA77BbjS
Lu1cUMdDm3fw8s38iLDxxw9/nQm43jTMoVElqEcQV+OKd3Q1eu7tNKGqqJfQIZ6L
caeNHMHoKN3Zo7d2u4zXEJS88EaL7YdAhRo3JW8ykOuSBDieE5YTNQtmEQxj96h/
1UGICIPeR+xuirGGnYj1iM+/XLRt8vF7+6QRwTdnl5bR/WK0fAdFiD4YYMHc1+MR
yQTmXDAv0Y58c9GzhZLIvk7Eq9l6uEGVA4pfSdfOjg+YOcZR9/+TNqw1+5zGEeIu
2lKGldaK7I/dMuy7y6JXvAPHhdmoncpp2eCEwnltXMlGvsUgkWMprXMQUiDBu+jU
+zUnqQBZS0k9v/anE1XmAxKO9qBTP4sIEHMWWxWIK6Tk6r50gW7cw3Y9oCbY1ch1
Hr7evPZ9qnUQk3XOdqo0Hvk7lzQl+ZLIOpT/lcV/oqhIHlgYUMfK8qDtfsy2R4kQ
z8wiD2yBQtsh+hW23gsucNOlxrAcS8/mt8vFXFgTXd9Qk5Ln+F4fW+ZSyMhgXWbH
zGcFB2b+gmYLMo2jqJTokDRmC247ZhzoM9xdGFWXc4ZokKVZ/h+VXbOZzIXLC8Pt
EoDCuF+CsxLddApfRADZQG8//cZQbc6nJ9VJbqXUnwTJWYNm4/F82wXjTWjx36vY
WJXJbGU9MGXEIt+xPCS4xXvPSuSszYVmOROFbOr4cF5224DzmPDYcyEjcvI4sfjM
CYoSHk4dQWqmU32TduxJ65uvjCoEeDKLDQ3ijsjNSmffOC2L8Pb2+SXNIAFg89Bf
/2mN+QBNjcXAefGN/6y9/nqrJ+mW2Tq6/3Pcjf2lxn/wDfArW+3lZTQ/Rz+HhM7U
PJSd+YAfLo8hb98inogo0+VuOpVTs0ENNq/+4M0CpGosArltOJz/vXnuvwXt148P
qmg/JomPG5RGWmzyPCjLrHKzfTn/fwM/4xx/9X8gnj9qS++3yH0gqIAis+L5LNfi
YZxtp+V9LlffNVt60/bdUdftNM6R2NYz1P5Tbbd6+Syy4Zs2YAogjWeH+IuUlotG
wzXTkAr2xSh6WUCtA2wzEVFknkPb+nlFJTpP/X1x8KDbIToq+8yKaGLrw3nUMSFN
qRyBOk1v6G8FU+vWesWXEB8GhNyh7qmH69AD3wOoWL/iwSdTmQ9GIV6RR6evosyf
s3710FvFV9RCb+y0vP2TegtMeD8o5BHrjd6yj71I+jJd1gcgdCplGO2MH3Cvl7/I
uMYSLo8hWuFDB6f9NG8S0PcHBRMYyfywZ8IisLDz49rsEw2cjHrko9RU5AsmlaIl
90+tPRChhzCNRtaAIq7SUe+1DyECM+CnvJHiIiguOCgFkbbhcdoI1c/w8f3HxLib
1lEhjjLijN3L1NlZ7Hj5VVDwZp+8dzlEmeR/WrWTFqIBpSnfmrDHgSwk4kciN503
uecPy/aN+aSmP/FdDCAc/UJ1063AmnKozYKhK/1MNnjILT8ZUJFb7P6++54yrdc/
UZABHL2njlS4aTIk2b9Epgn3wDGTpxi5R6d0ywG2ChR/4OYA4Dm3owajwJc7TcHc
QKgX+IxTTt3jLv+9Ab20RRIyMvTnlHYXeXaalxapAfc+evq/hRQ+khPg5pr1GV2f
su21QNjPcJ49Nhh1WXZeFJM57dAUmbiAL5nQP862zKjkAyerqqY39TWKaMl5lHzj
ZU7sMLo6SBwmR1qS3Vwr9ro/U39ov5NHWP/Tn7OF/a4QswxZO0BeR0OSvu62oqn8
L2ItjdajwGNJlr3/caB8cYYJ1sXjLGC9ZMaQecuOVM6ZM0gm2oO+xM8en30Jc9BL
miW6/U947QQEnNbeU6LaMwceLxJYt0bXjT/KliJ+ZCioxLLwXDTuPU4Nq4stV9Wh
jCW+p9s3wq8nTrYa5i6+1o3XQeRG1OWEEaVBfuIM6WgGimtT4Da7G61MyWW+wK2K
sJZoXQz/DJLgnUazY6Sb0rqRyFK8wEJP0tOJXHzXtkXkdv1xBd1GeQNHnBjq2R+K
LEk6xVmbot708/7TFQb3+B33WhdV/+toLAmtutHvo18ZL5CZymW7NwvrAS6wrUfk
sqVFu8w6lOK1UUnUP4mtLLkxTOZDC99FwnZjM777FUbmm4vif2Dpi1CrEESFc9IC
Dfmx4SP/49TsxGfyhObZj04HRlBN0hVNsPWSaVqayHlkGcSI+7gHmuIbQUZS2lm7
Q25sAPXyq3/9CtFi5yH/gka7My4sKfmJxUvCrA0FqQxf+DiAbN29ZmqIY8BSEMDA
7pR7bmVzY5HL+Umc2XyTbTiiAy4Ut4D/mknqOzX60jv6f0Uth4WUj8bSngVMzn/A
qbrc1feKkZJG+vyP16pVSj12D/sUTzzOelCjoAf1ItLhie1oN/IXXH/dK3CpP3EX
jb48+VcnMCNgyNdA6znStAu/il5ZXhIzgnG5JOFngil0VUsdLkGCCVJ30EhhkzQ2
s2kOM9gZgTkWhTBJpqF0E2pTU1aQ/ywkKDjcW70ac1auh8BuQhM77Suns35km2lO
E38RAKWCKaJCwV2bMf591WMdzdWINN9EKIZTfWGBV8UaI2zNqIQw0i/azSff/pfm
YTr1NjP763pXm5Gpq7GXi9T31lNvmsMfsmIkp6zJ3NbpdAKMmKGwgBpmCS6a+MuN
Yl81Tx9/5NIQqX/crQZ4wiJOqF5vsCngpWFOzJQxpT5jZoevSdQJ/P1fZPSENAPd
GVS7QAZAnJGBgl8YLtOdSKbHdsKY/KA0Ocg1t0Q3aHu15kY0bubqj7pHsfoGaZOn
dUb/beMSajXR/P4N2KgRv0N0VqZekWYBWdCvJhVbRt3+3se3/B54bj8ZK8zrS4dn
SjF/zz9F12beN/7PnoRaK0ezeVR5+AybSBq9wc9QjO+A+k5e54liC2Q+YVHQjy95
T1lMtPKmLYJSU71aH4Wo0FvZLj/WYiL4bD8osZpcriTbN4Ln0UZLLpXpwj0x6jvm
hHuObBON8t8qt+Vk29+icIhPbfr4Dx7dgZuLCAitC2uOCg0bcTO797ShZlJllk1d
uli0OEaG/mpIhbieEzGCWdjkVf6lKJJWQ7JliGPhHQlc1a7X3GLlAEVpFoQdB9H/
3gPj5+0yzV7i8fo/bU0cfBL7qA+uecLZ2cxvVlsFJ0m6FHIy9jB/s+PB5JN3bAMW
QEixzJ8DvmW+xXrvcdNVTBf2Uy1z7tv1PBgg+lYGYp3ANk4GfeLptt0o/Vj+1XG/
zgRbAGCIpc+n3A/QJENAyeilL9MFd//BeV1m0a+oQrZqgrVJ74RX4KoHfxMq+za3
Q8YtanjLRU0lcNFbv5e2NddlaaOVRtw8oEoj4K6zogWlnZNBTKHYfA16Y/MfuBI0
c6KozfNq7CyKvGOhDMXjAWBjCvxsQXvbn/EBU+3H7iJoouRz5ICHn6GfpMA8bLfg
5UZiIcbXArebK/mVAM6m+tSO5rn6Z78Vzwn/O2sOiY3gZwpnb91+A9NKNfzk5ASP
bgFAM/+NYAAGTB4wQtl/gGLd3bYidjcN7qoiZjMAKHSpVvpCLoEAavlWeh2cKBnn
Hr6LWceMeabl7SIzDkw0E68rCs9bmAt/cRgk5SOTTYh80GgBkBPsDaeCeD926K9u
A1gyeUo/7MEesm7zs0Qis0/GhBBwjEO15oZjEJxWTqiXJkzSQANGT4wWC5iGtPrC
IrTFu15Cd6noLcRhpMGtta1KyZXsxs+r2EI+uNDSNHuh6oR/8Nt1/QZ/MkgqO83B
r4wKSmR1E/pFnZzbumC4nI7jwuMAF7zNaqW9m+rtuczv7/YK8C4oisiOTPCp34ON
Z9SqhNAyKApabpo3Ng9WUVPdn7rSTfxbQjofjNHGnwpMcbsolBSaI3pXSJYEkfkY
2vqbs8VzkI1w0ZCgyQx9zOg0F1c7bTJaBz0lp61jt1YFw46oHMT+QhWpB5d93Y8T
GOScgpRDgN/HoisoOGSU4fnMoKrb9yEWWPAa1YZ5EWx96/kJ/oe0A+gEndkcLsOg
iNl4cJOirtBxRfVQ9MpHxmUfmr44bFuG5TULfYMUThMxAS+1RusTqaTXSjgorDd9
0z9IOKTIf35zlsD7Bt5kqZWBFXXGJHnSImdOg4HxaX960yhhjwRxA57CYFP3fPgB
WPv6lQcGeDv7GkLIyNVZwGr21yp8rBqhiCkinOd5EikDbsJVI2bZcx8iW0D1zuwQ
Gv9UMFDj8BppXbOVGgTiDkcffnriwW9TQ20xmMuFBItZtOJOQuIFVbUdtPnJhkj+
VIn9trmA285YFQMig1i38U+SKBbCYIRQXLuTABP7JnsTnnNAMBkUepD8j4VTNBT7
iWmP/hN+0aIGcrZ+GUp4/F/xdwvIS1ZVsQ1NxAEKoRENuwih0m1t5PdweWU3Z0ij
J/KLsDi0fhOwbTd6+YxPl9+LUFdcNFk1Dio62jon3OR43Zrhaqm1cu23W9cbGTpy
n4IftHJ/+hXtD2jGZA8FHDiYbAVBxvemycbwExn7WKyRy2B8wYFF4fJTYnYoHCEs
MHJjxCNWxuh1AyBbTgBd3ntJxVuECIZVisd1rESqdUYGfvEzAfAn/+ObHsEbstmy
jfF6CzwR7XsPJ/7ZtesMCHI0z2s+WZh9pk2Yvq3BiK78YOle2zk5f74n8KSisrBF
Lgzi9kB571jkx3QfM+5V38XaoI1VVenUUHJBwzsW3MdKBr5jHeyZ/YeAaji9JRGX
Fw9efS/W2al/qyGQhq5aa7UXGHYCcxxQvcjyz3QejuGsWGnjdtXXrfocXKnbnMIR
pzwR5LygAfFtnJf4W3e6e5b+qTbvce59EOP0bVijlqaqSD0ROGWR2OEAIb/ZhpD0
imqkK7BOBAU5MwyVbLtuW0Jr9aW3SkI80xV3fBR9AWv1JjKdE5hHE9D9YCzHVxW1
sIo6NLVAK5LMoc/ezj0Qw1IaspzZ5+sxOfNJYgKXl1lLa/hk9Hc0CljhmUUvl3HX
6NuvHb+Wpg2en2zb9LxcjJxt5Mn4orNAMYi+Q5UOX7nrwq72+KcI2XJ/rQs/mOtu
y488i53LMfCbcuF07mjxqD2LIfrM91uzd4NawjtHrHqDqcrScwyoHoW5fSmcxBXz
VFpPteAfm7FeuavBLZV3kK64Sg2U59BvFZy+xEobpQF929EFcfoaYwKp7hWfaP8b
bMlnlla/8YC7ydi0I0Cot8uu7DISdI/wNuaE+R/qrz9LHazWWf8rDyKuRSS36l05
yZzUcQvxRkAqLQFDhoyvKjUe543y4QBHAQKaWx4ClLEgTh7XJ51jv7uWg3S7YC/o
6+ymHDG9hMNmoRSrai3p5ine2Nc73Hx+FwUwe1tvAA87l6bAfmA4wqVw3jX1VXxH
2WrC7+oviW2ak0Rvze1zHQ7tQ1ZWm1lpPOxr87pYsRKkSXt1ll0RPnV+vmilXtSU
xo20yP8jBkyj1OJ0zpD7aKZs8gqGS4tjKDzF/IAd76KJUCgpVX7nqmpCtgAQ3XrS
9ViheZYPnJhoFhUVnfn9M1wiZsR6cVR5DSADG56O55zz94nx8kQ2o5m4xG42y5wc
rvN5hL7JYQ+gHQodA1X5LDr7Sx8OKKd4gKnPz4h4+2WJB8o0Yqs6Yjbcz9uxP10m
cTl0IeoUp9w9+se4870yMsb2Tdhd+rOAWpiAocX0NeS7HRiXF4lAVH27CiN5aUoB
Zk+H+06vi08G2FSm5n/PgI7ojTPLuMcgf2yPfiUix0Ojdj28kI6r9sEEgiCNrS8K
msotLy6QYOtIWsqc24AM/wjdhrVflVirKGtjbA22PL9XxxvcaAYYhForJXpsEXMr
6xRbVREu/T3Ce4Usjhs5a0Dkkj8Rq0DS+qU1BasJSVXOG5XqT6EePfiOqr4h5Gsd
QJpzzpe1olUWTN0jlgDb6TQwowKQ9XmSZwBVcW0Q6wKus32exMS8eUAQ/aryR9r7
iaL+//7si0Fs1mtHKFpMYUCNm71sHz0+Y0c3xoSqJ7U=
`pragma protect end_protected

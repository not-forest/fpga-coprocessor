// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
p0k2mC4ile7JAkpsNaQG/dDpcDrvaWx+Nk7kti3NIg19ZLJLmCdC4UJQfn/hi0ZPJVoUvbwyyEcB
gEw6vgJijH8bcOjYCIxy9VIzCt0so4G0Q/2rcblRUAipQldfA8LEz7xCF3YnSQkPb96gt/0l3/6s
ktBclOYvldFk5vayYUz92GQ4eztWR+agpvz/JVfXSpxYmXJOMjFhbPP/4LjHH+KSyfETIN9GDMQ3
q9e+QdM4ONmLdfgVEYiG7mh1RVTn6mfPOWrQWrH54ewjE+WNqbacNPOUzU+OQNmtHlH1YZDVgyOg
EL916hRpjE/bNjWxmPR1Bf8SZz7OxM54eHDAVg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 10864)
73LA0AASiYacQ+5oe5hqwseNBEtnNY2BKsagVEv58pPAKBDdqXjd18GMWuWbEHj6u3oPwh7Pehd0
/Sh1btT7dWUP58v5KxzddMccQR6+n+8l6D0Xy0NjC6QeUK22n9grgL3ZKiMj7/z8gIzL9smBlbEi
ZArTY7BvPWt6IcIQspGVMcSi2Sdeja6w8DKEHgpHK6fgFBmPKFhzXYmsgLr3qYrh8ye1b9gPl/fu
x6T/kURYNsdGNteMcDp0ihfInROUhaukrRN4edH4zVeEIbPEmrVvhwgrs0Uqvnk3VAE0xkyJcg5U
4IcloFVTiUcxzYxG4iDiCfLyvJSQJTsQ3ioM3FCK1JthCUCBJ8+N/W+gWlcJTs2q8NuefBhjZ0Eb
NglEsr9o8mfpkJCOraOdwsdLcfUhC50BnMv2v8GDSdd2mE1A2vxk+NmHZ5GWh+C6+QGJD0WtIVTv
8eGNBGKNPn8zUfx/Mw9vmSnzoOKTwhTXqcxOxkVk9CiZU+Md4oYP0tiNHwE1OUjOC7xxwj4nQ+92
iRNcgMUr+ycvOs67hkA5jt0KVxm26psOrxoL+bdxLfxFGPGM8Yhv6Ntt047oZWbfpViYqTpe7DmX
qQZXvLmFksagoOr43iLtjy5CukumN9Jj5ZAybntq5vb+UprDVlhuH5xAEjRR1Oxkvx0HAmYE0szF
zHGUXH/J8bsHkOQZ3HXQvaZJ+KhkD0jYv4ISaMpCKhCxJy1zAy1qUsqx2xZrCCTiirbu7vg/wFer
/4mAM05W72jr5IZs4gAidPMOfVIaA47dahdkyk+T6tgOERLwmlU4MKlct+gkXMVp+9EME9fw8Oz8
90MWrecCWst4/tqDAkfc9bUt4PSuTk0mHXUOuGZBlKwbqsHBdzoUbSWAlXCHprg+Hzm7BSdNfDf4
TpL9kG4Ms1hp4lJ9PVWIooRQXydP+4+5zfaMYPIo+8sZSoJbOTb5QTqBFnHrdpSLUROMdCOcz2q3
b9plN/ekpIbD9WxYVijtFp1QZWefbB0WZvkDeEo/HQF/TBPT/i/lz85EELYDURaOwzEaVVJ6T+C+
dwZGLj9D1hFQI5AZvrJRRxfWbWuPRg4f5Wfn/pdez+CY+WOLgN/I9jKi/Vde2LexS9LMN1BvVRnD
bdXnaV7O2wCA3436V4n+DSqHptV31yvdDNfwLQ7ohGZfKvkjiKVnds8lVDEo3Ic32oRXYIxWsf1v
P6L1QP10+NJJzS2Zv9b749nsFMaUs/jwChmhLdRLZDKEf75MtVAt6fsyASeqIh05rDHi1yWreIYF
Fv6FiWrUAKyzl9WRIUsJ+yo94mabpSoWXgOIhn2j/P3vV7FQk3pMgBDkOX9CR2epbt/TMot0yI96
YSCQYadHHod16BAleR7WRDbfDD4Wy2nlkmCEwQ5yCc/rc+5DEhyQ6FniNb9LyJ8qkbxe4IPwy1qJ
qxF9LfoV/c9IA0wOfk9Mk5Uf3u7foYaNaBudakxBSmR0ByQRM5llPs0+p7CtYQN12/FbF2r2xslb
6N9EjOXUOi9vSHoMvDvqZhhXr6BfewSRSZw7nbDSa97mdQHa1qWDNBxEexXQlwlyJfXy9PMdEbpw
L+TKIlS3wu7Lwi7K4aauSD3yr/MtQpJJ8AVUPBOYJVK4RJUpkuRbPhBZXt4z9o73Ie9sNt+Vh/1T
leJydvp1+7n+c5W+KIY8wvo2xVsXiYZ1eKnplWW/KCq6E2Gla/HSTqdJinvS5EirKUsqMBTrYeTL
ij7Hqsxilox1i5BFOOy+e9g29l/XmmdGhQMb5RKAqg6l9fDefIJWDBMPiNs2R+y+DKkIqZ9w+r4H
BYrdUZ/luo3bVeo1xdM4BcAwUE+RoghH0C4W8Pnjy2fMjT99OEmBukprqLLa34OPGAckx7Kamu6G
VCsaH/7U7rXtKlbBjnktO6mle+7niRcRgoUZMl1lYFDfPyQp25cIngtxfPGJicr6QV/UG6kQtWo4
KRz9uptDy0B5Rs84c3yTj0KQZk11DabEWZv+3AwevKiWdyjhtuH01UqXtMHc9CnJQMwuHWCbxHZF
ZhMQl/rp/HPWue5ItOTYMMb0QK9NaT8HpQMa2GzxCdSHDI7MK//ojbmwB1jBQlupTYi7dxNJGVr4
Rn69xI1eQdo24cqIWKFGFnboV7EzKn1rgUo90+hze4MDtxW0HD1kspqDlvFcCcJlXRp6EhyB0b+v
XDDy0ScPE/NKG7wziSJr1yj52oCbnuJmZUkdIlPsi63GhYQGTZLgftSpnK4gjWmt+qpxoP5a1bt9
toLTRlNphFyG3vnHW4YTH36+UdeWOgypPVnYdGz3kffi/CDxEFqzzrVKHXyKQkqrdRyQmx4EEzsK
rxugUca1WANKvUv1oBX/CcbiFxoDZ68deJgpxyFJ8F09USB3XSSTYF7bMbTx8yHXGXWNEcxe3N2U
NM9YdAaCn5wPYn4FPxu5yNpK8OcCCD15R8i7BaOwbxmzugYelAwIweofVMdOIZTgfm8Jes+iGJhu
8j/lDioQ8V7rix9BwpU/NFywTkNT/f4XAzFQa8GpXefTy8TM1zJwcvJfV2y4VCTPBKIvNs7a3LHp
8Prbt9VEM32Lju55tVHlWFiZ+1jzPuEMXX0OSP0pJcwACWpVr0SdgeEeWSzAVBS51Mlr04nof2HS
TzWUP28YWHtabq49AIPRezxreGF8Dm7KEy7zbW2AVRLx1UpzLKXGJD/WWcPE26KNzc6RMabJ1NCT
5jYAlyzKl5QndhsGIfdL0RuPDMw7QN7HywRMWMfMNays6yM/R/ebWdEu3zeuMeX1AyrJX/xh56Ve
HihT3kbePgY3EOaiOeNpCPChmgXEoBrFMVE9+77B7rJncCdpMPfrkE1rw8blUC9VVW8+L6vs3hzz
7ddXOOEl7Np1FBlZp+UH45dwIPWI3Qshw3QBjey0Zfpgvx1B9fb8jvhaE2zxVQ3IlOBXFT9g0wb9
dDlFpyf8EpTpNiNRzS/NS3gMy+wY695iBLjxXDacn5yy/6koPTXpyQpLg6iJkWMVtvt4QUBM2tpl
0P0FGHa9Muzrbd2UVGwJybCyF0NyqHstSTFDFklaqslla8URczmei2B0/JhG+mIs005zV6Bczyjn
h2I7ELHh1+Z114kmNGd3VGRKVt/BnA3XnJprguSl/s/2UpfrlaWnk1ngIN5IIUaLIQYHQNcf1n4d
VYIZLNCveCAiaWoC2R+RXarG26KdCIBGbpl8lkbo5blRilSp0eD4DnVbcvfvdCLaKxsmc92/v/vY
2FNZhfigIP4REWSYOcqWsT9vQAYaVSglv1lHilWqyjoheYeajzHghO8p2wFjLOVDi7fgPMFLh9TR
FnZ5WTcKsdoyVxhS7YeVrmJh7GQZRwKi0veDDb/iuiyfd/HKfQ6tbwT/F9edeMLEhaRs4TyF6J4b
LTVqc2ubKD7UIniNudBIAYpPX29+gM3gayTuUCbSckw1TpkwjcuRDEGdJ9AQcftesNFPYO+RQ4Yt
GNE7DIlHcffGwSna0BXnfhWQ8lZ8VrtVQVFdrcKtts6WVxcvr8PMynLJCSb+1DWdHgLGt6lA2n6J
lqoHNUaPy65/N801K+Cy439By0dyekwr51LRlzO5Y/T38hFuRXgiCu9YUMlgsJ18sy5QS7ig4w0j
OZQ3VTgEAu9XWm45diJyRGCKIK2lYDQps6nhN3i8Q9c2cSrboan96UcR3DjPDaMOpFi7cm+AtoiH
DNG0qTCmIqK5A1AcUSV6PliLAfZ6/uTRV1kn8BfDfN1XU1osFCDBXtF4+9S8tXEj+1ILCOoCGkmK
SHHXHp3Sn+3dIpETsB7tellFJi6sd8XwE569I2q5lSDd7GWqJSigRZl4/Vw1hTV2YqPqLMo1gUG7
/+3pNVkzVoHVXqUBUs1Rbk/acPzd29MORyEAVdtPBPsf3Ske634AkjLYMX906F5Y7x+8LQ3Bvwga
Nhxju4D0TGWtLugTY47c5g3Az+ajy17AZ+Nw2MfLmGL5qqK/VOd9E3iklOw/5CuN1h0f0mUpBBXl
d1Z8fS2k11oNdrinpy0lZdvLoQD+bfzxcpj+/SZU+BF8dZwl3tEtsdqrRtUdezxCad55u/36+Yr9
ZERWM0OYSWN+7x638WuN+mrT9Gy7o4w7GzJUkurZMq3jgaOuNrsCRVCnW5UnAYXeYo/Eu8HjuuRz
+TFpyBXd/LXJlSNseUkr816e+MgWMWc+6tYNLsFXyg3k0cO8DjQgqkeM31/Vrzraykw3EaSYhy8U
SjcsANbVDjpy7uqQYh1b3flCLTWG3kycVUj3sZWx4hggZUdADI+4LSJQEvM3fI6YDU0I6bw4YC5a
xALw+S4CAGsv+fSqFOL/FzPnkkkVSBPYPPvPvwUeB2+euVCPWssPjNqeFO4e/EsoyY6dTU4B0VVy
HiDhRa6EiHmk4NE8lwShjH3ApKCu3L9xCsaiAQLJVgXfy6uEy6dcVkPJAsvuvkK8UhjWihyU/Ilh
B0KFKOPNnnzzqY5V5e+Jre3jzViBoN45INjBBxH76E0VEZaHu+kMtAyXFqbOSG9ahxalyZvWIqHX
Gvf9hBkN1Lxr/ngYpvehx7geYXYhN7U8WragUba54dZcByLhCfxLUshgWzu1UcG5D0WC9qGEXXV7
lFrjX/fWXZUIKYvMmS3SFeizNuUdWJW9Y7W4V1cWD6lK1r6Ynap4NRlawh/5+vlUTh8gcDLoIVlC
h4d9plPrZzdkY/0RAma9LFj59V8rR95ViAd2LT0R6IgSedukuPAnR9vZTIDp+k+1lZF30hLFCC0c
6oOBcbTARTI+Gcv1FLbX8fOvt9+RiKl58EDhvqWXh0m3xFRrdmDOMYRrdVkzwROxn2OAkeJzYI5M
qwkYtU80Nu6F9YfYfES6i1+GrK0q9THPMsqC1o5qjMPyS0kkLr2OnqvOldQBlvIXVmlr5wuvIkgo
dbHy108v8mEUFFU7ml6KVM4ohOudioVOclPuYuzeTn3x5cTygak+DwWryJ0FfhwCNJhFqaLdDY7i
7oA89s+Gt+zq6hSgQTAaWWUcUMACQaPwLFio42qsc+4ghc54D0c7CDCkFKTmK6XnVUaIA31Mghsy
IgLUszIBqpanCMin6TTcnMm09O2LO1ZzSNmopTN6VYh2txqalf2iINoJi7XgcrzwVRwGOno2UpG2
KBsM3oNv9MFg1/w13/lbW2LJuiciqUBkoN73cYr/Uv0HAAGjG1SA+0d0iMIKt0WRPJbueHAjt6iZ
3ebT/q04/FAXgTRD9v+NFzZImWL/PRyUeRhOD3MjaxDDZsoAA0uXtI4o8cI4VGq384urhplqSL1/
Qoz8dQWwYS39oa9n6YcYDfrsFzGeLz/XOHGlyNHjY5U1XAHsiuCTPinyYzTNjyG3rkqJOB80IvQS
0luNYFUwdEovLLwE8PO2wplD3LBTrUXxZ/30G4t+2cp2XAZI2gxhvCyJ8Ps87sdovubod/lRzYVd
uPXxLcJIxjet3drFdeebyz9/lN/v4R+TmNEGt4MS/TZUbwlDiA94emBV+fgGrsDLEITZfv/qLdNg
sGfU6j4l4YqK2KOQelzNNjAGyY7uDss+blCGVD4tiCr268z6sUoD/EPlZ6FajyhCV49pz3SqJ/QJ
XgSqlm/7/D9f1FMZa2/1DBD1KTNfhzse+W0FZKdXM68bY/RWrN2xB69cZ3IGjQ2gbuADglf4n+nl
GmdLDdWcj23bEey0+oHoAQIEIx1NR+9xYrea08KiXqoN+B3iLkhK5MCxQ5AGMP/gy6TM+8SnmKaQ
4Ck+5lU/3FiV23UyDexYVN1jp7jo9D2Dvjn8pYiJ5JBlevr74K+9cfVLxmaSD9V0gLYwlinHgrPM
lyZsCe836PEOdqXx4dmsAhXgQUg5Km38R4YmS8pu1i0KPAhhUf0w7bk7q+GVtLPU1OESNa0/Gr03
aco5zK3LoDCIDTPou+jCWAfnjAQWSUdp648o31F95SBftYAuvH70wKYZwp7hGbIico08DkqvbWEY
XXlbPHnJVJ9zLR6yEGh3oPK67ZxfrKmJ3jcATaw0KY5qE9uPrlQM9LyEU+sYvwpSZYN6BxIXiWU8
W3CWJRSGJbkqa1vEN3/mjLDWIri5GTPNf2Bfiy9T+XqWJ58DOltsWNhO1v8G+RODn0dOzuejDIuA
TkRuNWEUG40Vw1vCQsxQ10v/e1/9YNXUwY31qU7lgeX+8rucBB8FzUcuuVLr6GtJQiPUWk2HnRY9
EqZbyEpWHvl/BW59bSMr4M1MJ8fvrYdY4pUrWoIjuoK0O2vpJepc9RIJgTntSHef/4n9dAgVAVSl
0/hBtHJ188AS6UPnX8wBCJ9POczx+yLx+vGg1sSfYfHmomkcO9AuBImTdlqu+DswhTLTWGbrO5KU
X2Gqxp2cyJaPlQan4KzyUrxpUVE8RUhjBQXyOxzHQTcMfPCbTWL1FbJetAc3ERX5he4XpzB9kzm+
MXlXRacJ8XJ18xKZ3VDGpWRexZjPqNeuWRodff6/4/qLKkBwpKKyCALP2A2jmsLihpKrQXu0ONXS
CDmy1jMch4U1hUC6qqdDdSRVqS4diM1+j6Z8D5DLToBDL5pRubLeKMT+ef7kDvNyBYXpr4OQZR5e
zzA4RAS3aFMyAvCKSEuR0neb9ofhWdagnVR40kEvwBkfWBJRuhNh4FX6iO0lMC6WasJwDPHNH6oL
YbmW3lcORTXnt70sSu2Unaror3L50CZwFans/keEbukqh/KPu4whJKgIq8CbRBFr4ek6uKGFX4Ld
nAjyCH4bdf7UnJ1MdZue/h277X1w++vP6t0QgOjad1EB70QO+l3umSuIc/bgKZ3fIFQxXqIRO3vX
sXrPdiNwPlSJgNrZgg+Tk8CuisuetLPaWFnN9/6VQT5pj35Ggt29/TbsvcDs+Cp3A6kuMjjHIgqY
I9K2WgXqJi9fgTrqWmKGLSmtQj2IjsLdvZAj5BB7xPSxw2cW/jucyJUkDWsQIpma0t5W+n0iiNzm
Rvjebqa4wHnQUi46IvvOtPs3wwsEx9Sp/eqzwQOX8jtY+HRm0YROUJWsz2usN7UDNo6J9SRq/dj6
uyai3R+iLJHC8/rR8kXMULA76ILYFnsUARqrz7QnZvBilF0QMBH1nlhlLHXqUMSknSzIsav/Ndro
U3RKEE0GFkPR/4UbZy0bUrcwaZCU9vwo3ZkG7K3ngWIg7+Wf2TZwPlvlRLLOM5WK+aa9MRWl4T3u
/Mp6Si4Lqt50sFc9+kmZ5lwXPZioZHAkjyp+6gSy6lHlVKpJUMnKJ2MzIUtnQaS9HO6vWPHJ/dWR
u5cweLFB0Q1S3Evl/0xme7KuHhU5bJtvFS7wucuYgE21UT70mHpcje/nd45LfTSE6Wn/8rirDE6J
qjsGz3HDF/JpAfwVX9eYEJEhIogSFOms/wad0S3hdV87r2+HTCtUNWaoXuTohDpnphq70vUowUcB
j4cflMSqaVgHxhZa2mE9R9U46nEwz5O4VvtRebuTsjK//njJ4XzeRz44EnbslJcGzF6khSOuWBFR
Q9TFxAMvu7/+V0wCRxpzhgWf9/l4sInO9Xnk8Ke7VXPQuxvahhPACryMbNtS6w7gn6xpaXK+Xo7K
b67SVze+5856mXobz0Q2AIaIEdL8J3UdTlhPqYLqPshkKScsTjJLa6HKGP5q/WEeBN/kmOjNMdqY
EC85Kx7qOuhSYhr3e4B+VrdxBeFn9pfOmT+jtfM8PiOSsRrscFDMQZGUDZsDM5Z1SpOqLlZdVwv5
Ov4jHc0IHzZsPFOywUgpji7HJEmsItzLjZpxng6G1R+OFwVH7A/8c1RPznzQzur5nVzN+pO5REYP
7skuCKLEstVHUFlVul4j2+UI/XT+DkrLOsEcn4IPGf/428zZz7Sy4lWtefhpKTz+JM/Kwi+foUOE
bWyutrPZtYbzLZwxhF+RhLbqppEq082s/nKHVNWzgfKkyzjAwmw5AXTinV6WCSigxRM1rMRBLVvS
o9X6sc90o5mXYPPbhWwQKJMCbjPakMr7Y5J54hS3VwNS8cVh1fGS3qWX7fi3adIcpVn+6CAowCVy
YmAxIhavpLMZpAYoWWVTFK6pqpw6O4bTZSCAadZ/Wv4yl6H09xNHp1WUCFJ3d2OeJbGzjjbShqI/
Ft/jMhpmSv11RK9tLytROD04eUoKCnlNP5PDruwKUABhFWyG0pztRoA+JMSOBltlWS8emMXPbi8K
9l4y46M6iz+9xC3vgVSabcDfKn3e3cCyBeBumWpRzIbB3AiH1hsZ9r6JAy4hg+oY8SUpAvL1eaCL
vmDUANuEhlian0nRz8kW3HM7DItjBL0EHSh+68CrBAN4gZfJvpkTQ26d7IzF6C0pAgRnjhOI71sV
yPxDeWQOkSZxSgnh9gYkKqnLVtStS2ilYEwIzsqZBm8gGJfqGl4pjReGH53CtZ1Dla/UK4w4Qc4G
C7YW4PkpGTiJlBC85jl5L6JVmYOsc/qlwtEHuQarHL4gMewEBKLtxU0ZaGwo0ur8ND3bhuw8RMZ9
jkBWtBExpIHCzfncOn5TCz9Fsu4aUtuKyFjQy384LOKgw7vC2QXIT5EpvNL3IA8X6+cfOvIgV81L
gBNmVZgiRtJsVT7DS4R592yVFQhi2GuW3TuhBtgQa1wTj4EQlO4Mq0scDMarkPzPWs2nDFHZA2FK
ty02x4k6yLolFtgJg40AHxmdA9BlfJGp79nydjEAZirs5y8qBZdUYrpTPaoWW80Tk/1ZJmxDWZKb
67aQkMzbuT54cUgc/w/dye9Qd4wV3ZBuYh8buxiXriwqObP16zgb43h7gy0ZiGAb4UAjfFS3Tfyq
C2sbHtG6WzZy3VjBRsKWpRFRcKV3G3us/87V4kNEplWZ2gC6AeexmxQXF125NMPu5adEaBhh7dkn
ufz/T+VyFzx+op8oxzCE0VrEkl3pV2OwhoPY5U0gkBEpEjU2birQFQnUpo3diTfzvJi+KHvYuMLh
p7AaQvthXoh0k5oTq+Y0TmGHNRw6Zj1RA08U6AXwdIa+JWg/VqPpLdzzpVlCq4LKjBJFjtjw4bLe
4ez9A3PnzBSFfNyXUrQ0OFf9B2zpjt+7NaHx1ohAfFZ84Q1pL8NIN5IHqc8AICNK8eEeTTr+f//d
Zw7sRcloiyTfU5bHtX4JiAYlfb3ka5/F5TtUt4KAQaG+Hz2FQp91jpMJVdA+Ipakg36Grab5XL/N
mOy4+a5denW0LOEjT9eQHAeMk6t3VcuEUR3D+TpBnjl3Q7knmByfl01R3NG9ObEKM1cA2qjuF8UY
9qbmq3CVV1dB4xQWGSEmBlkqW0usntBOpz1nUIMDbQMy58Ekf3plvhIbjSJ12Euq+vkNeUP9SYPC
AYWqQYB4+FY/NxliP2r4BnusTr2xwHu/B98wILjvPDX009ZESqAgCHoal3vRvt2F1W60LpqN5e48
VlKkq61Zm5i4CKwaJF3pc86adwFY0tDD34l0qERnaGPyaTPQepzZ4nh/p8qErf6rbLlaXMJdQO1r
i924pC2iRjak4iISNdNmMgXUiufnTYqSBIJ0RFE74z/Mq+YziaH5i9e8BeM9wjPRkL9/mBdCEkPq
7J/KbBMIHrKPa+Txhf1b5UhuE8GTccIhLiT+DLJlCCZCKbvQVVg2rqmtcQCVhqpwzksx1EOyBaqZ
S5eu30EEfwM8WcNyxmjPEHH6V+5+ckNWKJk/JBUrakbzgyo/8NansMJv/RBsHES1JXEZCww1vWiZ
5AcwDfPoV36b+4tHOKBrxBKuVYmF3gZbHUhzNrfa2rFZerJVbztHKGeTMCji3FlbbP+UcFbiVcju
lU2wL6ueui299F4//VwprUNrKrM52e90O5dq2ybaeGfEGIODJ6vxxLNNl4p8lrOrzZItLpUcP3VH
BhKqndXVtmBo7oa8vUGHSQy7wejIw9+xC7itc962XAWCH619fyyviHxyArMMFKNY2ucZUeP3Dju2
JVwm/fAHGQrYQh1iG0GbtrjUw2MBjrWFMwtYF1vyd0s+bY45FdF7lOh0OBV8O7jx7I3nl5MZHTw5
HPWjGTtSbHWHH2ldRNtWgtlggdewUf4wNkjfsGWKUye0rbEJUnMV8/5SRp8EoJxCNFjCX1rmGWP2
XbMTARDBEnqql93eLSx4322jm5MgTN7PpA1wfNqd7855pP7ZQ04qfvcgvGk+2spIDpZzJqJzIdY6
cnyxiJ5PLNCcYZ0hjq3JXbmfybMKTT4n7e+JjSuH+FmYXO2k/vS4g+N84yZmZaBuqaD3P1ETpmPd
nA+y3a+NROdyJXmF8kmtGUzdITZo6UOnOX8l0xKBPHqT/o+sV3+LmzTIZpxc5TNEvEFkh5wRmnMI
K3rmS4/7L+OTsYIzKE5+e4pYHA2ac1XjUqcrpVLY1tLyRGOPu9982fBGyELURdAr0NIDlkrm7z5O
vDCkEtRhptBshAPZ76WZ1ztHlRzrmWuLMniaq2gbMqWbtAMJ4GNHGnlYfh9QUIqULNlFzD84h/F9
8lOx8mosunjYNyJhkPGmDOw0DGheJxHiVKLhOfFUasptiwJH46gjN80s4GHraC2gJknoPMktL6Lp
rZGuaGZVjpfLsYf76FaSXzzV98D/eJH+3ihKzMHttRCIOPE1YxHRCDc3RDqfUunprTnZ3kTT8p4m
+YUmimvoEfHcQHgPCApRy/zMgHXzK0qLPQE0XskRr0NObSnZP+x/h5ykN0vPbWaw1udDXHJ0XXem
+O799uFNAWLowSNfVBmeY0MKihSXjgwH2ECBP6Rd5gIynFd2hfT65Mh2QkiAxW9tq5nHlP2bVVm2
fVcKQJYaRr7L34fGgE95aY+GJmswIYX1MWtwqHobbPu8d3+mKb5qKiLW0AH7EBPxbI/ATzD0WDOR
5/JaVtzYU4qzgv4nmA+uxx+6i3iHs2j+0JOk3Z8uANHH6P2ubp+fb4+wocAcqZyCsYD9OrjzPS5g
K7/NHsYNOV3dqT1dEn8ld9vB3jbTe0D6esPGRbXjHjk1ZNTIDis7uC2QryNwFvpyEXOyYORENl7s
DCyEoOAcH9d7MsC+LkwHdmK/mwa6WIJIR5eFveeCTyG9IXvwyZhJY8WPgb1ys0wO1SACEK3Ot1Ly
vMq8a3pahsqtXvE96u/v0nukHBgR6QIoH2JL0bE/23t7rUbDYujZTFkfUX5S7CfstQY/xIM0NVM9
xtgEF+GvRPosPzKeue6RjqhToFFAWyRx1HdZh1CfoJix6vJPmr+INk0wpHxDU9nTZBpMnOVIMrle
tF8nnNCprAe32ytvmj85hGj5QrVmh8qdiwT53Oy3U3xeN11SR9KNc+H18XZ7qcez+osD1DlmL8KV
D5pafC97xbT3AqTAiQjgGaXzcJ2JESbJPwsbhtm3UPxCx8LvsU+KkOtAizizaF99woinoBVuLdsH
SvlTNRtB20LHc2/yr0I+/G7JVvaWQB04gNlHB0El3xZwiizXUTDo8oguNaNyt57/NsYk63CisCYb
6XNjl13M/42Ifm8goNtItrqTED0CXmYnzmz8R+cmpzm25YQaFqirOODETzafCslm0pCC8wNU8Jcy
/MtB3iIbkF9OOmbV3rAAFfgS5X9C1S3tji0arCUD4zMS8sA2Xk60u91Vwr6EvRJ6GSlbjbPxQ6iQ
/wkNlmSTBOXF4CV+ogSugHEqvleC8bFudPkp24vJvCk1cSyznm+ik1q6WYogGeX40YAfQi4iI1bF
uXMuNQyJuFL4O5eKOJxmdHbOJWwzJGVH6IpmxS5YQuGG1STsh/V8S7dA+Q0Nu+HR903sO4OE0uz2
2V8MyaWvUJ93ZmdMeAFTn1TRMNXrLpnqvwRfEUyO88Jvdq/bcz1Vmy2wx/0sVkNj2Eev9qtp8dLU
PUTbm17MSWnIK7mm6lSPI5S9WTtJGXrosPgucdFyk80xeFCO94DQ+0zPnc5SPbyL3oyTbnpbt1Ml
jwH9MQfQY/7QCkQt5O/CIa0hVr5K8KMacWsRVZ2mVrNb5+Y1JtmrPN7sSgTlS642+L/QYqoE5C0F
n1O3XwqX/tv/Qne+t3rJAhGGFju/RZRlFS2uY3Dz3tNA4PUa4S9zDmkNCxLoQh4ZbUJoxsFE1G/Q
VIq4ZT6PCyglF7wA6ly4k6BBW+XSt683sJhJffzDwt3jbakfivNIIyY95whCZgDm5l9gIcjjswxc
ceN5YiLxFy+1xRWPL5odAlA50rBdnQ4NHTvm/oS1Ccu5E6zZcO9QkT3ox2lBxAvwAo/iMWp4Md6S
3sdRU4IgakNn2stUB9esZuM6wA85vTE0kIFMTRW9xhtJMS9TCp04efkeQj2XqBzYz70aJtYJ/XtW
p/j8v2+RVgMxu1x7ed1lOTt7klGjb9qVKn5gnXrQLtlf9wC1YQB2uTcu6x+01qhFZ76bci2zw+pm
J0+YdXuIYz02o9BL0uVmLmp1Gp9jFyWNd+AtIFa8XatAIC5M4k7qrdQGHEo3WwnLJ4DSI5DbaViN
PkjbZPSBGel3OXzoPqvRmsT+0vbnH3D+bVf7Z4RIvrmMGd2gzbgx6mEy+4/r54r2eC4tdHjod4/G
nWs1cYnMa04yMB5v6xCS4S/z6bINF0ZTh6YJqCmhpebHcDZ3DvSOAo3Wmi/dtpdQrv2xRcmT9eU4
zY7Vp+L5FdxM8vwT4zG5F0QMXR8ukL1LWjkiMb7dsuYGkMwi3kXasDiUvRf7i5ak1twg1frmv2fK
nur9yc/ONaHE/oGLdW3rVCRfSZlvx9KJ0LyzjFTTev0epBHZKjfJWFPvdIhKn0+HGn1oGHeuJy62
siDGuKJqVb50Olc6nuUMFz6rcmCKGpsaL7fiLkV8tmNcWewU76seZyrwITlGS6M6CK29CY1rryt/
deaQs5aow5ECSHGsRfhHqlngEmBojFQCDQMLHZYhSEtXoXh6nsOuoMq50FZQtVCpyVvDs+h8mdaC
vkyWTsvFwNUd319dIe4E3TssWPDHbTbAmr0xNfTUChuCWOzCvXs43kseIHP4DcZnfVJ6LEGoaHgY
Eskdh+5zSHNkAVHJCnupd0GDEAvcAT2tb90fscDoF+doBb4hAb+geT7QoYJ+PWRSaEu2SmEaaEOv
+vLTodmUCvvqtvnCpyeFnzpoyRq8wT6xAndgow0simnPowS5HGu/h9v+veji5Hqtf0NrSlsPqeEu
gqWnc4afD7DOEqPW3bdp+m05nHNztJD29buS+ERLJVcmqv3Bzi3ODT2bo4AIVylWUr9zQ/nC3EqJ
hDCxc9teN2Ni/lUat6PjxUawG+vi/jpzNBD5dhqa0dNqoDjIg4fVp9dknu9Zo7vJrBjn0eRv8ZD1
aD/QzQqQ8J5/v9O4w5nYMNG1Jv64B6xQe+nebb7Ly143spb7SWP3Lm3EvTG1SvuQwijxU3niwbri
+4T96QlPFLOws/D6kovlLE0wurv/ryRotMck5NIO3+yvP+5qpf78fcPgtmuiclHDu2ibvXZEO6zn
kMt0aFhbfxJ3QxmoIvcdihKaLBLlDAKntjjVco5BqGKhlG3ysfMxBA7l+5EDkZLsyeiqsVYrHcNq
NKuR6tJM3ltVqbhXNeAz4kI2EE0Xavui6V43+xLF+4wfaY9BUAdQGaOKWJ4Ll83VP9NlFJEZzyCQ
AxS/imiaMKywQY7vfkFV+5XW5iq5snfCEv1rVfs59f+ZvG1v7fByM6QPh9XaOGrz3yUrldDLtq5Q
oPDUNDiDym5Ucsob5ojWCiKpBIwawIhYaeUBUTwRVvIdz8EJR9QVvMzWNLU8SyWDnAdUj+GekHPM
xlMgQcMhu4rufITrjmGf4/18Lslob0122QOz2FAt5QJwFRGpKZUzBcBVQHFRhyMDYVxQh7a36GTi
pEOuq75uK12+krAUX3xPWKZ/TBAFJVLxp18dIrOT62D8LndOTaBE4ODuEyS+nXnl1s/cjV8ZsuOp
If7u3ZM+Cp+/13FuHPr23ZuodVKg2Kq+dFaLMfYD9nT7xVTUZrg5BFutAFxOT4jDP9WrqgXG+B7O
2iN4aIOVhNZ6ZH9lUGgf3z2Xhr5dXj0aRSvIgv0wDVNU+/na/nN1oMwULxcsmUovo1J3Jpd/qf6D
B2OcMmGaNx30kofXQNnvwTB0l954UUUuvVCv24VmUy7XZos+kYFt+isVTS46pp1s61/QkJugZ+XI
fuAYbSrsbakwfEMuCXFur6y2I2W0C2j1RDF6bDn9QwXuV9F3n8qqE/JC43dm9exlPgVjNURg9uBV
n3Jo8Nxy3KisI8lysQyFK33JkLUMJCGq74BF1oLfdlBBGV0n1/4E1BP5Bq/DQxylvkI3yDzn3JMo
Jx5EnPJal6KmG/cHqWRUa2/qFGXHAS8+u+WTsRkSUo50ro7eOV01kMIU14RmPk3+1PC4Cd5cNYQG
UWd6d+19x60EpHjAs9erMKFejtN4MNBo2yqLXfPX81FIrIT5dFJiXd2tCMwfztaszmRQt10qDd+/
FrfdKjvB8WH7I93pqHDm2udPcdVaI7uxxaWogVut3KLfTw==
`pragma protect end_protected

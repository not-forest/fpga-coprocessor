// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
RFOrCZdzVqNCvrK4TaCptKEiVrXRjoEcVT35MLlDAUohzGYr0CNCKhDm1mxJ4/Im
Tzz4k9jf+czuWng9fTES0qdajBk6TiIyXBSVIABkQLPoUfUfA8nkHRdfVugPDEEN
7TJJrWAr4APIH7PhtC0ippETJaNXaA3eZaZMXW1J+CASg7P8qcK1Q6QDQVZHZB1C
vAQc3twtMrZSlLAB2fT0+ngHVPEz7Iq6OsG0Nl55ytJ2EEa8IQt99AKvna/3NNbA
W8oNeWGZlYH0lk/HQtcGZm6xUz5kjZdXvzF5HtQl2jcBX3FnNIwu6GrqUJLdJi61
1M8avt0xXNXNrJo5kpxqhw==
//pragma protect end_key_block
//pragma protect digest_block
Kz2J2FmZR0PIXVR0bhfwSPAipB8=
//pragma protect end_digest_block
//pragma protect data_block
3UocfK7PkHqJFwfQvZ2Y7PnwQU4pYQrETPyc9FHdru3QamKs6LYy0YLBJ8H8txtW
X0AP9aQJvznmz7/k2SAtgJqLRfOAvNSH0rSpm0UcBpx+Zit5K/0+yWgK20JwKAzI
lKU5GWREYZE4NwbKq9EHWPAnzhKZaAAP/7PM/RjoYJX1Jk2oyT/Fy2mVX/a1UGLg
3GrNrK1KnsKyJ6iKQn4R+veEn+mEyy82jfhnX3RV7rct46nU1OxUZzXyx9QD7OHq
+p3sQW/u5WHvjDItmxDRv29YZ4FbRA5xcreZk3FX2me4iWhgyeWMu0zQVqNAY1N7
hc/hRTXCaF+kO3pvxhhrPc12YJnOeFSlostTUPJON/7lITYy/E2WUB4j/vaOyrR0
6KQAMW/0fM+A00TrjiPdQw0lwM17IVZ4IQ3Cg5u84+rFV27vmGQUK3Tu7LR/agSp
S/XyUkKx7DTA/Ac7tXK/U6gcYzJT/lzlDbJ5Fz0KyG6w2w6bg842NmNMw2zkvKsy
W9GzY8t34t7D7fRAdWEmt6q9A1uQGvpOZNWz5ooXJ86QaBHfAHE7l6PvuHf8jTl1
V0JzR2rfnchG3Jxfd4tnoTEIhHp/FJQrm1r8+/+kcmgkSqvxV6MHLIsr6cR37Qvi
qpJzr/SdefJDn3WVda2dEtWA3S7yBF5yFTx+BEWxWtFNFVrj1onEAgOYSMmT/YYi
oLqN7BJZhbQSPrmDun07PSv36FN9IEPGYjmzY12vUQxZNVI419Ps6FtzFOD9Zu7I
V9w0jyuxBsS7jUlIYXvTOO6W/eaOSZ7nLEUsJWpsoEygRFhSWZ3TlUAtj4gXA2oR
b/0gkXbRJxEEzXpG35CEbCCi4+vQLB3GD/DADrvTGfcgBl/zQ7g8pF19PY680atC
YUuqgyJyxcJURisa25uhAZAVOZUgpsx/q+eXoUjFKtmf2NPsEPY8OjBWW6UUl4ck
haV93Nuf3N+DyN4DODePXfY+GGkctmwFRhzZbGrooCV4PCzi6nk2nQtaPqZGuus8
Q6vy/0P/4T5dcg97d30ZENxeL9aUuzunckAm6/qlfv6Qfcpg+GNi/3luv/Rb58h7
l7cn8TswbQSStuvec6wyo2hXiqLFTBV4qYHMU0MDDjDlFiKpnbxNkLsPhy9jTdkr
XKFsm9EeTnejxr/6x6YXtX8Ls8jcGz8jNFZZ4ugbQ/vDIoHBeFEfPR2Kb5V9ENdE
6CRGKBReYUjAIU9BfWx1vRV1JiE7AfrBq5gdtkcCLucIgFr/IF2O6AOdQMRqSTPC
xPOvPpC5EiDdgNhbVcIOj393dWyWtBwch/7syoBSnX4tSwI84VE9G7h11/INHRPt
nhCtwwxM/cG7Lj23Gxl/UlwKjMQ5UVjOdHxmIwSJsYpw07eHoPMmqZzlqolaIwZu
AW1r5Y6ARfDO4sZgK4OAe97vh7F3VrLDtnoJR3FpcCn59BGn8Go2Rvb4GDdPm4za
6EdyrzEpKsMvRN8BCjP+xqlzB5CzpoMWxvApht2KWF6QhE/RMQDSxg5EdM+ntjrg
5ngE/Cj1GgQn3/+vkdWHU0cBfdr3wyO8ifneXtBaGyJwsfo7b0HVz2HOisbiud82
ljFU3hluBgfLZMWmCvIEzJ8M8SEPki2KJz3eSBARMvxw374O7GRQ32dYm1xnWwfq
aUCndzccKvrez85mfaV+TI6n7/yso/AQnHLw8vGZ2N1uwmdR/qmnmRagC8MkgrGG
b1qOETp6OPsQsDkzTtOEFd+sdGfmWygAh4VBF7u1STKR17zUEGkbbUKKF7T2e/qe
yP5/h98T1Jlfkgk2vkpjndO+BGjxNdw9iVDMTs+YAIae4wbTHGWy+m7UijrflfHw
6C7DgIpKERqUxIw8d4k3zbFU44LnbWgzqrgYpGengZcAoukPj1wagtQZ7LB4c9PT
NynwCcvfzBV5Nc7snbzinxNA8udp4Phvlo2qd4Egqash4bKRqH2ldiTiCc+sgyk6
SBkhs2hZsgRjqVaRhtbwIwqvXCufYx37w9IuDOJtv+WEMtny2CeEzgMGXkJSqnxw
l/nLU02uXPHP/PpJF3iMm/ipCNUmVRduHfC0AoocVmuwMr8tKhWHuUvpgmAPQTEw
0/pq+bYcWfcQrHWq+I+itGVzvhcfs4MUnX4ITH86QPUSaYfQyeGqCfCVo/bDaaPy
I4hSMGM+uvJaO7jVJjLXkgTUniKu9TXrIUSn6+JnnNNl8iJ7taB0KZ+M7f/DOj3q
LtJx5k8ji5hJaUqE2FgctrRyz2tXTnsCpqdfXrDpQhnC/JA9Gg2S1VTX05lmjela
PcHbUM8lJUN4vJG8/CvakmWNs6r2JIAv7/DCkHQaKmh3AbgN/Lmkdv8DYfzu959C
H2aiochHbU0F3OAHFMCVoHeSGgPWS0uZxQaQxtZh2olBpuaWM0MA81Ix/tkw5qAz
6qT6KE+a0CXx5cgn6jBVlagZ4zwIzL/7mmRD7JCUsHOF8fA8p1icvaXHVB4jcxvg
cI9MjdxEiyIX1um2sfjmcqQgCij8kHXkAxIzRBi1JmSlMTb5uqcFhuptVAP/GwQD
qbg+Ji6Wg0sKCnq5+S9xniA5FYqqZlizk1OzyuFfcvcYHqdsQAf0AYY3sSZf7lwm
StbpdHvsAFyH4cqovAqilpKVaXeONzV3KOu2rwsAc+gIfhmWnkH+wDO3BjhxbHV3
g/1IPUn1493XTYay/SlwFDGzkwIpGAlqVW05rPdjUqwolLKiBpb/Yr2NPDrC8bif
RL1mJpTLgX4lLTqBHPVM+ffTQJ4YBQXk1WV3AfdJZJUxAf7NIVj49lBK8v27KO60
u/dkKcHhfbP3HXOi63ozm5uNTwjM0/UNzSRNVvN0kyvETE75Fw6vARHhEHEzZXgA
BIUpb+omgjg1gfHT9tC51UdSWUeM+52r8tJi5sFA5GXF2AePcmrKK19nEzaFVfXf
tQabpriUFJR8l2dx/2IA5a76FEKf7ZM3ldz6mn6tnIhSJaIEPMXZPuqB9Wyr8SY7
RTKe9iXzyycYsvjfbGXWXa6QrDzkDMcrmV/bsW42FMJxSPy8ODofFZ78pmQcFZoZ
cmMbzV7DmGQRwEz8f68aFZ6DUs+rvxVUIP76zJITJABkuJdduvFuehRbSYkiINHU
vH9vHesktmWxOTwunUonORci++0GrrPuZRdIsS8uITEgBdOv63e9HmFLA9wYNdnK
Cd1A3xlGEHqcEXp4JkT56xTCkhX5UncDU6wwv38+IGtN3M7T5Xjr6ReH4is8U+yq
5+uvaE3XqUtCZcfVntPgHBcvfqz/UhwhV2gzGM1lzdxfMdt+vb7p6Hngm3jEIzEe
QHRrP14CNIrRvliKN6U7LjV0wGXuNs1ETgXb7Dpl+1zTjC+vLA3G2Fx9PMweJQhY
7vi7Pu0lbDsECbbQLWQEj5G2EXwj6/bdvuOx2dcY8tE0L+JFOzsPo71aJs8l70Ue
twlm1Y6xXwuGVPqY1C153BHQ6pDmWTIiUBVOb1SkYqv81WoOpHICDEc2hcOlDaVL
1AbywvgnlfKuTCQLScUFEs5I5+6mcHPleXLvkdsLLof5bYtLoYHDhLI3jADW4YpV
3b9kNXWmyUyZsxFaorIHD4rIK+oRqTEqk/imOI0wHKhGEJIQ8CXhdPdaR7eyhFnK
Cwb167CKipjpUJpYkeoObNMHOeP89kTe39CPALV2/FWp970Hd2xCe7Pjk03HS+0U
PRhpLjd7kj4EQGUBzODLS64Ow257/DNyZwPoAEj7JoimXjbO/DThdwElecw/4/MV
W1t/dwev/OWNa7oTkuy8qKWl7m8+QtVMPEU38HX7Lb668VeqkdMFdAqxxoFTKl/c
/qEjTtlHrHBG0ReJx2bPFO64lzBUDroyMbDJP7rO3gNcRHJrwFAYgBz4DY9DEtdg
EGeyE+aMV/510KQfY5C8SZlHEEuCb/hsW1NpsBT/KKIMvuawQXZufSNb3+i7tQUm
wrVqvNGcOuMkFh7Lohzu698TkjyWMzTi0e7f5KfUQwWOw13SqqCgb9E1YzQFcAwy
SRpZAYrELdCTKjwDUXxea9XfzfxKveQQPzMDoEY8QGGGlZRZVsIhqvhdqbMTtwLq
cknGiS+70QdYauNIvMMBzEkq1noPM7RzkUkL8SXWjRg3m6emWXJPG/UfFl90VMOv
uDgF4FLfOqC8r1yjpqCGDlXjOZntw3E/CYfcxwiVZ9yAHP6lytoDtP4Bjj79eDEa
NhDcTKa+mPwttkkU7VKKHxbr6dyg+xQz3b/b8nIRe0IC1u9luHo2pJ2ceEMXCpcE
Nzg9Tjjgr3Q1jrjlurpH1czNkieHmX8wnp4qLpbt1nA71055OYdZaElE1p+D6AGT
uSTHi2YN5Gk3qpGUJADwrvZR0cCsGNFlDbqGTRjjhYZDU/k0U9Ws3xTRJqP9bVza
CAnPJKe/eub5IalzQd3mQdc4xRFB9JSDjhXN5mAveduVrmMW1/TurxGAurMEBBRe
3z0gDQaHuDJFv/gWoEVyQbow+qnMUfBgiKauOQiOMIImmBPD396PBd4mc2qiEdz/
QuUTCTgLMpBb8LAs1ckHotdKixJqUe4sHXeTfGdVE8bNfVpK2o/wTw9drbKlPcul
TbAizeKYkGXhbRFZcUMNFJe9xgZfkfhTniDIzUDETG7vC7EyVwIpAj+HVdeQBUEp
RPfG+BKlw7GXQVmA9hxJIAygpffFhEjuqsIYDcScbk9oHp65eN7Qp8kIipCv3xw8
iAIO7dIJ4QTbKFNlI56OmsehoyBMqczwhy1s2jMe2WpVl0Hh/DNkStfZoPUk9tjm
csTWLqubXB7Y/5OByl8xEPR2SRlr8J1CI2Rgjl+CTHucvU+SxYrfiViaJwqioKYR
6zw2Wg7yW+lepD4zRO1lIP4DsVP5icUmfIZXPQ7SqAhRY2pqHepSOTABYS2c8DI4
zj5SHUVpycp8JydwHTyEb1eCoiGzsO2CZD8/kS0yIgTG0G0UEOJwFKI1NePrRue1
K5uej7bAHoYY8yFmJ2NCbXnxi2mPQhGKXhI41+eUcUj7wSCheWuHAWp+QhC7pCa6
qYpHneFpn4Gk5z2UF+Rso+3xhD/Uoe6VM4GO0tGjyCuh9Y8cyA4CYO7QfiEiTlkR
B8F10qKgJzKyZhFYlkczECatPYDHNKAmnifDqGJKlWFWlPRUM2P0K4GgPOl6uSRy
wy1AJhQyXIenbg/5sEVFWohks5nL/I29PVPplzesxathfalHVFE8Ioo04FYxw89F
A+hsQVz/FjfvkpnTvFbS11Q5KvXnqHm+XJH9n5JvI3RlArldWO5bH807hFYqfoCl
pJCPU6AtkfO2N8ZOWKKrwks7nCn9Npb/QH7bPdSX/X3go5R/AELWQKSJV2vPm9Rq
E/sCIo8mXzi7ak+3lK1+T5lqkujVumJPyCFMlpZX4cMTPwdExxwA8o8hP+GrT53A
kAt/nZ5G9srUdFRK/C5Otj3VOHcCzI7Bjt/60mEoVRcVqNhIfWr2h0Aq4aoLa8qV
FhUHgbHQaV315xihb5ChIpNEdXZ+5Ey7ATOTb6/iMkx8XCfswP7IIcExZNqxzKtd
Bxw/eNBVG8pFnBOOYvzk3iT7G0NJTe76S0sDggmiRd3fwUfjEtcuyLEpoIKemMIy
81f6q40H0JET0rn46H8DS+/zBivrUy/f/g01+nkzUc8DaGoesKHwUPujSldIbFtN
s2VpG13Tx/Zj1880lBze0c3ubsh3NB+FuJEFeFHvkD9FSHCeZVOPWkR5XE1ADvdv
wUhwTdr6u41LIc/SPIT4opG5axylQdyg++btXjKcOb7P7zRHOLwzHOskK8fgwmLx
RvylYR/UcVe+boNYYwYKwSQw8gjzmckSm+Qv6ETKw9Ak0CNBWSYsZ5YwoDcIXU6O
nH6wZdgarPCjm/Ll517jB3OZxm3zW/Xys2Dh1CL4iMaTgK/dHnnLduQIa6ldpoKT
t461YmTw3fprX7mxH8JNrnqmZ51I/Wy1R0Iyokyicn2Tz7HhYKL4tQPnqPnEqqVI
rqcjDX7fuQ4nLJAy+rS4BXBK+0l8Wy5GftbtrjLJ4iS+nD33G6Gprj37qX1WSV1U
x8VCtQLwCd/VArGcYU0v7Y0RQymXwOyUDhYYhXzcUB+ekTI6wOkAjwhZOni3Oba/
Mzi2KwIH1xTMh3lLiMVJDiVQjDIBGipSQEA1zilF7Sdvjblc6O/vUR2pJttIU25S
Sblg5AM+NFr51g6eL11HAa1se02uDVVdzmIGh71TcN5kPssGb3xoTjuUXMemfomf
htFKCWji4JaAdn3eQOjR11rYddQEFHWOXqJ5vrzi7aoZEOooxhaqMlOZWj2ru3bi
S/hx0UG/xttRmym0Q/kAoZejDvKZ6oUS2GZGg664W172PUrU67BiKJ2O1n2I2iJb
XmvlHwX3pfmg0Rn8xstWl4FmbA/NSfOW37yL9m7nG9/KGNzgj2cOglDm3LY2oZC/
U1HnqSXlbT3ImaAM1LLVIuBqDPbvGf/8oC/8W50hXNFhJaM2WBZEWuYqaKDWmDLm
lBPJu6lJRYDmVxMJF8cSaftBQP5iSQFVNcdfuObIwI1b6f1bC+uzqOd1LRrYaeK/
kjne6Gum4dAcwxHE4UfbApYfqi1gBddHL2lDsAGmD8urmu4qnMQa0giSZTc8qCwf
lcSm+WRPVkca1/9U/C8kgvS9FEDR9v4SPRClGq/7ty3sXRFq/D506YC8RVCibfpn
vDg631h8+MgFjUsJoEDWx0W+V3dl7ofm/tAsIeWwc2C2LNSP9YZH/gY0K3yEtgra
mn1kipttJq2dvMhHFwCuv16779Qh1KdhlHtnRrNkcRYRKIWY2rnEnR4B89bjiUvy
Vof+dmEar66dvJ9TeZyienFVBkJODbFTUoDhwxWewEAZC6IuF8DS/SsWrbfFrRaj
P/hN0gb4rCZGATKycWdEII+lMHHC8SCas3BJTUXgEdXzcllWFThuLHN5ASXcro35
oULBasxvoVmljNfuNm31YgQyJjUGSDTd55Y8RenT6ZLZ1kXREnEZwXs4W/7fdilV
qAkB5hijDgRRMAgNzDb/Of9O1dBdaPNZhjWnEHY+lHqZoopOXy3jkarVfAT5pbYP
qmNC+4d3aTrRsOLemHzPwjK5hXng6dq4ng8BhlaVOADbZRiM9ylfpjp3lbJuw57v
aK2NSvXgF0yYPNQVxqBxO/9B2uAd0Jmi3kuiqPVWzOhn8N0SxxYcRk6dZBH223EQ
RQx/GilpepY7ntQ666jQq0Q+OdOb1PGmIWaKHcy0hJMKuh7U4Yl8I0hTiXMXt81/
McNWCamHzfyDeXQMXyoOmlP2UYKZQp7D/5AkaeccVlxiCLeqqH7qA6rQRaO0vqF8
vv9M70P7OEh27+6ciXvEnBzgOBPeoKm2n+gNVnsem7n0gpsp0tuTNLFn8HJJSOdX
VYaiCQkmCftic1epR+3SBEpYOH7O3uwuFloNYh4zK+dchhmPRjBpmA2lOyglEJa2
uScHwptRGNhVK3dTe+mV8NZ3Ugy3IeTj1eVMV6bj/PHB+rFyoSN4JxsqJ2u8v6p6
x8AXqHSdqwYi67CRFtCnloIgYSh4Ts/4xxXoFTkW6nKw5uAYRcbrISwsDhaabVSb
DGr9QehjXmiEHPqdYt2FmcuK1EUArljASmeNTAbUADNP4gGJhjIiQfBQhgo076Dr
n2aCK0IXTlhXulUQmUZ9AbQCMILNkd7/rC2Dv7J+EkDCtYRB9SV0GUMnwLgWY67+
dPYNnKJwEdHoMF3TLRjVkzpUhi1pBm0k2jFiNC3aDNg3dftxtXFenRa7w77n0dJc
vLW/vrpozEMW5OWNp/PXPlQr7uiqEvz53kRFyDdWYc+suwws7TyFV/qRp9PykIu+
AgQQGTt/XHbRjaPLvP2PXUsXo8itlRN8Pc9Tb56argG4spnKtVBW6/18ii5amCZ1
eHic653XAScmeS10SGpdhYhBrpxP7lQQkKmtg/2gMHh2Xqmk8rZ7k+7MqA8r0BZB
w2hJZXmLlwzqs+xNtzbfjLUVUVyMSUFfxdXaSv7i3AbpG9x1pBvkqo5ST1wEBDUd
H9acuWIW4bAfTmlnT+quBrr6phyk568GtMYW+No9kfGI4eW7QQEspoGfthUsJORq
HY1XaL4cwAtdazb+/JSvExGIBu/LvsVwt+AoengW7Fu6TVE7ldHtOmR0sqY7ga8m
1YA+lbKBj7cYyEql+jd/u9vvj9wI6C61LOIFJZMBw/I6sKC/e692it4DheF+g5Dh
xysolRKM1DOkA3aSC53M8Qg/UziVudbv4GB0BCxVsTpWu8Ite/FM5FFUOQY+QfSj
sAu8dt1oiDJ98Q+ktcmmd3Ba7MprA2rRLncXve3mfhGB32AtETi080lqY24oRGQQ
SQhn2ZjUzKdRDQxmn3ineqvt3Ikk7zf6J4yCZoJdY8MLtp/yW5B7wkVhksFdE6y0
DC6d1TIHJGJuAVgSh7oS6+DU4Q+0YYOimApUivtMr+XEAt8s5siCuCpukE8IP3Nt
sJcmPTA9ErWTOrOeIBXFuGOABNe02GkzLPnfU9DRnwby8TYw6DsyHxjyPoiA4sMt
OT8PIAw2Ix5tZb5UKK1ZiWv5Co06T23ewdE2QbBW1p6o8oyMPVB+EjVItnkDTggS
ndJjOanU99G2j9qF5S3Yi6kVY5V5Qe/zPgo+qqRm5h0QY4KYmQNhxV0bLC+tk3Y1
jdSS2WkECkI6Uq1IJYEGWve33VtU+AIsnjKF+9hC0f3MPCqz7nW3BGyC1v0mBGpb
19bWaSKtn/ABcg1B45kBatyOclLP1/txS3MsmMrIBUByMfTUAJ4rHOigIT1tdagE
rfTCbm/wzuUU7yjeNZjcc6hiorq7rrqUVud1I7xYaFEjMiIFBz4ZoYA3j3GiUpJn
ZBpvX8XR+j90ThLF05Lptab3h/s44hGGxs++zYs+aYtfpqyfPH+jnTgJdvuhv3fk
nG7AhEZ2eSwX14hoCvDsksjh9Hmp0jwUeFTgqa2rbWIoSYevrMVAHbvrmaLvc0k3
c5WOPm1L8yudCHUhD6ADaU+A+z8Jw4A3CfsoesQBA6pr4PnGlRnJSPsShqs63dWH
gqDJWnasvXQcb43I9/5677yOUtxv0AgTXcMIhwjB3XIO2/yjceo88CVPX3HSVZkh
XrzagUnIPUXyiBBMN+FP16+YX2Frs1/txuEgWRUzJtqTO1d6iNpfLOh+FutEQnIw
FMyryqZLWe15Qa1uSyyLPdhfPXVW5a+QDuAFeaPTM7x4guQ0X5e/0A1D/r/K++I1
2GUuIH4DeWctQcPljBZoskQSv3IYw6GFUvcwqiq/262VW22FpiHrW3tDeeS2pow+
3GIn0ntoYImVqvqo51eQefsCet967Bzo023onizlMPcLF/dSXi3Ry8zuUmEfhJy4
yA1Zy6jh800PNqOn88RiOtyoR+hRa6RJfPpV3SGJ7ChYMutaFatQXh+OI7ZuIsAK
rVlDqUgBVEI3ISvj0pEG7TB9h8a1pwLWUFSOitwk8cSy1zCtptas6rt/wnmRT7Cd
R+i5+/KOdThfLh71Dz8BFC1tg24Q0sg9GzZu4Ns27SR5Kig1bHGp/DmfrxxAB2NL
03nrwI5dqWxpop1HZrk3vs4vF5puMNXYgawR8tabOh7043memPIj/Nv1vQrq3mJy
aKfCD25RikHS+dedTs03sgfri9q9t+lO7PCeAOY9n0t96u+P/eclesa2SL/hU+pd
2u0dl+sR9LeRcEi+tiox4Csyq1+Zdm5sKGpWkCRhneCv0bglyR99D4Zo69hM0rFB
+EXFYJItzCCP2Yioh0CofCnIb+4wR0BVhcJmqqIwoK4XnaBPazxq4yBrA+UNNPOv
uZ2M4qLSL3z30tBvQ9YjinzImupkzBedfYoiOIi5xr0f0Zi/1MKRjZAFXU8bp90W
arkxDoPoZfZZey3JpUpJ4Scui+TZ82kPyCOCtos2Uh81on10kWL23ktsZkr6eydy
iw7oY1b8C9I+C0VwQysWrAtpG5RXAEUZfJGOvX/de6FJgoK3CYj0c0s9OqBWc+LL
t4HN9FkoYoqEBOV72aE8RAzHMCmKFuUreoTVQcJnHYFV8bevZao9jKnFaXAjmBNX
lEB3O7j8w8vnkcrrVNnXrSoxfFi2dvzz8IRhcG22kyD0WNWYYsbXtQf64sHDxfpQ
HGWoWeiBC8lOgfjMQE0LlfY36LR4ht5HwuzZAQN6CzqAA3r0FSP0c6+AXVMASINW
yCyeMeeWYOk+m2VZCGYADoPSfR80u3q/RakdeC4j87blcHA+eenvpPW61rlWQ3U8
LlOZwjVaY7v3UxQvRTFvdGmYwo7xPTB82f4dc/IOfmd+ohQMy4/8yvh2P9LSqAKx
ddbybzcSxN1/shh3ZVYaNGg0eLNGSJ13E799gbm98BxMsxBIXYeiisN/5dsAdffY
q167XXh3V8SoVM9g1dQ/FNaQPeU6kd6+Cw3+hx/saRswp5RLc+vt9wJ677P/CnU+
Pq8c2mdygwIBRcMXGAKyjZfnTIQNFEqA6F5rrmcJj02nGDa2uqJYt5Acosxj/rtD
mH5pLf1jhFid6pXyrYU73aguKkvqNTXX5AK2id1tJfNf2FSDhtjr94v8l+21qssF
KowwFOVaSwmUMrFTweGCu347no8sjjALplaZObleBSHDb++QK3A+ho5QajUI/Cus
1rxadLxLh6LtexzIRNp5je54hYwhRALf69txHkn6kvNhQvLWqw05YkSB28BVZ6e4
P5S8Kz+gTUggbGpl2FwUsI+Rndjp1Ystt0FDkZ3BEJRit/GtVFtpgFD6X1EG6Ac6
nNFCnPH0qMbO4zGAokNVOFPzARjz+9iMvUbJDc2SVlzVb85QO6jSF513ffL4iMXg
35YXZXZp/Epffc5mP0E1piDMiufeZa8tDOPozkVYFfnvMXL1HoAYGN/MnOG6YrJQ
asLae0t9GqVdgjjCmVF4Nfg0yPSpRs6rQw2D7kFU10DIVhBNOLgpxdgPs55yjluQ
wp15GNBlstiCqn4WjJ04uUZ+X09KnjBbICI9o+xm/ymMwLMtYI+ngue5cgsWRLi+
R9IRXdAT6TrPOt+nPID8SBQNvvVOOE/kuGa6FpU+4XxpxZu5avqSk+waayE2BiAs
Z01fkG6Z01aWU8mzWeuKORd1a/ovCieilUIkC12vnwExOQwjJIBfKdCqIF1bnbln
+/AjdODXHz005mbY2AOEtHo9UqUkD88xLd4sL21Xf7FmYCs/6KlGEI6Rqlnqa303
336UVZ6MJ9BwRptYiXr6LyjwqaVXGIexR3k01NAdn7Rde1XLeXZJYr2ROjp/M1Ne
PZK+gZITK24CCHx0kBL+NAbpaBENNRtEzYZWxlPQCKFzEoEV4HE2I++oyyp0+PvW
xbspdoTopWKUw1zRnwkzc1O/N7VSAsiGsgUs19/E7kdRw6hWSnvIKNHZzPEXoN8q
sybM6Z6GM4vRqshQbvgtdLV56/265e4MQ7MMHMA64cwGqtlYo5inO5JpF5Qfbzbv
2tEbDczENM0Tep9vMqPLBSkGQbI3t/a7yr13RIw9ybjZptMRywhZ7dD32UVxOZ3s
meiopj6LuxUeFZl0KZ7J1fCAuXH7uBp669GxUGvJRycn3am/v8J1uK/F50QfH48w
TipEV4XeQFSGMPHufIQkBmKWlIDQ/z9G0TbUPXBRn7wqrWdCXeodAptQ2RRS7/Er
91tohvjptF5cJSnIAvCal7mGn72GxEuAyUjqS5xQ8zxMo1Mb84B82rcneMfxQJQS
8a1pNndyyTVG5IgX9T1GOqBrqa7yHY+CXjVxdHoxdXU0BHStEQzZ+zlOEtzQW5zX
sSbpjF60Ok/Wq4JazW5EnZejL83gz61OAvoS1nVRAEmrui1PGFUCohIRCqGJSsr9
4uEpkPJnmiNDxvXS8t7rGLOTieBP2+MY1+Qo8DrFP2iThBb+KBF0WDsGHYenrJc0
zlgFlOIVnZZTfAXvOTDlccQUUOcHuOefYSS8x5TVuSMSXXXg2ICoBfxfO+ZfA5mG
PQeylEgaZzyZtIrA+bXNTgnuB5dYCScgR8zHrJLmPkyJfn2Ymqv/hgnNXB0FUCxw
bsHomtQocBblpLX9v0lJZAEjIAnt/MBxdOlLMaCfu8Y42c6UyHUHwCBLfownuYYa
1L5B6zzoCTkWffvwo0eFg6j6vr/stP6QjYZwvwXyYBbHCjZc5k3Mfi9OzK8FpCjS
NAsiFyvYzqbzU7S9OZZCzhhoYkwtWOt1NFZwu1x7/TM55pgfyPWxQlc4zK50HlRo
jb9NbDJY6NzZ8zcLAwXv5UIVaBRZAQo4DhTLVMDoTddAmKKleZh705CRYOPvvJKD
zew08PRDVOgBEi9DYLB+B3847t9OqMwmzLGpAQbJ9WECAMxPy0sBI0s+uEmET7Zw
VUU+JxJftbTA4CUW+1SqVwtofwf+HFzNZ1PW7oPXrEZ8mxCN6XOySRuQ539uAzj+
pgtCj/y8cpGirdqgu+3gIzdp6wE+yBdbjZHIhxNHkP4sY3XilBq//I4EnDeHSUP3
nVcLlW6IEuOwabKD8nmtbbwtP27BxTAkv38t2a+8bITTmUUJ+MXk1nx9Tzrfa15L
O24X7FzKJU2nuLVo869ENKQ+8q6V57rmtIfVAi4IjR4hOkNXWiEkUy/WXu2puU99
LgZzyIb7AfxnmSDe+TGIef/ApQKQpF8ydHdEFJaJDZ2c1CXEMmKiPj8cWXp9SCXM
IOU19UiIyjBZCL2fpKxbZCGJerRrCKGYWQBBTxhkJbvnx42VylmPcsrN69GrJv1X
PzJbGEeV8QVhSJ+wPSK5WbH5ie7PlF1Qjc0jk6hXHNxf5NkcifDYsw7WwipXBInd
bTDa5MHh3JhIVRruc4O9LxQR0Yc4gMz5opyybPfS6C0YBiZ/YkkKL8hxJAuLjKfn
JqOOEidQ2qm90tdi6JRhzluOs3ZyBw7J5ULwwHpvFgKQMk3YIzxcpuNEDwGyVSPF
+VCu3agXvRJILmKTUD1wS/kW188HntNwPHHml6KE+tjAmaQlwAXb/bC9BUheaUlQ
7OXCRVVIwwQe9xB4aBObuvidMn70wc2tSoMfxTUSYQ7K/yShD5KwU239BmCucsbd
5wnwy3eVYCJhjec7fnhmtWNUcH89u7YmaUSsIpyX2Mpye3UhBMCzPIh+CksLzY1g
Pd+RDg0ss2iXhWlNnQ5TJ79vAwh2otTWATYqj2AbatXrQK/vGHaJ+eroAfUUNd4z
ooYxXnav4ChEu5ofFzWWkV6qqAjvqwOnmShTEMWJ6bcEFYevBA6Ji71bgB6EEoNM
1sSHU9jY/c6XuHpyNGTh/Ui+DhfIBUXs/qlKpTSC73Ite0BFcFEf4hJ92W/kOCyg
3rlHuXBYjX5tFXvPU8MV6grkqbYonBSZsspY4L3oLJFYFcEcw9bbKFNzGRh4PVp/
3LXczi+71bWH9d8GZPKfHiIQ1SJAGStmgiywA4/aMdaYxguF8epi/wddbzbod6DA
9Q6NZYFUkq+frw9QZDOvglC4LMkJQx9Be2Z1zG6VxwcPYK6iIIy71g/ZzhSMbSbc
M7A0qgaJMhXSjPFoSaUJVO99CTSqh6eTMZbRnbsdf5k8dVwmHvwCSoUU4dH44pQs
HXnkgTVdiphXaGsrvK/CglDFIqGOsphk9vi63T7+5vC2bG9ZqTPjWvj0+YuScoVg
GGMRyxkbQ9xvJJVfG2J/p6P8K3CT2cGgfulOCQPDFtHYRUSoNZtA56VGjRPPv2zh
zRVWmpSs7YfcvSeXRXAy0XVXB7CECRxKNC/xMTHUFKJkSIF/Vq+Hy+En7d55uWag
c4oN3pO6xUUx839BlJ1onR2lJUDwj0KFF56JbzWlfJn1U7I0mMk/s8l8cp0yspLu
dl8Waagvz3eu5xgv6aGSF4jlyJhMAH/ax0wq3UMMIG/kLb8XS5AyT7jAhD9g8fan
wdO/uTbV8lZ3bmbpwKwzOEI40oiwrpVJdTmdhK13yKTlo4NO7pPsCPeyN12AzOJc
mfz1K5JIqf2E6TCN8Y/5muPIloy7Ict5lDb6/N3E2NoGylxMq58JAJBXCsbOh22P
T0Df+dkc9JPIrnvpZ7X3V2dY0PDMtHq5/m637mTUFTd3cPhXWEsUYOS/BrMBDC/M
6Tk5b2IfwFBrhv1R+01n1dsThB0oP8ywUFnk54uiyDdR9N+DkQ1Y7vfmPOHeRQ7a
S6NQJgF7J1ddTz7Lb+Yo7SrkTvUriNzX/nqfZo3wKbFjwD/7hZNfUXO8oLcfZIRR
l8HEumIXxyDmYYDpLSXbl6NmzwmSuXsJ9p6YPISuJ4vv4dVN8A5FZHei1CVK780V
YLNznX+hXd0UrSqgzOM28nTN8x/dT3wNiUO85u3Bk+6aj2wxgfwkkSpF4mSfQcgQ
jtttCOV0yByq+gmw+9fwULE2PcTvkq152Vn18aH+sQIyKnJeMPOunK4afHRwfmJv
YlmWYtKEUVf5EJVnx5wEb2D9ycavx+JTinBlI+ncL7mxkY2CyLVOXvxHIojlsZkh
PsAaarh/8YQn431UDDhd/Ms8hS+RnGIM7EQ2fV3Onq9YUytXEBwkHB0XG2n+gYaN
6XBjnL/L5lXUufVaGHduqC8MXqGo8UNXLETiN4CvwynZr9omaCZxl6+3cDw1oKcx
d0fQ84hu6CChyyPkeQjm9mWhDhzPT5g6ejnzOcwt3hYz+B0hg29b8CNxNDzejhRF
O5ZrWloxPXrqAms2DRIQVztOTAvbgrUcqoWXlJMEcLRuWCNKrQjf+9nWW7+Q661w
6kaQxOLh6Kj1MV3zuddPitj7ky7PCR2+GoZEnS/L/sSQ3/PRI7HFOIY9DtfwTrri
YU3DgemIzVtnkdxh2HQyf2e8jMx9Ld6YLmtrncayqMfxxiaIz2k1eDIz3dG5onB1
hviHJ0HB4c6764Xb9pN9xOBDUTdReJxR5zKNnir2aelVfeqRPRmeE1JzqMkZ898k
hLetNJ/B6Qf+cQi7tj42G40rgFBR25ZyL92m7X1cfq810QJPOOaZBphK176lnh0s
Ig6EsIsQ/WIcHroLBkRBOVx0Z6wZNsB/mFCnXLaw7/ZAHJ4gCTUFXsIgHUW2XlZZ
TeLoW44/LJ+R7UU5FSehw1fCLOraqkzfVDvojjIeAdt0XSyZeR33yuW6HcRDS2q6
WlUtDPpWXc6kPVvMKVfnGRJ8H+kC60ie+sTuzTLDTkofP3ULs3yV9s5PZ7tgWvCz
72rpEt8ualehwwX4MOGr1m7zdjwkiuxxgFZw7fo8JE3q7MvdxE9XMIpzi/BzjY1E
C4GdZFWjpn3A7qpyeRQkD/kbV7i3y3LH5keauMUSXBvxwuS6As0pnPQQ1/04pW/X
kaj/cYNi2/BxchTXeL1x5tbHhADjnjm/pJMnSMSTC4Zmm6aMyyRdgPWnEgzbAUjB
WMxVVAC4nuQRQ3tAFvSGfmWdsITvkhRX3U34VIvWZiWD8G1cnlWwTCTbG5gcmUIA
b4mvYoPyG/1/ZftOzu4lbn+6SdgQ7LWPiKzsI2KreIZRDHqwt/IAGiTSbEtmfy88
v0GieSMSPeMQjQPBvU6PJskviLWhCOZZ/z4KUUinW6FRXP0W7cVRhBVI2xIs/qiV
63pp0F1CD/q5XPksL9v696EOztcqXLYeRUadzsr6OQinNF15wQTIny+0zBTpZtfc
uzwOy9UhYCj6OeICi30SSGiQZglyyD9aIw7aHm6XMHZRUKC+BaS+ng1aR8ubPWYa
4jiesgG6bIlKvz/5iP7vYCaY6+ssVzvwmJkjR0hPyzAreJdgNXCezeXKQG0sQMKY
6I06RHTgy9BfOsXzzO+4dOqpGT5P5+plzr9nwuVTQzu6iHwALc1/+NKo1JUsMEvQ
NYF0EVs1QbhvX9du8FFFRBINvbEv7Cg83snKaf7gnthNMV2p/C4kJ2WeA6mpT9pn
P0kHVxYmSK9dYRoEuysHogONTf9k/a+LsHBhqomuvocvF2Z58+7GhFNXXRr3MvNh
9WF+Lsb0IfwOIKAUuzQ67oNdKUfQa7r2CfQdDyhPcKSZNiDaQp/SOz8sJ6/r//Pn
d5BhzPyJtCwiS20Sh3HM4Sh/6dwILELcrG4rVBI8D1WfHiQbGYeTOZIDhUZPte1w
LMOHgOxftgySBzJAIUpDQs9UNKfjLJBO1rdiPAZ6k1Urybf0wko6l7tHXSQgoiAU
8W7BvuGAk7RxL9BIDodjvJ8txeIayStIqrcu02UQBwlqz56Q5cQvEPxti2lZ6q24
txmMJbdqE7YX8+Nehy3XM+Khj5FLj6t1hhvIknH0Udgs8YgI/M6KcvfuQL3+wSrw
BtiPKXEg/Zn2OW2pcVtfcpTeONWPWI3d1lQn7udQJRwGuN8Wa+a7jNW1qTaneqKY
eV3qm2S0D2dVHIE8b1eB919Th0QQ6p73d0FDl8nwhkYBbM0Xf7liHDUMK7UlqkAc
F6CwT6LjVfx+WP6heWscjBZz9SCXZ8WlmC1EdJ77vR0aoBNKOUMukGD+hQ0/0tU5
82KGiQW2w969w5+iZ/7Bxc/bXgprw1fAy89KCcGPz4RZQp/L+22GWfu0skGv2tEX
AeTmGPDxd+XIp8LCOgLP3oANyKu7RIqC5dt+C5dE0quG8QnTo/aVu1Q6cjYNWt9n
VoTyHmho9vnIWvusIi7XnG3hi4URBz9rgmgOWwGrK5QjmjQX24Cmd1S8EVLIY4qw
I5xumgwF+L1rx+yGQzIlLJz6UYtyxI8Ca9hZxXRBx9UozIp1MApR5jFp6Bg4+GX1
xIFiU+044z7YRzH0Gl4v5sjAlQoZbHrQH8DXtyU73jQiEUal1KHI7f8k2uxWmsB6
b7kJkYM16bl52JfkY4HYkzLU/09Ey50JdaX2FYv48IvP07Fand+p5hcBV2AfEmBg
HMJ0CHbk6lBtbvgkUb54j/IvyjwBIRM4X5SJ+4T0rhsfBbArmESe+w7QQOgYbtzO
z7HjsY7Lc/RlmtsZQ/pVsWR+xo87+I+iDIJbvtmOF3TGRyj9hrNgLn5Y7GOxXEtT
figsNtSbdrvitIWK0eNwIT7q+wj51aiMB78GNFt8OupyTrhCkErTwRjdovHowwaf
RJ46y0+cL0QBqXFkePwrOKnehYL+noB4B5u5mhfxCODkQkGp0PDz20ExLs6dmUJ6
6bmZKHUn1+OtZxVRzzYEisS5dFDqKzmWA+1s7SurmgCKQlMuQqXqvC/K8Q/QG2vs
v3M590mu7smRVVb6NWsmfx8eC6ucEYPBV8UpxPhB5QQa4JUQcbBGNGf+MA/zCngG
L42U5cssY7xCy/n7Sattozi3rWCYFpW2gxNSsyuacgunh0l9rsp/3WeeqGBZp+qI
1kHoL+8isznnq+3Fd2KjTSFfciOw1RXISY7P0s9q0qQNWzFr9GG8vvqNYAvDPvy0
ZcQ63SQddLG/io4pJtSK7LnOk07aZI9seiaYj8Q/b9WUrwxUSpAYfhJlrx3drM+P
+YG/+UTKe5WRJKMhPpTOYFOEfxQwfQ42cyhHny2ud2KW9lLpGJPDBMgMhL3AMpg9
pszZwe7DbjHVD2GTkLaepjOL3wn7UIIe5P3KVBf7rk3nNvldlwPawt4sZG6bnyHo
qdovL3xMpyU+IqHXuHYI0oCb9hAFUWCT7/scpthNuc4PLp459aFOI6lkpcDTLIsp
XhcWrjAivwL6DeLz3dv7zlcymw5A0bHV/jsA4F7+TF6vNq+lYnLsXZ6AygDa5e00
m2mqZWk4rWO7fJ1lftLSOMMunp3R/cD5zW+tyFxS58bIbprIuJ+dWp3bS5CUL5TU
k4OdCu2t7hdpTG6RmFl9dCWU6CT1GTdlsVgMMEM5JplFN8oPai6BetH7o82PFCmA
SqTbbWypxGNv2aaANlIBnnuUjGV3az2uNZEI3TJKswqVP9IKuXpI3Pjq2hvbB6Wu
YzhhtMGRhUPuh4qA6qiXAGBUf2R8WyBmZ5cEJOG0bu1V07c5FC12Z/x7ZW11ntTL
4zAJmv18TM8fZ/Eda20rzaToL97cc9l8JmPVflnDK0BV9QPf+PH1GhA9cqrAimwZ
pqetsT8ZmaRLCmDSWtJxopBZ19mr18jGTtwts+lDOF1NW//ew6KxX0Mc+hoQuVz0
xrrNmuMkPaz181G7wmzQ/Fi530KZkUqoARHqRGZGf87QAZGQCwL0KqrbyOVd5A+K
UQswCbF7EtMWQwcvzOxfNqDpIcPf4HJ/YaaiYFyMgilcKxx0pGf+naL/icbhLnK2
BzWp23lpMA+RLBDwXYq2Iq/xg1SSrwWWynLAxbaFltf3V0ZiW5OJljFam+2cNvr3
Jp4C47qzYTKpb4LkB9GfS3EQ3A+mIXOOvE4pgh0YcU+ceDctOZ7g/+mUUYOpOe0a
2BQnm7iGTiBcvZiuowJd6ZsM5QVNHNMpB0wo5gEMMtu+Ts8r5pYS7fCmdcRcFKCg
JnOWN4tfK7obrO86WDhQqftbIOvP6vWllxCUgvvZ980os/x8ayhqk1Kz8OISwSGB
UZhJ1xSEiIx6DgGbxGO8iDSS6DlmDGqQ8kEm1BWzGMxbaRO4tarKaHUQrd3IBk5r
6/ZzAxDc4VkrADNogPHkeFCXkrNHuTvRXjacAnJJf3IgzxjAhydfPjVBHXBYLLdq
FTHXHVsyVGYB2SeOUsUw3wEgSGrAFJo7Fwj91ywx3ypQa5SUu/MaPHPQ0hNivhlw
IUTiV0+Mbf41ghg7P9+DNjo/gixylkborqiJ+9PKEKfbU2o4CYdNQg8x0FpR+lHF
H5x0MmbzFBz4JY2JfCjTVRd2vxIfYRijVmyobu8c8DeIYBlEGbXoeQgheT8J8UNt
/7mVrsnsXVlw8O5096w5JUuKBrIGFWpC4iI2VJvmVGZheilgNDpamlQq3BcwKgFq
Qe3/byaDKSm5R31Ee1o9brmVNDIGuEbO//Vk16f9vn3UH9YXzSNAXfLyBmG8BPDg
ig3b+LInkWGW8YmeMy7JYJVCtMCksoECUHlVMZ8d7FTEjxxxTjEPVsuuXcIorrxU
UHzgzN6AboutAgvzv3v/QOjGwXxff8u/0ryxIuCQ4G+zYg9OCTYK6QZEtLkHKXgF
VfmthO1WkTRhqYX0u1WwxF2BPxtSJmNhwkdaIYEqzmyD2QU61fl/EVGZG5KC62xg
Z4+n6YDnbzJQgXTZuKQg+Rh4ldZxewu0G7+56ka1gSOsOwELNJ3WTn0p+Pz/zdQp
6j/Xzs0PBULC5OQtTKugbSHJT5uE2ohl7SQAMb21hbvdtiWBNQvbGgxZhb5L9nCs
wEMoPHCtgtYAgHB+2alYqBDaE1ESngrHh99s9+xMSuZurE9+Pwpaa0bZF7xxerfo
dAFmdlL54VSORLDJ237fhQz+O/QT6mRZoetfyHvtXy7X5s+dw+mcWi7Og4i2m1RY
QdutXYDzxjF6SAk9tP/P5KsolI+uEyzT5oPrGUQl8GYbjBgHAKBt2kNwrB4sd8h4
fV4Yr3KNKn7bEe6E/56mB9X2gzNnaln8NgvZUTfRayBz+g7L8VtNoRvSJf7XHWcC
+GUqJW8+N4lc27F4ac7hkCuPNSJqxXVb7BHuQdWEnKKzmOIGXeyCTgRN+OEY/pqy
G/J9K7Fi27hLKE/PE8edX+0H2AHAnanoq3KdWR9YkD9SgXcwOcCIMKA6+5faZVl7
JHGKeu9+5O4jJFbJxOgoKk0fH2f1uup8FGaGVBC5c7QKhtLoag3Bs0CTU/xo15in
gw+dx4Wsdjj8yWjQdpwS1uHAUwuZF936Pqah0B2ahVBGUMhi4UPllsKVB5gneaPZ
UbQgGp0hN6kNpoYPX+yjaJcoaykpONm8kQ3BEaAIrL/J8lmnIIUhErgw988Pc72u
z1bGVvEBjjr39gagvZsTGRJt6Cfzy+ANWZ9k8WvcAraGV5kmAN+eSWBKLls6i47O
JQ5KydahM9pEwbmxMeW/uPVQqmnklfCCFez6Isa0tqWq9ZKwDU6Wvhi3M7TDjJmw
6EZNe/g2GfqHmubikX/ixDQjRYBpfU4LpBxqbYG1zi0NFWfIxcaQ+jZggiAF9qJm
tEAIwM56qSMlUN9fBON0PSyLBuue6wtefR19vW2TnMrf2q4XIGe2qD0Q/Sy5jWDH
3jHv0zOwLDZ+lxfQozuNEljfhTm5himHy6ajZXqJhQjC4jx8WK2iJhGoYtgLkIuJ
AY6RVBYJuLxBq3sZ/ca8d4VFCan1PLhM5eWud3fKGLhsMeMvSTSzJA+Flmxc/mR5
afOYVmh+BB2uGUjyA7prCz+7UoM1nl6FMuLkfbrkMx43t97ahNoK3pJnuxarfXzv
3JaSr4xSeMyh4ECk7srQ+p42hEfMaw4AxhEElRxCT+Gov9b9Tm2DHEx8f+yy4jc7
4KlhVLg1KJ1aS5bpr0nIyB8kUz0J8NyoPSx4SklWRjKPUr3yu3r0DTOJwPn2l1QV
UsXaV1KSMPA7KNR3EogXQVgJ/xhyAN3uDudTlevprCd6fwaj4/arJvQDsVf3Oqte
e8goqJdPlVbM6Xr0dcsiLmW7HoQK+nCv8+iTKll15Xo6b4xG6z7gBReezLep35ZN
zYcxGAHzxlEbO0jJuQlW3eut83MIOIiOvd59foWnmTR6HLI9TfL2RhqeyJzCfEVT
ZOfHmWgP6iQRwevLfvzG8l6p49fnpzBpUVLOWbtbaNxEppe9p4WxyYORIq7FNBw/
78MZfR+vfgmn2Aiohue1BavUPgv8BI2iaDrWFxG1XlAY6TeUXHMQ9v8wh5ZcGW/w
9Xoy3t+yhiRroxjgf42+T10OdI6YioeDVnTIwDTHw+rqigHj5xL5BxdVii+Alj04
R2G4ZW3kz8PcsCfe14FAOZBMY2bLXFCF2uIBoAyfVB/egoFxhtFRR7KogcZKueYw
Q3X3JoUGr7CqEyS2X3hsKtJYRIWYd9rOD/HUh6a7Y64JoyZ0ARarcQHnT/hiOVLb
//pragma protect end_data_block
//pragma protect digest_block
btlqXwB9deqrrTEP4AkVi38PNNc=
//pragma protect end_digest_block
//pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
c35rnGiE38d184VGxE9g8yyTd1z4STsUSiFitBGYh2DhcoORfvqmeDWleKUdczuq
pWCsShmWfpAIdU57ffWx0zD+HeKkmiiW8pCYJaB8uruU+VP/VCIwebCpMq8FGKJa
8s6h7UWJOqr9Gyw4NG04PPQSQrGHCVPrGbPcYl2nwPA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 52432)
UZ5ulg+/EJROJHSbwQQKvF3M9DO+Vgg3SY2P0dVyGeQ6dT8/cRXnTiKNaVUkLa3U
xE/GuEfOOGGSn2YlrxLfGqrjakp69j6Yx4btlZWVKpfnvMGgq4L9E+iO93lS4tR/
Zfm5TxA/Shc0CjFiUxKzEM818eMaSQrb9SAdedgN8s15ASwLM5dNdGBuupm8MFrl
AIP23YTRt9fMBxA5SFiPdrFC8uYNURl1fypykx9bcUUGn5UWBKvyVSAnh69g2e0P
8sOsiim9IbZg9Y2qSofVJcLL2n/5k8kgrrYmQGvWUiBcyvcVjh3LJzJv/tBC+DIm
qbwIj/F2WWQlNczw8TiB6H/K9O40ZXLj8Ml0Nv7tgjhdMWThSHZ4R11DoVhYxFsP
/LDSYuqA47UfZee/JtSoshsF8B3E4B8MxQ0fixtirKHG6oIgYStxoOi/MZXOlKNw
CfU8j6zA+cLrqO4Eae6eAHGnwTUqPpBn4hxUTo3D2M7ad0AnArwaag+izjanjeEV
GgvYMHHFUAqgVZ8xLHB5SQpcN6cU7lr7np0uUBVOqrrIF9ZcZdAzjoN76sSXGDuz
p+Xp7aATUjvoo1LFk6NsgLrWOU/HHtklLdJNL4L6ejP7EZ23Fw9wGcOSlpETQ+NH
/GPWWCj5GKAus0eEcYvUGoFCoq8b142ftdt/hrqTJdL3NETsjciPk0hDVV6L9Sa+
EcfESDSbc93wK9koLMq0LDS6JcUUtbYBzatdXxxEAdnef5ZYWUg6TRJigD3FP0E/
t8zDRqmlXPg/5P7TpeQXqOXtbWJhT2Z50eJSAS0B/5VnnJogrr34je9qIco6ZYy0
TF1i9xLwHy8y+1BUVebhlL2rsa5l+8CWT9tr1Cm28EDHh5rdBj5qZ4LSkm/R/xBc
BR68ZOVChfmZhMPdl8rao8X6+nOPvFuhkixPBdsmg35e3bZBrCC+vEkVdqNXsIrz
ow1R5rEgCcH2nStBty/3K2ieGQ69uLMgcNMK29hZwzzMHQJyeiPG8zXUJgYJdTnK
u/a6ol7qNkghyHNWP6XX+oMZFIBplKi/T4LMzNSagPJpF3OJ/ZCY0B74jmU5OZEj
GFuuTUOQf0ZMXc7YIBf4JSASxcxKVn4mWdwuscXNb7OMs1+Mb6KJrr3j7TBpE/zj
ucf8dSNfCLJmtJHPj5P/JjgrPDdyYqcs0uDuLpeArxnt1Ee8amI2QRvq6364hOMo
Csd3pS3d8xNSaG/SlWpAS86PAadU6lobg5qd0U+g7B9nVgugr42QlmWjvtJa1arh
erNuuRB+qDk+kuPT4bAxWdnuMgoDQD+VVxxGX992b42lb6lGNIAoCuPOGG74AEEF
jqq87JSGtjYj73svwVqjdW7kC/jpkkru+Z/Ylhet7WjMXJnw8BnYbdRKT5LBZ/EJ
IiLgUzb02w1SIKvi69TM8tJOp+0eDdahuLtXCl3VU5c2ui8H3PwhVCjBMk7LGv18
3zYCfJG4BBENtfvXf0vKsYw/nSOqjz6b3S2Nf9vFkK5NtvFmC0brRcZmv2FMo1bF
oqI0i4Pra/IfTOT1rG9326LXg1okEwM58XdiWwKkX5Zl7qIMSHx13VuE1bMdswzE
4Id5OYocIpFyBwTdXmoXk+Qr+XAfb0zyV5Yb4frfh2VSvVkLjNa8nDkZR2hcOayQ
GHdIZnXM955BLdAHOMgx6iwaQl56OnwjJ8G/AWtXZ0unuevOSUKZDafh+uvMSrXg
LtEhB2mMz9sXIznLTT/cQxjmrasBxkeVY1P5oJr6XtdpudT/CMc1/WsY7/qLqU1q
8hNhwdxgeJcmXIWxexq2sWXfTueuNdKo2Ulpkuv7KabqZ7lwGat86hrz9PvO/8Ox
VI6th0Uc1pXlQLVD2eOz8AnIbuRCOpCekYEUb6DVepyeITxIlqynCeg4VF+9AyyL
zInFZOQOQOdsKJx9ZS3I1fntDnt70nOvQIMQavCYoytyeoqlOT6c8M5jIKo0tFGx
pSud91198RFMGqFO5fOxGV8JndSQmtdYWefO7c6LtozfQVMVNTxV/fENtICUy4yZ
XDivXhGaTNzKAx0QXWgHqAErU8fAk0v1P94DaYsLqnxRG3zo6in3Xw2V7jELqt4h
oMOEwWgO7WxTj+H/qXdcs+xWJRn82EXUiivNo89evrcG9W9RNXqvDmb/wqogcT/W
5IBT/bf208h7eObwo34T7SXwM9Rqvl0KunJxDkyrYIm2BCVM+6ncWIlUXihNcaE3
vk65w4CRmIPNxUNgjme9dpCxThegT1dbyaOvZ1sVsq/2rVYVISjcehMbPY4B8vAm
VxbJQiMrSrjrTuEGZs1u3kbItRiQVFx6+gzMnlE0btFh1gJ3cvmdDgK1PJVWdG9s
mKOg/HOXFrv3X9a01nbSn06jPCU/8CEU3iKnnG/RrVfCzu4iuO4P87HFSzHcGpX/
xjqwNmNKPgFAvFB9FOv+w41LbXFKlqEbjsmGYsa50h/I0LwQzVWDxnrsNCoiRj1o
osYv2Y0sE8jLZp5t6n1mKl1cLZ3Jl6U1agEy2kB+OjaESCwWO7OME+ZKMC9PEJpr
v80OwRsMh9swceFYmFQog2Zjw2OJkUSjyKkEsAji+otBIIYAVAgeVAPcc4a+sN89
m5DhjBrfDRSQD2XLNIZO3edEC0C0qLchobEV/mY7criZIeQSSX6GNwfZ+9W7rAX5
+/oc0QRulZS3H4IzQauKmPfMIgvvoHDo2SSrraVoIge2hsfY04DSJ3Pw2G3Vev1C
NK+SFKEfzyDRdZPQJ2zM/vRyYdzst2gPbPJNDiG4+m5koCbW8Wj2n44DfF0CrH2B
AUuovCf+Dj9wJ0BpnctHkSanGAFLu33ThQIvAh562U/PRzfuk9Y8XIUqhJWow9Yj
UleYJeVgFyr/VrhXfWSXQGD0thuncN7FzCA6E69gIlSw78z6x3JqnVzICWzaFfCc
55TUjQCFKMN3Q0DPz9gUOVcCtcbyf+LZi2CMxVIfayI0YIxgvYpLyIObaFBc6c1l
uvlVqx9hTz+PqKMmphJwLxShxYt2CekhHFjYUcR1iKKSwFXSyPJ/H3ln0ALeKZAO
IC8V5glUiimfO86W4qjeZHpsyIUEAReE+PsaKG7RpWsdiIGkMkDhUnHePLg22VTt
pzQzqzgqMzMpr0ZEyCmmPt2eClKtboGVHRTLfJJion8yoG4tRWGjVZj8jw+LQTOP
8TdV/IKwX9ff1EZnZ+gIRmpqEbZ5yxesO+v7sQfx7no51GrN5Ti3+6wNIMetuJHG
02DIjNXLzRF4QgZV4Z5V6ojzNESy+b6Q+KaSt/VxRwo26UhRFB6dStkwONrEkfNE
DxKx1l9qAlCTETFXYzDO+jgns8BOZi1Wd7THLnhhoZaCPF0qrc0/CsSbmyzFh0Y9
+hg3fmI9FyCK4DwWnxrXqgQNQvKK7m73u6wXGZ6ZpkGwGQxf30iyD3is52HX86f2
512B7s98FcO9pUFUEPUkzaBfHxhSpgmak7UMEmyHyY8GlgaBgXmn3EaMZigx5bXN
JR6hlwmjdwXsCvmm1zS/kaMVsEYtEkpRZfgSVZ2RXklE9xwaOhh43/fXw9ygD3BC
rfwR5coFOa3nVQblXMEKXyqP1hV/fAuTgaKat+xxzjwwCyVEwnaLQ1lXuUfQKg74
paBC5SPOxHqPjEQebDcupWBnJkB9jFxGaIRp0ShmwFtr0S+XlE/SOMOePxRYAvoD
217EzUriCMaQmI+fvefRCHLUFsvyHuq8MBeNtuvmuHxFs2rWxg2XftR3HvhmvfUk
nmwizo7BbHgXXHHiKyHeV0ivtUTL0EWCKJIFjBn3x6xYDbbePJd+oemLoSNNI0LV
TOioFhAz7zBVIi3XC8fdpUoK7SYo9LxlI4neM8JE82QLsHAnt93E5moUFnYZ+MJn
z2H+MpHPZOVQEFEnQhTN46rcSUA+nVMwV4BHmnx5+Of4AnpFUri93zjoxYcps4de
RGHKFy83I2bymwooKyRB+abiJSkFnzOII33oWaan2Yq2RnkV66bAhGfc5KAD9ty+
pg25nCpbYOhAXeVp5Q7nsZnrcXW9CzPVFH6DXOzPG4Zmac+x8nbGJ2mvWnSzRDlj
0Tbfl1WgYTQ0VT3ervpsf9emJty3xTHzJe5HhdQkoPr8mU8A8//BnmF62z7FBUm2
KFpvSRbr6Utfogwdjq2/V8c8rKy6jQHTZ55RXR8GRL/j9gxzhbOkKWnldHX52fgE
ifm4Cqvs23Pe8t0mxh8OEEZPTulcMyliU+95kAJioYX2rEBlSFMoRvZGIclIL0xn
eom32Kohdw49RgYyv0MAMcsKXgMDeBeW3TY/7UfwfW6n1yjwDBoMYJkbDF4YrSTB
6VJ0A8uTZ26tIAhFs4oZvIAvXh+W3Ubi+FrUEWVKLHFabLw6+6/Y7hxXgTTGriSc
UuVxrEyZqHKSsFblSWDYAp3f2eWzjFfUlaV5MRZqhhCCCLuT2Z8m5A8W21pL2LND
F4rRAWHHu9rcoWA+lNkmra99D25755yPVtGYaPlnJa6g+Mf7qfI5uHko9dOJFrOu
6cVx/0UypRfdfgL3efUXrgMYFK0Yq3FEK8JaJMCvmgWWoJ3QiUFsraahXrX/h/WT
VIG/4AjDs8kyi/W9gWI/3QGx1+sFDgnTexTBxARoc19pIplAfISRbtQXUtZPDzaM
q+m7NJ1TiB7VuDqlXIw97KFQKOzXVy/oTVyyCqz9NLQhEer+fJorLYE8j8iQ6wW4
Nf2YXONknsSl6WnKTwTEiQlF0Ranu6bZkTEvPE9qHLGM/TlApb3+7SJ4MTy5Aiow
wjkOYYXzPg9y6777/02/OWzRJV+pScDJufuz5gAykgvp2GYITfbpRX6DRGCHTbyt
RLapkmKxv5bIrwJXCBmmwrobh+jmMkPU3bVXgsoZ8gYCMvx6kL4mYyhxS+2E+MQT
O8W+G5ObemV7VGQoK+FzzeSZZYSEj5WjF4lNfAff/6Bxvdq+oES1biMDPcab/UKG
g5qqUGdt9SvWlpp1q1PGtZCIRvN1bT+MuSAqMPz4D/JM4u3A2i7qvBLrMU2c1lYM
apTce9xcnFPrQ5j1k2qiobouAmo60+bdqHx99+UdOvhfGEk0PMuTgWbnVADcqZbd
y/z45uYe4bfhBIWp+TIDdQ0Va4o7/KNPhP8jmjuiVKNBjEESLzqVm+2n7k8cw0Zf
V4SdSpusUfldMwyTxt+HYNoIK8OAp2CnvScupWeZPuhZRASjSpHjtS42FqsbW0Wo
XI/J9tcAyIio9/nIlKA6cjG0lFEUF33HUS0t/vwtjuhHX1EaGFhLYiigGjTMIYQE
Q1J/dyAlEkm7BI3LdIUN6Ff1JBGlE6fONYDXS9YLwJNr1IqxQ+sIPnssNS1TPtpi
rbpl1HACnC7V2g0yraOo8Tdt8OSUNywcWvwaWiS48Ybh5Elj0ZiqsQaJKIo3HpA7
v1qF/NzkqY2U39CBzgt9zmBqHfRTPAP4kYcC7mlGZisdSdvigH3JzedeAwvyLYYQ
eFLuFzj0HHIRSXZCXHgcU2UJXNPANAbfAceQN1S5FgNJg8w6uondnrnpuDCdzoMH
3Y4+S/X0QAhPdiGruvpSxkdP46PQFbZBgIktS/Xf2kYl6lwUELIkZbSmIBV/v/3c
9SozL7R/Juuq/dfBNQtGQtIMFGQuIUmxsKArk6j592D+JYqJnn50AQDTwONr5d4W
KdCDBYAIMzCXBOe9GaIUtUENiQuUp4timT/Mb1WtCPRw8tYG5Wd1Wajs0Q0UhlSS
hRiUB6xb8LmmvbskteW9YQAWY5W6FVvFdHnEcbZPIWBafp7ZgtS3yiYT3fyNez5t
7474XS8Wf0fhThbU79NH4Y2tIFOt6JsbIjbW1iQdbUv8wPyx6keXPyqchNillDku
hhDQSVHoius2BE+ntlsJGNLTzRuNnatIMzTKfslYSzYH/AYWmHKv20bSIZXWmDDX
nkADh3ijjqTNn1xQyXc8Ve/gXM2FObCtyZfMjpWZvlgHx6h3LV0hpTrdq588qGro
jYpQauAnUgQq43AtGYHDEFS5+cjBLrwMLG3/pTnDh1+1OH+hdhy/3vKcysp38NlV
+LpmVBsIK4qutOXLC7U+VEEir7Qa59ngsbwDzKKKDCtUcCXAPpyS1n8Fvx2yiLfy
r/V/L+s2Lt8qKE8THRkIbQW6hC8pK7EzvKcd6UVtCX2WedrjClfhR8B785u+OxxJ
krRHCEjlpDTFfMgYOQwlS1HYmHJVuTZY7rFQCdNzI3a9KceABpS79O6T73AOO6go
INc6IHiDmCRr5xSl0MmD+RbBM69xYPhweZMIUJy6k3y4+TXYSyOEOvsND87yHKVQ
VByCuEMiKwS8ZArzcBRn4je4f73utaNddvzNAWfytEO0GesxuR3IwYJTm9LVXTio
WhGvtJo3a5wj+WHM6kx6Jkay+u0XgvTe0OeFmTib/ow7WZ2PNDBR23JvirwQp2mV
QW8MXoFrBuwMeuzAy6th90qmUpCZWgrrfU9kqUnae7vweFJKD6bT39hWuTZ1XROM
q4YK5QwjxGqrN89D0CEt2obS0wxfJEThM1tPK5221OnDf6cGyJ/fTahP9fqfVE+u
IooGRn+i0HBTzfmbBzlV5DGJDPwVwpuRXbXQulyWcNDHQow/F+u2yHpKI1KI+Jq2
LDJ8GSBFpYyIeFpJOYtCG0AvPcqTg/XyKEtR6Psa+QV1bjyS5MBBJBX1sKbaWifH
Jzao1ivTLTV/IAm+cjC/Xo3u8OzViKVJW9ZzwYSqG9Imfj59Dfd2lDcU1fcanZ9u
KVTu4Pqt34+MhXjhbMQtnuLNx72Q//L4UQZ4ZT+W93kvRA9Xz6zNmogsfjAT/w9W
B/3ADf1PwAXxbgEzQHDLuolakOVMZ0SV+VSLs0V4jjXtukaC/UUWzqAu1ApFq/nW
+UPA3a1dSxLOg8KvBI357YmXgynNRj5NvEvrkRPu1jC5+t/zKB4BaMPAVpBLGB3g
pJtvSIATOQDT21ir4BYI7OMNp+PXsX5mzLJfaB5ozUrg/wTqGaLGqCzGTbwQNXtq
DOyHUsW0/F8oUrMXokKhMflCVVRMkzd5/XR5fn8MJMNxrZhMhQJDcLiKdCE8kpK4
TfD/XsSUT0VBOWBvPYY5lrgr/dxV4hCTm8Ocpjp4FTJht23/HcFqOCv6+6XpgE23
cKTOwoDLxl2L/gWBpyXoCQnFCx5gyQGvKvQW2zsmNF4i/dCtHf9VYHc8Qb+SZKho
3qhtIR/Sg5eqfKkYaP+n5DYjxe1SIhqnBzQEnTRGqUnKTxEdaOm3L92V25tZH6Qw
11KeDbLnCQAA8088W3p9siPYisuYdSQvLWyy1uVGVyf4xZ73PPf8/vebWLIBjcvb
MtRxSVAAWVwt9rDPZOvrjbQfQpi4eAOOvBK1tuZgC5mKG8v3tR4XK8xmyYvcasYD
fJKAST6KrusgWuMg2Ed64egCfMaZbQwImzqAezwcFW3tXG+lwuuYjEtxpVXpLAd4
ThTTZXzIpxbQQA+8mdTOxpiU0+xC4ik0fO9kCbItFfncMb5YUN1BAxA1KxNCY/jl
ao9+hibRynD4biDYey17GOtJ/j7sHeIV56EIgE0zkG5Rl0CeuZDIDHwN9RLT7yHy
RdKjQm33VBIcneojG4DGCDGzkyYa51CyXgPKYCnFYzzfkUvZ1s41MNKQ3IdNDJ2L
1ZouUUSA5A8SWV3gEtDUiQUEGL0nom/cUxVulpUO11wd2sgl8nU7CNHjPGrWjuGk
ozh5sSVxhS00oYA3YfwlpwwqjavSYSzuoT3lX1C+2WrObFp1hwUZDRA+n7UX377U
Ms3pnG2951a3n7T8r+m+FTR7WYudddmUXVEhxsU1fcpyCWFuc4X8vr7nD5iVSUYy
M7gPtx6HLJ+VKA87BwD/guGAxKN/ftNo2nVjODW+5XHoR/xGewyGIKYkhdQ7zOja
TWwMZYRZqS5wx/H4ddjYY3sDTALcvfPzNy6eZYvNSP4AgKrmP4Urk+ZV2fdM5svm
1A9+1EeXUk6R6XmL2z/kUG0EmZ6GyHD2X8L5xghr9ZiaUFZwK/s8O+ZRw/s2c5WG
KaUdkxSL1JUCCjAtYxpy7xP0eYJWpAZA/JaqU3DhseYR5g/THU9b79r7z+qXmopH
TB0uYKHw4wT5ddk0T2TsPfKvK1tf+DP6SMjSGkjvjsRo/i8tYpEPtaPZ1RyKhJ+Z
riJnMPSNX7AM3FnmlnvIdilhOLEtvFBoku8Np3+QxRSktbLelLZvGfxMeW6lrywZ
0WgWg2wBG/uM5vKmb6jPv5xGs4+bF6UUOV++mssXqBuzQidVcrQYSFlHfkBvoeVF
M40nfLjCr0PhyaW7JTa4SN/QuVbDmhHH7jMbZm2Z6kKhzsXTZmgTCNb3N7373XIL
3wkgcSRuE44UVrUUgTDRfwYxwyyKQOx76WBniaYjKwhEvkogK7UbLCJn9W5z1qsb
aG43C6ObVcD1dJEhxu62Qm9cN6JwTZ0sF+g7WfD/vc4rcbLzjrjdFxo+SZy1kETU
FvLgrIBOYrw4fqAwVcmOgCU7gRSyWnrHS+QovwjEbCY6v6F9IPX5VHPt7hdA5aC2
DKuq++cj55zxkejzP3cxFcbjsQeTRzmGB60rwnb3nG9G9tNHrNGg6W7+J9XnDLoy
8ofL7hiwt9c5Hy72kBdakyC8pWB1jHXQ6vxze0B+GkDkpjz1f1FFGbdQTVW5xlDu
8lLEzKKdJMlJiAIhet011Xq/nCgSegAs7v89iTeF7pmZsCO7ChCp6cUSJEF2kGRU
gN6eZCFOheKpZnEOuL2QyzKbLJLfuVlLt+JVeHsH/SI6RQgJfqb0BMEs1HwFrdA4
x26ZhK2VynkwvDb2Q580n3LKRmBpIxijkNhLlI1thR7PHGSJgkXUtZboJA44agx6
AD8xR7bvKNhek5n36l3pHUbS9mCVRdGhHYTMC7SZ2wjtWzwcN4bzMfxZrqygj5MB
kAVL8GKjKhlubRQ+m5TDPbzFi1WS4cy8JdLQ1ctQr1MA1SwyXl2J2Dvhy1Ekg4zn
Jkb3LawN14MGmaIbLfuTF0a+3XciBMGliqdjatufdFDzMcyFHz8Yc7pjnZUAHbh3
XNayoDdroR307wl2OQ1/bTIxWig0VFVuUU504ElUFklJRTbCLyKk6ckYYug3fzZH
YxbezGu6NS5E97jZEfiFv1DP+ClUGKTup1b3HmTUDamfiwy3GAEp4PPH0atslkJg
+XnVj1tI3CQOx1UBq332WoD6ANLUMcazp1u5rZxTXGTe+GNMGgkgb3wJkyKdJ9HT
XQjZT4jSf0qU6DxGOfg0VcJ2g6QgsLOEWZgKsyvyEpPVhxZfn8RjPkEbViPXiTRV
HtlNAj9wVSdN3WKOhVpcwT94cKXKlbAzCMFL949Nbmcc2H2OVJejP1bMGF5qBS1E
E/NgyGFBrUooo6LFnRgdhkAbGIJYny5iZ1leHFTLHEg4U6fjlw39/DlgJnGifTvD
DsJDDi6+Gn5uN0oISjQk56sBaYap978Bai/MNke+xXDfck/LFczj8boM8X1RVmPm
OTStZ3VLfN3GplsWUxwe7P0tiN6L5V7iNbsYyE6tRNwyQBANNDXNjaKPwCLIPVyh
gLaxu/O+qXssPaAZ17MZQoZn5fdmo8211wblJ2wmzfaGT0+LcozNZ0OQ66De02rC
FSxy5CB1k5DzImh5xTP1NVy8x+kX3wqsfILFpuzHYm+WKAJESIEC3aJe5NS696yn
+hJ1erLEJppOplGqCM+N3eSLjXC7obTRSSuT74Hsqk48mqS1/IDlu9eSv8TUyRF+
J7iqYEnSZdnecdsC8heksVQ+COh1A6GFODyjB4EMm/7oQh6chghMDyQvYPCTSnIZ
H4TaxRDd5YVHjTAGrLoIUQ0No6ELW05HZMNk3xKSVesnumrkju8kqjYP8Cgth7rW
v6tHBQYDfuDWjMeoCepZMZhnQqEPH/rcxL5xlByItxxduaHyKPJKw6qJpKCP65+U
sVRVD5CAgL7pOiEQjNmBHyUA4iWk4TUwwCywDMD5qALREtngIBJnvmB8oz46Xb6T
Ms7BKWvlqcFPthS7ZEYMK5h09/SNlqola6cn77p12mrYektN19vqYA+5UVakaJzD
wALb6YcsNVtWgTggCYoshP2tFtlgjWtx8Med6cI5FKIVwhI1AvI0Z6XMS24j9z3L
0KngXme2cKUDVYWrYQaFu++NWkRGm6ut2ye/n7Gu4BjFiLilgXyM9bUzTTjgQNxJ
GR7Yx1JwgHxV+PQPRQ2taDEEI5k48fwmzWLl6sB4XNqEP0I1vpmmSkSZOc5ciaEZ
OBIXh/fK3haN6FNKCjJ6N5QJz/HAUNGBMK4LFLQCtujYhsUoko0X4iLEuPwnNp5R
GNttcBFehRp7PYfS3cN/aetO4tpBfhU5+JccAV+XO/GFEV4TD2u+pl/jzPAof+67
HUAhf0OmWcxT3z9gPpUr19NFYLyQCh9C0N8f13mCo+b48DLQJATlmLf8G1qs2Kit
NC89A7eyYicAmfpJWWQlNgOGx8ZlrsdK7Y+EY3YqOKA8cB4fLsGdHlzQqhoPFJg3
raUQ62N3KM9m3EM14dalhG45m7BwCH6uYo+uH0xHdfN/JSd17Fwo39i099V9RheE
RVWByOJfPWNHxXfzvr5dHC5Dp90T9OFV4rJQ4/K6552l2CoPqV88xafIeQjJh0h8
QelEhNFI/3EmVxkFsrNpH7PJ/gTkMvn1rnFTPzmABCTVIISEvwJJ/f3ASAauDu3k
xxIvGi9/iddBYa6CQD4RqiKDAYc+uA3WLzKsdpt4FRN0Z4h13dGes7qqjWxtNm3k
okXpfvO1HEbDBjuPl24WIJdoEZhjXUuhED/Aiyg3Uc0t2qygVJ3iTzA9QHW2846r
FxKM7fGAeik93sbz78ig+KVKSh203jkteIsG5uemCZVLKUoryxk1QAarzGnxBYxk
aJLEJTmgFy/2tyerZdeyuANKZ2UdF899goJfJmKUY0ohLvTMJAlMYTItUj4cNlrs
lhzNZCnQ7CPaiteC9BWYBADPCAaKxvzgX2/u054VoBqtT7oP7vWCkEUXSRo29i8w
fOg7XLuRg788PZ24BSjBzXEysZSUL2x55+qpicrkJmhNy2cJBjx5EEWAvOBoP9lT
nVF5hoKP8JkX8d7CGrOH1oXTyW+5KNDgCD231dnZlfMPryqfcbSM+FDcSXZdPLIm
XUa2SUVXnRt48i7h5zKMB9tSOsDcKyZT4NGUQma/7TQQxSMFOdqlYUimOJ6fzviY
VImsI6gjeVPc7ScqtNDJGN/YUo4RiQHKiNoo2FrDxMf2rRffduBl1slIb5k+qoC/
i7agFs1xBTVEWta3+ZX4UszIzshNGdEn6yzii6BgoJev9oFCramumUCkhuHFzpmH
9QzXUZeXes9oFig7Y1bKwTc2a9UXOxh/XXe+n3tMlyx0nqY74VOgth/YJIgOzM2o
EerWTvoxY9pqElPYQrIGkDF/Ic4Aj0T7nYS73P2di8YXBOwj2KCz2QA+PqBwqXKd
BAUXu3e9jRFPCBVuVEu5sJNyARSfD8NVM5zN1XkoAUeNNbW1tFLkODdMmH0a5mt2
dvrl/9O7FlpF7n+us3hkoXQnczqVoagwI6wAczt2Vb37tjVz99NVXaQaoc13l2l9
oygV+RAlBccrrE5b+LpHm3NtER7x1CdiCRspcOpI8TlvF9AAKkGyW42hcs5TCghx
gtz/4Zr2qJkkhXrZZAUjH1slXBDeH14DlpoFFOpw7BIUjzTkQ/mdAWWGsWf8VGgm
1V4B5HFURXz5x61yz78AeF/DK3XAiSxkuCu948eqn9hWqE+Mnvh8ry+a3u/+4qAb
ebB5tJrel1ZSbJj8rqLfRLH87todOM4/pAy0wNnXse2vxoqAORJB+LXKNOjQcZAD
qbOc24Vww8VmpFSJslyL4kAl6gWB9rhg8lW3mQhMCtrrtCT6elXR7Gkfu1zj332C
I5s8sXeXTNZhhxLN3m5tg365eXStz84Hr7/XWPZkuMWchy0TblQ8/6vdTGAJyArx
GXG/stBkgFNt4TbNj34ZD+L2reKuz8ZWNXTNTtJ4mL8tcaYFqtwHzRTJcmKR4MnY
TPqFtpEckzLi5zOF+sO0LMtTUA/S7QbrWtT66SXWceLizZU98c9AysNTi/FAd3mx
4eD98PlbfmJjYxg3NZB1p26o4RM9U+RDgsUYb/e1g571WQeDdspOVR51xn0wV0yD
sLa9yyiuC43wJuX2Uv/o9owTi8I1qkKzx8Ba9wws0YcMOeejr4tnT+9Q1LfvhJPf
9zKfcG6cAYQ7IthFkHRjJjGL9w42TPDglFQ3ToSuo6TxqPW15EaaK92PJk5+Mvdi
6/sg7QvjSliUdQ2EbKgLeJusltNQyoqBw5jyuRLHDDD+2VVpuIsnf7z2FBD9IHUE
i7g2baKfyCiONxV0hcsdiwNB+e2cJEBTZgq1BbHTnrPTljc//2ffTI7/rdKwL1jB
vvqLtRDgHGK36o10qHifXajK6bnHsVG4y/Fy3ZusNRmMAtPLxN5TlliaVykt7SM1
YD6A/vc2aTtAlViLeWXs+IQ3HyCe70BXQ1Yt6fpeObdoxC6uM06BlANLKftU0WpF
oidaq4S2zqD/wP4TCOCxLYwI+h0Da+32Sz+js7+aMPpXXzAUSmfd6JzZSneoXxwR
wdML8C3wqaqY6ZJaQGsMg8+90PKxvmFM+xgoITghx4lf7xrZ4Hr8nJQS8S29i3+i
M+jievrtj3zz9XWkK3EhEDg7SybNsyaa9zD8QspcBZy1Vr4ILC8vJQ4pswgOCSWw
/ufFcuXg2o7nmWWGwBUxmnyVXyMZmP0R7+fMynocDnlsGf3kavzTKhI8K10UOUqv
hM5k8v7kQZEZx9D1BOSzNhAv9L+gefoKi5qxQE7hwWsJa1kAQ94ZqtZAMNj7p5oa
x+OEAUfsVtd6FpUf1jYbTfKC9/TCFd5p65BW9NscZLkc2smuImWV1LbzTO2p4yry
ldTD9N3ED3UX9EuAJfmXRBvNppWSmjc7OBZTKhgZeECPh3D/RnOL5EPTIp+pYAnF
dY4zZD+0DwnX+gB0cUTBM+TiwFT9e0Sr2xhkKpqR4758GGm2lrmJEkB6zXSCkXe5
HUJUhrF+pkzMdt1NolbKQW4wdSirWYpcuPhjeAlb1R4zNaj7kxJaeHbxWVvMFhRc
Ey963VgEsh53x6VUxF2SgvgpsxAlGahwaPUkyobQekK9OUyYXCE1d7oDh5attQ2p
vSy94j9z0VmBXDBusgiMrnbrMT3R2crdxo/l1OXqyB8BiEReOwsh2wgbn1if1Lba
WreLmcdG5jAyEqYMUOuKU7lBRD1u7s+grChOnlqKTsNHRQGG2/bPUCA7zAAD6lGn
E68SvVWJqgiIvFsBAUMe6ExYrpGJVkvO2nYxW9jUUy9QuSju5RSEBA/GM5DuqoGj
x6gZ/GQ8FInKB1hWJCpGMFhhCvalTkoj7O1wPKgaoGB21aNSD9NN5VIut7piimQT
5hWoAHvbQzuLaBUMUzrZ4+wnD2GH1ClJjNGn4dAcAIEAiwzaZTv5zDxnKzzDxbj/
sR7V32+ceqdy6MGMGb4ME6cKP+GTlNdCjS7bbU4IP1WHtbbyDUz8RxvnfZneKKyQ
6ksWNIIsblyN6q5+LRt5Nu1ZiDMEW7BTPfjBIDqtRsljFHfBFTz4qN2IpKgozNrv
Q7jOFOjjdgyTyM4pXVNzQyBmA8P/aBf/ViRlBuJd+9Vbv2vPFoaryZv9DcUNMrD5
dKFmHFid3wxeu5kzmMPRz8YMCJvUiM3rFYhrmIhSwpAuJMofm7W2Xppfad+DMVdu
kh7rO1TQ5FRTIiQ7XN5M4VBmmuwc4eUSExgRxQdplNIqJ2sSubUM4eax0L8+gKMT
CIQ4higB3QMoyiL4HIIZ0N8sXAooM2IJI+DGQnte/74Qtc40mJZHhJ1fc5UI6yKR
u7cS+l53GNRz7J1PeIFLYRJ+YngCF+Cb1L2PEEtfD6ztpzdSwFYGe3PyK9IQv0Hn
yt/ONzwhc2o65lJgrmzRJwYDw3l+YW1f/xywA6FJfsZ1S2UmdTrfGrSxTOv8ZMFD
zHamRRL5L1YJMAxTw40YIVJ9TLrZlJNj4TfeupjVNiVKd3mbzlmvqpB/uo336xLm
t52tAoAc4r0HXLKKDRV9EvBrOdAVJfQs+9oLbcNwBrBfA3fwATjLbPhnlADnGyYS
ER6Wvo3mVjoGLLgIyzXYc94vXrUmDoAs4xK8wy7v2UYnJXO8HWEXLfUFfU+tMQ2H
So9YkvZ82JLOpa1nqrK93Otg0eFkStu92R+Dn0b6hrgp53PJZIcR2gCK0onx/gIH
qXYR0JbP7IpuYZikWRlEtyX6hS6oZet1oc9XmO/vNBKtoMP+9d8WtD/7C4a3FucT
kXGTdfleCMR2ESnAPN+1wOczcQfTLHWVGJoPi5NgWw2OK45jkxt8hpi3o5Ox/L+U
GAQ5xpF6Y6or2obssppdKeAuTweahB3ji+8fyEkk83Cnck2sX5ldVMebSTyfYfXH
HaxWUPdraCNB5OMBUGBaWmdWvWaqG75uG1OhzLKpMySB223eIJt/2/6+g6h6PXS4
WWKyzxSGxuakVovyM5kHHjDRlir3k4vo7Ukes0mjLpzSQi6Wv8T7N98lltftrBOr
w6j5J4h9haUO01IICDFTh5SJFrkw/BuqGPQNC4U3em4WJ8W/JnfQxzRO+3DZhfch
107WlNoqbv/Y//I1ZDn1SriGKfbfr1+abJFmC1baAV8+pz3LURXycwX3PM3Yb9Al
wISeO8fXu3EuJwihW2hVy6xOfRwPNnwYJpWqaFgCks5OV9YcyC4Xm3HsqHOE5JCD
cqJbpge9O+Tt3uUevBF5lqHcdmjqeCWUajB/rp/F1Ubmudgri0Gyi8wFerPwXYoH
+940OpJ1eKGkEs63sw0b3qZTA7YJNXX7WunCx8oTAlLO/wCOLcY75bELSDxh6AdC
UUHTodiQV1uWJfy13/o6wQroincfGyA0EGTMmhaucShLQhhcM7Iz5Fpr8P4EmDyY
9OcUZkpYo37AKzj44fbMSRAg+TUJNaOZK4DVfXGs7YTkEwLHTvz4O0jnXDzQUz3J
6n8GP9PyI+dkfqfatJWg+jmvz4pVep3DIOdS2X0ZPLV5D6vGJUZmPgg68GwwjRFJ
YPYWPXbUlEvBqVQYVNSQbWCZOegVfDscnwV72vqgEa8oePsr3eZ/rahqDnmLngEI
88LVqBKME/5pFFeZku2BJ/GDehogj0DguEtq3V4571QcyBI0ordlVLZ9V5JdFmnn
85y5aN8fG1kt1BxktD5m9Hy6tZt/BORY4C6ooWv9n5lPNkhysnaD9c24b4LFktBi
lE95Zj6dTr/MvBvNpfb+XjIwZIKRrw7jSmB5pexDAmQ12B1TWmXSYDKmGmu53rAH
nj9VlmIO4mbx2Y1m194riKzg4aKD1XqMLm50DeWxGo5ejJVrAw8KNRGzSv6n2LP6
0OC8fZ+r5LDKkQex0/ymhmoS5s/ek8mSUHxHO2J57jx4kHj841DZDaY94Tb7YAzv
+JlHl/Ga8ymnRcOPrBQbPBhV/ioRq8EVUf5ZKngqu4GvUGk04IOoeGa5uMOSj9Bp
fyUmHAFmidrHFQP3bnTzMNhR4FnfSxwwjkETGLIWD5gNZAGT0vP7zTQdWhdoIg+p
pPnAByPGQMBfozMdoZwSnfd4Zc311Yr1X/ChesMIsmzM4G5aAcCHhbMLVDSuh+5Y
35TZuYqVaTIkFVk3g6rgHhR29MTBSqnOAbeqWIo+wTV4ZPtw7W8hJAQujy3LbzwE
Z1cHGmxU9LMVNlnEvBOIs1Y2kMoAfFDLIt9j44l+zp1UswYXkIfs16Z6u5HMO2bY
JKyy072Tb4mvwP128ZFJBrPyS/yCNTfGtOD8OlTZa51/98bPmHToIkqM1bGmqO5U
xkrCqef9gA9K1FKXfmyKZsPc99kBonbK+CgGMB9dYqKJLO8ok0jMRQOEo01n5rwZ
653kPGbea3QLoME38OxvaRz6N6UxmXXwNU+3VP5R1FZ2AJWmlNswoEVyJg8FDN99
FIonizunxjmXzlMU3pLkyqUDS1pO3vcY3V6SZLfKentk8ORggLOw7b7ukQKw44Fz
yc7eeqH6oDBZFS3J6Vmqu9zhIgdQWUxbzB42NDCFKOavTzrtEbAnyqY4XOwSMDC9
r1Xzc8+TPkK7FBTuB8n6i8Rzbes6RW89ZzMMcdp1FXKpJArudVCNxuAvaLiQPRam
DR7kYyZ8COjnsiyvs4ATErzFjQFdU95OjABpFaOc8QHV3SNlfs5iLV+Fvvc6kLo+
ZeL8COCz+HpERub4l41rZtW0Ee40mSHODpDqzOqxRMBqqsVzUOGG8rpVYSG1HbSr
yJvKbThwTaQEqDSFCntajQrI4k6npq7SoqCo+GQmdp9RnQrNMioYshuOxkyOGjoF
j6U0lkgdoiAq4g9x2VqLyJURyzlHzWEfJn5GjQVHCcpuxNEXPZJv5ysRJhiJpqFl
KkVN8NTzh4t/lpg5vQDPdv2k+Wi2qh8cmOb4eAOK175rh1U/ci2IOs/PdrZbFnh9
Zm3ek5iYJDYoQgqSWb6WBOyK7COIAabZAiHrM/A0gBH5c/cQeWvXomonvSEkYmcu
Fr0X2AdCfsXJqCj3CzvoNjGfPK37lD8FpRGXYOmx4at6MLhlymgjWFW0Cp15xEre
fKqnsJYr/RKpJNUZRmtnvef22GU6Lw16b+wbe8Wx7UeB3ozKxUQJjfdcVkUzY66Z
YXA1INSN3CJoaJXd1K6SAogfWqM1yMURXVxMHXqwgH6MSdN/IAl0yoCnwK7zBWcX
cein49D2PLrZ1pZwd+5hra+phpOR4Aj0yKT/JH3s+JWSdjAkbpoXtNNMgtl8h3Sq
Z5BmMBJL+RcRjSOis1R/yItUkTcRmLaNXS9WPNTE+r++CHZQoEuOaUywD+/bCjZV
lL3mZaELZo3ESv0bNuEFMH0v3UvetE6ND2JaiaxWrH7BXB0ipHods09KVn5aJJBm
5b1r2HhzNR2WmxCNVw8uWJeWFGzi3G1J/riWjUcWXMyEcYuaOa1kHazdQzIP8acB
Gj68/3MIYAuYfTfGFK9gUYPz1X7ZpEqTLzJBeR0ymTmxf7Pk7SFG+VA2it81zvbT
g4MePQUUTRAWvZ+H3NVTdYxLouNcm5OMwXGV/9oAYsucWDgCTLazcryIcflrhdQ7
Z6VkeVd20snywjzSBv6MEeopPOvmi/oH6g3r/rSBBqlybzbr0W70WiMvAB43zPPl
ehPOy09L8KF4sofqbvCfMZ/zu92vuquRPDj+wP7fenbipRH+RwsQgBx6U+C8BW40
dNzzlMDZYHgzxXiaNW1QPcynw7g1bvO+oXIz61LdCAgLlkSnWDPoFtgpdLKBkAeu
ep0jRs93Y5IADjvlQ+xyHeDCq4oCvMxiif8rO77DoDcAdfwWkCuE4a9iejvWZSX7
ceoJYbnv9txNAlS8YC0HprGirXYH4ReVsfh468UlysiZs9xyfeKPBnx20zI7J+LE
T+SVYIKPOz2YJGhkR3ZsS/J3yCvsZayh5KqHAIVXcm1Pzl5gtVqMWGV820wrA8Zv
5DTk7EuE5RZel/s5F9o3b1OUyvxsio2S4Pg9eWEr9L+A0rch2hfnboBCN5iKwGFG
40d45WT6MQpQA+h/sv1xAE7ENP9t+YWq894j0bXOrz9GNSwno6+zYEf1Y0OlPn/R
U4GLXFJqfPE70XKCv9hWIq0pPyaUuDWIaZ49SIbLQoAH05GVZsfai83+Xvul5ecT
mT+z6qSCF+4deUDuziJGq9bPyyLtWqOoRZw4aJYk5PILqm5GrV5dj7In615B6vM8
3QGXGYiWNwSTXbAJ2Qluo5OvMatOSDKk/q1AFfl3di663+JpdWSr/FcgXKeIXVKF
1oAh/pUn8XyNRvk9QDSFUcgRHVIuvrqL//XbTCFBx5aeoQbjNntD9EBBI2bWCC29
pytqZbDUHgZ1sHzBJ8MhZfpDV2umcnHwesgB2XsmKclj9e91VWqbO8q43PBUmY1g
iWJzUHParzs6oJwsrFHC0uuj8erzgg/RLZakE0cQyniu5iIANYuFF5EWHQ9qSBZh
yymQ0KH7bqedpYed7d2W7qZH9qqxxhsldMrlzERg1spkvWGRo3NLnIpPI84xh3xf
ggIi8g7w3U7v/W9JGEZKihVWaI2EHNcT+dcLQF8IM+UgQ8rFtZJyKwHv+cakIAdi
RYD2p60bRWbUUKGTLr2wUe/lzASy/jh4go1NG3XvHdyxwaiItdBjJP+nHoJuAO17
OJQrZykuZ2nlDizCUPj6BdmAxK0l9g4FXEu90C9NiqaB4lFWQ3ADLbkSLyNoOCdX
8M/3WplmcZiImuqevPkyP9JOXzrxg3WFlfgmw+Q10vBv+8uNIZM4yECnvk+UDZMg
ptUeGvpXG6yFjkZ6b4JdNloyfJzSAOx1d6Kn0XqCZXPIm3HvEMferYIQ36OMsD8r
wnyJM6qGeuY6/Qt0fcY6QROuKaP+76vu/JdCYt7MTFfqPHDqZix2iwWgXeHU1Nj+
ie4B/UhYzFl4bLuFPeEDaY6aJ2xlHJq4cp17At6A274vHoC7PuHHgkguuDhlBqKa
O0PKFj1ILUUuamsed8AGbpttYggaBP3i2mPZu5AH3KHq+i86O4l8n1geIPB3UYAR
immqwPpMazs1mM6oFHtPykHIlms46pzB53+e7jkz6XgYBg0mBq/KE6u5cINep7Of
J53BB1O8N8nzvTNAJdWu5hEy47pMUynnWGvMMOYcDDU7KVTf1pyIC/ZJcNWb9FuG
PNVfe8AzHZ51veT7XyuagN9hJZUiYtKmdo0VI3eaT/oGvnuB8YAWyT5egIRA3bH3
eXUPpyzmSkJaVCQzF6ggtH1la4SzDYNg8jAuh+OQriOBU5b02IehDc04FKARQ5mF
mqL3MmXbeXo2R84+x4lgIDzTI6wz+EoX7J3vOd7iSeCkicQbFYtKx56OtqXfN42r
CERGhpnH6hGCytmKZxmGm60reB5cYjzREg7no6zbI3WkggqZIm2IZizpGZx3SC8C
nKCx83/29IW89tibzvzYZ4lSkTXYekr6ET01/Dve5V5xMNxZ2a/6JjbPEQM9E3ck
fLnGc2wKHbLczd2pYWnWEYwCekUmgCFom6WisKIlHZKFkU362k+4KMNctnSWTWj3
85EGTb+e9aVNtKVlbSgHAjpvDqjpyYr2HQkR2ZjyIqRnHtLVcpmkWbQvghwKuzd9
JRXRwC9kdP516Gjbi0WGH/5/GY2UKwRQPCQc+fQeXW96++BL+W2wHVZnHXPd9NWt
XE3eIND976D3LTT8HSPjgf7HeToBdJfKYIX6hxFK1K8Ei3AfR3OAfJV2cmuSm6v8
kcv3pP1tX0nzlYIq571Lon4v+Kty2yiXnUdP/8m44qNsxd6N/Y2DEQMrgs5TR37u
TFoIlXFlrpLUDyqW9yQWW749yxyMJueifdTAUV6x7vnHJTMNpHUtxKfr9LGqZNqI
NF6V89MNbqK+jkY9oMF7UeQxFwpOZC4nkJQDFU1OyBIAfd4dZWasZHMqaC7kR98/
WXR6cU/aRQ4mbF/EXkd2q+DQLitU7EnL4je2uixtWYGQm7q7F+nM4kY/6OWty6sX
dp8TN2ZGGbnabH4eu4mPPieuZwNItJ0FUbcCaLh/c90j9b1kRlpJQ2VDW+lvCA+K
GhiVt1iZm/iJ58OJ6euQxpEhGVnlvq+SApgnokJaP62TtqFBKwQszLa4yZ730DMD
uKbM1Addr8OcpIG1B2xZmaX1cztXcxoAzD/RcEabUZFz2x7pTgYdx3cfG/Li7RiW
UP7HcTZJG97S6MX8NDF7ffsS1eD4CgpkMq3XxVRcpa2Kthvmr4XxQNQwnoBJNbPM
Pj8sUaIvh5lYBDoR8tNqLJCMmGT2nwj0K6mcl46MECkxXQEzZrQbQ4YlOETJISo/
2/etgAyTp/9yVdR9cGPQzAd3YmuqftiSkMB7b7X7DU6NbzbSEJPgbxxBTJWRwQPs
gw760tc7GHv6NcQWFheNHkwKdJer4LF10X3qcifUN4JACcbtVmbmRULgddTujSXG
2Utsz+Z/NKcuzMO0MmZXxuFjDHr2+2f5WaJt/SKTuqUIzWxm7olFGUPDqMqEHFor
ZsC0hBzeXrB72aiRDyX4QZ79SsRFrXAhahZQDcYn/5llFo+IXmCBvjnzDvmBd/nZ
esjlXXX91cSMRTL1X9fjvky0FTrh/TGl07MkNNCWrEkmCZUEJvkXTEcdWbS+MPQ1
mfSuDiwxrI6yRKmKks+ehc0I3cy5ldHig0cTKeDKtthCb94AevFhxg+/O5PvB2/U
swh8wmZJUEDdWbpLVUngHj0oHdG+SItFRC00Bn9jNo4s08hTfrNVpCEd2WaAyh31
ebVwCcUxnrWXwpYTE1Hv0JaYCkampiNFV8yGQWTcjiF+qzxSoLPt5MTBofTKGLKE
Oa3QIQgwKRZKNn8U02qaXYd9r/jkazjzCGfAdkODFe1345kdBiosU5z+isBmEm3e
2VVDJAIMx9IvkEzxC1GwD8r5t/nWruES3AgSh67W5yGslH0TMAxvnwdkBuyQEBLK
qXK4/ZzGBW8rKfDQlb03rpjASQauOiRgMiuNsrVsTq1xPloywjrBc9RSGjb2LK8y
UNfKigFHBe0Pl5O3WsGT1XabJNAjo9zpg7QV+y4krP6EhZtjj2ercLK2qEIrwVuw
Ji+f5R2s6ruynEU+OV5zwvylB2amzWqk1jTLATezxsuDQl0n2P29ID6ca/TzIS7z
BQ91pPWw2ckYTB+5E5RrSYpejBY/wkaeqrUXQqKBjeXUjj2p5Sw0bhn7gA2pgmwV
qIZSdC8YaikhnUwfbNynrVx6YvZ3RyaAbjtvxy9WHmFT5+iZR/BgXBhnpGZicNL5
3l/SAj+ST1KBVVPZ9e8+7tl4YPccnwcnPl6G7VDCwx+I9WzBZ2oxFNMon7AE+bwV
44R6Si3ax4UVaeL61F2wBMT7X6Avk2lKnZMeasDHFlx4UHXZRNwyDg6/b29inz5V
U1Ylm3BR7IUpvr7HX4Y8qEQpp1eziLk4TZegrLTWlZST7b5zjO6IFy+RfZgZtew9
QBJ/ERamZze2wgbQ7Sq/A2FJaf6VcqX3NTBFq9gqR8vb8c6IFs8sm21RaozVtyfA
dXn2ZPjBtOOrZthrnY8WqjpvInxvLALkx9QRP7U1sAzVhddoqbFxMZEYg//bG2b2
JtFhChvjWq1q4oyj2WWJf1Z9J7NRktipWOfgdIpRL+6GDrEU9UhCWqP5rIJKwuwB
jNAWu4z+Ugors/wvnRyKlzbvzzBQJlxQjApLk8ZWliKiyNnB72rVNgLGbw4wDXY3
G+BRwNhiqSAe4EY+JtCzAHbnN2TXE5Y3Ty/31kqemJMMoomtTtTWf9JOH/h/gJQz
fbhtR0t1RykjKhKvZ0o0R5V8E+zbW35KPSV9ipUdy+DniLOrg1AjQT3MPDbq8GWH
WNAazr3G3fcwEnmfyzEsqTN3lqF1J4SkUNv+nrgCttN8w7Ba066fraPDvSpF/yA0
r/lbZEUyOOZjKNjyTErXU7bvNEPBWUJOQeR8k3In42UjT7ctfiTdC+syEZxcs2pY
KkCubDpS5lFhIxVabPFCebAN4Z/1M0KlGIlAgLwHbiig4/CrdN3awXEoifyXZPhT
HB/7Pmr0eiHHQ41KlXEebLXcXTaMZNtIU+O1Oc+4Sw2gNmu59KrrMXxSNkj23Zkq
vFUAqJcLOYV1Tb1dF85RJ1Gonq1bf7wMQTcHicBmO7bN6uWQxNqvb+/qNDiECB+6
2L3yEbYkMjga4ntcrm8ht2nu5bdy9MtsUC3d43mby5WDsLFpbm+Tiv2dc/n69sm5
43ptpQOajL1BudI4wUeFdX5vSJsiwXJxlIsmXQ/jANcUJi7QrmFrDAMVsS4eLNQi
Lbs1vpWVWE9PshYsfov3aJj9KMaSQHfhji2P81Sf1fGDEjfjELNR8vA3scLI4inO
7exBGXzFAsirH+kmRMt4kFplPUfIuGE2MAi0CTuFDnjSeZvZR/Hc5XeR67VULcy9
zHkRSg/pbVrBYaWV+WgE++iss3nbX09K89ZAw8bqGtZG7Cbet0FfgHF50nv+/EtI
D/tYpVD2/euh0WDHkmiokVkkkxQGDgOLVKZH7rbNMw1UDDjr23X5I2SU8avvvniA
q6NYH6PzjCo1VZ3H5iBAqOiIP1pbT5fHWlKSeei5FKEorAhcqDrvqyJ179AGpYTb
4v10j9HT63IJXs6dI0bfCALAlbdMwtgYvbhGxTXKM/FJywoTR388usxJuz9YWbTr
8bC19cTe15TMkNKwdVaUyVn2nLx1dETyucMiUE1vtKaC0iTSrbSTanAk+1aJUWny
GXHGY1C9LJ5CEWAzI0CzxTbPxmv5ZWXKCsoCdxtVT8VL6qjX0U1I+yjSaR8zBalE
sgGhkcMenXCKAioCthfvfy2JE7i1bUTVnZxBoGjm7sfDCbj3ZykV03xadgsqaj4G
IYxQmRaqpdGGUvBi8KlSlvKDTrje6N5yE0uQPkfPo2H9miFJ6KEglPyifzqBM+ox
ifu/9pUalInZ+pZO1DPhGIA/XwIsrFCaOp+r4wyfENlvIieYIVgnUNbGL6cMmxEa
lDAvFyaVolDnP5ctV2lG4lOsDjJU6sT3AV3fq0MAFAPvQghGlt8Gy4rsIjYH7fvm
JdnslB5R2d1nETPhOWab4GGQ6FFaIlYOnBx3tlHlH7PtiwvTKyVXmMs9ubWMZBW4
krC/+ffHbrOPs9kYhFH9bYtT8KKbOqvYSWeeBVu8jsjYqCMNt+gC5nAcDkwzMhIW
cTe56ncMc/48BY468PMEn/btQ63Lzt2XYB0GoS2xLAZjMVN7wB3ygHLjQJg2Z/D2
UXcchIMtmr2sAbmFFvGzSEB99ACFmzpvche43IYtkHKAII+Utmp0PQ+loUttFZUc
0Lqu4Q+PN7tlfoNre552bK86XC6w3e3hvBg8M4/WQRFiE6+21rKxbGyw0YNaArCO
gPY1y0QsFU/hd8PFKnbYWaktCZg9PJHWh7mL9yvsfH6O4ai7m4DB/90ixQOeP9FE
+V71odu9TTyO6Aq+b82x4Fo0vmVO4ZzK+lGnVCm/uD9iQVc4pV0M6+hs5hC/xioT
/FBhWHy9+tWu0x6d8N2gEn+2kd55OruiMRZZ2njxL48Zx6mgtaLN4uvsveHsPPcW
2YhhgYk7Ey9SVXCFNwfB+sMf9UugfhCYPGf6PNLfCFHaYd13fOh4gX4WKLD6Wc/I
/4DADgtKNWACdekvtQR23n/xpqhNapj3mvLRYhP0bv/KPaHeKJqzHF8wAUjGLxAb
wtwqMuyt0InYhw4lwmqDnX31/mAofTlxNACthcSicrKTv5O8/AzuTTfIqgoviXTX
j+FoeuD375SU5pQ3382l+0DEVfp4YaDmKhDUsKCn3baSXIr6TzkUbw+LHQdenILX
mHGDGwpsXMe237jNHeQRqCMpi3VSj5/JYE+SRa3GMHsiRfyNgDz6K13NcOH6FEBh
Ukx5jotMXw8rN3jV7Zfj7PeVYLNTY7ih8yjnFsEG8Gr8IiMzp34uaGLs/kj+mclO
DBWtqVkHwapzyioaGJdq1xfc0LkBaREmVYkBlLaR2KP5kfcBV8rmsm0JujdflzFl
OKODFOBQtnojuDXeyeyvhvY9mBByO51i8EgX1VJ3hezpfFR9Xpgc2BtvhLAXsmbq
w0w42IOXRJHVOjMBXLzUEndIzBTnOS4r5u3cP08w2obhuuiJ1pmg29DNCBCd2N0D
XewOKuHIcYpEjAhhQDxsrmaJfc2oTFmG+1VfjMWM2++L75KmgtLvtLw64a3YhVKF
6YHclpqmBByoPFQISE7SC2BbncbffM3k/owscaGpH0EytCwx9i+fJ60Moe2MO6Pa
w1gAw/NLE91A7s9KuHzLGwU6D7AfvWSqPh0jY3hYd/WkjIXFX/i4aOnlLsKBuxpB
kbUa1cXBjWZgh2mTf8vAEEJMitWhNVaQANFlFM2bQfa+aBEuVZ3MfIhd/0YYdqUM
J+sdtZDd1guco4mIhhH3MGQpsa7f960cNeTsiYSNNArSzpLXHz+7nVP2H6dO62Zj
FY1Pu59Uu6w2qPpb11HkHqokEkwkp8fMRo0rcpNXicp2mtQeVCGJgK193DVWIcbh
C4L/v62wEwixMppXociIj7FWTAFfSVyvRYZulhX5cCXd+KGBkRJWrbuMvClHxTo9
g0wAsaf2X0Z/oVIdt5tvtzql9LTbRGTVU+XZ0rDtX8renrNjbpHBOYBTz1lXqk+X
2XFGwRb62Jio2w0tEUekPzWGPDyKMo/ZZ2XcN1YSLwTt6O1NsLdphk9Gx2tn6SK6
+RPQsV8h/SzRd1/h27lHFtpAUwgT1vw0Q3tvyts7DNs6mQymptdpVGN/wM8konJ8
u9Y28JO5Q+glJEynLN6vcFvWa/x7kyOLwOilexUi8pFojdFBVqqMQUbKF4SgQa+w
YkqnftRp77hZjrBwEGUfvDhzYn5wRiRFEQalVA/lfJtGBIf0VLYA0+4Uo/Oqr+lU
XJvnPiHzMYxYyjR5re/+LbG8y8YzDeOV7XdHKjoSoPHKC0WdYtH1Sa7dJ7n/AcSl
W1cesYHgDo7PHP50dO3PWS2fjyKJQhm3v0Upn2xe8JjxQM3vTbnQ8QKaZ0eQ79n+
SyfWewxVaCJ6YfAO6UZoVhdxkpvLA153fStqTeNgac62b36EnvRohW0tjBh0E2Ww
Pxmh/KWSrx0dyT0qmPjjM643/LvAUOfE77IAfUvQor/YVEE3yhh8soYqSSRAtZ16
WAedXOWL3SsQtUKnG2X2BdGY95dVJpAw7HD4g2+BXqP8ixx8rKhLPjlutyyEhpVG
7X+Ia5zpfbiZY9k3OVYXppvjsTz7rGZ/WrAdws4iikXMfXtiExxLBfZgg3UXMAk2
cLmvq/Zybx4vkGefLHjDgrTPL8voLLn+xcUoVbjhtzpAt5R0lAnC/FtyN/0qqguo
gNP02JnaDScttiwOuBrTYJJl4PCVUWXw4jRPBmHzwkOmCWzrzWeO3NpauomES+Uq
byNiGnXBWq0NDkqWA7r1d755tYBfdSlMiIK5+yT4Zy/HX0aNog6EC8W4r3fIvVs6
p12hOq+53pugymLB5TUvnzn5IirMKJIyN6PBdeW8Ol/ZvlEGH/02fVo3jWZDhHbB
jbAlRjFrWx2SvK7f64vyNPHGLRn2Qgsi+SQfb0FT80khzQf/OMXbGy7efZlsH3eJ
0LI5ECQr8pn2Uy2pNZsV76J9aogn62xEA0uQgKDjMZtL+AsR6Sl885ZzVpg8UilC
WG9YpbGehu2aHx635/4a+oYWgGzQdFVqmVHyCG/QEjCig8sy9O3vgFIjoQJu/4wf
yyTL5151knn0TXBhhD6g2g3RUS0B/jd46k9I1lEKhiIUbjQaC+F/gAo1IsgivgcG
haAJz63+z/V7InfmfkJQWSQASclRz1ed4U2hfM1HN2qBzcAe6g6CF9iQlW1KpdF2
1WuCjZSeCoRu6LR3xvHliTWy1NI0jUxVTGC/IlK5KCG0jYAcBkwLgiIwOJOxIHCG
sD/KgsCN7mb3PavxfY9hX1XYaOv2Joh4ViXpZzFwW0bnpBow+qfZI4Etvg95i5t+
5xRo5dF3y5hwdiSWUGuSp3KX1mNLkHrItSDRFwXDBISIMsk4pk+2WnEdsWa4WShs
fm9OPHIzIK7SKhU6nTBAgWX3K5V5nJalVk6q48pCmyc07k1aMhIA2V2GTay/CAUQ
YTa/RMJmYrWmF1e0/txP4tXEwQVXNZ1wtRUhHhz/3SXu6dZsk+tsmQlhNUQxVWcV
+/kJ7jO5Bb/oDjvRfMMifwGTBMASRXKFIv7EAq4tf2ttXZXhHxC7LVNAXjY7+Gq6
/mSRykn8pei0N7AF4lX0O0+3kKKGfuGRQ0nsZRSfHC5o4H+71QRpMsuGHcYevL7T
ondmv6SsKDUd81CVdRJgtMb8KJMA5j2XKh5tuBSs1MfiIc3/oUDqwBhVep2xxHbW
eZ3rq7wqUWlCx3g0TGDHB04EeKyRUAr8ruvDRheTD/Rg6vJswr+ZtQWN0ELnpILq
DB837+W8BP7gr/BJxLSlpvYN4V0/zXF6kViyGORh6YaYZ6e5t3oQ5/ZnywX7mux8
t4txE1DBj/m5b45H3RQkduWN895ONiXaRR4wQLU1jwzPVfuv1lPNYf6BbH3RwZUw
usOA/0JphGwPhAKnjACFnzmzmwWgsDCX+AJpCxWWqTZWFreqEqB9k1dUTigiwj2N
/RW2wVlWQBbibh2VQWMybYJ6ClKT7+lAsjY/wyqwQZtt3JxKcz52jzHqktVRNxhp
Sj25xCb5xEiJuLHqBeDEc0w36CAWae8+t18e6DOVV9AqXNIYz1p6xyIfifdOteXU
WKWExZFcRzmwBYWUQdSXTqYeJmfGRq3OkJAvvoSVCBMXrXmhu+2UNwED4cQ72sb2
HDrrreoSxGCoKtvJeq8BTJ5exmPBRrZ/x0mje1Osclgb+aE9D8RDj8sFpVsWXsbz
Z3Ln+TZZlykYppEWGLkbwk+sU2NOhoEdcNt7zfFX2VBRl+XqbVwc+45GVwNEW2p1
qPo3Ob+F/MrzU3oNOigIJSeMB9ZX60/sH9W6PmmJA8OmoFimx358yvJKNFSZc+6U
Ut667SVeeXjq2/ec+AQaIhbhArdbdCrb5n0virDpmt9FAmnUg8f5y9+9DPin7H14
dk9AUDZG0pSHwqRrQusZ09eWrJ3ZGt7KbWnA6tLke4PwYucbOf9PZOhOqLYvG8xA
qmrfGvMJHRWEdWg0ODW5nXnYjfmhJxsvVqIiuHo3XobP10IJDdL2poAyIAzga3Yo
sRlnmjiZxbcIj6Zxx5KR77S4UjNg/d3L4lSw1//F2OXHcASOtPR+qhZqQpkOd3gV
0HCWGMOEHmUfHdP6wKSKQU1h/IffyUef0KWJltuyRlTyXceeNm+lZtZfqk/++dTc
rVArz/nLU9E4ypGpBstJL/K0GghYZ/BEKUPMi+GUugZhmSQIDLqhIEL45IbolMoZ
zxSAMmyeld2dEWZ0ygIZ8C8Xy3pvAs3iXZJImKTmnY9ErqmLJRzZMevdNZUnH1Bu
zw0rn+ALheKpXVvz2dlbsJ0/30tYcjXG+CIvHKN4fccQklGe2EkH4UcN8cBHk2Mp
JgwaBproCGUSeLG7IVdqtZyuD3faPERwDEkoqfdu4RIUbi54KU+TYvv80moZaQiG
kBV26RaRej+G/ghlBv0u9YihePapDLCFlJ5h/jh3AZ/OCZRNRHYYkjd7tljJtlGD
7ler+7qI3Hl1ZQxarK3CzVNfL5XpEoFvZ77SWQ1tfpQ8iUyuUwpgT8TVOIwdhjBH
2fT/WfBsqo3ob4a2JOUm0wTqZ/1ucG6ktORlmw0Q2C679Brq+XSBYi99PJYwNMkw
Cs9i5ynuizZ7hnXokJP2+X0ijPySeOeVjTVIJobQ2msPKkfTL+cs6T4gx9I75KYQ
XKXOfe1QToMfPGxl4q16ltHF4mHnCRrqmvt8qlitKtaI1sTfYZR+xc2xtjeqY8uk
mg7ORqgo+imktSrH9nGKz9DM8Y6MvuALgcsUSLJ/rwZ8FzZZJesWGL0Mt9P+uaIK
9tStMM6n8Ens46tkgn6MfTC4uEt6nG9ABBlXBpSnsBatewX9b6BK7fYY4Lw/yXlk
ihG0iytVv+8bSAPAeOe6arF3L/TYkg/PKQJXx/3q1IHNsrqZYtzYIdpZ30lFAVJT
s5YVyfCDhuTJBo8bKH9ZKxPBDMqaXjfmy8j5hP5969eFo2Upps/yW4h7mgVHRjQn
NLBPE5SpvYHk2t2Wu2sUUx/fK5ClZfNoLH8ljha9PIOgjIAw+4VK6sMok1yox8GM
iVwImNat/MxwID5y2uytmcBUWrTVX6FA7+QmiRuLiEVRFCPWrSPWxVHzz3xyT+6S
C3A0O68ndP/okDxw4SxQ4xWetis6nL9dzBxuB6gGLrJYmelTfTNcdQ4OH3BvYHBI
kxUxWhnxWnpKATLO25UxXfiKjeNo4QxGXStlDd98P9XTyaqrLTnhaYyZLXyCvRCo
TYQv5hQkiT5gDNp0CoVgxgx6Z4/H9XxjWBnOFxTffU+5ZMqpyCk+22UIggJbUrdg
hlDEeIXeQ/WTOt53T9Q262Qg7ieAO5v5jLDBr8+495XBZPlHFP2HA/5WqPVsK8WM
0GVgwsAIjBehtYdW0go/6JM9LB/FbJCBFATn4gpbitc38HP105Xf73LrX1khXGKt
M1sAZGYzvrwthOYd8ztsJShCpJIFfcov5HH7lBdXgtd/ORxxiwOLq1Bnum8cZVkd
3a79HfZhqhqvQzevgzEb+OG/w1a8K+ZYLbriziv0ztBoYO764wUw6QRwNV6CreRi
eLCRk5ov3RnLbSfIbgjHfhanqaehSx/Brje+EWUICs3km7WqhWM/RcGSX6icQjTX
yPCNnwBewDIvx4/YAUTQjOWJ7R/WegfjLpBDj2SeLClAzfuPM36oe2/HfqQKnbSQ
BCQcw/+ipn+bllNJ8X4opNG7hfka3FKj/LjvkXcruc1MCN15JcKa+4MMoaJKjJNm
3yCGRCK12cgCpEUxCN7rKnN1o0EUBAvNLZKjQj0tL4Yw6yAv3PyYw+MU6SGRcC1H
LSr5rBhFC2INAOmUwI/u3cEUyyGyvaO0n7CBZMKshJ3nn49sFkzzVyDSZpiOmpCM
t1JG7iAMmw9JPRwHAA7xJn+5GcYUa3FJTeS1N2lG17JynIyhu48Qg3mVl485n//V
4cdQryfgIRcFpZ3PBm6/VSoRJpIcO2BtZSplBpBQy2XBGRDnzqS17eqpUOnUgN4g
Py314CuB3iMqbNxXlhUGaT9k0zdp5bg4QzNTi65CG8/X+9V5XfYie4QlNgV0mPOf
3zXddkM9gnXugZZG4fxCyErA6nXvo3stJlkxMWkyOia7FkizUcjvOndBwD8HJmDI
8m22d372QpjchwLeeNSAXAih6Unp4dzUvEiVlmQ8gLOBp1bp5eX5zl2+EYXIiODT
SA3ty+pt6viEu+xVLhumZ9DOsR5jVGnw3edQWhS3ZavZ4ketYFppdkHjoekvUEJ7
xl6yXRmIVLcZQ5W8RVbvLtQ0quVphppP/r5fwd7hGCHGiaePB8zKYrGsHjAbNtJR
Z1QvmPu8HmbBXN/N+XMuyoox6yERVuasPD4oyDkMPemI0TVcFT/B61jq9zXWu8HC
LaKmWDMqlJnjm+VV7ucTnurJ53eSUDyeCzyY1paA4rE4jtNuRRqNmnUS2m3HrMoe
2fNSxwDcQCmImPFYE3GQfwyicZrW4TTpah77JmyG/WRsHDdUyjC8HhIz7dZyhajP
6oSy6S2Q0LIcy9oUeDt1PL18GYvMmoVASHbJG60MMzVmLYT2VrYrEF8DMo0Xn1JG
7K4HNMjeltNEVfHpkWJ+i4MkIesEdT4osKZXyBrKnBSCR/RbKsZxLT1FGhVmzg0d
7Q4ldelydU+4Vmt8VYltRnLs/VLQvYAeeGnkgAbkLnS2kqI8JtTBIG205UyUl5qu
5YOiQKYNRZLZ9e6Vduei74gLz71Dd3sgeqRxZNNNnL9WRF6ryL5cCzxpPv4d+877
iphnzHGqoe7Vvwp6CMkaMOgpkMDjT84LUp81UoIJmpUbxFQtFxjWdoBbmGEKjbWm
QDwOoXBqpHwSKYAU2uAGvedVvreMBLDHJSPmzMRP6TavZNgXG38HRX0MQiK+/Rzr
t+vYf38xBM9sY9leRn3QxIH2EjwkTO1P77HbN/VGYHFPKoW80Q9SofK9FgsYQ4/C
GjPn16pEH9KuTNdlmbTgUjhJQt3F2/r/ryNdmgqXcOxx9dnX6GRWp38n5uL4go6H
Op0yK6MffOIr01fw/uRpNGyt/T1sr+8DvWeo04s2iuCsLLmX8R6s1fJv5J0mfTOJ
mnnbi/KpvyydaK3OXbh+PguvRVhdRBssH6NSlCHwOMZowTb0AMI+P7gubpDZpu+W
QDpAESAd5oD8TmTbxd3eOQQ54iSl+vxQMXMn+MLtoMtNeAfmggXqu2xVmX7LnD5h
Ta9sbMpkdXMhVdZYxuqOJVIjYkkbXbGwVHhLGXfHZdDKBu/tQp2jExqELY9ai0Vd
p6XmPgsL4AgQkqWNL7qXdHLKvuvC3n6qGmVBJOnnZK3/yHQo3BwSHd3nyJXdKWXO
ldKzJDer8VywCG3sXGqvj6hROI3iEWq1OzWgUsQod+u0dxpuUyABQBhddMzK6yt4
WeKqllnZXcCsIHm/Kp5PwNF2ac5/edln+Uj+3HoI0wWF7rTXUlnzQazqCzA8aZ5M
CboMSybbjQmnZAv7Uyk87CeYy0sTy2lw9l7AmfpBh8wsl3a5GvNGIeasu0OUAqun
1pxR1L0oP8aF9oo2L1dDKfeeEXS7XYUDmbQkDVy4f7ljcNJBMEYGL5DQKkAgNdFA
hUqdQH2OdpSc6P5mwx1hdn955kNDDzLptnR/SrY4zNpCsLyLvaPc1qRZSfgiemb3
o0ZTVC3NU8nq9vNzGMgj2RAdgodjDU0rX0ZtB9f/lZsQEzYjozs95bLZbyuK09n+
G5Ut7xBJpgF/OO5BQy4fUapcmAodmATvEX2FE+hgvqtscac/i3lmS3i8kugMBJ/y
k1ujTwWjKy/tmjIsaBB3SCdBJXXE8xhr3idy4leVMk6SRnF6gbT/iSRmPlauOyP/
jvybmHFA/PyEZnvjrohYA3x/fp41aGMNZHJQmkjckc8ShqHYUJMBXw3B1KS2btAY
hPLRq2+hriPn2xaQ0oflSsuN+vVONy1z50wCowzj/rVyd5MGHee3tDi7XAk72Ps1
zlHxSAe4xpOIKk4aR1jZZ5ZnEn18MfUJW+PBuSS/0ubqzH+45Li+wFW0kI8UPr40
pgJbGH8gMb+ArC2xv1FaJs2xjKvwQ2vp13RwW4HTLy525b7skqJe4+IIMYgYDllf
H5Pq8f+7Jmkzmy9CASMXEpNJKQqKdCiPkJLHy3dm2bO1aBOaREJSBFDkFEALgcko
LAKi0UZIjJmo6a0s8xxtvNCIUsHQUUC4wUSHWSpXCFpKXf/4Vqd1N5ArmjagtKhe
vEvJY9mZpArKCLNfCHPZgt9WGuG0Jft2geEtuQVGHMpcvYIM6A+LYBptHp99y5TD
Lb4cwUlFbCb7E2ovZXiX26J+TmPrgJR4hUQseY2quTrdjSKDmo1smXpYdBqKze7U
FYyUleTlU77PMskX6rwATD+Xa1ff3VG+pgrocWn+Kz1pWZ+WOwwoSSdjPDVAhIMh
IQLilwPZ1/Y47YiArC2TrIk3Kbfh1flA7YVr6QwrUhkhT3n8BcnY+rGgMRZ9lUeI
v5Z1ZHzekgPGdDaYAhn63S2QzfbmEFSXHZEGNLa8PkWdxWAxK7z+ed4nGqvVUfPG
9bM/Epwuqi0QYJzr7XshNaJ/MpZG/Xjxc2/+LbWaT61Oejaxyk6/UBZ2vj2WNqwm
BSiY1W0Au6vp96I8UQ/AW12JqG/bzPD6Ga4voeqwpZF+IYLbe9Z4GB6LO7AqPpNa
7X1sPJL2MzFtaWI0aM4XEevu1kggdRfBvXIB4tE+Ou+RIR4LIHMPCVnm4izbjNi1
d7vTv1K+HNbFFGQBJP5vwqd5M9BDoEd9nSBhgpJX6AssHaTK7LgwzYEWyiXnFemB
p6pMNu3o/6rzTEWU1BKdx4vTr9r/HbQ4Hswbxd/CVAawyuaNrt0w9MtTtLPpbUzn
YkhCrcBarl5hdSLvj0fRbKy2OyqmiL0j0nxyUgOTi0X25RbQmwt1tMdFHRu9CWW2
w0+YETcT9fzyezr+4nLPMDBy8eGtP3Fjgq5+/z6S6xO//ggfhvrSzpxxo/H/+2ou
I5oUYidIY4HSuWuRifbmqFl3n0JpUC8mn/P8I9Xq1+d9ZmWPTF1EzOJ6FxrK4b2B
AzZE1MGouwYchHVZBIgAHKLMzYNXGYQnpZnuIxSCMTlpF2dpUs6ntgzfI/9Nf8ek
Kv+Fy7ArO1HJRZm049NsjfeK42ihU+AvOC8sAqxDqWTHdxOReEvWNJXosZNSvZYo
WcOXFGXqXFHZkHokCvhCvEAVtO03xFeuELDh1jpAE5jIA5Sthy9is1mDwv9koGZv
JCJXi0SJ8FLWgU48+B0CFnEeWT03sj1L6kgLSin8zdSCqMZTrhi9VtW0Z2S/B6qY
+N8hrHwSa7amuqWY+czA9a8aEponsge5VCb3WA11TV3Mr4W46hoxfsvH1DSMxQjP
svXyG8reePQDWO00Jsfb7Yx00sBVzb1tZxR2gs9s49vAkRjie9HntCxhmljElLTF
PXgJh9edX/HklRYMfrmJd1EmTwtw+Ze2BAfCah0cH6SzeDrTK4s+WtDal42PrZ5G
bBh3kcBtDUPc959MQQbCtOPoaA49zbOo+ll8ZiPJNhF4FnoQJstzllyTVhLNHy38
AiVaITXzSMWEW/KMMazw299UubYANV5W4ZuuooO8qYRPUNvNlOg5hcR+2qiWKQHM
Z9s1NreAuYxu9ECsLv0QfWCMkILMjX8RNaN0qGi71BvaBQ25dVUkcEKjP08xLM2L
fpHju1f8w0vIgY40Dm+IJXOY9KiL91ogb4VzHPM3GMyQ8QtxRfu1wBxCA2HbRjfR
Is1qO0Aub+RZxRbEubXLkaXD4kbKCwoVdI66DtuKSordo1WPw4XhPVFMT358B++n
dOlh1z3a2PRlfZqCuQcGLMAGu8SI1zgA3CmDAYV518AabFp4iQz3WaSU9As3ofp1
R2KJ31Do/COoy3/JpPvqeFpSmDCQFWvNSbdK8JD1tARyqPoyW8i3Rdi6oOLnm3Ba
E1Rdko7yS1N2ozl7V3eXY+ZL6nwO9rTKnLlGIZbZL/z2bzqMJptoO+1mKuFyuzmU
mMddbdAJJyzKmFiXy1FO5JaJkTwJe1nmCFvm/28F+MyPKWQJp9xNjEpkPuUjSIcs
OPFDCD0U2H0geTNJbkDSynaVvI+u0FP+PQ2M5BnNsngilq1Iy2PyJYeFprAcX4fg
PJuQu7UE3xEoVjTrxQRM4tufyV8DjCNsK5IcWYT3yI4wtjbeoqN3fibUIC39DBrG
EESzwgGgtmtqX1OhiALGD2SH7KSGcZ/e16a7mlfCE6A3luF2i4lZF6VqdqLl0xH4
TVoZSZEtSMB7Ejh8brRFaAPbBMvu5tck0NNcKoYOD2BMhHnm6qIYXAa/p5mLGrez
lDg4U5eqqZo4ysOWlmCvjdSS6FgNiFXPUJIx6ZXMEhSlogMjcDgYsMpsnHGpQlJv
FXeyeJAzcivivxe1xSLVmRgHpoQG2ST3cTIXEFoZ8cfbgermDMItOh9Dxchl0qE0
uZsa9gpBoruyHCfp/A92MHTz6wyhBdwsLg5e81szlPUpRLL5dPzwSQ0tCMdUdkb2
MId00M+Q94lncjssu4WQwqMObqKF2qDFpu0UNo5W5V8uTRdlujawxAJW4x2IiaoN
33ZZDgx+0Ro0UJWViWuT/c8cJA7iDtpqQABpwjDYh5xJpYkKhstuY4fS/1vSZqpB
YFMLtgSxOYt750EoQJqazb2UF47UA7pRX1R4pOvdq+MHTjQggHo/LpHEYsukWgOP
ZtiAeKvQaSCxCGZPEVcKDNZcYCa4+xtDDdPC9/U2fgt7W9HlAIqT8J372sg0X6pL
UVV5HxV0xuNU2xGC+6KEwNjYcJVNIGBT6NQqTrajmTTnHuiHKcj0wIMJbMcvsFez
tTagwEMOhmYO2dbUtMNI4nlFGqtZGbpXLuJSoDpePQAJELMuz9FRjOUAChMpBwVa
PMv359XhI4BzZtfDruIBNnxKhCsPV1J1PT89eloPyI+fnBSrs3aTjxg1Zg6aY1u3
QBRVsxj5vcDYa2pADzGc8Vglp0gqOQTV0bFzqTZCzlhUYJf8oEd2lni7gphPNDvn
7l8MRlm3hJvAFzoMYx6+zuGwbIVkyGtj6U+Sw1SU0fdeC1tuaCPd7JM1GNGC0uAc
8htQ5I0Tr+xyOlTDUFE9a0KdZoAZQ5JN0z503+F89mU5sE7/VfZUtAn1uIdZK6G4
tSTmLGm0QZ0/7ILB2sBImtRQNfVWNyXJCJNvtHZ/HbMJPa8c++Y8S2ViSBvcG1SC
SizAhDfkb0emEPNBsBoed1/JshUyNydvFuHt8slBsoj4w54hSs/bjCHF06UagDb4
T4EEyEjDNQO+QPbkG+nQBOnP22WSAL2yh0meGL4yIp0V3nG7pgvYCJNBztnuh3r8
CFJ5kpmh52c4tDwup4mm5C4bHS1nUOF01uan44erm8NJMb2TyLKp8qEZF1vKkSla
ts+7kL+ncmM2vnJ9RAAueKItxHmaxQiWqT3Yrw1usSZpPkDKFs7ddg2LDt9BuDRu
roOXfQm2/R9PwsAIrqby8wYi1ptuIFIGH8j20YOtjqMb9mpO4BvpdtmcdWi4ZbHj
xmZM2UbUv/brRJ2ChnBf145tSOw3oBdpaVHFj085S36E8jZpsxibi4zeSRrQ9LgE
Vb4RROoq11gadjXZ5AnKPEeYFULx75EBXCdSx+4whKSs+qxO2pQztjaEEYNFOO3n
7YYcMQ7/LfRXbi9TtoJ0fLsK7ObYUw7j/k6N47ZsXOWYyf4p5r9gzMKfisEkq8Vo
jZ30AG9G57IzurUM7ga3Yq1Fs6Nln69XyRpF2cMRa85fxhaYd9wLp8orR/WyGt2L
51WK09MrpsI/bUI01UtenBwwxXS6F5kVH2bgQWWgK9Eu5z8GmMWhyCA/nwgCqwOt
Ki4YaAMjh8uBL0/uR0rlA5UVlwWROor2oO9Z2O+gUxqnWA5gis2LqhJgGVx7J7Is
nxcwNim+AuIqGKpb7eaPj3l6EpTu7xDqVs5viaZR4BMxO5DI7qek6JNtqJDqtlHn
CY70e8MNZz2M/0rd5gso7Njildohy1/CPJqssZ8QWRfFpu+vvDKoRgKlJ/v0w7Z/
Al1htEPp1RMiVvmCSEK8b3oppYEorKypEdQ6wsvAnMdoHOjlduexLP1sCo9UazD3
yDAi32kmjteFBFovA+KSVSD5YOV6QC1upEaRxuSEIIk4vN1ZdwAAOnkeSkJq6Vc2
tI9hxsrzlWg1/CxE8GoUl6Tjt5ZigYvWm0DC+tDc2XmdO7EznDE+2/Pdo9/M6Tu+
7yGAG7yn4AI7UWu528pbalErIsVFEJ6GaAFyi3PmEAOcpTidwpxZeXNIUJ1nuTSh
9L0TRH9kWU0CKZa4dyoiyodaqseHfDc/kJoAjYyhk8QdEyXaUt8bNWv9hJFAXyUa
h8ysUZCYixHeibvNw3QTxK1J2Ginp67JNTVGQyPbLg/OC4UGmQC3AP4HLAC2leQn
X3z28TegA/0j8OSQrVtyZwYkC0Q3RcsYvJc+k5R4OUe8Cyc+m7WtXTnThC+ItlSH
gGdNfiWwPYIo7Y1tVKR4ISwN4onoOc03Vs4VcaleGv2ETJF3jPSyU2ElixlynGh2
ESQTgpqZmLARp/Ajq7WYluuZst5bhUI0wdvykjVQ7hINsqSiwiyo49/cpLEcomKL
ihQSi7zJAwutvKGLnTlfWE3o+VwpbBlWc/BKecU5t+jNx7MF0mTZ31KJC66ACqLv
nVM/aHwLquiUYWz7AO8Rz5aMoNq37BwYsjvy516o77R1V/817QhMUss43Lw9u+yK
e6iQ5fm6kEdDbGOCJBwOYaClpizOD8q04Dgr5DGHaL1gDmYjUUdZNCRwwY4iE7r1
fsf3V89z2Sn8Vw5WZyZkBptOVafUL3p6d+YZxYXo8gHtv+t6kTX0L7X+r9sdP6qG
pN2HNktyjckjYkGZTmd16L2uLJ4XfVUxUh/EfuG+QHl1/cGmhv1OeD/HcpU1r+D0
RZHHMAQapYd9d/DQNNzdWNYpyxBdWC8DtthI5w9k88pXS4C07Giq4ULKtz70FvVP
y8zzduHTS3EiALtf0Rp/X9x+Sf1Jowwvhh16J0ZiXQKWnMOHdJLOdZTneI/3AP0L
LcGyzEMcl9/kkQBvj9wWXRizUR9mjD4MUgkMK1LKMm/06lQSeF/4YXA6yVPqOAD5
Br6TSZjMzCVteFRER/AI1//J9hk8J+5BIt+ahwGtrzBv2DqQ1FvvJO9sIOuvvHQC
/+LaPgpdAfeqWefdTmDzW76mre702SQiRyTrpAZXz4CT7Om67pL46g0OYA0GKSBs
gEA1CMDFmmB1mxPk0guQUgUjt4Ud4gMokjuEMcrEfVD1FadRBq3LAR+vL6v50qPp
iLQvbiXtc2OuNH0rBL2OJGL4iNOWbqeh9sNuvSnzhk8yw8gsZJUu+SE+SF5sw1q4
AVuS50nnPAPhaHClSjM0TkPnh4jYRgOsqthQ++LxPzc0jGux59IF6Ml/UrfyvBYs
wxQfe3ZEpO+xIJ4ogzYltd75zed1RgzGQQskqt4w384Fki8a1ugM2pqGrsZyTxio
Z3ijVvKjCGyI+fMQVWk+l5A8tIUnCcR9Sl2/mnC1IEvla200bJB658oXUy+y703I
oxmDLs2vYVRiArTb2AN9ef5Z0HgQP/srRBsL6GE8Q9B6DtrgJsQ9xREvYSXTFimQ
SbPfX1DWlA8F9cPXKMN1m7YzN78mTfn5yyV1/37ZRiEt+MmbhURsFWFOUA1270Hv
pegtsZbfHoJ2bXRwFmTEYfEtIN9MZFHkjewf09hvkNgH4k98S8JJJsrHG+oC8rha
pKovfzPyW10HVAYhLvJkBZJT5zwpHmUyuh5BCx+b7OVJnmNuZEJrWXe7Ymyd8V48
UPppCynRix/74h9KDWl520mXNqUPAs58i2XZjYzZbVcW9QmTe9G3jY7DnuOkLcDL
qMB63kP+wZOQTrXnx5ZPkTjnRySzzoqS7xiuKf02f12XgW9Ba5W9ZLTRx+OcVWVU
240w4xoudpOIBw9XV+cNvniQcTiub9NAMduwXit619y9+bWpKPdF9R3CAvzMVPw4
Z2btU8C/R/sVfOP2m9sKQiVbPpt8AbSbhCLWBsc7t/zWtI15Qer88AHjqiIu84WT
7sKvVM2LfBIfuB8tavSTxjQxgm+YWe7VYDtBjHVHJxUffrawRRzcVLSKqh2pcT1K
5vx2gJRhTGs/gqOKuvl1xG2wlToN/zXVqmo7zIhVcNIkyv08bhy035TAhOjWC5zY
nzaRAmd2WXwXIhV7jxSu/4CQoV6O5d1ZL3plXnYTAc8tIq+x4P03/p5JJWzINnz9
F1CZnnhWUt51YoWaVimOm2OPg402sefJAoup18d+iB6fgGUexvCIOLD86iOGX3eC
UYr7zPfrzq3erD4O9rj1S1P6k2N2/vxypCYUZESk29XsJ8J5tIwL8RrrhBxwSn6G
XRfwzZ0fv/0HsqlSA/07ihs81OazTDl5XIc4ZjOHctMJ7aDpi/78gY89WyeEI2Ni
0vGN34vHbus34WZg6ML9Zf/+aDfY7+K9pO9/ufKuELDpY0oxd+2JvhUlGI6YHO9Q
NTdVw8D9JS8FSxWerCzuHoKieynGyEfn3EwjnJYkY2pDUCNSCvrFhN55dA1lQfZ1
aQqN6KrklFy0aPlIwDZU6iLrUqLUjEy1fHOXBa+nXD400bQzfr7uPko6P0zhb2Bd
zGDapN3qc8l/fif1OuK3tXioYTZ3Nkks7beWPvxl1McoaSppjTcBC4h97zi2OtNQ
/FqQ85fV2xsdXjg/tZ944zgmOwrz8CPXh23XWtfOAlbCLGbJn4luqhGavmtk6QwT
g/5QRcV6Vfr+YlKa9pINiV6843h6scUa0LBn/pa05RTNLty0WXeRNI14wfQUMr+P
1LayL8OkcTm8Q7wj+ENLBxGfgfiAXXPDCzo/QX/KAJCrS/7GA8UdeNGbrWmzNTGp
MCJWmqhDxu1+PdlCefFnrnkknnwaxQ1L9vuF2HJ9ZTWN8PXxjER5fJeyXq8Mtm9v
xZJtlSLTi+Ph0vI6mYs54VKpDhIDPp64d6MwMP/X8e/wYw9ifIODncAFcFPExEO3
jkmfgVi9XwD+0uWlBb925YPVymZ21cTMl/zE/NEKTSUUH4OvbUUkZNP3TDOBFjFu
yoIGw8t34zP9e9sR538zjN22Yfkm8moiw5BoIQxorpGh1gA0+UGEdpBYNQoBd4xo
xlr8Qu9ueqmQQrRq9HHAbENDCe5A3JD2hKsWR4xm9OF2NAXENW6dRX7nS4Pfi93h
3Eof+MgdHq09e14YyNjLFQpIXFTVSXcdXmF3I+T3F1Wwq4pb6bHN62u1XFFqtc0W
RjBUuSueYzdZBapcZNnxue0oYyVnLrmRbJaQJL33WVQlssj5eL59MqpuumBLNYav
Ncer4M436W+qXorBe0ZYnWECZ0e6UYepKuX7Q0tILuAkw8RgHWOL5imVWMZKiMQi
PzeRzJ8q0/hMGWJQNy5bbiFfHC1OwfJRRasogde19BzwS8ZShOdNPR+Y20zqyTfI
B9d8h90IuE6CNW1/XrfYvayStd0wM0nWCmWewqhVMCz5AXbnPyzTl0zKASo5OHuB
ssjjYyXMfsgUXU+2M2RvzmOIovGHgl1Shyfb/DqC+lHBxtRazQr0vhHN+20DGgjJ
Of2rS5JkzvUv309V9u38PpJv5qxh+bN/xc4i3rOC5NuetoF2X3IYXsYjnG7gbo/h
UbljZn3jh25G26qi1I7DzOC1nccMFDryd19JGFOqO4lGxcvFRHIUPiKvvcl/glUl
JRnH+K6+B0D2ooU5/ibWQ4u7AHvs3jaF1lPQlnW8FiedKsGq7eZAG0ITqdUgB90z
kFi21qBPXLRQTYkZ6+p55uGQUmA+hYPq/FzlphVfBNponPBFlib4UI+WgHZZqamr
3TfstYSqEpImepLUeIe9Lcs9z5lCmr2MO5GxKuOY9Pk8OTXhaINVvkqL3gulEKuL
Q67CQgpRPHntiPaJSkqw732H41hAhlpiL7qSjq+1A+ipQEa4o6hNwkxu9lLYz6fk
sl8iG61Y/sc6DF0ZlXe/LXc3FkGuziqwXsui7y6M9yg8SHf+oz6lcXGKbbt4yhnW
eOxIviFXVpR10D7Y59CuoUsFDsufgmSKn7zMek7HBlTaQhNyXoIuQoVPj6rIY+/7
d1fo0T17YqGjNz4nsN3xb4EpEPa8jtSZYY9UKs2wa13KBhytPxhlhHZ5DOgA0VDn
Nl+vRXKzg6wrUqaZ2dDQ8FUrmd9RCSb6I21+tHT8d1yfjravo7VHMyarx6S3mbW4
CTXN14QehCR362Ujj0J/lw0IEFsNYVgDUC4jAldQbebXB/UftlUjNt/fxv4oPQXS
oIGipBRj2YPvDoTDWBDICorWY8/s1OGpWoxyT1yOhBnAnRPunFHNL+KDO35nGu7w
a4n2rnXDfQTRJVVUIW2a6LbuZTIuS4P2N/YIcNnaicaXw7g2ZlDtL+ptAzXUKjbF
8OKYcbvecasDZH8vVHBkuLDhLSqiGymsUlfBmdSIFP1INyCqCQb8VzEOMt1ga0QJ
LCmPOJtpvBm+mtHa8ZCxaNl63c+Zclmb6pWW1eii0vLvUiYORvkoq4XGFV5Kc+Yd
sVdlWibDmZVu0sEuPxGkn+xOiu4nO+ah3ky46JVMZC+BteF3ZrwjfkPahX9mmnUp
yEizQSYaK2eNrxYdLa+4xIbGpDaNIKiuWw7pgfvfI5Y+zEk9aLUFv1LLrRpRC3kr
hU/+wEZMePF8xQJabmqD0dC7FTGDSBH6H51AVqiYbebqlxTocdhvtGZsNrBxRMNW
VtRAWQhz/nsBM/ryYfB4XDds0H6IC1h19HspP6/WNzc67QtwE7MwzUeOUBuSwnY2
Pc2tk35JwMOjR6uHdh1iKvTIukQP3lJEvaM4LC38vATO9bh5+KdKZ5FtZfo/haCo
b51EPJtOII5SMBrgF43VTHPViIRT+Oi0imqBF4JshjFeLRV8Hjxin6XpN5T2QN3A
rco+BL3lAkJfpKga3tBWOnmoZgrMDWZoeuD3LvpSY9XPf9IdihNBU5Z0eTV5taPL
qKTTmc0TR4hE22x2PWVjIvy70Fc4OoWdD7Ne99o+t2oxa8DNnixqLMOi0087/k2E
xFLTpBxttwLpbKzbIk7KceJsJyPIfK0z0xnqwuQjABjqPTW9paC+zGayADxpP9Y6
LY6Ms2uZk3PsB+XbauyZ7DqMLnUgWkbMkGejRZFGCPB/I+OXBCkvYBbrZ3t9WDxy
Q+CWpNhLEVWMGnmi6y5Omi0WJZE4kOI+Sm2LjUwlAWJw8X2Zjoyn0Iw+klLUH5dn
gHoFNvTAfWsDxxHBEulXhSUxgjji5sRCZgApZ3ZgZJpEPGe5j6vfbA8DJEV85SFA
YLJsuFzu/v0Tp0VNGwdSbwEmdwjlPtSfgz4ptGLkDBV7yjFmPS8Kyo5znEyNFbQh
VLjR5UHH8RehF6evcwCcwsUZhN/YuLioUO3ZLKXDqj3OoP+7Plml9JKfPbLvbS5Y
u0tkiQ6fz1qQu0JZlg8mv5KFWt7D5tAtbTxlfXLRC+gDFxH2OF1KhaykFkfPV0sv
UKtj8GrKCHwPRuzEYdUnjypCZ+YyxAF5Eu5WL4y8d67dchUM8ZMbI4463ntWE790
fDvJheJTXSYW4TwRrEf3dblHiq0vbOy0Q4l9j6F52E7kVdzvbx0OhPq+TXGrgnXz
j8fTqUYhEn281eb/L8aN7mvZNV2+/qjtIa7nWY3Rrzf8dlBlg2DcrYnMOjOgfATg
TH012ejdYwypVijYEQjdr+/9tx4NqizEypTZL1yGEC8dcFYA6AADvJv0zFATZGEi
JM2OPrjUa5MXHeI4SKT1Hf3EN8cbO6P/aIqxfWFHA20ttSJDQ8UrVqTvZR2fo+Im
E8mZ8Urk2WABjbEjo8isId93r96Cv3PEesGjWyGTOWGWFADIbsZTp1DzAobfTEHX
fX8hWyOuQOgiS15a8ioBOv//ESt7pYc2NyZp3wVhivSpcb/ZIBz6yL5iVvDiSkLW
+WPmV+Wrt1aqliJPDeWNpREmFaZ+cSrzLJzps26zgE8SrKFeFdFft544IZZcKaqw
RCcQ8jVDWMN5/uSMzBW8Gn2lbEplwhKT2JhxN2ZkRCTwMkU+OUdMh7pio3lbd9OJ
WxPA5qro4sePQQ5TqDlnXfByUzyaJIJB4I1zeMjTyHGA/KM1AdKEsSC/vp4BQtYJ
uAB0az7FZVUm/Tc/Gc/VvxQaE9R3rskIgCl9at4355NNkmDW/CETFFIHuFwz/i9g
YrHtKjfoZKI6uMVl8/94stREZOmCqwnMDtv0Jeyq7xd8lPtegNz3uAa7xXkE0IfT
6IFSrxEOazJZg6VZZXLCrfsIF+4RhRABXk8yVV+Z2A207hw+yCMb+d3ta0MpaujX
45T3A9+B8kKrbTlFFs28IUzXTFTl3VSsBgaPq9uzurFoLp+HlkGezOUK52E/r3Hd
0ILojpiYwLeqovrrb0KZcbozNSDRoqOQXsFXltqOfh4JQlOBxWZMFlrxFaCqb2Bt
3Dz+GaPK/hU6F2RWNwLuJik6apwp8R9mf5JIutmcEcu+11PwNquYbX7rPa/jhvfg
G5EStZeRw9EuK4fozCRzmwnz3mIYW7Hz6CNnw0sGsiJiYxRBfPPiUJuYSLEpsJD+
XhR3bkQegXVqhjtnH5hL821Fj8np/MXH5dUlat9ajNO9hC3eBTs1etc22xxeXPz/
5njBlmYwwPP6NGTdhmXrj0lmuItLLweSlF5Mg/nnWBPbkq6SYL9TM8tFgDRgAeV7
AddHXyQrm04lHekD4Wr38nqZGmL9PQj4w641EU8wOrqFv9iVltC2+DCNipwqnmHn
n+LU/eCK0j4C3Ykd1z08xFSr0Sp/MEhqPjLsbtXO7lThzTmgSG2fZ59g16D6HsIf
zbstOEFdK12uWJrY/t3sbSoefMlbooqNslXFVF2HJph59xgyGrqt+uKSe8PCjJz2
+VilKeRXoC1AxBddoO6RdCnm4tf4UQ58qsYR11bggpYsaVp7bx/aDBFusRrCe9su
0hfsdda6LixIRvcs/lng1yncMz3RgSaGuDEmLJ+x37SXiBhh4mC1gREws255GjEs
qvj467H/S4yR6cmUfBsOIaa8nPklRMN0p6SJGLGzK9BmyxPWE1TW1BZiWlLPzX9F
7NI1ljGgtErQWSZWxYghMSFIt28TnAYvOIj7hJ5rIgjOycMXY4HnH7C3AqV1nqm2
vZHDS/jpax55jOCde/5JH3UhE9h7GTVqqylN2xW16/wXFSCn+sF4aGrHReHVm2Ty
8jCUYIXBGXoi+P9+MUuIsCuw9cpegyg9HU6fzG8iauUQs6JfpHYRK7g29Qjg2FnU
HQg4Ni2vfAYeEHb3e8l3GTJj9yOibtd1uD1xWyyxxFwZggRKESjtJcF79UPVTN8a
5u6CD3fKgycbWpsgqcIRpefz8jxN/48MlWtJgqDO17elA9kz84K2Nj54VVAY7gh0
2aNVDBI6AI+iopdRc9IEGqAwQDUkuSGK4gcR485FEJvTQJIJEgG2dN1GE0WBEF8B
sh/ZTipuVxEe7u80Wj122bD1+b0t7d6T3eAOYzM0zudiQxk94R1y3gPRTRIqJR7L
TRi8jHKUxAn/6OqY60YIYjTopDn/VyMIO9DKRK+Q3MLP6/DpcCCv5yxvGTIx1uPt
q/X+7E37iuDgHmtXpnfhwBvwfa7paFc9fwq7gAIgrgYs310kAB1blboCcMZYvzq8
mGXiYEfOk00i00Gg9GthzFQcLAz6XxuwbyBi8msEh0lLeW1gSRrK20CianqPVfnG
8o2uLtANeWty8hKUHLCwyS4Tm70o3DJjKwj6U0o8N+O6rxO2l+aoy2gcjM3IS3K0
uFgnT6XFyoXatWNwe4wbnK1FYcVHbYWs+xE8ONRw7tNvZxUhZuTZQp1v3cDiOqWw
9xEhtB5ZNNKiAuCM2MTyO5UsKZuNW/m2e3V6nROHd0VSoftBqopgs8xWJzuthKVE
pI0Z3CN3EmybDOaHVXaWIcX5HFtSzYVa64A9P502281i3j7bqcdxQm6ebo3MnFE0
jECwze82eALp1SpdptkEebW99e0DN6NbeBdmpPjUwUoyQCgPCQf0R56hSgePYbfJ
HyoIjkh5GFU1njNKgd2hlZhrAG0vLHEj2ypx7eBYdF1LrV9G3I9FOvaHMsR2CZpV
9froISreDc/Sep8aj2ckBuJePFr+JU8kKx0inI3xzSVFfirMXwF6ZaTEHshRX/EG
n5NhRjsiWymIITzcTVmZpZbRcbr/A78aEV+ZdyCx/JJko4OgvcXWnaMpM5Widtw2
5zxf9GJVlXcDtHNjIVon+TiYTQgE1YFrMoM3Wi9vQSW7IqCof0RTycoFZkCePIla
JA6kINyKaSRqzBnCYkW9kUzw6TYhaNhItzX3ZJ86IPoMzavqAd7D7CGEPu3B/bOY
PuDmSWZn8C5UdfT5pvOShrcOLNvbP/CktrQp3388w7NrRfz4Fl0LehTO/Uthzocp
5t49i8qFztgwfcanEgvexsXZwJQ+vv2KwNcRISa7nq4T2rnqotwq3QqpStvpBONX
G2B7fz+28hTOcylAmEddKcDgBoxX9L3FludSUDleSKk9A6RZyKaR3FmIIMJQHTkk
J5kPXibLqdlteegAEqR5Oncz08bNr3LQbyL139jhsTrITCTHIIRDsmNLWPW21dee
NFiHP0sOIKhHtfd+MU29YFGeAAajI52Iiw/rpXMDkYzpehmT/onsQ5APNyqCOvNV
ai0llAbZ7NeyKmqLXqmnXvdnjzWSwOYr4LNxFo05Ib5jfFOTzy5wxwyQELg1gDCX
p4gT5PDiOFgpE5EH1qoTU1VghsZBOyPQ48W4a0rLAIzj+m8T8plrjWjghcYD/Wz8
yg2EU1PcWYeYW78IfinkLfb54cFd4ln9jxUOuskolMptBxPJvin4tbfkkOJJORKL
xF2U2m6/P0KP8wTvsEsKb4zlVUsotgsUBZtYo4Sk438yFwjaMmwwD9tOuloqQ8jb
hkCEWKAeG02D8rC2FIhoQlrP/WWp1ZVrPSYOQJQas+ik8MQbHc58eHoZ4znjHwpW
exgqDi/KtumXzJpm8c8CZAD5WstOiBDOYetGatBOg4butawSHLaiiWRNjdCcLQ9h
3P46P6UfVm6bZjpQ67kp+xS+iCoUgHBR7nuatV39XRDOL6TSMdbqrGU/fLpJQ1KP
CizJV5WxWZ8qTsC6pVYhp/GrUBjU/MDJ6rtaRfyCsQmZDPei0pyIXpchB2HfCr1l
+mt8oLkg8KsXLEMiyROTyMdtJ5Ni8qBKxez56qLJ5yzY7DTh6X4QbP0f0t2dKh+U
qXeYzAM4rUdHp6cYw74H713eH7Yup50efdiJvRYspXtbEeOlPuPN0Y1V7XKX0psj
PIfcnpPYfgBQdt4R3cylYkQ3+D2zYAgRs/uO8r7R6hdHRBAgQ9LQn6lOkBJ7oZXE
JgLTqnUlcAx2mpumH1lc1DOpZuotM54wPWPPD7LBJTYRS5BFMt4Fk0grWjH1Fp8a
EF4YJOqCrP3MJCp8EhlnLf3x1/ZexrOK8uhsr/Xrq3AaaFp8mVFQYIxh74Yleuu7
VlWTC+1fdUVw1FypEyYbRqoOA9hYSqZM6xlS/PRmrcDv6dngElrSRRfZOjn7A/LG
FrLr3/Lu48DI3pArTpVvKURDpYCjtSk5mIt2X7qQRs0jxEvKj+Vwcnmn+9AOrmS6
1QmLmUliM55c6Qzc+NNCms/dx9JRgZDAgAbWynINSQ+5+Uuxn/yNrOyjVq68GmBl
cEGLpTjq81pw+BBRFcewN3nXwnTMZdbhvS2G2awIsPVIJi00EhNv5KXuahR8viSS
9riTczui0ScIBaxNNgaBD1XsbMgQY2k53KVB4TefMmFznv66Fvwokp+UNqjlJALD
Tq/AdYPUqUDNJCJIlb7yQi50FESGA8UzkCMOK94pFdykkRqzk/AdZ1qIdS+/CKzT
gzmSI7SI8Tt62s/s2SchQfoNlGhQCAFFN3WCnnrez5STCh450VGdig0C8LR0IMmd
7Yczjj4ZU5M1oAHp0szdQUSWqJ3TMnijxBSt5MLi8SXRQKPtXZl9ye4FJ77SxUrr
zzTIXpKLbm/hF1vkj3ike3vXzVGc5gkQsXztauykA5AbVNDQ/+RtbfnOp9hsZisg
30S1F8Q77cVkgpw4lR259A3BRdCs55TzZTQCyL309R/iPjBZBuM41TNBC4eAhWVg
u0v230RrMDf2+CaQcAEGCJ9Z2CBeVUMC6oXrIw9qW256wGPJJ5wce1zRvQWrglfl
WzEgP2p+YgDfUZB0F0Orh93uLRR7CS870B2hGcUVyhLmEYyG5UM28wqDhYzDxKss
80mn0lfkn7R/EMc1K9ESHl3OsYyqyIQAgXpYzCdwEBoX6jKDQRtO1gma8Kp+vLlr
AT4FmIzA7g6MjLlPZs2wmuBCKUpPGarnt6jJki8LeNG/t9gLpcEjPWv4oxrB3GPN
GlX1JpSXXwinYcQG8llV5qiyHGPjR205Yi+mPDvw2BPx8UoeS/2TJfw9mqJIn+Kc
yqI2w27461LVybErt1FRpbrxAaPaDPX0qBM9OKHhhi4Smc3RGX13R+3fzRRyIxvx
oj/WM7zHvcVAZcCLAsJr9B/TQfMfmKwub2nsOS1UUCneLTHrXQp2HiKsx3oQNkEb
1yUP2buW5tqlcsISXc/NO5pn7+m9qMKDEbscBmaIURDtCa9WwHGjYOYCQWbyfdL2
+xCGcbBSubPudk0I97C4kMr6EPE3yFvLgHBh86rTb4Ewo5aynscuQjLnfirmT3ff
2CrKHLLNumDmOp1PHRCxaPbVvQgM69KjYA/zDZD+2z0iMfyzi+00LwncW1KGzFip
O9rACISIAOPcqeymGm9kxl8uzFYEWvm4kZPkqG4iGS9gvHa4QtBP2e+I6gV9CV7d
o52/cDqZsn8kPJq8hHkJyuHIMDKjZq+mnMOn1UR+IhC7k4SIckYTDfSBOh8lzF8G
lcrCY2W7DZnuJpgEtr1q4BtpjkksL3Hgf0R+eOupIJc/MTuyOkU/Y88XYXtqcxJ2
uPuz5hl1VpZAWA2bK8d1fT21gtx2NGlrLLH8lJaIzAHoLxtjSm1km1WV7YH6i7aZ
iDmbCQxETbgexPL6BKJgL7luJcV6CG+qZkOtEThzQ82yNlzvNkAvFmQVucWMuNp8
jMLTFuSUKdcGH5ydLieUaVkfCumJYPqyWrvm5EDayC0C9hhA9V9fcUovOCnBR0+G
GEyVm/LgvZIUg24yjgvQb6PBMXUSIEOHBDZLQl4KQuRw4uPCEdmiUvLGmRQl9Vln
aipnbfOfGDI9dss0xSTpCkcUllcY9VvZNhmbxHWBt6Mc+ktiaEgmal/HFlObMlH0
v3BQoVt0cfICR3MiM18PXH1ZtbjpnbJ87952e3ENwZRzicTY7kir9gNmugTgs26l
VSPphWvgzP0/lfrZAoRbdgPpH4ushZzXMGy/EWolX3Im7d7mpoaaAwFoRn4ND4Xd
LkVOuU5ABi6osnVKX3cN7oCby0bF12h4pheH6efCMtSowLUJYRkKGyTEMtZIv0Zf
Z+9erpsGgsJJ0qhiRFDBGBQMoplNmt/1UjmNudCEty1rQEqfMSddwTN3qsoZExVu
V0BddQiKXYTzBtmHgV5aNlM07KvNBVi8LoGqjwkiATDs+PTGj4yNHdCnYCf9WoNw
OZDFJhtNylkKzbmrlQqH7qisjyETABaDNCyE0oM9PpX6lAU8o5rkHNGs2MUNCx17
4e6U7RuGG9hoYdrinS+RICTEv8JqT56uoko84FSaPCLU4YvgcF6Kg1y9pTIAdPQs
12UwD3Rzc/hw+SUTURO2qcDD1kctKngww2NPb6WFbUa4XaLWYEmx6GF9EvWeovPu
uC3FqTU+1E3wFIzinNvH99Iqt30/+Wlxes3wPBcyAyiThxdnLroVgqZM2jL34JWy
/jfOQBoqAxckC4JzgP0Fp9h7eFguDadX6N/31E9/sgY8rRaWlF+X4AJLsXOdOXVJ
UY/H5MZbyPEo3Y1fTSnQ2PzWUsb9Of8hYnLeVXsWg7FzJHLR0XjCle0bMDhrkMn3
Cwn4yAT6RUSTXJsoc1dr/0b+Rp3z5uVjxokCWH5QAFHxCkC3DzquB5T2o6+Rahbk
+RVgqqJqK1dmwv/Yk870oZ/NFt950GcqBDoHt++hlllYtl0r08r38O6IbbTFwY8N
okB2Fifrz/uDrwhK1p5h+Kivc4UvSjWStIIPhIz1rrC7fd2TToSPIrLbcrNZH3B5
XNIXaN5qUkD37/bL/t/uNmuN6fWumhw+ZxglEqKzJhwnVJ1CPbGGo2wXM+L2yk6q
X8B0Kyu9aTCblgPNw8vjLEb95V2xjbnVKG4g5sp56FVhyAoVX2isnLGqorn3nQht
xoXCR8KFKRXMVjml1XdM4f+Lpj9jK47cA3J/FIHo+eBdI1H/e9XMiENeBpAg0e65
fTKOr7LcBLvzq1LeA0IQTUsFrJYXCyTYV+TsrpQLxxZXbKLm9j0kJihVrdqDzqX6
QHRXKzeZA4Fk/Nn56kJ3O1pwJ+esDtzAmHpKREBEkqQiursrwlNeXnMXxzbYNVd6
4hzHzSp8sQoecZpU4E1sRsgjkAE9voWldFYJkySpZAOeoqeTwRwnCkNhIWLK4i8t
ElkVgNm3ME5x46iePmpV/KMURRkYJsFPUJcsXrNK18HlqW8m6Cj0bHBOveGKSGQd
dZzJb3jYAdMUj0uwnZ5UjQQKwrv4KiAXTYxioetriL8NMZZmpWLkVd46MOc1UVP/
4OLx+PMfVwNbUWiYGM9cD5trYzWhPnvqGHV4O+etMG8HmMoaAFoGXj/KHEpXQfl+
v51vLfAjJ5BhoVD+H2h7ZtoxpPqAne6ikxf1EX+aPuVhmQ9HU6sCCNt68pC1oVY2
uoN8FBOnQT/SUZ/j96r+NRlLxv8LqWsSE2Agvf+GpG3DNyE95/Vtu4Rsc6oP26RN
7t0bFZ4qHCRpokR/fnH+E3w0ply/3CWc2OrrbN2DHGp3CKgXbW3bNAybRUjTWprQ
Lo4+A/Js4YQHkGn139iv9EGONokjVNorJtJN1sxq9BmgF4tKPrwCD1+X2i3ScdJH
cw1jNGg9AbEFYdYsOXgQkErc7EYMYF7MG3hKniEo4Ah7tdZe7M48ohUYS/us1JKJ
oZ/q687ntBbMxGO8feZ5ZA4lJRM5EstI+Rjp2iJ1egfoUsL+N629Mi4zeJCvPsvA
mpa128OuIpu8wdOIHBsQYga+p6CGaLFVFX3vkITlSLuXcnLLGsGCAVoxd1lmpvtG
0Qh+HcIehvkBkKpqdh8rBy+WBYsFxZjwVN5RcPQnoSzwK0odOP7VJ8N+E6tboR4T
zk6IFoyIJfRoeGGoo4WWqmmpnNiYDdMqgibM2iqvkvCRqJcWdJ1kKrGXr7ixxYtc
tp7OJu5qXKfKoos7mUDUxwG5xJ201AUE7m+1d3QM4AEg9qFFImgCpKs9eOuWZxJ5
wJ9KXxU1RTBHeC8mtfZ2YhUxINQuOtOAF99yZXUIEj1RtfY46omhty2iAtNc4JXk
3+39PktxIfwK/iBqdjxzChRIMjXzxjsZLEDVkTXwpxIEtdzPg96Avc5i7m66pdqK
BnRnSTNYjOSAItIq8xCgwQalZnHpzbPxBNY74ZwHrt6ytxWYOe1XV+TcJzUV1zoA
5/U1CnD4uW66ZSCywL4bQBfnj85bW68mQKHhKEg2fs07gSb4/2N0JDpTq/+C2qYY
nbhxyZ2c/qZIhMUZ8UOJaa08mB1Nitbt6NWKFcgGrEIRaJ29WzVJ+6udvIVI9ahf
CaOL39aucc5KIBoflPe5LtWIxtK096MGHr0PRZcawnvm4GCwiMX80ft0yR4hcFVS
3RBtcjZQAA/o5YT3miHFgPFS+sAveXRtkpxF6VAF6Rp1w8x4XN8IXGRRSn397A0Y
kdHdpcTpAbAYgHLOBxh3W8vnRv+Ei45SLwad63vFD7HJHQSn1JqU4L7nGgXoH8bX
RFvWCnSOn44cI4nsVVlpj3u7TrugbWlGKx8IX77MqCQ+/EdiYPZNegvPj6lrGPRM
1UCw0NEjRtNtwLe5M2pSK1KP6SHOx+HgJNx0VvmXXsVQw5PXtKGU8C97XvgdyvKZ
4Tn1tEihe92YBukIkpZEoiu1fc7r5XujacZS+CBJLp3KixV0OoupXIQxNyESGtEp
HE1O/pVzUO8vA3XqCOb3r2gi0yLD2t/kP/BzuCeR22f89ZnTzYJi6iHgyVB2URwI
SzMtM+562ROZtfjLc729cUiaevmE0Il7goSzavaiT6SetDRJyMdAreBuUycuOflL
5luLAWjQKP2ozDSh91gwlYrFmCShaW/G7FWmeoGfur8TJBqxARV0YkHUJ+L08dkw
JXdUb4nf8O+/NkBG3s64gqdXGOaoUFydR2l/bplWHsZZ21mkIzovwmMlfm8hVrql
vcSQS33jrCS0aNUS3ymyqykM+3IgGN9/jj93JiknHSWYL/OI69MsaaCxqXeH+Oz7
0yMXZyrZI5klm4MDTVDl2UHgG26XDzWzDvqX69FGgCbNvh64maqtsEls0VRWs83I
Ii0gxojYnL3v6k2Ac3GHC15makV08fkA76nisHetkHGkJzj3ArmiX/TY+gRMFmZE
ThCViYgBLgX4jh2hXrN2eIyNIsLL4SRjH8Ym1m+KN4jPBmHSTHPMR2GV99IiQrEJ
iaiPMWVG3OvkVziL+Dx77aE2wTka0O13FAkn+yA0Fra2pN3rA9ULfLpbgDw+Gy99
amhRjDtBLqWRRN7gMbqzalxPtwJtpndgcezQXORQjTfdP8L95o2u/NcUOs/ugXgt
+XgEUGfdOBPmbgu4wUPtNdwJs4U/v0h/RvdxC5TbUEUq2xEX+VKggNb6hEW2AqMJ
dmAd72cj7yX9tA1R5CDj6u99N+qQ+F7rLdxIC5DGbLZKV4Bte/UIvsluR7Ua0Jvp
+/74qKKNGAhV+rr8tzr/rJ8pHBASHEIJ0GGmX+HpD4R4ce+xsIDhqGx2C38gjueh
BO31sUbQyAgqqGn3IwE05UTTS1bdOeHsYgDuKIhO+PsEnbBYKGWSFmOE3AmCeOEJ
JXvqlawvTFmqzWD8ntE41XgPNMurnh9ZVSc5nd2N2f4QEkHSKAa0cQg499zBuDw4
4Cjw1tZDUuKVxvn+qsr0a2T8cDtCeedBGPii2/gBUN8ozLmCrwps2uSK27gzxeS9
HzdF9cM0kfgyzuHoIqaH6MVo1fipifARmdz7FGzqxR6bcekHkJO/+Ms1YXlTyFx+
J0I7UC+2TF++lFaO7soubf8YhV2QKDMemKVOCCgTEveamd98E5bkyzkIgx67Tlx9
wWSQc7Caacy0LF5IAmNgfNNIGCotnB9SA76KPNNBh4skCRUGgk9Uwe2xjkTIgd4w
+jJbrsq71PDQtmDY+WJzKjOf3xeE5lON+cbWZXs9/iXcf1mRizaYPPR0jnK9vL+7
C6nNtbkXavExYogt11qtqSNq6mwv69lrhdox1GyEPAJFvpDuDJtbSJFEyMDqDgx7
HNgnaDNDk0smhDwJnnZuQoBtBJJ8khlgkF7n+6xJ2BG1DxiyTnBIb3LZuCrP6HsY
gSbn0o8mbnBbgqrHny655vFPAlVMDrPSbPyVpih7sYvwalQh+z8lcyLwGqwWW3c9
hbvwa7BfURa1gEZ9HWsR52MSd6tzfVE68+VllnExihTa4G9vVxWfzqh66qMkrPYz
tsy55UvL3u1BWdwfKCUD3Gc5DM9ekovGlgK6Ihzs4qWt94yrc+0RR64BS3uXP0+Z
zW41cVgD2f0DMYBQ3gXloe7RpakerfycvhPcsxwAX/1IieSu8jZiw7U3es+42jO+
0Cg6x3WK843JvbLDweYe48IRq1LkgPxiZgLFm2X8V+wg1pFCOPdpcRG/+aD9yxwx
8TRDt99Y1bk31IA/f09mnedV7Ty8LlbWXBkfNAya5JnsyejBA6draNoEilsjjpX9
sRwd6/Crmn46stisHtvt9EvTM9xANEGRyK5SxvLgaybeL9ra9aXUWTbIXohhyPkP
Jtqs8J2bgF9eir7DT2FdMRowZR2yHARlHNazRDxPZKpx5yiah+kjhbIK//Q3a8bb
Oewuf6c8kyq/9raZuYgjFVKER+p2TUYMYtc4Fy7QVpQEAhTHv2ozpbmPwss1Ikwn
OpiLCptJs+klPLwdXq4+Si6NGWP4UvDrsXpVCld6+P19a1bSg8aBsLhJ3z5pO6bG
vsSj8bMZmPhtDfruxLe/KIZyPMLnfCtuYhN8tQDKSVcEHhTYcE2QGswbTNTdF1Ks
DSQ9iJSA3a0/aAR+rXuaHEU3b+L8xfJPqkMicDi9bhcDnfsCoOofNUwrf3H9UWXE
3Fd6oHNFcXUfbqCaPEP+YItMFTg3GHFXynEvhQYEqKezXrcq/O3N4F8+C+1doUJD
sJXjqRJyReycVkkEI2vtLUv8XR0a+YtkREQH1tMByXGn9TYt8hA3+N8SgDt4kc+I
c2bikmAnUqok26mcumsEnIzh71LsVVA5UhIFMuefdNJntfokB3rG57JchFrnhlK7
IkZo7CRkKTRYfsdJGMIhCa/pM83uFZ9jsC+ocxMDKHKFNYSOcu+H3WAAlAH6m6j+
1DsfAPInhCZ1FJuJcKnfv0ls9qLfuwGjHhQSeMYjbnzM8GglyL0flfbr8DRQRJo4
DSD189QnvXdCul8tq3NJwHyanAkNfEcp372soL4A4vr1aykNfWAwk6JgoRRPCoXq
QCsCkTpmtkk31Ip7s38gZrKnrVas862xE/zG4T7QpkafGYhS+Cn/GGSlN9mDla5Q
kGrc6jPfsAbm1n4eUIRUfu/5PWpmRPBp5bOWaGtivis10e/xYK3/d8rvyCk60P14
WH2m4HNdi0ccPWG6AQ8woRVY1cZHQPEBtdWB6kmc0HDIQBEyjcXw4VT+vfLkbFZt
Kp5r2emB5gWNWqFuQzV2tof9inKU2sjj3MdRNEWjN1o691AhlLczcrRCXTm5as9T
DQ1TZmtFSZqKq2zVwOmTV18XZjCOYqdRJiWVmG4iDZVU/iAD2vqpoQ3Se19XIUIz
Lofyhfjaz+zG1hICLEK/zbO4CSuliNsL9Yo24SlLPlZ30Ru0gGwq74hDq0oBxmL/
ufK+4Dis2qsS6DR62YOF6L+yVg284in1EQzULyXKHjxooWIfOboz4dqpYK0KbK6i
ZnY9kxV+O1p1sy0/WEX1uq8C/0p3cZAq+rK3yrkcXOB+o3cGW2ZM6aaonKAmLdtZ
I5g8nrjvHGuCXhg0B1r6ebgfoxTvW6M/D6XshRRPr2qXKzsXHu9k/eMe1UplmzKN
jYUcHFnGxQjj1PwfLdy/ZQDYScsVlbgIl9/ZmDQe3KjDEdRbTdpRRFv+CWo9++3I
LN+WkiWZ5jVX/m2bjuAYEV/qX8fVf28+WAXpnkz0mUy3P/1XIr3SoS/1SIQ+T6Vy
IQPn/KNPGH3q1xr0iMmFvYOgNvGomYdWFLk1dxSmmabiPhS7LMtC/rqH+7Xd1Gnz
swYClas39lFqOenLGX0IEuT9cxtijnR0l9aETkgw7TYuogC6feEsA4KFl1KXIkG6
1X9B/rXgLuEvRClblfbDVzme7kZ0MsQ0SYHCJ4Ltc0/ZHkFXLs2Mmg0pN50f4c1Y
EAfr5Q99MIzT6Yt4YSV6EAr3C6GMOXz+nXUuJweFyPHvZsYof7r0rRlsE+qdOkxN
Kpq0g70N4vI4Y1cT8RM6s5NQmHfqSj0lAOfZb8rgbsKkIdzN1GoIDSEw1+HHgbUs
fBNJDW+gMj0j9hVyEIJa1g5ZGajyVSe2Oh6x/1wHGTe0mB/sDlcTz4rP2R0QdIlS
M8IsbYnzZs35im11rXhnLM87HCDbeguZpwRb2jHoD15jkPm5usICHc/lkq2OcbEt
k4T7h5o13dx9PDMNysaOMtJ+/KETKLVIsmf8zJWn+RQU7VtL/5fpjG1SNqGPIJSl
sEiwqD6AcfSGKYgIcQAMi3Tjr7SWkVxjzrO63vNPJ+HCr573h/kZE0h5JLNhDhOf
j4QgBksZtwx4cbjFRRmRgEYdDPLxw0K3/4EVLujPl8E4g6AtLVnBPYIA5JMt1e0q
YsF6PbrwXArOL/shSmFydk/liY93WkxugFDscvMD5gCHMa28DjdEnWS0dNEFy6TX
E5ftZ6fzQcu1O+6K4dvW7ga//vjHRfNZ7NQUKwgG3hQyBi93mkpfJ74EVnWReKh6
xUetWMQcoV9ok3MMOK3WS0A8WgHtgUeFnxPcuYAfG/MREsO/b46qmIFH6A1INsj9
000n6bGaiwRk30bPwGy9bxeV1nXdEsX43PbL1oLiSDU9nEWZx14hF4ivDyiZTsVc
6dDBt4z6RJ6dSP1EIgDs6BmLELXTuUwLAsS67D8zBmxWXHNOZadOm677VbY8lK9K
V6isuMMA0062vMBBRW6bqJB3OdZCVv0HC9aPF9hHxhwJJXsG6D1yU2A7CnyTRMaA
TAen/SIVUr0P6CIpPsvK8zQ7fa+IZVYid/+H/a6hIadTOwp3AW4lqXR0PhDW+ty6
OByd5duEZ84QXWs+/wnPnWpEOHYEvw8B8WyL8tSPlVNV1bXi7KsjSq3VT5WrYHlS
F4ygfoZvjFa0pd6T3lDRtGDhpAw9VmG9qbRjXg8MdGt6ZNxAPJPtX0OC0l/mmDYB
cBNf0fK4EBxucVY/zvqlxXUExqqzTnCKoh43gQVf3mJb3niYOiX1Z7uzl9JDlxqZ
ZGYijwMJXGwVdd7vgPrE0dYLwzn7F6XTOAsLoQ/ElSUU/+VNs/2Td2GzHMiIwqHP
7tPDjtVi/WBTWRLx2rroq0NkfVHxuv7QSlDbGiNjcy6F1Pt289NWMYvb5WAAzIGe
47GBGId9fC0Q178yV54ahc5+9JjgDdX7FMBq7HLrIrOD2jJjPq1u/ZY7hghroTMs
E1ZY+my2U+Hi3bcK6ey3tZdy5GInhy8OLYKkrZUhFvA+10xqE2kAMd866U2zomrV
UQQng5TKR9p3DqSfzcW4sfI/WxY0/9rLUroBlffms6seLJEFI7HkHHnQMMOpGiUL
CuBK+JZo7arP6TvcCa35GcgHdmHRWpHRlpWB6BBYxQRLxim/FmZfu1S1nQUJ9rSJ
RhKYd1GZyksfE823YuEnmjgGDFwMknxVWk6WIO7jQ+aK8RKATiZPvY/LM6NXWiF3
gZSdnWrSkJOu/cm0EP1x6ZJ+5t73UKmGGMzHN8c/ij9Tl2BHvi0HRgvnqVUnm+Sm
bzJT5K3zQ8S9GNbgY27A+EFFZKhnWCPNUVln+UhvxQpMJoEXvMQCtBlKk7Oe3HRz
N6H/G/+hi7xmzZxpS+i08Zp02s2SLY7qAS0FTU5wO3VOhtCUBFhVMZWxXyHaUcod
jqyTOa1GiF0LMBw1cVSl54uM/myb9hcaca4Z7nfPmeLDiAodcgv/IZYQD4YHNphf
A1bLUV+eZWy1W8CGx2FdVuwQbqaA6tesNg/VsoIGuP9/pH7X/V95ah5GqJK7j6/B
ikvcEw/+SM/dIUykiFHOcTdZByi9RCEkF+n8HClmDVT6RdO82VzeVyZvxwn2FfrK
Nz5PaHCzpJ6QdZvixszPZgr7OgLmT61mDFL3WBadD3cs/1hqWzvKRQ9h2bY1wCKl
pjDsCRvO4Xdxplm7IQFJHJ9DcZtpq1CoXuAO/BiG4eBBWQF1AUTSIEWFdORvM/u7
RBvi6XcK0TGQrVhL8YxTSCDk7bQNMSf+d+HovLmQpstjznA+I5L0bMBeY9Z8/wSW
VMkV3sPA4Frokqffn5lTyrkQXCmziiXgvUcdwbcO6mdwTkEi4zvHO+Di2dyZJZ73
u+cp6BLh+DVbjEczhK5Wsy4tk5TBPTFjlZVv9S1cGZcxCIXpiW+Q3aVdh529UN79
zHHE04gP33mjJQLs2GjprmAQ7KYGsWSJvhn1qKWwALuwWst6LOWusEZ2dG6laX+B
80IvGo2hlkwCErPXWqFTJAgJ3sG5Ib+vQNKjj7GurDdz086l+CK1TImmtM2P0Jvb
oPcs9aPY/umC1cvkjuCpLzINhlcA35m3c4AbtIu6ZMd8dAG+fgp4t54/UZDlOjge
jl5cnY2D9+t2uGGCYit0/9lJmmk0GV6I8YLcJPlDQ7wonP+TvNST0pTXYCbY8sm1
QGUt3m9i84/9PKdMM6CTHpSHsvyXSmZNK6p7wsxx18ooVfdj2wktfk6d3yzE6rxu
555Ttz4y2C5y3uWEIgUH/OsOLrUiCXgUAsbvYgUxPKUhmf20oRCFKJznxBHyzRVf
J+2bavSnBb3pK7n7WLo/6X75SF9+iZC6oN8S/CkPAsQokRhCWrCXojmu6GH0SgZz
vWB9o7h9hJREEylo5OlXaVyTvYz+2Z0UX4w1tNXLWlrLYi84VBpw7i8UOBfLCkDw
LemYbUtspw0fDM/QNLJqLrQKdNcI7bzXn5lN5gi2qk3wyANITFcH32QzeJ+BkQCe
HBQE8fV6l9jIeREnDmICra8Pz7tSHPYJbioGvxDQLVXTvyu7A0BIEj7efeRvHICf
EbO/rZaZYqDL/Bu8cUCNucNAeLRRagbnT2pOP8IQ1fLSxxhX2Xpib6JVYcCxU1JX
VLHJ/CyGdHM6Pcp71OR5oCvoi+SqbHHogc/lW5NJbYTqWGIoO0/O1cokaiV0E73P
NFGKl/PmhdBBC/AR4JJBhYQKnpL0OeO+3WPFNTyKf+olemG7ty/uCWsFARO3fkMd
r3FW+HOcV2ROch25bYscwWt0w/AtfJ0XSMz8z2vgY1dLKwuYm0iohdPdEt0bAnVL
yuHFSqppLDxmHfjC9P32NtK/zSGCIIy+UZLkGgf7a8nMlcMcte6IoNQW27ay1vhW
bna4pX3jHNCW/EhDm1FTKUHd8BKbRMs8hkoMlUhntclNcjqgtwQ1ncS3T1XEkQnD
8rRYdDCSazC9PVUH9yQHV+isXQ1lic8XXNSzwTTPYPtWAelk9mY/QWF3NLpR8VNH
bnaj5EsR++B/+7b0RsGDJ1V6eS/+ChCXNI/YaU0FWpsEGGAthVZHsMP/akgLKfvA
EoClt/ydkK2xAoHFsPZk8S11KRITXH8+n/d+5keSH9z3kmFetYWpqh5Q6FRc3Fhy
scbgdtowy8yM9Y5FDTagPMeSa9Stfbwf0X7BD9hqoswPcyQpEy9RCSJTjI91AdDe
ZhMqbWRj88wNpOSsQUz8dihDGSRywiHxjr/PtVYXL+77ozKUPt7KCS89gaDZkQLv
BA7tuzTWey+zFqgfwny5YheTNZXhRZBGp/zz2vy+WUdjxvDtAwRlmLMq7dYv1l4B
cThTbo71D9kg8FaRCCrYV/6iNsuLNxjkY8/xGhlZc2HUrk8uX5n9TKLeSXN7vpFv
dvOlB22bR2KnyLGk5/QSwqwuoNCmAafocfs5dVmhUH07wp9Di8RntEu+aa2z04qb
ecaY7EUCrL0jmqDTOZF3QofkwaVGC3+D/MISW2blZceQuNiSe3ueM2KHrEKAk9Ap
El9MFutu52DypQ+pORwcFdRPpAfDngamDGmE3fvSzUsi3Q+JB/R0aCHn4W/NVHTW
jDDMuEBIPcslui7eDmMHRf6yLodR5UOfoxKJosNZH5dfMH6YUtf9BaJr89yJifja
4IGJxppTe8eKy7Q7ui1nV2SlO3eDHtck/ZGY8ZXWf4Ravue99yPLd4PovhMU0oas
hhPf6XIQNYK5oDJTmeyqJO6m8qQxfH7PrOmOSbQba14CZIjlgFRIANce53YXd+us
3trNiI8Hsj1snEawlnedCp2gKm4EYmpTWbrXZdptr5m2HpZ+61EY33Zo/6u/lcxZ
6QRQJalbGa+hOHmORThGPaTMRcZQzLbxd6K7zQCIb1JxixGpN7jiNVyd88tP/ULq
iaTViFW/7ZC1pHlxNwh274vCYyWW5IKc1vNfftOEjVUm17ramif7f/+7NQ5kdPGC
3LCs1RwXLeZ4O9PMBdVEoWM/sYNQ5lV2ZMHs3yrTzKyHIynG/Aem2QLOdcgd5QSN
rwcB7+WG6xNVEKp895U50/HlviUYqFQk+IuRNkqJETL05p1VxhucuCHgeUrtKFna
960N5fPTgo/HP2b4QNzqAS5dJ+NWigPkHPOq6+vvJBC75y3c4V2d0+XL+4Df6w2d
j/+JsHXCp6uS4dF+bhJGWiiThiyurVCWPenswt0GTjnwAfKfVjXYatqtezMkO1JV
Zlx3hbVmxVxlyoHuYQ1l76G/Nj1NfQsAPW2Bx0vrAvb3ysj/9NkrFzfWiKfgPcWN
CZmMANSdshROCu+6FnAdBQgmyH8lxqy+8HrUPQiPJbGSzEQtrluDuru5cRAf5Ehd
pKxRsrtjCH8lj3oN3+x7crTfexuOwX6pIJotoOrDef71P5P5zGFKs5OsTJViEf/p
WAk4/NntqG+hhRfn0c++YTkX9J4TonmxDSBWmU5dtYr0wgI7d75rO3/zfbduz2MH
V3ilVYmWoXWswSyZYyQB/qq0X1/drp34Dz9JKt/6VtX3Se6ZrC6cQrJ2tyJZMjvZ
jEISxolz9cQtKE/jF5IolYABJReQF2jWGKo5b02ouH8MFTDCl/wU7VXgI/Bm0/ii
rQx9Qee5p/T64q+romcvOab3jbdrjcZ6lzSF7TslcrxleE7MUH9ffQe+5y0QmwQU
jTvAJqXLV7s0Ndnm3HZJNPWpiBWbA58rbWmHysCO3H3Ob28AVzSnLnL7FW0WPCUi
jbbV3nlqspVc0HqUq14Wf5wmJ4QXUBNCcGFizXghFTqq6EaSPucA0qTkvAgnSipO
XfzytlV+yNPHRLaMvTcdIeEcWA+aDlY4w5eNpfJgGeuFqhK/4mu2HgRf5+JOPirF
pMmHUxn14a4NQIDqnwhtDS+BUqcd3nER9bhYPNMmnkdP/2Nyj0sE3m8Tpa/ZoVsl
fJfhSrQc1sVlV2eVzA2HgT3YWGylFqlKqOeA8jlk/Bb92J46cjhO2LKXYd3FsDUF
voS+DTIP0IaiY1TuwsQ/w+2YUNHlIxnmeeBBF3Zg3KZRu4uykU/3ax6VHHs7FgGq
ud3RNLfE3T7pCHmgYTgSbjKjSvWa2Gc6nWUEKsJefmLB3zE8ZEetj5qscBF1HdZh
j5y6kE9yMdCDn9j31/yzhRGc5N7zEPmUcujIDm7vWMavVdkW8nXVA2JC0f9Dy4Zc
2wMz7dNF+9oqksVUf0kgczAf3zYp8WmqlTVKmSEuQs0H/6YjcoL9PNou+H01lbsp
zMxtHamTy1nxfGPkTMhtMZ3It4uGnWDEQGH6X9EDTXSkEbCuj2m09PkHrRE5ND2k
zmlUFpeUWVULATN9dbsymuKH+Kl8IMgkXbuDL/CakpivRvY5lP/iZtWW+7Vz+Ymk
+rCalTDnMQyjIOzsIjrj/XGjrxZXjGqK5trkE7G/GPoXTisNXoL2tWBLMTKFzrlb
apC/c/lTjnbB5oJJ5J5kGcDkPadNi0FxORieDQnNngi1/xuTbc81VTuIcsZxaxH/
LTHUsTHp1QjDJHc4r4m63PNuxmK5wJCW+IRTBJ/0qg0EUQv+lUlJ1VhyC0HfH3OM
BDSwKAEJU6LoUkyfmqgAitw+JsyTtRxbCObWBBGSm2KEw4VyeGGJ+f5/qQi50HTk
slX2Y1dnPxjR0f9/BKzVtmvYHxW4iNWmz/IkYqDwjGJT2SXrj8yEDkFWTH5T10SF
lYqSqJFdiln+T+pHibKlix+vDrPeZ8vqXoyXRQ3Gg1oufaXCg2QTub+l3/TgjJwi
G13MYqN9RlkLwF5GUVsYLOordKRFA9HjWNzbP9nvQMlUcRMsU41ieZlgSite82mb
SMrDve0eBDp0e2yOl5ZCsJSre89ZDhA8iH9xoBKXmN16XT9o03gG161RYFsT0yKb
FXjb0xfEhp3tuKsY+ThlY6blrbj/qnkUKO6971z5mRrprGZwUv/M1MsepDcSSEXz
T6cBnYdpr1Syi1HbQQCazzYt5D/bTxf1TpxFSNMkT5lwoWOtjozX3Fjd5UDDcsER
QA5suD9NcHirWECzMq7q3OHkkHuwSEG+Gc3nSHHDg2qAE4BGfCG4RnwmIlFARNVK
3Jxn5wlx87wcZtc+e4wMs+jkwb8MGvjgjFsmuMSBR+lvulKH0mcMfy0dA09ekZJe
vNaCizpqn9vBvGCD0dNFNv622ehqsGQK1speJ2UsQJCAYSzzLW0AqvLvzjD/R2JZ
5j6PTIAlwWSJUilUpSDbVO5fPrd5V22EZ4UGJEGcRtLG2rvR4BokGADp8Rr8aEQE
HKavjn3lsinH+EhnlrdTOPFohC3bu7iLxq3wGr/GZMSm/mWHAayRFwLcDkNE7US0
YTXpz552LUyejJk59VT/P7GQz02sxOIGCnXxx32DVgLs5yeIJqlAVw2wDsXc25hj
mtsTN+Tu/nhTt2eEUDB7ut60TaGPThF2XdeilHzqmdPy62UhQpj0jwSVygDV1d57
08asoWaAFGul+oX5lz3aFVNDisqVYgbxvs9yuQNB8hQhfRMGR+dO5fLD3SE3JguA
glVxGuJzUupi7evw/d46jCNDqnfVnkgizg/XLyGbz+6BxPH6BtXsW+aQ4BphbCd+
ieEtZT8YUEC1V3j8J6Ug+56SzhMemezT9OxJGT7uYeyZJfHIcvDHSDxLPFncgNj3
IAjun5gbBKH16+lV6kx+WhNI6Ybb/zd5vB2cepHBN+JBsYlNpwBUPmNRIzW/LdW3
xgSqJn2F1T/ET3TiOrgYSDf/CzfJyulTD4XG0ZrjOPhbPsMSSe7gRrZR7uBgOioB
GdxhUn7tjytsjIIh+BVkfBMJyaBc2NMXV/ZjiBMvPdPTaK57qCYTi7NVPnm2ccGN
EcKyqJwMCTSlnc44yhWfG17m9RWcQwnwnZNzWGJ6zqlHa5ByUi1J3REAcom82kIb
FL0UHJFB/VDfPOvTq/VYErQOMv75I5TYEYILgl2Gy1IfhjpLovmIdp3NyG3JCxd9
PecbDX0vodZBuCGP+bb+rH++CtM8LLDQHS9M6g75z6EBkQk38boF5zXbIoRWLWQo
yhEzzQdZfdcS6jPJbqzvCjyY7n/b+7RYgCXuZ+BBQTl6finCfvjli17XgKTjpCxR
6boUMiIGo8kx99PTugUah+68BOZLyIfyAa9IY7J3FsjLySeO7YGCRtQGrB7CZAwa
L8671pdh/ILjz/J1ru9jJmm8lrxTUDdG78kVF2pfUi40J29qOcP72MMV6dq3t1qH
CYBfJzkcW3IpBWFD8enwjrDLpG38qSnT/SsAPsjcyll+WRMjdnPOrGScv+3GL+5W
92K/z493WDIEg1fjJaBX8zgoBqr37eUQn+0R8ED6ldtru4bkjrqajz3kid5aE5IT
k9Z3qRPVUZQ82VuyksZE21uIqZPOk1s7+sb1hk4PkjmMRR36+wQREIU8WI2rPt+f
YNEC/BCcLHLiWqf6t7FMYPylXSIiPxpSqWdgY7sgFt/TFcbWfMDnjWdape+4Afhu
lDR77kmYogIjMsOrJNkcXXsldOWbg+LsgG5+dvBl7b0qU2qUfEncxJTRgIK9vVnH
UeezesD+BWN2sb/Emfxc23CJjSdFVQnwuEujJWzWTH8TBWWflZ3bNiVqCpVoiAri
6/FMaTAJrc+52O1JNdfBj/KbDhI7GwLiGygqFTXqlIv4ffTZnUqLUTKaZjNLZ/Xv
MP7ONRu4Xl6vIF9JHky4epPVTWRW+FuCHnfmvbMgI71FDAuF9+28iacJZUGluGOy
92Mv6ik20mX0OQ4HPdTfb56Upai9HbT6xYS9Zrctk9Fd8FJynwLDnuyPAb7LRYl2
X232x18EairfCYbpehOMY3p/2YhTMXrxvQ6x66XKn7vigUI/7O7x9TIw5zciU8T+
eOdlD18U51xrchNu6+kZJDyzlqOv+t+VwZ95PSIa3cxHvTyDWnF8hohRZFyFMOmI
xhF6mZFuT9dFTB9gfDEuJsFFOIFWZ0DfPgvgOOv0e7Yfal9j8vMkYeqMkE11vlbF
sAUP2F5u4ilIOjHB1pOrgvuew1YVuxLnB2wDjRoe8JJbyhXVJkqmPNcSN+ElW61c
SmTJEy/ssrIXm/sC41/21I3hVlCktoOJb6DQtn62bB14GfUt4/x1674+/Ne/E6nl
ZfmCNqWsQkL2O5oxJS8LSC3gaYvHZWyLuKI/4FT8Gda9829brDPxLYhxyIc0MRJK
7kBPjuvs3Cj/W7kzGwrSzghEDQk2Lf0QBl9Oj5T85/pA4fUvl3CXRu0nOQgVlvo7
juKU+s/GLZfZl4U9vWR9+q7/ZiGDjfNt/T0mo5fFYNbKNvZ04KMbfbbOrX5iB6QO
f2HpBT5bEqW2dNp954jRFXII7/m7Hhyn2jxi0mwMfpSKq+jmNhYg9X42egB7N6e2
8ze6JI/qvN8yeh2vhhdtlg5s0LC283fSC9HeAi0vSFtVxG/ionz8MvHGreb179Vm
DhrLg6zRAAR8Z0vAbbEdJUDzij1GGWf6wFQnBTTIIBxfYbbjBRg8UJUWQor57vdG
BJoQldkNZvBUdMNYef6wWW930JxlgvgwtZ4Pfxdn8ypdsg03/g2ueg6gaCBv6qdt
RRFRa8oqXj21fEMC54C2zVaS90EUsmlyXvaMrQezqTfNCk+2caPd07JTYFvQoBAV
vdDpzrEeZ9MKn58HUn7nnKW7ucG625tG/OElzMqsACJzEzd3q/6FsPbvJBYO2a+9
vMK02q7zG0+ilA8zDt/g3nFP8oZkp7XrNFNfTkVoLspgVK5gXhPy2DdEyAKroCUt
T9FPmQwVPQcjqT32QQ8DUYQZpFqoYqo7F+DZJHrIAmCj55A7VfY94K//usRi4d63
0OfM2eFVr/lN4xrLtZI9lTVLxnG9aT/DanfGf9WaBlFQbdpj4T8WnROq4VJgolFE
FwrPN23YFZniYg8RYUKhMMbQH2cNdxYtkVftzyLh/HOi86uOiHMCvMvNyPUQ00RW
McO+vujbm6IxGcQCxSgYj1cJxzLwW5B8TIvEypnQSOy03PNFpuyQbwmcWzzj4Ckb
I+B9pGb57YONuf0jy8uvuLCmeGDMbTohIlMyGFwcPYGoQ6ymSWkZ1Q47ztBM7hGH
vqw6l3zcSXTZsjDf4LaWKn94eZXIk91UZh+//b5z2dlmKJ/L4/BxD3PAX3q0TFWh
IcF75O8P65a40kyPSQMQgrIZg1kSAba4u35YK3s4sC39T/hYx5z8hW9LSi0TY6XS
Knc/dM6s90TLH15jG3DNeGugv9zvcrd4TnB0ya8ETgU4fCUgsq0B20lieb0b5/tL
4lEvaCll3g9ibuzSK/CUqRmOOZX1zPl1Hzsa48pg1uUQpANcoFCuVpytYE1hBF8b
3rOouFCX+XfDs3QwloS4rc5ontfIqUKL8MyF9XCF9VOY0HVBRZ+DgNn+AzAJhkY6
yCfS4Oi5JwrBry/S58Stxs3sWd5IjVZWEip2fXhIFIQot+KfqBF0IhmHosskaFYF
/AdSKiLNReR2iDVN2ShQRnZgofln8T8YsXU1jtqiK+YW3x7mUPV/Kwzr2B9nrukD
T/xYHWktLHTYG5LNJRvJpz/F39gXeTHu/X3YbsTGEWfNQ6/7ZDNfjJTNfwBgnGJ9
VyNvbsbtoOhMF76FTpD0gFPiTTj+j+TDgfQtz+xQUj++1DMYBRbKWF+8xENbGsMk
uGx0CGUJd6THIgWumfsfIjnT+3yGofVJnwTInnoLwTMUlUf3yxs72SqzfpRktkFp
4MP4+zFI0T6wIH2EjfYyAJeoIFxbnnxn3s3tmT7Kxwxj6UOLDoB/1lwo/rktr50W
9VU6ULmg1a8yw5tfIazM5BuaNnVCmas59NSuCPc1K4wXW/FwjlRX/3f+dgp2SmY/
QKAKC6xiBEvs/bzP2xifTbfsbQ4z09vBzW9Q4jmbyZKLcb5MdcA51Dltxd5znPl9
6SDyzj/j9unSI67mmbXGn4FWFLiNvlfZijnjOMn+tFl7gZ9unLEcHTuWBQM2QozQ
TlhgLJim1YMBKlnIAPjVOnBYjKkcC9Ae6VCmFH/u37P6COO65fwsivTmTZW8Tovl
khbBCReiTusrj1sdifEmPJCzqrIcYTXXIkJVJyjzsD69LO7/GiHX6yhd/6j41n3f
b14WPTdpM7LQVJ5ofUOp/pkde4nFAWLnjGrWpZLZ/omX0ZePZurC2uYhf+Wfd+zb
BsIiTVBBYi+oPYpKnq1eX1NcfuXM7KpWCLK1HX7k/LvAWWXrehgQmh1jelnAxxfV
RwY3kLR5OFYiMKB4I7bTVj18usEyRe+6rRt9CGALN4hoGYxF3XLf5+AQZxyfwztl
ZC4mYFFp9HNgH+BE03nLSUu7pncF2xA3Zc+s8c8VB5T6XxpSjZ6BQegEzE+9R+gx
1MhX6y78TfJ1qyjNE+bfR8S0KfZXqbi8XotYY4jHKNeI6ITdHiH/rojCtEk7skTj
iJ1mwlxuVDeYWWzRF3G6SHy231Y/ILeSQrJDlx8pV9yw9VhNwy237RIvFGhjei6Z
eptJbEoq3S25I8I4egjXSn4jSc5z31iJpn68oGg4OU9v33jySlDkTT+LtN6nhhmD
Chgj8MuBmQ4SR2X5b4ii2pXW2ZvJybYYH9NkVUcAa1CbuGOlA10SFvmqsXiwQbfW
zqw3xq5a8+kbC9aOI7yV77mN1xmc4w/Md7w2wUCvxahG92PDpN914q06PhfR5ThR
sfW4+NQqoKIzsnbHBgVgflvBkuqVI/VuqfyPPNKkiXftMTpljy2ZZ7VNrySzh5VK
yqsDzWfiiU7IrpAQtKHGgT53q81YhOCxgBC391OOrT2wQmVnjBDn5YXSaIwSpZyO
pGCfCu2eE1Pq2xruk2VoneWLgoY8qtYKCGlF23tDfX8d1L7JE0T92l1UxHAXiKOl
Yp1Tnv7UuhnJXW/C95gUe+KRfR47W1TePJG5jSk7T9ry/etqzZHtqX7h2Y44RbCL
g2sF0CsKocuEYE4Kj7CjNrHdMVAltMyS0a8bPnfPgSZJBscmfxwuEMi28tY3t72j
5f3Zfx5IxuQbuDPQBd0JXyyLk87QAEMNPQc+698QCU9gi5x7yfPN/ICbb9uu+a0a
kxGTO5Y/SuFS2E/QG1HwcOXEV7WhG4MkwBdL1HZBhrh9GzZNpnbKXaYtABNMR17R
oPVXUkO5IBJy/Mefyo6/NL0mH5SmM389bxmsg4bSzPePAWyMcpe19UiZVDGyAaQ+
PapNeYxTXlOxSDGfvu3YDDmLHIX1wIrIDE3kKiY6hiUG3lsP6rIJTbQ9j6Clby/x
7xJESFEuUSHuAOFc1qiqEmbodQgx09/7Jz6YxorASTDrjlPvDP3qm+RB0BvR9bC8
163G3ewV45fsav8wbaHfPGqfb7JK5ShuhiuXTawf1kpSsZHN/JMztJ1q1+/oKjAN
VzkWmqDJSgaq3ijjcwtgUYuFYV9Vx1Y+iEskixkz+ez1OWQxX/EPzAqrnjhH9bBT
Mi3Xcvqok9Va/B2xaJsRGwxG0+rT1AwAYManw++Pn2Sdz1G/fIc7FwbvTN4K0f3T
9jJt3JNiqUdDyfHeoDYCaniwKy13hbfC8FAs783ElvRJ3Jn+LtHDJZD9pHWOdncC
CXPZVrS9PSZJ3+TJgWqD5K/6+3FXppMPOIeZqWktWUxfzBlW0RHUJtAPNY3BMwee
553xEF36fdQKjoTPS6+yKo5pLF+j+510GW+fRKdpcTGkeS3+kCeJLEld2hj6uz+p
CzU4b+Ba2KysIzP4VwPNrZQVBomaMNoDzBHCCqqRAXvwV63R/C2l/lpgPXD2BQBW
N5pn168xsxODJ6nAkboLBoBM9OgQyodRVYDwwD/vyzcqNvV3ifpW0iUBt/oswONb
0B7hv2c+D2OV9Q+iOt8yBnwRvu0w8FvlzrVfdPUVJ5IjUxaBgbzwTw39AdbuwxY4
xuSLMBrgdFqUbRgNULIYhWQjU3Wfsx1bnFodlHOdG0AjVqvY/CDAlo1Rh8BlmFxF
8o0gCjJSTToCYkk4TUgn5mZipeybC3ud+t5rIlLU0OV3zNHU+KItz0GPg2yQBBvw
w1RaKvkBQ3HK+z4eoYu1y2Sh0vwusNYxPT7pPBemI5UyTXJLHtXoeM7umt1cepnb
amdkv5XcdyXkJMgydcnpbJscVeuBkjmB+G0UXrm1Q/OZzWWU1/1q4FCJKR1aRgVT
dDI6ExBSZ1Fl9gVakeJCXk7HlJL1bKs9LU8a+pkYoRkD2cG258uNmv/BLIVWm5W6
ivfOxS+5S5PsawAP/wqNrL1yLfAvk037DjXxtHqrq8y8tJBM8WwhMa7D2txTS2Ik
5uD5pSUoycoKSVlbANgVScJMAO99I1cSzsrf4exzgzN01DBqIUW3W6Kw0UsniezV
A5LbZ48+++Avt9sG6zWiXv1PlPyZ4LfhUEAshyZiixF4H4tcw+wA0NNrW9197f/y
ellTavjJtOhZUWZssUBB/UfzbEFEuqW2LY3CmukTO1Y0rZpjUiPSCkKo/nJUrtR/
2fj+rq3dJtMp8o7Ab+9DrGVV0mrV/2L3NTGw1VVwIJfXH7GCGzrCGMco6GSGImb6
p5rMDKI5zvJMBoTXPkgDyGNwyyc5HCB1lgnfOzk8k53mWk1EfP0c7zp9WOxJyFgv
LjLAk5ybDydXERhh9LLEl/ezSPhvixzv4k1Mt3ZDO57mHqpn4SA9ejK6OZWaleUC
5zXFF0eMHUuGKNXn+9RUXbGom3CoYvBnIUpI/G6eWoio3+qt5UiR/BIEQoav6L2C
l66XXYnRKEEW5IBB6fM2FLNaCymiSVe3lNZbPZQBbjRQ4nlSMnNNNE+JJkN4zU2x
5tofzRWkKSC5du9jMMrjSDKXdjZg94hIBzGF5KuJP/FpYeWt9krYE0fge/ZsK3Tf
TUEFJOJXsIhp5KUJYGQDCtf2Nqo/A5usxp7rsi8y+zNXW3PwtbqiILo8js8FTBg3
ZloIOyAfryeuW1f6Y+LTcRmX9i9J/qJbkUscIOpMX6Ebtj667aibLYQs9KB2+4f2
GLXzdHKt6D+HqJ90GWwEQGK5F1hcPr5CbD8vSPvQL+DpyV5MYSpPNSUqAAlFuE7t
8laj3aB9Kp4H5EInVJC8RYQJpA/aC9o1j5JvwXoOxuhMDJgW+DpOXrmThU+MFE5U
+F7ocAA18P7SM+GvKcF98Bfb9eR+3tOdckrEqePB4XVbpnEGW7UOWTrtA6bJ7lFJ
b9S+PRu4HNmzULVrQ6h39LKKfWUcmfRhRIIx/DtC0lW0AwcnRGmqLbA+7h1rIQ3j
onV3q0O++TL5XcGbMfNnQhUPABrS+F/IRGMTI2JVXNo4V6w6OWanVEA2OhVYNc4z
ZWBOUNSTLXD8wMsXXVsWBuJMfrm01fST+zYASec6sRs8bHZNhl9F6ngLAvSn2NVw
uvwBSanAMU3vj9A62xJoG+8O4PwyYU7o40pH+HV7p7gSkgQiZCqFM1t+9Y+2ESI8
6mFXUazfnPIJBtRzQjHl5m+H1jXsJgZlxc96iyM2Y6NzlLrANBmnTZQPj7g6AENW
iHG27jKxht5ZEaeKI9bjlAGV2mmT8uuz/dZ/bayPqeDk+NzhlmONFrAyDdVNMiYN
tyc09h8Jdyw0N+za+HgNqbtDxnDlYG/DnXaAQDYjyn2FJag9g7Pubih/0p1reMWX
C0P72jIMuZ2e/5Ej181FZa5E7+ETtNciJXtAP6JPRZE2fXv5sqEIXMQHx2SnLtwP
uCyd2jYDRX1h6HCMXE63vomZHHoV1hesv+EfhwNs8ooi1gfB6YQEiIe9/h/urXcg
iIa5VJHuKJCwfRqTDDXjGzwT1DIAVKAbOTpd61yH3eHO7BgAm2fGzfffV4IkIl+d
KNVdbFTy0U75Qiud84jfKl4v9RJdHOFut6SG5cZ78Zt3vTw/vYRSF3abn/5NE2CL
NvP4J9EbBW0K049ngj6MX1erbmDEW148Ht8a2PmGgD03uionBFDFCzDFOLWIsu/R
S5hNb+2F81ZcuUAeyHMW4idAzEPl6E0oDuDLRCf0zrw5Z5Fk8Gv1QYpyUAmuJOzl
GXh4SNCgGyROV/VfbnXg5IZ8Fkw4Zjwy7iEB8q2B43KxV2bMO3mFtQYOusWybASV
6dyaw7Oafu92IZPpshYhx53Rk8r/WPa0Qcn3LQKeiRQ6K6yHCSYKT52RCON5isdp
q995A4s6aRbJGyGeKEW/wT/T16I5f55zvAA/IHWRpn1AkqXRY2OHg0lbludFi1Bx
V0rDp9jAZElFH1C/Rn6Ps0gwrkmNn03VH9VSj4T/UPCo/aZpmWNpz5A2AFgCGFFp
4qwhiutGnj7uP45/7U019OYSXGmjEcFJLy7uKHo/thilBCtIB4d/yScvvoksbOxV
D3g1Bi1pMQ/kbqBcmtep8QngxSk6Wa77zLdt5o3n3w8MdKO3EcEvlJmQsdbTdpIb
n2TcxPIAY8j6o+WmKV+pdN0rDnX1Fe9+i1BcaJRbwmLNdkSEOTtcIBqZS4NFLcBV
z8KRcm0y2sI4Pvv1HtYzf9aGrSGRW2G90OE9harpteorJcB7BoGwNzsnWSBO0ZoB
rwtiS0yVQA7JKix4DBFkJE/U6L86aLdIDtfI20aorArYx14QavuI6tHaShk086pJ
vd1p/gcsYqsrTBAubNj8hTZ0Pc8yO9d/3DGOpUn8kjLhKa+QkXtNmscjZO1VfWlA
vjMFshEE2n+grM353cqbLU+PcYdab9dVJ07tcCU5mcxTRPQaYOn46vKFl1WcW5rW
lYV6Y3YIOHPYwXvLDDVs2Uk87KuY+4yZIiVrzN13Qvw3m4cB0SKfa3xhP+w2t/e6
oxiaEY69AJu64+A3ARex1fWvcGmGe/BCyU+jojn/iZairFS2sJtXE6X5AUbcJ+Rh
yjM4MB9ie7eWfb6T1efy5g7M+VtJVj6yHEn47gi+g4IyH6oMHYX/9Arm7pxW01Qe
ISLf3RY3bXSFlQVV76ZW65/OuQJIAiTWJiPzuZ58YOIMacdhg8TkGHEUg7QV8LnC
fNG02wGvMgGO4WO08MaBA0jmLZhDBnXCt3YL5K3cz1jAk/2slB0sPziNUnuIbzzk
ukKKUAhJHEXFLxGC86ld4M+JtTWfBTT9o7QyvAEStUNv1EoDCVaX/pJr3FjQ2HMJ
ET4SfOH7ouJ95TLva/gSTu2XWFKKhLF62nQ4CR8DDyPTt9FbjUemqJZ2Evy+reEm
OUT7q23BMa58KcvwaeOym6EbwIm4Ygj1nvwYfGExz4GAP8jj7XxrKSb5xq2fBwo9
okuw+gi43k0h4dJcGjamp2Cx7Et0dfuAPFc1a8qajhqiMR1vXrgHW+4Q8l4zbdVL
jCuem9ZS/F2F9lk2Eo1psw5HF2ZMQbrRMt/4VWtwH7/WgVhZE90Q09cc44vFwdS5
r+c3rjA1EsvO5jXAL4YeJOCYe8IlKFYOldqX6Ga8F/BGG/p6fNTOCV0ZU5FXHGZS
QhIuSoJP+5ksNBEX00WzlyowEGScHXlTWIgJ6eaG10hbGRcyp3krvy6NEMivSAdX
LlY1BcC6gkC4fcTkc5t5dzsbPCQgtPSPe5pcexbkpQVz9n1xnefarm/+SpyyqrEY
zQSG5lnm4IkGx+VJrhdIj5ezA+Y4teaLlu5ynyvjr/8fzoCH+qPsGwBvWsy0Cm1z
GNAlihVgKEx4eQrET5w18vD1cxWv1PsIBncPKnBgrnIY7BVI8hbRHFfHkdN1r6bB
MiWLOFJUo2FCBKJbleSOhe8bpxqmSTlgj79+e1U9jRJLbZO/TcHhHeIq5bi59rrJ
Z9YR4d4vOQfjPF/IIMFlrACcRwQ4Pfcsz9VoAS+ZY6lHyh+WLNY1ytYB4nNI+LBV
YqkoFj03FsRF24xAiWmZYTFrq4BnpbtjylZ7cYesx1JXoE453V9U2IgXQueq+Bjk
RGS56xURfCYmZlmqz5+ArS7MaDUypBEpOCgojFZNoPpjvMznDAPvv5E71W6gU9PT
wEahFdpZBAmCFng7+MEKZG19w9sEN9lxNIzwbzYyFMX5HWrMLfDr+rCT8Y7b1Lkk
2xK/yBTKCFwbzZJCWbpPIgunpOhjAMjcBC4ypJyY4qx3sWbq7nAOSpB5l7OrWvGT
rZHRVnJyQJ6Y2fIumu02ghgDaT+KUiJ8+KMW2OEZETP9Yt8EuOWg4a7lPz1ABPTY
3fRw88VpH3UAZ6R1mfX5mJYyQMpj4FbfWoct2po7oIyBA9j+0X+l/q1p91grJLGC
3Fjq6sdcfWcpZgzaBclukrHGzyGw2vaAHiySf5Jgr/OaZT8PiHlUKTDSAALB4XdP
Y9n646kiH680O841oLbYcnFZpJYywY0sm5C7aSD3yWGtJCGgrROc7nm1W8WXTQZ7
GKiXzkkEznSepyNpSGVIbmCy/yq4YzziI47+il8KFuWzRXZYwxaL/KI0l1XpC9sI
yPGFD8mEjp8xqL9wLF00ruBQr96fepoUF8anrTTOHuC0EE0KYMpfeeB8xP+qR4IJ
XVbQnf0e2miGTYTUJTTOpbDV6dtX8HQp5dgjh7Mu8CW1OMqG7ISVDUnoRs90/Ta6
UMbV4Piy4+otz9pczTgkmDoQtO3y6Pcin4rVY11p0+Avw0L5Ml6s6f/U6zop3znq
EoIIbgLAJKr42+GjbgyUxfHkHFvPYXiscILwF2qLuHLIkR+uZWl/Rmwk6gNmwg9P
7VKizJgxVM55LEZ1bkGGVX/fu1+ZVl/3YfeLLcnUf5UmKI9SknIfDYPgFPiiwbRl
Ii3m1q73FHXYvCZWNQQF/EqLz7K+55O5vhHRQl/AzFxc40mVGzlUTnmAi9LLl1Gg
qbE1A3NjbyfsRiF1Ec+IfuIlKbAVi4/xogo+stHnQ4Uz7Xrni3WkbJmPx+/GWAfb
VyFZp0AP7+vB+gcaJ/aPP39qIx9CCnzf8mPi102w+4uApcefaAacxkU1LWd661ro
cMhdrW6V1PWxStSj0scKanta5/7KweUxmLAIZeLA2vGJ4/kJ18i4utj7xngfKy0L
/ngdEj0EGJ5W2UiFZNzFd/viION4u9p7QOceJ9s3D0DsYkqUfkygXqnHjJO7xerj
CIjbVplDuSHYXSzUCpgxJA==
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
CxJgXjQHj1jEndtn/7ZoO4TfrlEh7MiYh7u2UqJ2vRPNVuryxq627Skms9Zfatw2jrgDnYUfMwd3
N5MwVbdFl2gWvbvmplZN3gP04vSoIli6FIGeSiH6ngGwNn+n+U6PAwasYeIJtXLOllSJnCEbifl1
LUHpkkSgzPBlApNRWnfsyzLMhRJsU7ocCzemfGnzJEm8X4EtbWHpHgCeVyhmsNmoUbMbdHfzhdz/
2dBy9wI0R7+kTgU2t+qzaKJx9fJPfr9UA6icP0VpPGnTlL9u0AsdMCLHAS+WkYqI8wZoq9ESVNsd
S2DNip9UyOURUKsCbnDqwBb/T+W7j2fWRdOnTA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 52352)
YIwDvKpmQZ3ajHEQzxfpMIOHjhV+u6rU9/doaVyaoduDPQGlc/Aczs05q79CDk85p8AbTvLFNM9p
wVC4Z/8G/3M+scxUBE7CQGG8sGjF1jyx8V6ZLiap8pZLrQ+U04kQSW9bazt6nKzUMA7zysCJf0mw
UxMCpFGhdqE78nLofSYEZqcSx27c+uZ3yW7i2F9ZN9lbWVR9+sQXrC0r00Bx2zsj6V7kiYTXWXH3
9WWwuT3aPYIQ0TXEPWAqyevoDgs44+guQdLp2I0kF4AeN5HdsJO3sQHWZXq7o6K5b2OHVQsBKZT2
H1z1r/4pQTIy1ggWT0ohDqh4RVZggMb5GDMRAibQoyb0jKVY1jb6O3IVY0DfOtjDChYMLqRWLe2w
NfXiBF1ihsX2JJG3/EV8x8ZxGHSKjVOuZ4iY7WCwJc6i+QhC+luBSWkDBw28Qfu65v5EW3omnTv0
fJomoBfJVdP0xobbo1XboMNazvQOzALJOdANFR94GGGhezMnBnkeHQt1CNdyFgCVhXw2bTqsHcH3
/uPZrUljcDR6fM0r4lhYraJ/4vBlio042Ij1pKH0du2dPzr/NWSFnXCmBEF9+3T8bHo11SjC9E9x
1E3PQyjXPozLox6hrmSSkz8gVfCIIWvXctAmHVnMC7Hj9P8I2F7HiVC2ZpnjuulLzj2Ybdkyd2u2
XaDPek7T7ISR5tFDVOk1E/CU2rJczdH2rTGmtUlDCgBdIfFCVZdYsAd2rlVDFxc3qWD+Sam21dSy
pkulVk5piI6kP31bvR12rF2AY+i6pgP6u9XUUifdwa0IUT7Sr9T6FN9THPp/2T4aRfv7Z8nN114z
WVC6INuP72c5z/gpIqn7r79/RzDSMA5KG+B9RlSMjrYD02B1kGJXpB5SFp8RtH85kWFUGaMYXJRh
+LJLh5zH7WM3MolSNdlGg3JG9JYfao620bPg/hz9cgim7UJcf/Y1WJ/d/8obJMONPPqzuUD2nRfr
WdizYpJy2iM5dja1tHhY66Y2uduZVZ4AABgmnP3I+eAifzz5iKe3j+2bwFK5/4hfk62TD4K1v5ah
dEsvBEE0bXctbnPwm1kX+AFvwWhAiL7TOLIOnyeBT3wrRqlrEs5Lzx1Xhn75SLJvhMGwmZHi8Lsw
d3zI1MYhlBxOCet/MeAG+ETNr0fFPM/rtu7q523BJ0NuU2f1yQINrCKSIq7WcD8v3rSNA7wELxrj
1FjiljkIjmxIR6N5Y+CPbIrnR+Dbp28OsE0L/kbRDGXgYbYkCk/05fJ2QOCJ1Kpj78lNE3pAHYh1
sj5Qx8eHPZcYfwoveQtZ9XQnpWrfcaB/FZjr72xYj9YqnUg7S5vWaoaVFwa53V2oE32F/xFyU/4k
wZxHdvrPQRfGuQktn/jS2pDy2zejxjijF6u8VHc+6eJLD4SLChi9ouZqDgJ5Fz6TlEbtuOOe2WL+
uGKJwCXQB6xx9w19lGmMP7ijr9QIP5qupyvlmbQV8xcwAPxjAAqvIcKzsSQHnFljuVrS1C1PzaIM
Au1euS+gFGqi0fpswGOBQ2DmkGmfgvwJ0fJwOnmQtuPm1qy/eW5AVJLdqiIMkPHW5yT5d47ysjMh
bCSnGCcBGhTGOLYHSdgpRLzsOitBVLrYT/cc2e3Z4UPyIVreFRqzKwJNL6+JeFBkMuAKb8ZGf8rZ
yhl+hd3A4BOJmC+9J5le/BJFU4jc0mxJcnklmfUS12FjwgsbmbvalBaN21jtnaOWik5xKiQ2wMPC
TVfg7ClSQbD5V8nalRgA3181ZX/VwAbss5V9ZjifnB50RipAh9rMrBlAFIKej7qC9NkEZxYCVXsp
9wEyraJ5sKwcS4+Kia2GEzrRML8TPgb/Pn6tHptAMc898OVmycjtsQuDsy7GGYnF9k1Lio9zaw69
U3vOp0acvRXNMUkPOEGhDNesGrYfXdr6Oxmdi8Pc1COEaypwX5KALd3mD89ghSn0MriWSWMqmLfW
NpkyT78SM+BP7OGd+vZ43UwnvHsFQRRfr2WE24un/5onH9wa8LBN6ynxuvUjrVAqD9Vb7ABhChJz
Zi+rbHodMlL7dSEJqBK9zu89dHKsmTlEYosliFcRCW+OqJt3OW9CX6g5amHZK9R/rBFZdhSKfwEe
i97fc9LMoSS/kjqLKCVVO3416GsO/wL8BnLl77LT+JBS4JQpHVbG8sDCOjGfuvYoOvVdc+SDtHBQ
WDYb3SfZNacx+Sv2rheBUjSjmsudmw1v6F4fM3i4+do89MudHqNDwcNgEJPJDKqG36y+1Ymqa27f
+2dnT25RUw/zjysbKKEhyAxP5ysmd8m0Cx2h/yUQ9CsV9l3lQSbeRv8YEHWRSOXDHxUeBt6ORwYQ
WSuFmxv6z7yArNA6RdhTWGKgIDpnq6QAhy+ErvHWFd3Q/p8G/F8Zphucq4ATUtnbfzDYBtLEQvBN
TseG4pRN9d4AL3yS/qnTegHyvZ3znAnuzLEbK1LMQyBHH40/aZVgCZESJjt1/NclCCU/ocD9yPVT
yTeb4Rykg+MpwTEQDizPiS95RtOn6OA+axtOc7LZsr0YV1FTIk5NseviBBO7OkTkCao4/VOA2wJt
N8psd48VfVZK24MoNiiTiGc/pWnltjZ0knEFz2SOH8fyKyxaib1wHIP6lyITULwz73wjuvXmdLce
XM3LR00BA1r+kXCd1EENYN4n/7hBuxQjLzvXfnSufh0+GPCW3+J+2nHyE295ReYwaxdAg2/CeeH2
iZo4O/i1MXAd+hhUemJCGcL0tlPD25cUvT8ubXrTfOVs7uxrvXzC/52otUAydDrosHNG8EzAq5Q9
npp5L40jMmib9hkSpADfnU/tZnboJbKGY5v8ljrT4mwMG6jCS3jqIHMmnOoJKYWV2nrSp3wvXBRD
2TqEoX0xg/eiZfoAEsbiOiSMBRoibGV90A4DXcOnrT9kJp+wIdvKzggncslMrWJUzYLaMN2aZeP8
HakWXIIjKgEEnW2Petid5zWp+6/zOp591m42YPHcBJ99FO2mw4egLHxvRuz1Wu1cxjh693P3us70
8xZpVuUg8MNvNScj5afFvlpGJyrwURH80gPh411bZjkWJiFXxSV9RCsvUE4yI470BNVyRsIKrEI8
rCfX9Ol52/i7WAStai5giMIrgQUxplbVr1wVOu6q9bDzLdUGPfctsYyzT6FfHffo2txpOoOet0aw
yQWq8WmLYatSC5Nx2geVgpL1UEbOmyBlNw4GCWvLGjdCH+FgSg/n15QijyRxBKKdKRC0gGgCul6i
GOyx5dMvFZAJMEY2NiCg5HGf7rVYnbUMYwIikqc6liMs37Xew4E6HfNLX6+AeSmFp/svbDXLYK49
i73W4mXWl7XhriL7FD0TBaKjUMrKufDMc4SzX+rZplQOl75fqSaY8LsSMvbUvSdHwZPmX7p4F8lZ
idl/TRmX5IRiboxrMXYb03HSwgyR7W/eC8FXd48r0TXHc4UKLIwJ8FPugLpnNQsL410h2J6Iz9dv
q/niP1EoKlkFWD8ZaHzfeoMKAX1DYDsFreaHK2ifn12RqWbrBKlLbTHWZmUhYgI4bi0X1CWF8M2m
vYODqLFvDKmVvE61fo5WyODPZ8j+v2QA8lg55NR8uD2EJ55/Z7NK+U0sGEa3J0YEBlTdOTNma6E4
NBtvJe96T5/Y69+WRAPNN/W6Se0NhnyyNbZcVKwEWUeAwdSgwolmb406Ef4W2dt8qZF4Zoez+3Ak
KTV62bUgjo80u4IKVTykugFV9s8klwrt5d9ByI7zS/6PXusFJDgnnMtqL1evrXnHzsx3+qS5g+rS
FRiiFJlARha6y4PUmVNexJocFrBVrQsowZNOmGIB5Y7gTKg0Nc/TZ/k/QtR1XAo/0vG4xCW23OW/
0GOndZXrO3/3OgkMFo0ULoObsiNkkJvteTeuo+Qh+Dz9El6Y8NPaawfo3snSyn9b/GxjaOrNpvkv
/gWLqT2auvpEiA/saVOlBi4C/b79dlNLp1cITxdIAQHfXBH4HYZK/bJMiN4b5iKywuFChRB6ApWE
pGfvOjviw/wV2SXiKzSCfSp5ryvC4fu20KcW54NMvcTEWGODIUoND7ItU+vb4MJZjGaM1aKzEQBN
M8hknQ82HlrSaSxh6Fkd9e8q4FSp2F04XzyXg2vjOIVQtVNcuKpPw42Z/KEsjA25u0WEGZbJLOd4
7yWiYlnzchg8D+Ys6jrkOhmcDTk43sMvGF620YEs05289mnE1TDw4VamhxAE0tN0pNTn3w7xU4tw
kiVElSWdtKKDuN30DK9/+WyV7tk7cs1oKnraKWyKTWWOBfoXKX4+vxjsk4gDH3FMHczJRY1/kwYp
EF4Xtu3Zq/GhQYofhsYYVHiSoXe55yY+UAkgWcGc+SzcNIpJLIAZIULAGdwpa+M4XKNhgP78oX3e
4VUR0fHRamESJQ/yPN0uxS17fcsOHgR15ygAqfQD9roJTAuAUmvbm5DtOesQ5M1sXsatGMVllE9l
cvgp+yCo2JoOjLAMVSdFrSGcBcL9/kuKgVqteM4lPwYehQgT3Iv+T7pA83LeU4238CP0VjV784hS
ybgDwHy9FjznHGwwR/C8YBIJo55Q0UE/QpQjPD2Yg81ybW/fOFSXANctQTEgyn1Cjc5FKr7K4dD0
YfxcCZ8UEPVEg5Sf4NP4mg3Z/z+yN63ok3uorObrUAGBwKIVR8PnsaEUuqqxx6dqLWQAady2exc3
M1T662XuK4DzTz9IDemSV86qNGiVrIgvnhU+EjoZxFQtJ8eYEiNIcYYUk1WOvvaoP2mNcgJ2t+M3
vNh9gKdtqiq9Pimh6gKbtzjLK3BxdJD2iu9X0VVEkdJmzbSfV8qzhIzd74u+Hi+K3u5cA1P2vVk5
7b9tswzk/NmMYnq5TP7j66f0g19jFvAGJ8mkY7rrRxM94j8bjB/RbOyqJW63oUBf8vgXISRVYajF
1EkWlq7QjOFNh2ZQSBjWAgLtggWhUHGcf14224cqfIvOFml9fnd0dyuImBELYjibGGslqoX2gaF9
IQpHvq7+ep9dIVcWmlSxV5Wus5rxqvhndH7Y9YhyZFlVYgbaVdex8xJGz4M4ExOVtDRzB+9YZfmG
wCKhbZ/+BVatbPBXSc1hrXaO2j4o9QpoQixpgc6oTfvnRNoXFOKfY9qbgIAkXZHwKg2jOhdHpedZ
MY4mBNCADavDCv09DBjAd9khEYGx9z9bYtlEx2FLvXHAmvrKia5C197ljc4gZrmWEaHYocPRVNWl
tWbj4TAaCzzOkcNEZicoL9sl4VXFkcZrTNuDMEpUwRktvYUKyEzcKe0uAT34KqT8qqjJDLW08/Yb
nAyNCpHP0KZltMIpK02L00YjPXxsnAznv3tlIqf82HiJjunRm2QoX/B2SSN+PEuYyysjLUAbXnEe
aAT6f1RgTTl68G7IA4V+u2Zw8SnrN3AuFkT+zyMFh57YJJNYB2VJDoKKtTksGp3lywoE3VHYjHnI
J0wKutlfqC3ghHN4CG0eDoIImbmhgK7mCunFOq050Occdo9ICZz8HOlwBuIe2azGXDYm6K9jMwi9
B+L71Onrd5Aw/AJMUFdnrxcknNPoRX7PwYseZC/2zglirjiys7SJLni0ArYJ/6hCtTs1oteuRHFP
DITCvFxYw/aEDUJubXSR8h22QdMa+bxO73kkKmpOSg+Dszf3PAQYPDiIKP4Y0BwsFY+NAuYWtRHU
Otv6k3FYqxkWNgvTM1V1vb3jSD6sggDeVXw6n6VT5FvPFj3ZQjDtOiUovAO/SDzgEX6gI/oSTGBv
mEHbciM0WgOma7CXKMkUd0+p8nfW+wby4p66SGrNTwHjGe6rDCbUAScZWcmSXYmgZBuxY9535iZv
Z0EHPF+A/DG2hnOPo8jOkRZ+PJiio62Q9E/JxNlIqMYqR+baJ24d+K9/JItI+XHV9rUFoVBhNDjO
+qrfDVIiS8vqkMNBv8cZq/XkDzLzyHpaNop8j5lV6dif1VGsArPJmRlXZkcrPXGndHUMP3OoIUBO
mCmLJ6lSZVy7zYxlQ/GPTaDk7srE/UI6ReBc1lgR0vZser9mAmcApt6sjwE+wyMAtwHxsjZcPw6g
jyNZnQgvFjz5EveQaZZa8jSsa7wGJJgkfqlafiTkBqJe8QGgST/MH5FQChOL0cbXqtrO35M8CaYt
gQ2mZV6Y6xZgfSGOFVrzORAqQXCBqoAlQwNSxbsmbR/gIzQx8IfJH65wISoNZkS/GGGsfPANzdBE
Avx+G9O/3HYVFeg2/S9RHtYtC9+OFQCPj3dxQOlm5GaOJPGKdVPQaidjWtffK8xAlWxErVPw3FSo
8GC/BtpjbUJ1HRla6uM74YtbJX2O/vIQhPnikjwC2Hkoi83Px2Kvt2RXYUI4m017bEycteNavLtB
3KSmQtDmMpaEymMPgMfhaUlh9fV1echfZF2eDK11V+d8uZeRktquVPobcB82Kevq30J3Lx8m2xdT
qqzUxz8ypVMfkuRI/TjAbIEEjngzp0vkzUlEYTyVdxIFtZCPIpd2CI7sbJ3ZIb/fNrqV1nxEVACW
iSgpFwHnjt6ESgveoR68W+fobTN8iHgQxFyh+cggaNUzi0c+GNhDqtFKslG8ZE/15TUZ0ri04EK2
eOF7hOlaotKofLc89lh4NX8QlseVnEqqRhZmRKMrCKwEL7HGHSbfFr2Q3EXBfxlv4sEZ9E0N0zcq
NMqVp0bMGxXB/m1x8RqLacp/4Pbl9cHWBYPY/bj21Kk+BzIofmn3ssMui93c/llectoGHskKQX+k
xAwHdXzMq7sjMw3nkgKn3xM4JpO0jJOP6wXyLBX5rrwzogzF2PddRH8eiXRLzF5j+p/RbOUW2nYx
g83DsttHbupUU+ft1BAT17IYvRI33F1zK1tPz7mGJ7RfgTc7J8hFUDjzWudq9nFgMvxw2Xyj6fkb
oVm0/Kbv4gxoiKvMYPV4bD3qBn5+wLoig7gB5HUHMKWyx9h8Y3HbiFwKp7IWSNzf6x5dCh8QJMt7
jGFXXXvNnf9mWHpr6ymd0inv1pcUP+Ob3AFuTHuAzLPcyFXlrQArHsZKquQfQYnYun7BpEf0qgch
Gxz2OBKVJzEfMtfO0KzCpPlAZkXiNQRDNHBtEFAFzg6Ij3m/pOoo0NzIEzVUk4rqD/QiYSD29FYa
5vo/GO3FtaGDovbcS91eFTYAuD4FQ5Gn9p69FZSMxojh9M4AZ/z1NuX8gkmZwCjsxyNjANgtdqH7
vnLtkqLSSLBM5inB259x6KqZBhqpWKQI9Nqu/+1Hua0Pv/UcJN4H4n46qVzMxw1lJ6Mgsrew/fCR
/CZHjS815dE0Bsz5hzUK6NXzmfukC5OEIJjhKlFLmEndfkCkyZpR8dE+yND4MAJ+LAwCQBdBWM06
McJmzSrvPKOYy3O4meIDhNOfdQNbIYKqbfHHsg52cGnyY3AD4lrm3uKBP7eplD7qgUseqHhfDSf5
cBpciEXQlWTD6P9teoJZuY/VWWfvf/W/64oQwDCI84skAHrVAJ6xVsKgmKh1jqAgpGzHI1P0wYMB
SvMOP9pf4NFlY9tp5vVbH209C13oW7ujgh/I0zEyrbxiQT2duJtcPk60U3qvNGQXyxQQB98B9GkA
jx+nCljAhuIILl23rzOAU891/wJ2UoF5SvsB6Iv2AdVCp5sO3OsVsT7z6cbkQLXo/FmRGtZ2Rkka
+wYE5u6mZ5WrDV7JylDaxrGPmDs6k0dIxsPmzYP4LImF5Kc0Zec+q5WxzPFFU7F5a2qiOOFyWbnT
kwKdjEEmuhNlCYTX0EkSuS9ieGVHBARBX9n2iNz7sUSslzq95CgRztbZvfX8Xhzxwx6BKRqoqKM5
3E4ixUfw4oBI33bJhTbPkbJ1FZPlOFkR7+mVtuu1Dj1CpK+gZLG6GBlZQi8Ib1FDuVIyB1yT6nWL
KDNQvO6PV3MwtYyXQlV7MsDCi3BgYhnTgSgdlVO3gWYDJFfwlhplLDAUYbhlnXSN8XeKD9TQbwy0
zf8YrWzH8fZJ20L66vnSpzIGG7KYs5y32oxJ8cdM3U8nC2e4Fm9RG6SabGy7tF/KdUqfeH5hBavi
mGFpXbmMdm89O+v96VzJFnsLHoku2mo9ew1TWdPGNtdGJjJH/WSWmrDi2hZCw3m4zb4CnVqkuKO6
SLdXx8oVjZAMKkTUpImSJ4lnLUtu6LH4RgAV+BHE2sF+t6e5RJWox0dEG4i+W/FBqJuO6upm65R/
HQIN4noRWMLnCYDEjwSre7jl+fo99ou+wl2iFLV73HivA14FBy/RlAXQwr+2BAPh4bVg5l2F/lSk
DgjCD/MU1+moGw2X5S7l17WCkPnkfgSW74HHO6q2wuTzVfwwaddl9rmidSYoJwiYqEEsZexEQnWV
yR+uv3EBzoYhNGl5uGWifDhsH7FOdX9U/gCUzqNJWOuMUIX7KeWjQ++SmDgiRyfZ0EraVdmJlfBd
cqhqE7NF80Zq7tqH0TUS2+z33xmUvytMh6VAsrgcZuOV/H0FJkno2Uea25ugu92J1hqcRqekTd57
S6weriKAWHKnUgYr4VM1MnI1cheQx1ci+ckZaxCn8GjygdOFKLvI3doJh48s5mDF3zhIpiUia4+4
Bp2jjibdoQ9To3YTwG/S/HrBLB/F/dUFDARNBiOvYon6ciziYXepsEkR/DDkbnLbaQQZBCtQb3Yv
ylSzoROj6XAsbbz+6w+2asIkRKQS6beS48HuX06EEH9pnxQcXpBQ5CVqYv8PJyciRNFkxMw6uXtq
1w20bTMurXIy9NvJwtSgc/6gBjtgY2peZb2823EG86n5TrOVFkbYwllPusYFtFabaEkke0jTdDjw
dsOIaHBi+MGz6ERc2+bfvsPxqgNqhwG/gsLViw/OvEpTRO9IiGDd11mgfTCZwBnHFD9PAJP48vvH
G8KRnnZuP7SN6jmqFxPK3FHIoMZb5tvTTodI0wXrm2vqhOdlR6wf3lgZh/5vWvCsBwTAIt0Ho8O9
99sKJjOuodEgfOV/fo3WzVpws8c6mM6sMYdxHhl6RenOtjnD6UkS1+pyueeUHBOQMPUR6drId3AA
Ilt3tl90rCZ/dLfwMiXtdo2e42mKCIy77dBAziat8hXmtTNcXQy2mHbwCjblj+yukZgxlaIhHJ8n
77tr0Tbh2xJUEbHX6LPdHC/x17uMHr41gslWHIUzaosLDDJmoWxmvKCUN7d3YjjvCCRomvsNbmoQ
9aBrxzkeB3DU8urdw3rEv0Fh40hjhSpmKVQKK5zQDrv5RrN0SAX1woPljBaqX7odvWv8VWjT1tj6
GaQ4D+GD7lRNwRDPLf15KjxhVccOX1ARBTyjo/Iya7f7gRFbcbfxChcHkfiT0ZFU60VyyeNkJHRe
9hys7l6GWKWSXxCUdbmmZNuK0+XI7mCqKTKV1hSWGvRIKyb3PmcAcOeorB1PHCFm85lDX4lMedcR
g2oAYvnhWoL6d60pkGhWqPi+sDuEiWQ967z9gBD5sidjf66D5eOXmXTGTwKjdncyYWIWaARUh+eP
NaAdjX2ugd4IMAoz5RvelOWXUWtCU0iRpQxWvv8i45r5GLXaPIxm2G7ukFwN/eTWOuj+fIRvLGUM
EwKIGjKiBTv9VG/UKhp2hak/NSs6rVFuX7M/EhIJJcQHZ/U5rYBmxOJsPbthKUQeyyUYAZBHQpwt
6ucBRhz5dy35kIhVngbzpBBAK4Ifmsf1fbJQRz+tdX74UJ2M2duJOiM12fFZON0gpGnl4cqmsqb2
KOe5Sq6MhWM5upGYgB5/nxPd/aWFXzD5oT7QkfSYcNBS4KlF5qpOuEKZwYUWYjR0idkXMMlKTGGw
NRx322+6EpStm5jPw/y8XoHrDqemTawhN0rWKuo0wGm2kRL8DEKTbZLEZP7EghoENn5+UYFF3EBQ
I1I0Xb1kofMdk7equiXt63KGu1HKsoiS35rk/LiouGecO+8kbiQ1633IAqvPCigE1+H5cW69+Gc3
e5SDap3S+caa5vXVo80OtywAGkjHrClnpTDiJEbFCY44jJTQPtrM5xtBBTdba06wOvyRlf70bGKf
8PtkLcUsvyEZDPChACIsZLJ05oxejSW3SsndmLuWHZHRopne2On0vqL0V0VBo2xZT6+vCugwu8+M
mgJyeXhU/F3NrnYJ3JS0RM+bZSmddm6jPDYu55pORhA29pBe7KCsVvaGcTlZNRD7Qj2rNjMvMa4n
qoGmAK7XT/+Wh6wyaAV5/DES3AYvXCC6VFu0329u6pocpANVX+DhZCPzX1/Ev3xkjPvatTxInBJb
0Hpbza6qZtWs7r/hbijAbgLz78wfEx7LHpUzHnERbOXQdWG4alJWU7tCbotsnuSB8//VW4Ra19tB
8ATndeojt5VjunWPq3ud6YVjx+nFB7seWPTetYAXwNvgbl5Ga6uf2ooPYuqXIxkgF90RP4MZXH25
YT4dph4l492ZuisshiYZHBlPG+T7K2XFubDWRyz5XTktSbP8gRxbLqBtKjF/ZoBupw4UX3g2V6sx
M3kyMtJJiqy3Pt29/CgTT9P+qP7KOad0pAqFj70nEL97mFXGqTU666Hbt7Vo4G4F3CeVW8hmx+C7
ryMDeCGGY2INCc9YJuSrNKCvcuQQCtiRXzsNmwVGdNyHk6J0wuDTcD9GK32SwULYSarbf5orkOws
NktjAsPSb2Vpd4ORg6qg6JBNdo98nghbEQIFf9U/g4eexOuG6w5TdF44YKPlNUNpoIIKjkSS1r6y
3KuuY6Kgzjg3jjwPWwm5joNKghM5O7OET/G/BH42hkpZqPCIF1ilI51Xl+7XHSDefSZiopoffP//
1HYbSQGIswIXIXq+RyIwovtEveQqw+lItQ1TQ2JNHqoZMR1BuC/KDun2pKtBmdwawkbzk3T7b/nS
oNdWNNmVAmYaFColoxGtT+a906ddv2IW0fSGYTwZcMVj3QSjydHg7nlhvhkJaV20wetprAIhtXop
opuq8yPND3QWrY1fynSwdzSUsNC4SDtci5//SIGsqwuQhbhtFiOQxaSyMRYcyzO+ms1Lvmq2lxV5
/xZ4zonEynxQiHVqMGoDB7fpYkJQR/XWfA/LcTErKxqFr2J79bd32+PFQonTMB/nE78A4tOG8VzA
99LJrsBuHP0I22E0dro6M5xUsuqBTl9V8JgchxEWCVGxcvVXsgevKW1CcW9kc73M6d/p7mwh5qfN
lfN/gh1eDFa4UQ3bJ1PrTCZmeNIPeAtUDx5zbMpwZglPUn/iPkjfOr9CBIwqHAfrk7ASX6qqIegE
Kw80y9+oSS6E/tMj92m6N2mVlj1slB+8zkBAL2o5FjtJEYLJlydZkt9XTnXdLaw5AqMpOIyFl/vX
UxWdOaNsiw17519Xuj1B0kDKT46X1u6+KmnPplznqtUNa7BK/KLDNtcTtUtah4qtKC7OBaElbeLT
/JLoZo7K1DIGaCUOUx3ZGDcP4MZKKAM9dJkWnFZr9i8InQzY53tRB7H+hAvHle+x/P3O2WLVLRel
KBZ7uSR/syED7qVEfsKTMQGwQuQJMFPlhXaTq5yofrUlwNdHGCtumAxyIJUt7A1iX4ut1hkCyetf
SrksaU+N3Qh01m8wWaNmS5EN2rpZqHuLWz/mCu0zCp8agqQPW6eiOQrqBPj74RlewwFI2ZlX9+mw
cTYKu4SY/9J6RSZbhvLK84ysmNUN9y4cSjBm3DNbYG8vkF/iFgs5nfFdEI+2WjikSiktsQkfn1rs
5KbtWZOyRNQrJguc334pkeYbieeE3joxsRdGDxHalLiUoTTDSmx2wIyau0ATUreC/TvocypsF+UK
y8begFCoHJ7Z2y46aYNCsFjH3FLKP5kgw/juxLjgf5v8WowIrPwm6HEd9Pbu5u7lyCzzZOrjh1aV
qou3RTbwZI+pHFoiaOYlx7Ow6z9ZiySu4HZQQbiV8ELYXzJOcX51BWt7RnNlpYrksAia48Phc8x/
bCDjK7Iq/0i+Zfoz989+LZaXzBypbkjjZVgRmhQiOXuIWkqQMA1vqGZ8LP+e0hNIsJSK7Fgkbt8u
FZPT13XhuRfgPlx4A6MLrGhzCnTiGvCgMyFdUY2PHlVpg5Kn/fihi1a+kDUjWRUqautRMgMyi7f5
j6+RwrwOUGSiQwr4Gua09+TFTOEtwXzdK9TRplxsnEG26w8841V/L+6SrVtLvJTS+tTATIfWSSut
6cdT1ix18DuZxhRDw+ClbXBAKqmB45dobdjrTZuI4jypei1L9SpznOoSrF7ZqoUrwtbbqoKNbI5c
mTd4stJbE6vlqejPoj8R6DL0LT95D/dKEmgi8mHf9Hv5yCzO4yAvz3FTH5/Ijk54bMD4KJLByAKt
75cnzrYkamnYIr+Tr9FJl0w1NL3igVHdZmKr84wvoIaBdqAWuh51MKVeWnjrW5+qbzP8OBi1RLA5
x3/18BoypPSZGyjKmVodk5diALmLRQsP3EjmWY7mwytT4kK/LmHgYqgPCR6fsWI5x7FinvN5yQt7
w/wVNUkQjXqQEwnC5qLw5bqAnshqqsRh1V0VJVCZ18W91FYvAA7rs2T7jq8uiOXzmLeuuWnj4Pru
aj29cOSVmk18i9fhEJl/XZInrROQ+30e5RxOYwEZ2aCv4LqjUOXhdpv+EXAyXo8gXAWHlH3HTWrZ
IlXDud+dizUcZQPf0uK3MnBqoq5hvjWDPOzcfVqG3z8pFUIFTES2MjRigMsblMskHA58Mb0Sbnuo
J69TQRaBBWYqxEaS7H4uxYP6HWCfrL3FCbYV2iWg1ZOBtToacvp4vXCG0OmB/4fEdM3/GkRX0C7p
hR2zF8gJEutIhQ6/7+8OgNlu0O0AaEMiEAkvAjmU1MKrQuGN0mr+UCd/Q8oT3FCjtr7Xv3ClDaMt
ZVyBaYR8hn04KTvSKto0mIxUMbsTyp/rp04qeQRN8JpWF7QitKjdHmzdtLt36WcfmWdW9rYo12OL
+AoxtyfVGphKJew/8TaNydNdIOC1ES9x65lelPQzKChu/gyEWKWKuFD/Y/2VU23Ac8lf/P1/hKMC
7KoxFPCZmjexE1seYk/4LLANsBgeOOUMVrcJlLfELqovIwyXVgDUkVHnEgABvmtKbLWhSXagFuNm
huyJmBMm1l7ejOOod2wWc1W73302Lm5M3oxlWwM1ti2tTDtKcWrdlxa2NsRSmLnnxGNf2Xp5id5x
BLVasEVcHtwhVfAWQrP6yIWiaWBbVG2EjjGnJCB9JIaBCHDvNWuRbw8qkOO+1lUxSICICt8BJZe5
JgSA7ZA/nsZ+yipPbebEFJ//28lB6wkS2Dv1bFhlI42g99VMC2rg7PU2h+Z+T3Ftz+bNSMuuRIfT
2IoiCSQK9dqBcCJSKpjSx3alI8rYIBPBbLQiScY5ACvEBcOYXReB/ugTOOAbyaKoFfyROhQeYnIk
YRSGj+lkizckwjmAmy12MeOU0oa6YqPL9s5iZ3QFARAuWxwAbuT03ERvB3owWmcOlH+4qivntsv3
jEXOhp13Z67UwtmQGFqyX6SD5FhsKMVg/Gm/SYBQWC74ea6M0qOL/rW5UndYECQIyWCmzPV8CMR0
bRcg805OW5pWctx5nGHP6ZqnELaRfJiC32Jz1m1hU071W521zly0usKnbN3Q485Qhleoe4o/0ENT
ioe66PdO7I5vSh5X7VoQWVbLBNb4nkUvdvdp9fok4fYcgiKAngG/auM+rqupuD/alSBd2HtS24Kc
0GC/vIHG0FvhIUXXQexFh40xRku4jaoHug7JgTWF/fPYntuZiB1M5pCbV53Kjb9kCgIXtz6l6IT6
wNKeGkB4droY/1jZljNcY7B6vaan7wM3si+nsDm7OwyGMKo4cH3E/JxFC5AB/o/FEwlKrUdkOc4N
WY8l+Vuya84XYk/yQdvuycLBusk3Kzhf4Iqffevq7fqCJjye7411x9PQMHJsJ5Rz890gJ9iRFDBL
h3qQM/Nf4dZ9YNq2EGrwc27KDpkZdB3U/wsf+I7pYcHthRpHzFs+cKMbnbW883zJH9Nyzqf2RZrR
hNig7AMQQDCR33eZiETVGN4mkME6TmAVKzqVoMEzUYJQP9XqkrtVH21uWYmB9CQOLDYzDz6Z7lsp
EOrc3ymBY0+1/qpKBRVkm2vH6aRfK4YozsqhBX1qayvl9eZ1Z1RTHCzuG3xq9bHHl+1mPMTX6OZw
Hs+mC14WdaIUQxekxXzqd+DOYHc9RlI1RKmVjq176+8uAJdX6gjKXj5gSG+roVcJboyYk+C8m/F8
WKUTvHyeg15b42x6whSgw9drF1l8+4qlXRqE9mpSO6Q0fy7wEmX8SDF/k/PUGOMuOWYNzIHFUiuS
KG7KRsPs1iaY2cDvIJEVr/NLEiF89KVgdkX28uNfV6afCULXrK0vpQSY+5DgxyNiY7IEq5qmEKo9
6PTIRJH/AKRdxzErPGkYjD6/Wg9OIvYQDRTSvcC/YWsk/EYRsp+Afcw3m8jPrQr0nXz/alN3cMxc
xiYKRyh3ErjYXiA+42wakbvVmJr7jxOCugWa0EUDy272N/P2UneHlf8exSlUqMF30YBE1FR+d/Gz
jZiwf+kMtmRFmGKw3P3Gnmy3NPXCdoEiWGZNImTDhhUKnvZsqgpaI7jAtf9kUbAzmbw/wkQ3ntLX
cDcrE0q44rr+vIP4SkSdF2IVg5jzxpiY6eVvcF0GSoLbZq0DWjL0ZStRVFZaOqkihgBBxq/k2EQ2
j4anmiHGcvtQbCHtN0r0No0u5KAGAgglAWva5eWGhzXq40LhKuXNVQONUBwpDb7LA7bN5qFGZcHk
7aTzZcTzjVRIRBsjE5cDLCGijP+MY5/9mOt9BNP41Q0oeEgfbz2FDaE52nJp5JgirFBxYC2yo84P
RBq617jbNgyzkDv6WUe7UKq0L2kMw4ten92+mwdDAOWiCXQkMu6nTdAr9rXSpr55BHnCpbWdWZLl
qzC7ka0fe/tsRtcd0h4YAeXaMyTZy9zq7RreS7o+C+NYXHFMfcdBLlIwpsi5Eb9B/QRqw2V9Yn/M
9LVCjqZ0XRwCi3/G2Dw6iWqMEr9xEUNCxL6WC3CVdTJw6B8cyiB5IByEIxqBXHRd4t+ldAAmMKaf
0sY3ll3hCG/5oi7TBYOp2vWzxnzh8aTV+/a4vOGQy/5R8K3rWF3/NE4pVhYHtkLBuYJzc+l+P28x
hW75Uv6mHWPDo4MEXNbpj+8o2sdBBmaVJVzad+8yNHeA5Lz3DB9pz5eC3yvfDy1aa9jvW5gSj3Vf
uLR8JZXjDJpPCUpJfVC00eF8RIYQ8Ede4Dhk3idf6FfwG0FAYyTBWYyXwyk16ShUx5n6xWz6ekgY
8Idf+DdUOwHzevS7SsMcf5dCTssy7rGxzOiAGY3t3pwtQVYTwjS42vFOZD76m87CY65TZWhmC4nT
7fjzI1+XC360uct4h8/5cD4uJjvCV7zYXnKdN1PQSpOwQv9x+J3v4yAQ5syGYDGlNYdEt7uG5QyF
5nlhGoWrELx88k6UlAw+UyjsS/eZ4EVq17NVpHR2HENnUzna13nCzRKzMMtumVUCeMtxpXNBjIbP
alihDX6YpOTomdmg1EVc8FMV41LCImEow1f4Dq6hpXE3eAF5GEv0gCtePjcVajrOQSNGJpe2HhUB
4ZbOpkKCawWUdp33Sy4NV4EMNCFTFV0ONUBrgagJsnNK25yYMcoYwQzbczuVlrmIONIoEKEJO985
Q4Fwh+vHL4mQCJxJwy+YJa2wwFhyyTupuER4mnGH73YlRM5TTWUwOvBdhAU37MTr3bEpdW4XMbQG
AI2ywBm5WRXQwO1UoscF/aYdWipMguvo1V/N0+KMD9mPNEZmPxn9q6Hti6VSXIOSoNi0G5JY+23n
DauV/vXdKx29bv0oHa9VcesTJTL6rRXNXJAtKKp+jTtHEAW1cYjUymDVjIixm3xS1bbvikY6C6WB
zfCJO7Kwbzw0WZkWzjujv5Qt6v6GsniVTPmpJWHhGvOEsCmIXdncTXZ4+c+S79vAngn5LEUtF0z1
bXHNVcX+F/29e5A3TfdN6YCTQa2VfyxJBcHPQCsIyj8Y7VFVdTAU3HFgwm1+SDTPCkh+tJpZL6mq
pefR4LFsSycHu0t96BhBAv0Ww5UQY2HmVbkofD26nXTbsaK0AhewpvHLpilzaEkArDyucbgTfiYN
PnK3epT9Wa07i3NXjpqnRwdM7fdDwKotmVyNYtWEojeVs4u293sPAtRPj3aoPMxRrlcE13/aFXRr
wC/0ZewiIuS1s4n30cZSI5wUw9ojy6b3sPLD55m2yUe9LtY48Dw9VAbbrhhqMy4ToOCntld735Bj
4tW/DIRV6rajor3ZHccLFVbFT4xrkeDgmCG7v8GyB3oAIVgUM4ZwGa98pruI++rsLNnpIDTC7Ufu
rD04zxJAxB8Z+usNbHN5+Dgdk9tdtxoP1gN9R89dT3xs0VLZbZ9J3NEYYbhjuLk62RgI9FPDAcDd
wIdskME6/inAxDabDuIoWGVVdbFIqLain2P7Az9hV1EDw4grpj0c3jJZsdi39Ru/OEcmi/AqLLC2
wuKuguwwXoR27/Qe8R2I+rQy3t07M/oQte66lbGfFkfLcZmZpRbhBLie7N8RHIA2OD35LkY6URIs
Em1cZPlt7Y5oED5HFfqSHKYh8dikhBvZC8Rv/6MgCl9h3ajNdZHldxQf1uLcAw3OWzG92T+9dEgJ
ffwHz61SHxt2LgG9cqSJrm8o/I+An3Q5UsP0hyyCe41OJndCSn73Hkj0lZzzZxdd0LvZHwcQd+dG
V+lfwya6TpIQCcIQEsxXbmNgurSbs8vlA4Cgoij3gtcIrWfDjD69vONzhxnKW2tjoAmm6xaFyADE
fRDl6udOFsFzw7FBpU4iVX+B7bSSVtvLfdBr4a5n8b9g4oH34eoQmpcodIp0PND3EV57jwtuMvOn
uqRKowaY2XmmFmm5GggUFY2ubmTIloC5vH4ErmLxr/+6d4BoccidpOSgHPeiy2r2Nr0Nz5zNMffn
Mg+3OCuYdKPSzUXdx5d1ThlbOUr2/JTWDeHZ6uTtrBD7UWFnzS8dWbnyeSwdHFQ3vHRxdhq0DKoa
8z58A86IHjb90Vw/iRWX8tHdtYi8hr67j8fibPgDYSHguyoUHy3AXQ/qv1/blNUBiNbqft+mMhJU
E6AawVip1Pp+ShSuMWnYl2lYrw2XrWO6NUgLbr4+LHwpkKYShuC5zmu+8vbpxT1oZ0PyjkD3YLpM
25bsiKEAtCmX9CSwioIzwYoGcraVgEaB5+A2Yfam72oK+8X4GJImDPQAM5bojhMOFpCpgEcCdGpp
+y9pCeDqjzK3zL1gT729Yyuy8oqh2BnEZjcN51yOtfwLDEwLKIg8UWdDwzxBs89fvWzG2j50fUcZ
1UWZ98Mlq8MTdlrBxh6pDNZfLcLkFjukcLmOeCTj0rpRXzhli/MgNWLwSi58gvpp3LUXOl3qxy9h
an81m6Wxya4bcVE5tTcqUAGazVsFiq1qI5X7hlGN8Puduc9Xf5UbYbdGhk3tzyFb+22gQYoMTrHr
SYgUiS8+Jt+PsA5yebUrLjOCPENPdMQ2c0R1vhPYFR2KoJfYZ6XW+DL+elTkB4g/IRLdspE+I/xq
0fvN7fI41JvqzPS+iGu6wyrR12gZRdF3o970A5IWiqyzpa2BGhCk3QlK/+dkID3n2mRQyDCx9xTw
1Dt4lft4no66IkxxRvQhga1jRpRHv/Rej4YNv4Mw0FbjXY2PIJBhsu1FM/B89aQ2hs4lGytakede
iXwM9jWzSnzGQClFcikEQlMuxS27/ZDNAHQ3c6Dtt9aoiWgZwOarkF3yGP5dVShU3ZGH0lrnUN/2
VzZb4iwpdhyoc+8NNaDd0jKUBujF08bxFJiq9HSwqdLFCCeCFzBxxf5X1wtWBTv0y65TaufEI+kQ
Be6f66xUiWnQ65dGRRQujGwKGerKTaGiVbvuBeTBclu5JN4RytonGkNnqDXPFHsSZlay5VeK6ihp
mrsDtBlnNI4TGLdZdzBbtLkiHVxLItGg2QilvP2WVQ1470jx5NfAc3qXxmg75Y0jCWS2qF03aMR8
o06cfJLIBBQh++Sc6SgTkd20PTAc8Xg2ZkaRgE/FJvtrpXG7jdH6PmfsdNyZ1oEBCiYJLRPwELF8
Jxud/9GRFRKwGMZ96G3D2chQGZUcMedalZFV7WX+ITikRkhJwHn8MJ5hNNqXh0nJioLC5BOFLicD
uBSJmzgatjICyoLUfGVelQIGwxWfLfG+dlsJnZdm4+O9sSBJCC9QKZzxkCeoXNBGlU/7e+2mSWfT
fAUjUK9vDolg6t1ZGxOCmTmf8FXCkQU4CiymjqJT5I8WdvACobNE7io1Vdef0xTMdMDrA4U55Nz9
3DajxX0VZIq39fK4dahEGPafGAWL8noFy8BNERAJXn9J6lBCFMvyToPvmhYrsmgCVVMo4CvdRXe+
xkyMuS8fuwxwPr+0IVYByZpDARxf3rFeh53KfpjpnHZLrE6aaiJgehN7WgL8Ulnys1v19E5f0nn6
KKi2dERWGGf+mqdykX1OCA/gOXSsKdBHudqX/FfTHpFR7n3zuiHKWV1numvDiBdalAP2kBKveODf
v/xnx2vD2vafjc94f93YBS8sykzWNW0D2ezb7qhamfW0U8+WtucHKJXEV7E5ArPp/1pQPnUai0s9
jqg8YDE0wA8xdjOdajtNpGLTU0nYbT8lXEYH1j5cVW8U1e/UKQWgnqKO16wP9tmu0rbi2JMcfAcD
6NR42xRymJ5RRb6J6S93vl1WADqWn+HCAl+6bPWH0HdCerJ1Qf9po48tdwjw6VjV9/GEbD2egRMS
52JyXVcHYoEIGQpeme4yRJ5mNaANHv1ldTaVfoSHOdoFiWYGHHNnt2s/mbxDYBcGktliapPNJn6Z
xQX8TNyWVM9f0Yb20ENRES354RA7X6eg5jDtiGg5MR/xTjPADk+11lnBygWoaC6VLK7yrptUn6vK
Ty3ebEa4DrY3sEyfaQtBYqZktx6ZJVEWWKgmtqTgZJDuXJZ8nolOmpUhqFU0JJYgPPz6dVtY2Hd4
aiBX4jcT4jWvlwevF10FykTRiN1zhqewvXNlwc+ly2k3iIBZsUYgVgsWyzNLGeq51ErMBcU16jAM
DMXKF9fS1iM7ADoiN5N2BgNJ9wZcAfGNO8bunCVZQaJTkxRt9O/yxqluXHJCJwp6xcR2TDdUIi0i
G35YyPDS7QvkHHccXPnpN/UdD7YPCIGAmvTp00TbXoNUaqeJtRjvDSujp4H4mLzByGiRIxdHG5/j
8qdn9kdMN0/0c9+gB1gh+vl6SuTXsregDcXx0fcN5O0KrjRmkOVHTcoqbClE3P76Yfwn7zP5TZgF
f4oyM1hAQxMY1i1elnDk/I0CkQWFu4gZgbV7J3CsPD/29DX6X7HxNKj0w3c6anL6mgw/vHFVHAAB
SUxrqJeeTT3MuNpqU8q7x03A8Qw9+GERcXrk68FzzTLVRsQLOtSPdQNg198RGfjAgISTzd7Iz2Uj
jsPb0hHRM1hHQkw3sOpKETDVMe0/EvMHxzRo9qTsst0cBfmQgQ/+mObKEzNmPKSllAhV75wT6qvG
UNWDVGPrDPSJZlSdCbeRzPHpmchSGAH7DPwY6WTpBNnmpmgIEZowgMwnNFk4zvW2E4BaC4GU1pbe
S3h8KGjH6i5y+6ufoEIourDN/I+Bajr+K6r3K9Q+P0fMfVejx+XM1RutkzV/pjxGbRbcH7RipuiA
Zi6XdasjzaC5y4iJ6/Dw5e+uMkfLvhExq6BF/Fr63usvgcjf0jqX1jPebyrPxL7Agq/EfH/YkOsM
R9A2bcB+YgPuP0coq8aLcoXs7EYJQvtFCAUHz1lyJpwu1V85AFaiHOa5NsNPMAUR3g3UVqJWeWNL
+WVrV8UzqCnexEQ7vvV4p2ZUiniw1hImpUT8Lu+XWY5vFxcDWc4J+SBLJf5BywouWEHHM8puFU3o
2uCD2vHXSAyyjUIfldkYsNOlUgPV2RWdbRguer5mHkwRSrLqxpOjNBZt0aCyTsSXjQlIQvV1zZpV
OqLpEaKgniwaR/SMD4YDGFeLhh5/E51AXaHs6TxZZEjXFeN5CJCiatyrzBHdWvnY+EFYQ6XEuqdQ
rk/WqnDTQNrBQKehO2BknU0Q9kq8e3vojp/lb2IP/uZiGyvKCb2P8gyOaI/LS8r1EBrONAdTP/Ls
LGZmXGaWGquTrkIaYhsR/EsvmO85QEU6Vrta6rJJCadRaa7FeZXjLGTGy7heqQBj8iAjwksyaCni
1DqKtyym6bJUfw6HMHaCLrbjUWE3I4XHTT3KEsWM2TL7g7Kl3bN/yjKIz2di7X/fRDarWpnYcUIT
yXts1rrIY398dUYDJ+Q4LHf2s+SkDsAA6oFc7QIo7LAcgxvAWN1j5f462ZIaYaOYIvb7wJVEi1Zj
vTKSur6hcAnZEiZttt1tti0ymEoCi71yM0EUZjsnoeOoFv6pHzUWxivF+1oLt871u1XYPjq+xhnd
J8URl0HaDM0shyxQlX5Q8w0Uqy6jiGqedskX7dJinx4Jo3I3cl3siN7uerxQethsizhLyvj0fdfV
OVGKkPvUI1VXE1XNWb3nS8rKgSGeSkEvFV0jKySSO6jwANBkVdjt/bCmJl27ZGX8G4ojCRoWrg2z
SdtzuoT1SiOTpCG+xbjnfMZiJmwatvvW8wPvGM1omqsyK7UIAwpQnN0mDAwcyULeQB1olSFdUORN
H+MtxnO5SxQKTGAeUXMIOqdkLHTiLjiSNS0O9LclYCvNXDHexVV6Lwv6ve2rfsy8XI1pbFj2SH0E
RuZrQMqiYgTiFLD4E2iJv1mkjYjX7RqBwOW9tQ1xBw2mlTh+R/Xp6WopjtUC6kYYXpRThLRsipnz
dbdGuUwPvSi/YNLyQGDpp1ppKi7G1bZlPoaT1k/HlzkdUCZRq31tYHeBG/hf7Tc4mWDq102CO5ox
RRh1t5Dk0qtJiARYd6mlvPh6YxQWhcT0unYOfXWnuB4DeRxgh2YTK0ogzjNgWw3P+0Vj8HShrhOY
3pofP+yDA9Tg4vJHgMkqOgsRRTVfl3ZsUZRvp/gvNPTdo05V2lqA7Rh/7GV7XiQc5U7ykH3sGdph
dHVBLlMLxyV0HXRiT5Tnx+2CLTBsrIDYffdqMIEpbKkvY8KwHtNIfDXGzRn6XVeooUU5AMf0tGfM
buFv6ZS7QBgNeDKQ/bOa6VRfDMbwCzFjBsV5k+An3mx3619o33BtqWsHDyFiimo303Vu/JDuQklc
Caiii7b3XZlHMpOYuh+zPhTzgJwuhhaposw12zMdnuoT1czKlZSbQuQV4fi7TYYGPgQG6btLJZUw
Xpj2hDMTWopxRJuwPGF8Vp/O+9Pu+PJUkHFiQc6b03za3sPokpNo3SD8TCmDvRit98bg0tmVfoh9
H0NOnb24Hg2Wk3CiZAS9939xXuxf20/2dnBTv6K8VbsH48+GzHitkxhUSUz1p78GRpdsI1V0T920
zc0nyzlteG7cjCSIuywG9DEkVRVJkgVYhz3ZcKvwsS9d22cNs+Tylyou+fxKt/Hw20yBEOz4eZjd
8e6fogIebTC/ZqKgiKS9YEGL3mYO8xXK/xkcYTNf9EU6YKSub2j1lFG4NsxJkGj85m/ZbfWhE6C3
QFD7amW/mFT/zYtmTNOKNLAIhiZMcRE6ut9nVfNo6qg1JLsz+79n7jHDw5JeDysEoe641IA3nBI7
Gh+rfs6FB58X2xrmKXzdQk6WD3M6dMy6X3MfBPeJ2188F6SQ64E4Acf1hpD6vRh/1Pw/ApIUnPQH
zqdhvKCI3x5k3WGKkwzwVqYhBpDOMS5BjDuugRA2rE/AWSVwbNnYc6X/rJxp2HOTYSO528vieMsQ
Ubi7oCvb4usdKtPkA7kF9ehU4yKflruEm14owbXboSK/bFOgMH7JJHHEnwkhd/knPEyC4M5aDSby
S/0+JOnNhnBDl2n/Tc84CPAPZjvlxnIQTgfpF5IMgR+aeshgc+aDqx3h0zQdA+Tx3XnLTRjDgwEe
mzzdNO3O702U/oVcy458KvEHySamrnE4V6z1r7QDGPwAM8GYUGj6t9xgfc4LzjbpBlJYQ7mxHV4T
CHeoUX0hbzlnxHoP2rWfTcGZCKhPWi1A3t/dpmPNkU8NmOMhaoblyVHgsHJEVsgA5Oxp8vv4Td5N
avRiaNa4QPNwWLGjmpRhZn0vOi7z+SUyXC5/8908yELzf32rPWr/ICzCdSsZhyvOHGdZsN/2Yxey
67ixK1fXa1XfbHW0MXO9s0lnt7KBEYuBjJvsf8ce4NrPnQkiUWI8CO99vjnYb6tvbNpm2muxE7uE
owrTPYQ2cpcRUinfuHfeO3/HQDVMRVATMcbgT9CPqP7lvpyojQFjBqcutf2oz0h3Lj13hA5LGCa8
jJL2WiGc3zJctEv2L7nb9nacxEG6wzT8qFgPMzOGJ/yhrYN6IEpbsSR/g/ufjwS5fCXxiktgML4L
vy07tMa/k8e133Ep0/uxAUB9MY4h44yYirCvqGoTw0qdNhbUCEOWw62uyB+RwoX40vxkEtkzkRkR
sS+T8u5YMIY5waZ0MC8mh7K0DO8+x8uYvInYKmUvuh1kAJd6qLpyfg3uSi8nwp8++st9cCOT0XBx
hBp9QrjAf5hQ02oFNfbwrkDmASve6ExxXGRCEwXJ+0SvfsrExmTALCEe6tBsvFLRviHe7KMPItSf
Vo4iGaCZ2bXAUmfKgmKUhOBgRXefNgogTIsTP+UQn6qDdPuJHEusUGs7AtXfP2X18rSLLO5fSbTS
kfhyZbUEF6PJS2dc2R4VWpBQu6A22ervv+W5H61bf037GmnaWffdcoZaZq3hUxB/6Ph1SsDoPtLj
TREyymR1EO5tWI4cqpTNNejWMk+cbengLxJoHoBASdDdT5WhkZR7CRH3yuz2vQOcZ3sTJSY2X3yK
rOIh0csuYXcWbcqlMlFtVQ63KXcczAg8ehu9Dh8jqgkkP4snKfHsrHgTBSYcOC9vdXC5pp52Po/f
1FKPmw6k9i9IMLMSqC11rcZt+gaSHp8exx9VjpHovol59JZwTPGYD/AP70AlApfrwbecmzXs6Gh1
tw4CSTYhluUHNS8XL2mAFDNe/+PFkLs3FC+JDoZ45ftVXpUkrzT6QiHEFP1pfULxB3epQ74wB0jx
YPt5w2PA61TsVAHgCUsY1c+Vm9dIRMTgLRkSaInMq4oi/Y4uVyjZ+Zc+joySrlFvrgBhCrZJKyUS
7SEb5yqz/imF960lr0bx6YDj5mdhZfD3tDogXSvOAFzVTBYjw5xjT1UwIA6X0vfdRYfZ2ZL2HH2d
CAah6Mw/EY5yDb91ThvBL6tll1hf7PgpLXsfg7GMnhsnXPydcMzIkAjuO7iDtjkiVM2cTIWJjMtO
ngegHCONmL31c2fvFtuwrzC2fUc8K4h6j7JRfOhIJiFOo8e8SlKvOnDM52/jQKEacJ2NQGSDyooC
8pLWMK6RfYfX0yyQekJ8M7HdLv0aLpcHl75KD9RWzsztzEpGBqZQkvioeQVh+xWPqRtAD6BYcZM0
ZlqpQd1eEImNUF+xKF8rp1RnV+6Dg9A7kx4jHsToXwcrz57h9SyjxkzfGoQYO28mWvvwwGlDo24x
TB+b+JgDSSCJkAZOTc2az+A5sTZp7e+v3uk05dPqOGQjB4PiyrNSxRsUaS/IhLHBVYedbIHczQWT
JjrF786fjN7bp2Qf2WD44vJNZpFxqVyYBy2ie8Sh80/3twgOj9qR3e0hEV2mxwGAqc/U/lgtoW09
QfUgpCOFy+nhCNFHT84YeeTzfAamjcg5SPjd5DGMPLeVPUJR2nU+MS27qqqoLuL9g3JRuf1X9CNW
U7+FNQJaPDzM0g9vF+gHH7xDUa5iglTv0QhaMBPsWp/oxAL9+WOFH1xXwpHwHFYzSfI3eGmiFZNE
E+FUZcmbREfyvw5/60Iy62FvgLiQPCQQU1KeEw/LhfHr0d9clVX01kboWFfhT29WReEIETCm8RNt
QZrkatU/92s9A8YFp19g2JE0QZl+gVUkw/xhXqlHvUxczRgStqgycobgHIGBvlXLEGtphsFeHPwt
tyx3DEui5+DxtkFNb5xZ5ysZ1p+chrMpgpac2WNW9QXJRc58TYgT8XK1ie/1FtCln8JptjH0gxu2
oj57hfPf7rQAXxZoNBLBwurdHrfmsaN5qkllBB+/fWgAn85jXRrBaVRadro+xiygA1z7T2TbUUom
ccQZ2M24+vWDZ/hQVRzaGSUBwADr9hQtBRFrLHa7zLpMByaQsoObjaLv2zDIw47mBZM2qmKKFWBo
dqH/1jL/YD254SsxW6oQbOIreGanEREsD0c1mxutnDOPaearCEo9goYdBu11nYqUG+dMM9zyKP72
pdR9YehRRyuW93kBB8VrQpOFMubObg2LUdYupIv+fV3JbEH9rMNaml3R7KUrS4Z9LYIn/crGZY3O
9bT1yAqBfcvuXMTgHbkqHrq9utMHs1u+2lp8LebptlFK4tWJSynqYG4mgt208gI1IVimxe0fIIS3
gpJZNS3HmnXP4Iq03PF4ee6Vdce7YhOXzj+8QX6kQgAxRkIRnxxl8Ushx0fthc65nIP5LnkeYXTF
hKHphhY19yzeqY5Zu39ue/loDtG0MWFWrs4s81anrEKw+GPK3ImYau4S5JV7zHJxW4YjxW765WS4
aBYTe6zjWPMVu1/7ShpG850BIE8SDsHYQnWJ9PE4fwVuJL9cRAHMND9LC9j6Qkse/Kn29wU2+G5S
9TmiO/9R/UmNJNHnEpJ4eeSMT0ZLHWI/HiQfIHIpBJatbu7tW0jiLFUoHNeA1Le8ERYLx2KDoxy+
XMAvlq9KQnBrC+p9MJGi00OCz/LjEUo1f9iwdhnkt6aWTronZ8Rw+H0WGxjZUKh3GeaZ7pWMsqts
NGeN5mln/vA7nZtuZf4UsfzjlrnTsMfB6vWNihRT97bdSBDOYdRGPxOTYRkSIdATR7Mm3TGc++vE
/JU1FWDf5p6nK90KJGa7TaXB39wH10UvN5D5cDjV25N5btIbKoiPeZRNnrtmYMnY/Xww6rVIz+PJ
qS6oOu48ydEM0M/FCTvs72VbwkXBfrcm2+qX2dEV4hPYnaOUCQ4N7W1GYA4KTFeCZ+YFaXpZFOUM
YlvUCTnCiPmXp3mTZm+kopprLjC5Tv+DP1jnSCL4hpXTKSsW2OcYTzEwGD3geutfUgZ8fMO8ZT6b
z6BTUMJeOx15zeawxiMR1VOz0WHrv0gGt7c5lGYMgTUadTR0OcQr5tFLAV2hingL+LhGWDaaCvLw
sC3S5mXlZIkOrN7C/mH+S/1pVa7t1ofrfdlTEAn5iJcFOvpiERLicErUY70b/MuagZJFAYSgpNjT
OThUgUUbfAuM/huxziTJt59qONsxZbjzO4G7MvF6lAeVQXes3vF9Uoth7ocRNWDo11/FcGxuyW7F
iXX9IjAUpnCwNt0JHDAYHewCyV7vtRgLwP0+FXymhmE16nmPVjj8dxcNrp/jQIU3RtWV1d62Iziu
T1R49P6mcGvSIv0Q/L3uEe9tOR/xMSvtyhKluKvGikmNTy+QN5YYgdslIh2sltxfQbexiM5GahrV
ok6CpO9xd0tHEDQYt9xMvC5dFJtG9ILrpFr140jFViycOHQuwS1kP5wpgK4th9KevWjFq9776rOz
KaF793XhjFqnl1HkIRDFLg4dvPymGzy8nyVNleLZI0UcmmEYNX8E1eBTxAI3tBbQtLd1EI2wtHpU
svnnoSs9TjsDHI7A+Jg3qfzFt/pmh3g+Vn66PLE2Hs5uvIyU4GeCzz4/pcZliAONODzK4ohIZrvN
A9d3YMb17mj5U4MWOzd7xv350PTRd7KpjSQeTlDIvZ7BHTk+G7AUKRo7MJ6/s0ItjWiH3qiZtUPq
vKUi4dd1obmqngwFEB9htJBEp/UhfImnCF1H74Xlv17ttGSuJygJjZ02u3AQN75rOpXFhfJMVd2e
vhOf9Cze3clePAyPKLeP1qIkuPfGOaP88s7n/nEIx0szc0q6QfS4iOZa/HxB1kwhbhFZKFBhh6qi
di5eHtQpDiTvqDqi6ZIT+7ePzLdmooojqixPIkkEKbYChKrxG0urmUq+tabzeJHEfaKXpwZ2t8FQ
l5cvm4e1lkfr7QVBL74L8ApTroRiecM4CzC+utctTDQMwMJllkq8ELEj5HQ+9sQCSxpbYKa0LfcO
fqgwpMvb2t8GJvCTk4L8+2duPQwb9IlVOBGgqpLRYQWBfsn4bClSzZU68xXy4JTKOhKS3uS6VoPC
4DmuWbqr19fvLoeAeaCll4MFMkQr2JR/S0ENyVzR9X3Ixnx9I6ibHghuDRtCfIT3ONCTmQA0HuRQ
8fcxD2js0568WXbj9zCIFsj8kjVXQ7P/6M1aPzGbQeBw/sV6F3ytv/bdP8UM/awOtZzd53P2euFa
9eTrjdfKd2pSf4GmKQRvpufCJhH8BD4Sw+nm1TeXYC7SDBUDPcmvKj5AOb11LtEElZqejgjEprJ8
Hw+eM2YoCBcviPAHNMmmwA2cJ2PuzTfHpeto1m5ka93h1KI1cIhilT3YiIWnd+bQC4T+qTX9BJzw
H/7YtZ5jsPu4JRvEp+TcN3DeRLON7dx7mn8MdV1SbyT71FaQokTsN6vTMOQK4Rh7UZER0K/LqyFA
ckjTvrVfRA3ocaXHimgd8rRFPqT2uSSW6XqeF/W42Z5XtgN8YDoQXInp8dAEoPwQA1055ftcN+R7
Md62zqIq70cpKPxlUJsSepE2ZWw0TmaTj9EvW/McV0Iw804wY1Ni8u1TsJ7C1QZNrBjMVtFaXUNW
aAxDA0TuZOMVhprXSffzRkR8lFr3R+/deWwulSj2mKE1KtPbXI67qM5IGwu1zQKq6Rsy6jL4niCU
o1Q+Ux7p4lNeRWBu1VLvlClk0h/dHZHWgg1dS/D36lY6fdxQk+LcJUgh7pQE7lw1UjY2WSWq6g6q
XQfG74RAGamF8xidWHRiRndoJcv+9I4Eut3bVgtNN9V8djmVzldDO2fqCNMtjrVyD3lx/PvYNZpI
HdjtX0w+6mG7+XbuvSLJUA3jHnCU7Dr5SllUZxsDxl8Vw+NwRohxyvz7q2faXG2yKf6sbYTZ1XWA
Uvfhvll2JcnJBOo7wvYxJUFYKFGPxhAVEx6x9pJOl4YO05S9pOqAiOLCkOOjNJBrV6YT/xGV8JLm
QTVary4syHs5y2+uU9S32MoCGzAFM/1mW+iJle8EmLn/mtkA88z+vObH1aMMlXbuUmgbEPOPdFCK
gWBYcGE8Fz/EyvN90oPzoPeGj+wXFNtZB9/8AlIHXa48ly9RnVuZWAFQW7YVFUF6KgNZ+L66oMPp
jAbWW4nuhY0iazj82ST2HsDkIey2nCl5XR7BDri0FnOyLb69/6MO/i3h6VMCwD6h+PIybqXLJfbh
csABqPoP4myjxhgXrmImJ9PIMCZHBV5EpQXgl8UMPA4zpN21pGi1VoVHuuHYyCOsK6SbfB9LI5wm
RuA0ul9iU/WIz/9cfx9NB3tm619KI0Yog2wyu4d9yZZjlUNZSr75CrEwOKeBxVDvIJQf757fJPF3
gg6SLB55DM0PmnWiDKAj/SmEnyVJyZR2oAhV+jGD3cOiq3y4GCiOHarjpS5zjsi4ET2UmYoTzD9w
jQH1dZRqSIF8HjVKCkhcmJUQ+HUndDsmRfXv3PLX4E9VcOG/LDShQivasQzyZ5rxDzqYannjZbiw
ItrgTrwBfbn4AzKj9zgC0j6y8sFHvL43clSGncGECGH/mtY56na5kuPhqgHsNwAH1vY5Rn0HYhGe
f53J0JW6NzjJJBCpjLeY+9zr//LHh+VFJ4VsnDlhZvHkWnXvvRV/KXHtkOOhRx0ue9IisoDp0J9O
cTkizgdj5UJhpAHmxAgImjJQu6tv65+gi9ldWzf0lk27dH0Hx0ZqmtGokK1iVmCPeNcFTBM5E+no
fXD9zkIwijxPA/INhnIIeTKmwZXQ/kA7djA/h5KgpaX6bl/f0AzUl0548XhQuLe4s3StMeYkJYhH
QnV9q74HsoiCn40QqDsa2JzXgV24wGzM1hOpt8ZSqCpnaV8bnTqMKB2WuvRrVJWklHHclEGo/gIm
tpCbcizQRIbaEsSrAdbIoZLBHXpMhkAfiny0nQwdVbuidd1sfwLEFM2mi0X9n6xpdEAQqpZPfNLe
QA+KHCUe5mf2ZvL9xC4bvhizPKOcGZr5vUzplKEnA9su10GuzxVuY+Yx5/65XFzMzxr73+z3YERE
i7VnEx22y25gq9xt31G1bTWFP8vYgKiAXb5cbpPaX7lFcl4nyHZoxtMm2Muuf1L9iS2pmY2AjV9p
CSUwVQoA4TbVZwSpDgvU2ff5rhet6ZbKk/qv8BR6tIfh3M5o/pFr4oyS76QK8xJ4X9yabTq9MTSQ
Zn5gNC2q241jkTgMEV0rBR0xs90nBtp3FHPXsu5MLhkpUtJXnRJ1WsNojF9mAlGqtfHOytN+zZvA
f5O0t+Tglwl+cgeC2hnGfa41WJPZOOCm5QY+DoWtZouJRnDEa8AH+G8NEoKq5/PlO2csH87qUolC
XIOETmeYh0U2AE7Ltc7BTceVILKBOFhzmEkxcD/u+j/vv2rrjZwJGWNLJrAutp15FPOBdS7VwuKd
sL7KB+VLtofUNja4Fq8UNO73Ka2G+TeDnGV/w9HPwS4udJA1mLymsd3+lZYJeRcludAzLS8MiEpq
XsAP3w5V51VrIX7PdCAGayv4HkCKmb6Gg+6hFzowwj0UlKODos5kSRFzQRlfhMIgbEdyClJi7WCf
JebgvAuBTKDsGU5qkkDQUIVOQrfLVuMS3X5gOolseZKndzmDNDu09N8pecnmU770DLyl85+eO+8+
6PcHeAbO3dq5/JD0rJL+9/zu2ScqkcBcMmx2VC7Q37yHT6cczz2UUAn3ZrRPEirqNdi6MwG1DdRL
17p9gPBcgnSZe+a2nC5GHexL7v8XoL7kby3LZj6+P1oAoCciVuOtrVvYthXH0IoSFWfpnZrZVFAD
5MeLapjcZqWg1s6Mcz+TWEyF8J0JNlWAj8+0m/3wMd9R+3FSp0Em2fAv5DtbJCk42R+3aoK6aDpe
vl7upDbPixYpWPE75D7HtyF6sfv4CnX/MJKwaXQeFsIfFI0OsurCMxJ9xzbK5SlLcx0tM6yXJTZ1
gdM48vuwrxgfJVeHhCHeTxEJe30+pWobki3R/mQrvXscSU2XUkTuFbfQua9mu2o5RUkqV7W9a3rC
b849okLTUuXy5HW+XPwGaigvTKevD04eLN7xAD1+yim0ieuymRx09x+KZhjLsfWhYpkW4NsOIx9v
0URJllIlaheEjvSdR6lwdQhiTD/dA5VBqadN4ZJt2bxIYjyW3HtHc/I+OVvhHo+TiOh8KR3/Gwk6
+DFZpcO2EIx7l40AntGxT6oAKwAExVbrrhn93jLQox2WfV3GkcftKp+ZD+c0JS8T8yG0ShcbawQK
s6MdTRBGPvwW9MZxYVckS5TuV+LhJeNbdBq5qqwBcOmdM5NDI0+dmz2vDl++NBvyRVDc2oLdcKq5
eeGNLG6OzPoDbK/O7NLbNIru6XoPtJlo7AddWPLIuaLvBeW7mbUgiMJRgG1YG6nY3AhlipqSq+6e
/+uiYNOF0aaD0MtyqWd8vgZHyfMcXb6Facg3S4CQinOPiexelbanWvhkKlsM9IrAs9NW7Pf0UW0g
jeEQIMK/QjZ8B97cJtLnoUHxQSdDCTCGyDaBYOAxQD1gf0dvA8NHHY1MgPBJ5cX9o4KG2qfZ72Q+
XDzhp9d+U5RcGny+YpqMmlTsEtk6GoqWR+6yy+6+p0mmb1htn2SOOxjqQh1WuWMi1zzoYbT6V3aT
FG//e3ylJz8qmfV7/+CTkx0V+HBm2qzloGcGhLC2j9kwoF9TKS0uSQFk/BxpekxrEhukUSITMUzR
csgJ4lL+zgSc8ApMrC8mpJBHkVjHH17JkHVl7LR+Jw0xHOKT6FYRw+VGARwJCMM1h2uuOUjs4E/J
CYD02dOC13ah9wklnjJwaTutePN8+HQbmVhC93XYPQZ5TDf6//Xvxqoo/ijdF0g05zEcFO3aAFwS
NVudBMmYWzWf0RPxj9prBBl7YmaA7dhgrgfhcnBsHESjbvgVnUwTzBzcPqBnDC3ePwxSP3dXxKiU
nEa4LrnkpP+03Q7lUgDvvKjCldvDK1hO8gRwmkTw3N9pm2QJKlHGypIF1XmF6i5N3fFiVaWo22af
7fo/KbhJdPX7VvojU9kI+FbbVL3AM35290JJDJVdui+Pk07oC5keMt7KQbBL5lcVkDyoKqDQ1D1l
XvUl1FYY1hdjq49DT8Bb7T9rNwj04rECrBAQFiY16wHmBW0sTdcDOWrJ3zWbKwFLbrdbU89x7J5/
cFIrmrdRG+62wvhZ80+m6fq0WpAcDvILOdo0HF+PFSzeLeUAQTE4BvXHO3DRqgHioiIMrkUQv+tC
Iae3d6vzipYcpdvKMbs7hdXg+SFcdCrM9mYExgVY9KF5z28o/APSa3LrNr1qwjSY0GuLiCrdvaST
ceaVEoyXAehJQCpqtdHVenSkNl2u1ZlUhYxqgTesKOR0iABY6zd2EPWqzipIu68fNbG1FoaFge3A
RwSZgoZAPG/Yxc+b/x11wIthbDmf/uwxRJZsNVlKpKWialpuH0lzLuRBlgfBKoRnewBitNmatYQx
a+4vaLEoWEmSgGP+szs19R0zy8IwpjyAQ+QYIPAS5iqa3i5b4II/fKmHBTqzjMXkZKcqGxHIxrk2
zlBW1ZglAtdlQ+Rcs30ifbYo5iOw2TI5rQqQqp0xkhxnXb9j+7ySDnz4RpaCbe69kFfxkbedt87W
OATU/oRp81j/+9WOL1gqJVnJwpyvDvHbZGBtP86jKOy58QVHSCgGrWx+ILO+Jmd099IpLeeEcsAc
SEixiNdAx8ytQznSmC4+fCznxuYSlmKMyXeSlnPeDaaEro4wCxOVqcnpA6e4TRkHcnvVwpmbUH0f
Njh1B7MCR5meCBktapum8FzJA85lCGwtiyJb8WZRdk6fgva5yvvnJFJ7JgixZXvHmABLMud4vr1N
nj6WYzcQg3ZNfmW7EvVivmf+gltqOqY+mQBu684ka3vUoqERlw1b3KqYN2SDBlHLMOCYiMvln6Pf
7nweGaDRlK8fe0nw09NU/L0RnSygD0CpcDL9fKcFl31WtDFHr435sbZARDPTOZ1G8CNlrrFAu1ng
nk2nuSBRfYddziz9D/XhRwACPwpM1/Vx/1dDEW70Bg3rRmEt4ufMPdpsc8fgr6vgoTFUPVqXJ0an
TW7TJ4Z1meDuGgI1SGu625jXRX/AT8u2Lj/wAFk19nv/N4c+lZKMYlWZrUhvFkLWXbqochJ07YDN
L1ItrPyudWeyZGvcOAWYKHsGHHOb1HyGNVv27bNhyKv8LGfCxzYsoZwaFPOAagH3HsD1mpDFaW3U
32yIdnWt7m8BE8Adws4iesj64I9SS9zmmkYL5/ToonZrXR6OG9IhEMH0Zf5wZeSzBXTKB/7RrOOt
UF/3qZwv7Jp3WFIUtgGxC6/CVDK3DIo5StFvol52RPayIfNtgZGH23TTLMXTE3QopKZ9aW1Dcd4E
HYfiiUBAz9h7r1YvjIp68/FCkjr08o7LwLDWikUdfLzQYW8uZsXNBOtKplFVbTd+dlPMtiCsDpo3
0xP9KGzoEuc4Pvj/RGi3gAmC0Bdh+SczVJiwIwbQXnIY9IF2u1mVwRI1ZEYLSpkrBVCndQlx+pao
Yb1Z7XLYaMUJSLeHAYgkWe35Chofjxglqkrk/xqE5bIT3I1U3B4TJT0PAXeC4sANIa4rgmDqv3OG
c392tLefcnqi3iLsnf1ultevIR13DM0IhPrkMy6ETlz6nC7gTodSwrCbI1c9t806mvrRHPetJh1O
3hM6gfV3DgeQdm2nS2O+Ee0bmLRjjGyatrSCy0jSjdlk6EGHh/TBo0xfe911lOu8HoCnglBmuRXo
Q7IWSepvqKzkc0SRu2Lme2s5GX3eQQO6hJBfa6mLTpM/A6WOXLZUzXWOhRZVVUfOozxZGvAEu56R
ZB/ItAT03tFIHkKwAoQlHtIf01aspdLhk8n8WRF/tfPaCgi9V2r+ugU6IdSaOYh2FbsbTxO71noJ
T1S+zk/C9pMNjZs69ikoR1oZ/3Z8YtVSU8B6x7tE8lIxk1rEJlPWe2Ffb9RZmIL6P1YMm2Tg9TsO
uByfZWXHMaisaDwWgFaZkZin3SqEVhZmctqK7T6EZKeGCnWwzzYXipz5WcRIVTNe+fKKDrsEc97C
EgEBdZWeyySOvmQptOaLaskE0SXD3N+h6+o5+j2TQkGrCbAYpI0zvnI4r70efFUeJrTM4w7shPlc
Fr0IeWtu3CSzK1YQSm7Up3E4uQGxrBCqNMnL0CMH7HBTIIbY3tYvqp/5xZurtSKuvgwPWKf4HJlT
ll4XlrFnTDfX5YrTrm9Ej/izzwW+lMAuFjsM2ixZ8GT50n7wq+NCdqAnxnv41IvCEdNNx8D5JfYH
hG/ZIXdP3xZlQt8JgN53lN93yYJm8+hegkR14mllp5QbX72vhQNw7Q8xIjZ+LMn1auSwuMEnxYqk
wux1Dt328XCVuNwn+bi5k+ZewC8srqtUDeBF8WUYcOPpjGVFuOpICDlpABCXHoeNyCHB7Hw0Az2d
b9tp8fjrZ2vFgtZQYFZp758gqFqRxV23ZSZle6g9P0X2rH3DWTjYKgQERPWXZgsFljy9hTXd+AbU
WEeUI3GAcuw229s1zmucF1owkQpL5LbSo883c5+lKozFNdX3eU6BjKpjEiH3kAALiTXCXJFt14NU
vp3kYwdG53DtT0xqdcbPs/DNWnXpNG2hiy7D6CZapSdE0hpXalVRvH/kx0cTC4eVm49bx8YldbOG
+TAh5KhRKk/Q3KpOLF4Yz3fL2238i1WPD3JaqbUw2N2xVfjNB/0FzIYNBzPKSO4EDQ+WRtGDZ+8q
DTVO3LmxGGTZdo7VonqfYzE9C44vE6eK6agc71KPfHv9c/j/i8vgMZ+//tSj3n9CAvLuUvFYsyUj
15F+j+pcTVmyFCYD3PFIVKx4+yL4wsan3ZdIvkGtmKEHaYXWVrgmvCdxpHvBulh1V9rgg4AmqsMS
XQN1I62RRfeE/j3nYlsn9ttHV6SYtPE0JeWJXe+BDiI895hP9b4qNpMRA84gmxYAE9YPdoTMfpJ5
G8/5YXPPm0nmZ4rdxzZ8oYj+/nPwyCfhoKhIpiwP//L9FAA0a32ifW7L3D5h8D/kQGpCmfR6OcD5
SUTlJOY27yA66HFVHY7GszSDJr4IkIAnJM94pUZYVLSDJTBK/ny648oiKcnvg6V1zKe8M1dUhxLy
7GvbE6aEmvEs3LgTeDJ6HVpi55QQmGRHIos4s0495h6SFMrfWnKxxqn6Mp4apHp6TFOQxhGgrMNv
vCNjsHlbpVbNuNaVvjkKCwABhHHiqOwazo9//tvZzy24zvYzUEzPdgdwGntsYl7WLtl2AEtmGOd7
Sjh9jpcu6gxWa+dS2c6ihNMswI4H9HQJRapSOzGEcBUzqXLbxGU6tUvMZnFKcOeGAMqavCWPRqCe
bjIbygzhvRlnTRzf4ySLJuMSpqh5BQ5vwv+LWWxUeSumOMkqWCuo7Wsmk8osW3z26xMJwyWXF0bu
+CHvtJuvUUFrkFmilP54/WZcsh5qVjbun7wzZp+vlu/KCqavDrlRJW0Z8JjcC14L76u++E0HNbxB
jjygTjTw4Yd9VRW7BHdtqz3GOl4/lYtaowjpWt2EoBCyh++tkml7N/x5rqrXFLmBWWJScRXvhcNw
RG64AcRFBbOiac5SXMdTmm315nibFxcXP/VHVosfvd1iKa4USBgEItVrjDKbrCXi/y9CEms6SSi+
ICJ1V3ZuZUgLa4hg9Wz06cjCqAOiEzGoGkX22rCKdC1Ht9yrDor50CXL/INN1MeA3+6SGI3fpNDN
lfG9IYJh0OZ2quTOhBUm1YJ4xPHq3kvPlRXfq8DXkXbwjhPAwagqchmxeU4EIxmolEixNwT/QdUY
hzcJ2WT3exHklryVC1PUKMe+Go/1DLDB+4n285JgncCMDS0lGAmlH47P5fB5lIAOtllbq4d/Vgeu
DqrsskSwbznPv0VPLhjcIVJwtS8ASTAPcQ/CglRq3D0AtThbESs6ZsbLD9VKxGpkgVtHreX1oqy8
CNfs9DX3lkmDh6XWn+B5DJoHSNUwBxVB3V9Cz7sGdvV1xPwJfsQMOGDa/TGSdESfvvMZSeyxjbNc
sS+7SgmfnC5NpOQkIPa9kDTMJOzHx6BnjSyMCiZ8qoSPJViMPNEOSOgIlyQkTPnbCDPI4Q+KSo+V
bJRL06gS9iWduVjIb+wVPTYxWqOxnr3MAHx0pagMmshQZUYsaGRMXSMMVE7JwePWc2PsZhZ1wi54
cceFWbdHwe8DVYU2u2NeNTBLRg7DPaJtYMsiqqtFL2xFucIRIGe6ANAdwTkzjp+AzfXclWYPEt3v
GRnXih6S3ijcQ/zthPSn4NUdx9yE1R+M5MmC6s0oY3fCgzlc9b+NxYU3BZ4G8olkyrTorrV+/osz
upASXTilg6AzbzxyB6lAVgsE82llprtTQ7VpWtZjIfsu+LjsaNZJGQQcHTMSgXCV1ETPfYWHZoEk
XZuz8mEpGq9T/cXlDQmactP5EslYmjHw+QpOTCtnBuAheqFh9uW4XT6paD56TBlUuAq2qH7wTH/r
a7fFCnsiaSd01o/AchZfbtWqAyZaokD6O/AQMrQFXqyH4tq6i9KuQYQhz1rCBb3BXCXq0ao3cGmC
wJ20e/qsihBzQFwLAUqFL75BbEz8Ihe4ul3FzUUFWL46S2zVFwRZ8+JxkIfWIegifsdjCLACa/5+
brmh+g6Gy7Hkbpkh9TlfI9nUVc1TD+nlZ8LWvP58GBxh+Ft7UZY84g8xuCqMP0PDMc3dgAgAZNuJ
U4uZVnWXOJXyHdcGUmeos9zOQAuqTBSrnW/EuUJ2zo9QTLyF3dZohD5XX1bvzf2jfjbr7fQWngxo
HJz6N7U7LuGZPAMLE34pU8+wkgjM8n55VIjm3HsfQ48YhCUEvGbtM1LUJm43ESsFt6M7Y9g7rWv2
vhEjt3fWC+YDxqKpx6PTNAtx/YxY6jnm/ncUISE8jMQxKsX65I36kXH8O898PzynxgvrIUx4Ccm2
4YYd0LGC9AtMLTihaC1aTyxrKAfcSdpYrzDQ7PjQuKPKMeY+mQjO+1F3SxxeUwVPVZ+29TWqo/Pe
7hNdlnrfWC0cC07ZmxUrIyOxHPS18NQjjHKJNdGjAgxrFJ7STprwmQhaFpa121P8gwtVJ+IPrLMe
nFY0ATx+nJ58F2a7npzx1FtEjU6f03u1v3gF2oXywt2XGIaxBiAMMD/C4zoZMNMzzi3SndYi1SVo
IORSD4iKMEEAl3kRs3VyYXgQwTLy/OTNSABoaqTwZPqKN7poyWxX7FEOtrdumWRIl75gBezvx8Lu
2578szk5GgVjmyqL/ZAn14Eyprth183cPPDyZTS775pRTkrLmIYbQCfDSMGbxD4IWbUwILZiyk38
NcZL8c2TpBzmHPB+9DOMcBUh8phrus/8FI3fm0cPvcxljMAAIT753s7lWjgdka+6EP7/R2elyC6C
HgNaTvhKMW1uuLmkW7gkwdCjU9DqrSbCSE3fMUQ7FgG9UIDYp8qwq01x8W3oQFzssEWtiDNl50WY
J4588GnQt7zFHWDF79wcpbT1IefYftJRm5A+C0RdZ6hSDmii0FrnYWsQH9KbfaUUkkFaMp4VaoZW
ifxbf2iQwGIPZOldYsSIATko8CNFxOV0y73Ib2y7GusZjd+cdvgbLgY8vr2q5LQbKLX1GPqBZiiS
PYlOi8EDmM8vjES37IwhGEu87/Mr9Dq7qc54OXPTBD41VrW+pDzZVpupC2bWwk8alKgmjS3goH06
UZOn8a4Kwuo+cgEAHMFfdKxCdXqWSh2VY9CIVze/QwFmq9B89s41uMH+8Ug9JfK9srARTSpUlXGg
B0cVhDvdAXJUYrsWv1q6yt4PElzGqerPxC+k3L6LGevZLg9ep/GAby6GEGAkNYfp9wWbvhVS96Vs
SBEugssOzZh8e3g1PW51FRejF5uvguVifSa9vb3+rXPIh9M75YoNKOQl/ZMsz9xLGypRDHP4fKuT
FiltUtEw9MGr8CilOIpf9tUbZ/HtDgsJZrkPHI0JPpMbilzO3+5JvEVR6zp0ynYOFUsUCaOt2+Mw
6BB8kBf68HvNePx6VaVC9TKihstrfi7RnyAoQ/1Lw5sqUyQ5gp+UVqRLTG7WybGdkpn5X+t+p/IX
05RMW5hd3oM9u2x5CECqPpPW2hue6diksKBpfDeB2HXZ3z9lLyKS2AxWOOsgPAL3AiSdrHdZyECP
mzvhFyjBYgWHE60sGjyYsOnUDAAO228UStc7uteucaweoVvYTibYcUD8clP6VaanY7k0wx5FRKUc
WpUbWHTAf/g9+wjOr5NiAL6nOREeqi71BlHzK2ZfbfK5MFmDPhDW1DJi4GOpRYFt0UHyde2bOCi4
FrBNeePGqi+Q5j2VIQ4/xdR1th1YXet3Y5JukKATe50kA41g3FHufeb0OZwcyIYzdUnU4jBBnIXI
7C/Vf6W15M3pjekP9tluVUEDuLOFqBqvH8ycuk7qqJ6KhDUygJCm9E8xJYZ1w1rQdBZ0mBcSWeR8
cdvCWgLbJDaiyzboZeqE52owwObrpug4CF9I1Fui9u7DmWUrMhUxBiJKl/3lXMc6BrN7gF1UJEbN
5CEgmQcocnjS8T6C2ndv+RNMm9V3OJ/IGDfz8vfudYPGdS9Z+iULBSElXRuxXynv1xvGTqCo87Gm
GYVp4V8ExBZ/dD3uI3zbOlY5XDBv3Lu4CQvyo0sdiqK2RwR0um8kG6Lz9dOmknGQzOdndB/f7whc
FLxWgCGQ8FlkrmNPpj11YPFaZQEj8SUGoAsmD9md3XqnsIEOnsUabAzjv5ulCvRNUyYfzui87xz7
ClQuUXUH/Chx0Fge7VqzXIdExtvLYRnwKKjyqu6X4KbQYPGpdGI5ZXqrjIJDH3LDPNKlqHlud7Rk
/nQ2w64nvZQ17J3Xz23gBElHDByLC8WIRdWGsfPi9cmZHbGtDB7lEEjg2VAm72447BO1fiBmfCV9
fTLzMci9Yi5aiTEoQ+wuZVu5vU+gybq0crJcuXOVbUaJX/FxDyq9fDvsU1my3t+054kHPSIf/4ti
A4em1l0Qhmg+3HfvEvcyHIRIiftLe7C9y0/hE8B1YJW9vMilD3pXLo3xlx98g/cr06ZU9MWRpLrA
ybmz4HNROqETxMK1bVlcdEVd3eu1x03SIDhUT4naBTXDWHEHrjVvBywfQeBsYajC9bUVm9WjGdmM
Qmud4G1Hc16LTn7JdkZLPFRu/SNvExtud54/JxQaheDJFZUAovb5N8bkJUgigJn/EhU5u63J4ah9
2O8KhAeEmLf9ryPjU2OyLb2mgYhfjVZqSfj6TEtBAqdIjiki2mTF1m2rvNh9PBZTSA3Klnb2AeKJ
a0MdFMmvwRn17NU+/ObcAR9kZVO6WZnrI2n6mO1gRlLn8ZADDXP5YsiCcRxcWv5qHi/z95YGUuHc
vUzQBqvbrwG+AyFKzb3Z5DhQsF6tyzm9XdwReL/seiWUB3eQbFvegndfwwW29L9eNxdLu03Mng+j
/tyM8jOeef/w3uKxRA5ivUPDykNdwYGg6OnS9UG5c/+Ssy8M9sgKhqiLoACMWMzDGmto8LSBlUTC
Gv9IKEMsHI7ZAMiAjc79c+0Iqs8IJ07UHU2U+8XNnhEWnxuiBbDpDiqtMmdED42cTC+tV8G34lFF
mA6DaYDmDKAwAVlmK/U/bghHMJ+ELxIQQ9G1Z+bI++8YvucD/Welozh9MjbSVnkAXP8l1nwneiM4
USQewc6m32qTmmkg92DLDlQzBZEETz7Nwm9MXXoP2PlApxIEnjFpPPl87L3Dzgf0RvDWD99CVNFf
NnsNWuKNlU+MxzWSLZC7TGIInw6AzeCkkmZo7RHZA3LL0wUnMr/RXp1IB0VJDozoUdIG2SDpm1JX
fccaN2WMctBuQLn1fXreWlN3Pq+2bK1ksSUmkqMXMG2dLu9q8Co56rW3f8+lS/xAw+P4p/OmsUyS
2bW2UG9Qr/XpQmRhR3FMh1Do3NLxOp7yZO/Zw8/JH9FO/HMKCpwK4mxERUdewHLpJsfpSuwu+MxT
4tkIe3zvMx2w5jlRUZYH7l6O0KcJGP4i20xI3VVEwzpiLRu+dcUww1FknwdHAD4eUubRGmbTn+YY
aJ92h7+P20QpH4qdBycwUu9phI0Fr9MEX81FXwY76EDR+C9G+7Qw50/TIejlfiQRmvv8azKGWKSS
BzkwUTFdfy0tjxq+NL3y59F7iAGAVrhEeVKBAKtzbRnoWnOxaaH+ddrXIoKRivogVZuPuO3+OcUK
midtSjrv6uwpY+AXc4Q2g4UIkrwyeHhouMOaN77XEwmxhDsP37rJBP20otPvCsg7cc2gBPHp6C/Z
qbWRPSUyb2x3A/RsmhgiRvbXqQ6CqXMHJO94bErVS04rjbIghUfEKtlIOMo8E+bZZ+mnm6VCIEfG
l4xioDkcJFAgJUqBjmXsWKOQQLCvxzGiENbn81DYDdMt3sm781NjL+BWAJ3DZBPshq7mZPJHm7My
83sU8inhycM2diaJW05RSIh9Q2RZUxQEytQiSAj8WW9uqIyVPe7eARZv19BFIkFHB2GLyuOn9/9z
Asb3j9vVykD/V6JWpvFhslAdz8i2TqRQLDuDXcILJ0WCr0WzkfMKojj9gdnTdJ18T9m7Z1knD/ls
kjJ14o5+TdfIdd1eVjnNlPyiHgRUYNXux3VY03ClwLspPwLqJqg9Qy+4+x/ZsOgIJ1lXpYQ1VSGj
8fttGIUhs6GfThSZh2GdlBTjLeLwcqqdJ6M8h/mHzitwVkR78WaB+Kr3RNWewCFjPp29UFEaA0xH
e3+2j154PQnKPawsh9rHwRUtOgQEM6usNpIvzeeVlRoQEyZTKBligiccKkVoTAl1WKoHo0YgrqGG
iuLbGyQ5Wkp47nuAydUB1uByyaKGahzbFMXynyJ17ow/BzNjqDwmkPJlWnKhOEn6dpNFU4hoOMMf
pxpK78+2jTy9C2meW8wcqiePsxbib6ZmIlCqS3lDtm1ztQKSwEsw8nDtC+9tDkPz4YsUnDDBqRCn
iFoPkyZnreLIOZa5woOV7L/htBaQK1TyaNCOBK5Qf274JJ9rhVn87hxg+/ebQTXhbDkZLQIPMA5R
YgsO+/uNGmeYwQ96rA/LIH5nTpzWbuNHDUK8IyPjZlfw+9q0bDD8OPonA0gZP9B6ujSBtW4CqbDI
xTOYMujzgFgi16Di/7CIi4NZlCOgvsDOb3Ov8xNdLvnQQIOVzpFNlquIv9MbK8O+XJh0uozKk41A
QXiFYOB8HC7yvbAEnenCmaWrIRTFbsvTFSVyyLnf+Q0NttzJS+yrbE/F7zXYzcei9xnI2KXkG9BB
r1/N4RquHG3o4KmPLh1nkpjXyQ5qAQaIw8IrCYnoDTpXHpZA6mchvGtSYaSuB0XSE3hD/rt6Gdqw
wrGrXO6tfW3VemzFV7mTENv5eCRiiicmi/cNhejvSwcCECoZOvU7OMtAvM/QPlCVY5RLAuoiZ8uR
/MPV3OlgmjiUiGBNcezRvmLKdYXVum9WbW7A8MhPo00j4WCCyU+uMACsaSji8VchxNQLsWkTG/Tl
XaktOf/JgaNjwmfKcxnIXFo0ueVTuUJsbg5bandI35fU29a30GWl2j7ashSXyoxFzX0PIza/2MR8
1uql8EjOODFKlWGSgrnv42CmgB2jeYRM7XzC5rjwDPbsHkcL1rnl4BrYF1xmJZomqjF/i8XV+of1
/aSjJsEsSaAhuJFtPR1/T2QeJoivz5v+gdtjrg/n7BHxgfCLBEhmVpUyIt5DKCunZ6hrn6c6yX+Z
APr1lXxhRVAwIRe43WMpUbwBtqFNaEHTPFOcI0tpYvoAg5QHhHoKVSKc2IFRVJF4CJ8WaeiX8qR5
2UYp6/xaXZmDN1hyNCMftI1OhcUkOOeJlivcOWR++uUBXZQcJPxY+BOc61Ez4XSvNnjzE+lnbGWg
6d24Ix6HYNCthyTb8qb1xjmNEi5SF1i/v15QVcy4M3lu5C/IQiba7bt2WFFf+xY3Yg+HP1v9bebc
SnD3CS72wbNR06C8DCpaeNiUSwwZN+DESHuoG5YycGu0VV2tmkNQVCUrZXy/76hlA8fGO6OK9B4z
uZqIhVJQKTNfDckeV2YN+zhDdGFLqKEp79wBnxAmDM8qvge0yJhs3DsO1Q7pG2oeRE0nYXQW640E
BFEjEmYD+NZ/nR77jRtP1tPom6bDyNX4yEMd60tR8AO7AXKVxn+jGF6P40SSUZ+scrnyol3P/FyR
dVKnOwRzZy7RLRPxqhjTswUbFR1YzqpHEaRi6VDL0nyk1fZPxf3OQaVshbx2FVP31ZorGw3e0dTL
E0gZ7+/3SSwt7U8EoURKEswFrF5ynp3pZbF8KQQwd8QdmCYi8fhTnr6eikYfxXcH/YxtqLnJLbs0
EWu+2ImJnd5lpoyJU/LpAFw1P3U+IdvHor7Mrr1jWOwoEosrKUmrKYytwVFticvA2KnzLFLi6+8L
/t22dz8sKRPejtV7NukUBp3Qgfi5xEiEirlC/WwFKF2rhx55PTWDbLGn/pjdXnMG/+lzpsf++yxe
+3vISqZWMOUxuz7WrcCr125Y8HpZhae+eTVEZUbwcacVDHL4KxzVSHxo4ZVa/RD25EUCPyyv2GZK
TrwW5yj6DT3kQ942taHV6G7GhPVLhFkUNY+c9bBO4MezSo5zJ4zouL7HmuShw721O8MzlMVI+qfG
muha6sFqUJUTG5bwuZV6OQ2bfBhFjkZf2atmOXWpBg6++V6c14n7qQd0V/+ySHwGCKhAx64S+A+j
gJf78bS5tZnWJs9QdcEhddgZSbaHSO5kI8UGnFUl6is4IONEq+9rp78m/I5iY307A6Llg8wwjoxv
eJObYMZarmNp6O5QKrQfreicnVa9YIPzq+w3vI5w4rvnhC8BZs9PVTrnZM/AT4GilefZqN7cmLVg
olocZzfRpgB7DvqKSooEiVvsHJLHjoqwEEQKQ/HDVAx1s+5SokN4xnTIR9upzGZsDV20UrgIeyp8
DyejFAv2ise0/Cu06q8N9RebzA034UEiyqvkOrW4nXYUOh36Cwx0UYfGHaBA6hBirS9kmsTUn0bx
RMTM0CH+J4wt7R4gQ7yWVaV6T+VEcSYpHHTbUeZL/J6n5s9drslmxgw4dOR6DN2V7qpXobYMk7vD
F43LRJZpnGIoML1M0/LNPEHeDJ54PWfEDnRXdNUYU5JtvzDL1WtOYPKZWwSsuQEl6ROYUEVDgt0u
EoqK6kOUbNJIKMUraAWFPmhXnPKueO1wkPSrfNah80V/kTbyJNaV0WFWxdZC8UBPRfcMm3poZqGa
dCW188J9qyOcocaTGek/g7o1L7AsS84XhZzZpg4RlylWgem5IhpfOROjk3/ypKvzPGLxvDA54SZV
X/K0hJ24WdIZlqDTTn2S31CkZBlKgGFwlNcrdO3h5xfnAKGChaiEb8J/Xl+l8n6UJw61A4G6wDmT
4ysFYlueDdeIHF32SqTjDdTtEI7zM+Kru7gOkB6DqDQ9+RRX8fx4nFES71sXzMPwKA/mYjlngzSz
UMiyitK63vzB+93kTjCI0nqghqUn1Ukd9IGksGAD2CrGEVY5EtkUi5eZfqRxLo5Awd2eBrTr2ecj
1XXfgWNldagzFRz/AHGBkAX2FOhtpf1CF+ylvpQmP5YfBPmp05CGU3JjBUMn5ymRplmFh+M4aa0q
5WrR9uevVSuHhn6AUTRgDGoiJjkSZkHIgB6XgiryVO/bfF3cjm49EFKBUSH3AhsKGqvPfvK3ux69
gui6vf/9L+EzGFz+pIPwu29U7SB6GAKf9SNRdb38iQxNLgqiZG/hj3KItG3wOBTEddqbzZ/pj7Vg
p01gD842sbjw5NF8dEFjpb2sRE4ETS+UWZPStnUFnd8pZGQayOfvj/vJCfYPa/jJvTKR/mGMMCA5
OvvKAiIh39dfY6EGtSKe/QgHzqpmbYVH+4sYT8wIFyWfsfqfQOGH3EZK1W7Ax06MEy8jLxjHK60D
xz9LEQYANv657sxlcPg8yDhu8XsVw8nerPkc75qZe0i08vryC8w6A8DkgqcbtCLIBNs8VO/TbO5H
hm008mO8r6UzKI1FEUtuJ2iFM5nTpT5Ugh9lPqXzFcQBI3CpTUq/1Vos251z/m2JAkn5GgPusTDA
JD65eHMJYWiZW2jn7db0ylPW7rbtxno0NKEtmf+zQy7jPXMmeQYmwnDdxanGNs+tMmIVw3ZRd/IB
kM2QV125A+KyIMCfB9alUI1wOh5TVBvEEo5lBbjzL5qRsoHacXGm5LqDHDGNmMTaoJieAURydQ2y
l+91k17gLQTHuTs3RDZJeOaU31Je9yPHz/ObPKSIqhVFL4XhD1f+a/9h3cKuGEqtOp+LLDKozfSN
JTcJuGAwhMHOAgupuJInLtM/f5rCNM9UYJ7ytFnw9AGOYAmX0RfkgHInvT+gzN9pBumAmqfok81c
NtHOKA8e3kgx6yNdrxGU5tzRsrZmW00OrxlUkhw7ixO37/BBp9ouN3OZIFu7OfCLn2/GlNNSZmOu
0c0vaQeX4kEd9jXjPBg+DlTZwYsB5Mc/amuZjkdwyxQiTtIr2FY8AhGYNSSiO/vm/ozPZ9KsGVzW
Yy7wh+u3MqoxEtnph9OvJ9wLUU7CYhpEd2AFBeiqnYUVaqMYKJNKsKGrMIshd+sV49GuH1VV5ufy
9pe6zzV/Y7KblJOB4/mgUWTzKqJ/7PTvPHDqhYmmzM2KEN7rnf5VK+GWy5O1O72hAklxqX4siMy+
ILU+KUHpeEy6kNhpwvjAvfEgoyu8NDe7Cx5CSNJ/JCT8xtJtA4mip0vJEqvna2G+yljAuZ9BlR/I
pt1MjwWX4iIHuFWb0ikA3mLg67/DUHoKXsQsqqX/GuNWFaW9Y6x3lYZYp/h/YkIbM6nf2gzvVQmJ
W27Sqa2UnDLaBiNlRLADtJ9ma7YnwOCnsImLU8DVwbA1SS2HaHd6rW4hmyZ/SDf2yE8//wUaGDI9
UGzHEqz9FbbCb1S846Zdq5hBxKIUx0T6fZISK31qvuC18FDZF2dlHpsVgMEXAaQErF3BzUobtRRg
DHf5ts7aIQB353cQkXcDQvLc1lGntoc15ON1v2jyMWZUoEo88Ex8CS2b4E/H5WIKVFoQCaRz9arv
HNOGi7lwIyLiHCi4ngdOUfCuAWBhr4PhsD5MUdZU/VXmaoh0ddEvsLnYAgftbNkx8Z4J8uudwaMV
uEUoxBgq4fZt3jSt0+8EI/hf6R+fO+CNDJmSOwf3eDBuhVAuLKBAr7dH2bPq43YDHXZxxrjJyu29
zgi6zyLnWK4DHjM4xwpjMFIt6KF4lsTwZdeuBVS7MJ/aDMoDDXj3rVWhnCfdH714i2rYxCZ9y0Vk
H55JdeP1ryHXDEM6UIiL/qmfl9gmqcRM/2Cgm70QoadM6A90DhlqBxZPMTCFkmQd4ivahU9vUUCm
WNpqIAqX+3+D9E6te9ljIe8//KU2EXGrN5Ut0Yh6e6kuU3ckCJhkmzZSLfkTgzaa6sI5wjQTTuRE
qryMJAsdaGePh/dGczphlJykhG8F/SHXMt1L/bxWw86tLBVYje+qgWI41zYEwALVtYSWlJwIkM0d
1R6NrtmbpYBjolthPhEG/3L3CkE0+FwYQhOlBtIay0033q7PeWkC676/abORoqLs5W252pQKleeR
KF0iW2JTlesh0ReZVa8cNxV1CNMUtnETAPQlC5vWR6bOGeg7Fjal75b9vMeqciPTx2auW0BFcMkZ
x1WRiFP36uCz33Z5d1nbvfP2LGkpt8Y50MQmxu9W9mEtnGJvOA+fgfuNcGNVWrU5kNM8JXa2n5TO
+zRMTmvVX6dscZLnx50luTQgbMBfwRv13qB2iDvgDCgimXWsmF++L6eqGegszmv31I/o+AOyRFBA
c9aqO/MSw3DXPz7i91bO1AaJm22kpk/5XXR20Ue6DbTnUc4ueIwCKz+kL6Z7Ht+xoayNzA/immjK
Ve/Jkar88D9CABs9KY+ZdUCrLHrvrtfT7DPBWYmGbjTKEWS6PH3/vEVPcVwWV1ND6RbgkNBTTrgG
pPEmnO4hevg6792Cn416bK5h5RIJEYi+RxjVaMGeoZfj58togNF4T8SC0KOlFSRhrO9ARUueogfr
u7vA1RCdu2wk0cKHIOxa2MaiFEPlJAm1l34aJ7DBrCaFYjsCt2Y/3/yWLRGCkFnce3Mln22VcGqG
eRknE3sFTcrr/uHr1gSRkEaFvMx2g/X1+Kd5v4YBXjzkw4kCF02aBsF2rD2WIK3/u0paiF+751F2
Esgr2WmJeG1vIfchoF7EoDGH0T4y3Iq1dmzItYvvF+JngXsw91FzN2JiKf5PIlSK93anMDFTDnFb
Cefd7FBouX3rP9682srk0hMCVm7cFVKqVl1jFJzFnnjpZ6kPpa0Rw0K7wIw58Qpnz74lybNMSa15
gzao905ornJbcw+bruv5YIO1C4a9uicgd9Le031SLG36X/XoHqsqUMktbhLGevQ05h4hMf8xXzu1
nU/7I1uKRys7dVCRZ/IkpCkfFpHkXAUWpkhEGj/TsA5kRw8JKjxHSILW73JN5UJVO2OmYyiQ23np
ATN252az/qw88/SfyAwuCOUSDelnHip4T8g6DxJTUy8dUHDj77fbYfHQjXrf87AbgZUA4pxXhriA
DMBvpGCfG9/s512w65/piJcJ6BoDyQZX/iBtDlVDELWVTZPmZyJaFgPiDPlPsXoMQ7eYbkr4gDoY
L5cijLIq+wC3EPTMzUNPxHt8nHV7eKEiLWGmGpb9xDHL6PDGB9TCZs3ZR1XHytxfmNzCYEAZ015E
R0VN+iZtNslm0LqsPMwY6+1Io4+gn3EJ44f6UL1wS1cFIUfHHQD9PR54W39m4lBCbXyMJwWrF/4g
WZHiJmARUDbhXe39vWlm9qTRugzC2jjgzu4CzCROwROSYxln8pFgGa9AihBPXQXCGh/k/TvD5jQq
suBCbk4tpy9BBOMfAnW/yZt135PSnVW/FEAurICcfkAIKGj1HwYgwRaf88C3tLJ7kshBwPJ8NL8f
cqBejWIqm6vyB6ZSYX1oueWrqCkw4LhrmNTmEZFQAARxIfPDcCicZoRNUEsOOMlx3TKnjdfVX8Hs
nuedjltxuvnMpw0nmKv1XpGEvyXZ5B5cjQeM4egiRqsp7CbRvFMqP9GS3triA3i8lwyq6N8+pg4J
TxXf7pb5zoaeMbdmPNK1XeXE4WF3J1/+uUSFC7m7tX9SaJyKIp3IVWCCihLfvRul5Tv8kkFAI+2y
3tuftMyCDfFh3dFp7VtmK5EQG2nQbTOPhqMU5NUq0Lq34Wnd3L3M/IyfO87rdmhpaU4q4Gk2avnW
4Rfp1YJWf/LUmIkjJcjRzm7cG5RwE42QPJqn5xT3O1AcRVCYVPrqw59v0DnGeeFUzuTQsah7Uru5
Sp/YoyczCJpRc4Ye31tVuVUZBdgS1vrI6e/pWbHmDrBHZHvkJedj/l/jRQy3cXbvKbyhQYUDJzZ5
GDNPoBoKtgG04VH8s7PGmwVZoJAzEkd14dguwF5y3X8pTEf0/T1B5itqmWfXsEkOaXHPpVesCEJM
JYHSdspgDA3w3aQ4UlW0WAEQ4tjV0Jd4pptZ5gHXPldqOrjoiDOq1U2sA6quPDHvHqhZOTYZStYe
J0tdXQ9jH8Sn9j8+6vNVpMg8TJDeHlBVA/lzk0yM4CDiOldQIZPU4DI/2woTuW5XKYY1n+U8m4fB
wKu1Q+WcNTcsZkaSPKBi1tzGfX28DpnkLPPMtixS/mrKxLMCiX9fL2peNd+Z5AUCf4FJWWwYRB5z
P6VivFG6C5aofWDFl0PJYNstQlOlKLR0gy1BaVgvJBV8rIo6kXe81ruLUJ/x3Ma1zyRd7i2GSjco
R79JLG/EzuLQWfEIQp41Cv2c9ug4oquemzQBLeMYdAB0+znNltefwS4eRBa5AZA8GCHEz1oPhMUE
QT7xLPBZWUMZN/gDiQMou/J1MABUaEG7wSfcXzwatvkvmX9S4hokCQ/GPd9LdPVvCqOu1tppHXq8
IFu0wIr1l4+G+19xAa0WRdSqbN02dqkB+bZRoaymtseyXNDRkhQatIsuFFPlqX3BIOnIVHiazm4Q
SjEI7OFtSvyuzzSYdEKkEjLLKsLEfjyd3VumqUSxHiabsZdEM3c6r2gKQdP+hdu1LEefwyoDgQNC
q3VcyN2NU6eI8VUS3qtuWyMi8D8Cz8URuMswLIiKRmTtxee8YTIjfbHrslpTGS8QiH3U1zp4wtQZ
UX+35iC5NO7v8ZV6LLY+84mk1dnk8HHDjuVazh/ZhkmZVDh7gyk0rAyoQdJNfM3Rmk0qy3NdwNWF
aWgTXtpK56lHBdeM5ARJaik9AVUldRPDOcaxjlhw2eXh1edfriQZCfthkac1LVwA//eKj1dxKJFj
Dc6hkQ888tDKu/BBGUvAkZ7+gNMnipp4PP4ojFlTobX2E7OFbHXZBltA+d46so8f3tnqUkXlOyh2
pjtOCNteJ2QNHicRLvxf3QG58Ccg9rU2KdGtkXLStzofRSJtnsYzRqNEpK51DMtB5GSX8gBoIYj8
Ovaj3GIcvE3RwoTfUDK6VB8typ01W1jtbbdV9v5iT5LRb/lfNwx/R2q9LbgDxkdhwfgSJExPM6p9
hFX/IDS/UqaBipTL7qUhL/dyVT5GB2KaTOJFIct5gykC8Mt5wSadvBanMo/cjsJFA5iBPhBnwasp
/QJ0QE0/0INOV0Qu3Hz5VgHorLE3quhq8OArPBQB3RMQuCr1hZDMleYlKYevc0do1X8d2STQpOID
WbYExmwDvzV2WNGPdgfrIZEwEweTAEkdWZmGXpnBTf9wCsh0aSpIv7o1KaeEYxF4vv7atnT2g0PX
JLUwODiArcoRgkaidWXB6vxkXKjdEtaAFDYN/+zPfN4p97IoPIerqHTcL0ITYZQcGylKneV72BoQ
4HYKyvwsoruo2mIpgbteZTQEIZ/6S2boN7JTBhdybeT0FDRRsC/HTJYS+MWbQTKH5vzn8XlqMIqb
CFbhB7r/OFQY5SNtEEvqCxLUl/BdTMkABfPYS3oX7KGxhz2rUGNPv0smuwEVB99bT/HktcYysg8o
zRb7WvsG6ze5P5jjdT7WOg7iWamDl0WN3VN4q80ZSLEf5FnYNkYDKIUifKx/4bHYuz9wt28fmE9y
GO4Ubu1xNtsYC/ZDxCg/O66NJL+W6zmD+M5sGwbSIm9s1f8FdJMXdRpH2QqHtMZ00iZA5PAt9oRp
R16CD5RRj0HvrZLmZAlhOdMZ0UQ2aUd86gJ0KcpN1yTSxO+nYgagQI8v/cH003QB916Gg/NJk9SG
tuOau/Ay2aDSVYgLKIXdMcNNtagDepR2TF5/VSm1p1dRuNaf3cm7F3vhqXK4OGk07v8/o+fo/U5P
V4gMPJvNTDvcbPlX8Q/dUNGicg47Sh1SSQwNRreechh4bo21NVQexBjwFkO2SAWXceLcMEP08iCL
Cn7QL8iGFUi+1a9we3VNycXC10hq0u7xa/mmr/sCq4izE2mqYq404ApZlZ2OlNYfgKvBCEKKzVbr
OCvJnu6NL2K10VTVkDkQMaoPfZc2kSgWEhNBaegLMV8OMD97aVtnyiwxOA/HRF57yCYXxNdQNiOy
rAlvYxTntQKT9SDnLkrlpDGjirA/qbT/QJIxhCwxKZigzlKMw+Ip1C+KxJ1U5Cjp4FAxkedvMW+d
mTGrx46wCWvN6b5tidSxJlktUalrCpT6xoHglEC2KnYQAuham6nuIJM5mBsxpwrvWNKWOieqzbRO
/6jnNCCl76w+HANA+qbe2/vR1mGMHMvURFZzXXCovinS6Zwom7+csh/SOeFZifzEdjDg4grmhn1B
udcylwexcIoAC0eR6GB07nkBfj33ZwlfW9taNlVoL3h2RN/iaILTGXxqGuGVkmPy32KywMsVXwLx
FHjDnKJgoTi20sfmQf+9FtoSuLYRsi/V41h9UgHc20w2DnZDRgueS0lPc3HaONf2TVPrmGAZaGIi
vb+8cmImNPrO4PaS9cQESRcPDrowUuixmS7Chs+sLLklaj5YP8rIZg5eysRNWX+hMkpv3WXjZVIQ
T0bl2v3gzrGmHB7nqn3fHJPIQ53oXnNXy+X6qGP44tUuRJHTauMcxhTUqxmSB3SmexMqOAAQzgiN
GobKtUxbPxt5O+ogsEOPI6sdNTa4iYjx7Zbp5gzSqfZVWeyKzWNrUjx4whA+lCvnE9e/g2ijimBp
Nt6+eGwzlj/OVmKXxpddpunkLZfkM5nwaoIM1j+P1PJgvi2KwAahmQedXGpUMCuGsEO4IHEIQGH/
7fYBMj/BlPuqX1AxAy5x0LFZkpClGX/1xWwXCRB7wYPjjc5yzGFpNo5zj3xYgXO25lPC4l57OHH0
BZvh9MkgOKusnAjWxOA4uYYf6xMSWJRsVJw1+FUCwWFS6IWKmSXI8t87dgBo7x3ZR3PBn8l5pX/7
baUqdMVJKHjkHp01kK8VaNNMlH/9BjRAMmVYejRQfcgjbqPRKm89c/OZ7NHB6yZF9OIPullRfhLR
DGjnavzSXtOD00+lc0kNGStNMj31e28b20yOzgJFgN/to9/F0xieJBF5LOMMVc2qh7iavbt9IRDX
P0VLspqqDRQagiJleeUXzujmZYnskJI2wmPuFxEoEXxAOUjUXvT+sqpshS+7+TJknmDCBmmr6oD/
izYvQxJFHX0ySWq9oR7/ML4/UzucbVMrRiaKIAfBIdZolkx/n41t+HESfPdf4Zqw/19F8uPRO0lS
Ntg5gn1Dod3MdagUFf+wCZEUE0FPzbZo/Elh9CL4cerdPtIviBreFnYaqlxSOGCJK7TEhzhPEimN
jpKFS+BxS+6/Qahafh1wMwfkAdMoDyhTYsYDkyboGmSfhrV7CVSj5d0cFgex0wg1RjTsqke4RWME
5FchyG0GqHM9PajYz40pwsqJmO117P1hTJObMLl/3w3bJJZqFZ8uqsfflbxFAFD2uq68q9p7+z2M
C30RWjdSLJ3jUMhItJOX2Ko0z7FDXXo99ZwpqXW+nDZ1kR3V//wd0uUodroc77R593S1gstU1DK1
o/dJPCzHpgS0e20tjfpGYwK1WOnL13VPPW9F/8zOqK5f2yNVArmpUpAHe0PAlw8OoWzuDr5DxEhk
VOM7Z9UfL/bf3cGcZ5J6O+WMtrqQajR2UVb3umGXLm4qlRTdbeFrL2LA64E4b2iFTRAmxqDdqdjh
wCoUw4bM1JZYdxFlbhR/O/VGnyUKZ96iPfPIbsZUmz036H4e101dJ6KVZLj5xyrN3uX68pu0yuS4
El8ZnWdhiH9t3ERDO/r7RRvV6K5wqns/erc15pUbbQ/UNbsBDOXgtpYc64k/zAewvr1IKNm3yMIQ
HPSdsGwzJnvQcwmOiIMQnEXuHXVqb5UeXcBb5whw2hpLGaX6BupgiYhI7TXXqI69QbU7YfklJlYz
r94/PYjFSSd7qZU3zRkaiVH4cJsBc7/GC0MW8FBIEDJGFi2vmN90osPko/nX0cdycnSgLVBDynEe
RkuvhEGch7ngf68w6Wd0maSUJCpeyfKE5fNSv1dw08ndW1tP0Vnhlr+xt55Xraam3yXtSJkpUm8c
dLTDbVIZzcExffSXZsy2AUQm/rC2fbwSk9ksLY7DLby60bVBYHhl8DXZl21P2DTl/mluKOdMCQxW
CIfS1RAv3da0Pu5Q3IpqxYK3KMxJgFM4OV8aeQl+j3KMMkRM8e114+3YstMqat4mmy+Ct4t5XGV6
Q2JwD19OvdW8xxIhYihUXXQas668MAT8ozFKMnb3j+MsEwPVGI/cEVTb+hUI1/CRftWXp7uNw3i7
2PfaASQ1GbIpQ7A+rmeveXDASchHXQZXScTmRo4EEgpCcDLOit63ULe1tVq6FJYJSzwNtk3Pqk70
Sq7uAneluvqEd1ZisLxN4KVorzti1UxhiOnjq39sepwUXCmoe9xm/XayMuY4zrV2rWqzgT+RKGky
39Vl3M5EX8NbV74f/hnYEOPF1qZOOvaNn7NzA646rFBf5STJxddo679FcI93+Squ9BOkl0GLYqvR
u9X2f2i38wdZvnR4PdKH2+q62SVgbMbcsgI6SxLZAL1hfZjIuhTmJD2hDAJ5Ugc1xoo8INU8AWVu
iayDZeoaHPif3v+4bWfLaoFoNBJFwsk9w4e4WDsf8uyZRi+DitwEe7hI7TumQe6Ywtbn4Mkuo99z
Cpo3yZAO7ijxVD99eLQWzPVxAXpc9fLP5uy4ebax3oB3LqoWm3DaGdufVX3IeQMPb2eD/yPBSsAl
bGKE9oFWihKczXEeAZSYphbvuzqU6UY1xrgT+TO7UniI5NO+DllgaUfjGFvqbO2q/Ljpw0leWyuY
obkPss26zSpw8iNN7cb7wjxsZ2dvjHGQmv1h9RB5VSaljEtKmSidtaBq89/jnVDQPzWaViJpz2hj
Tswqf9uCtRaZn6nV5mHZ8mxsjPnYwKWtJ79lGljwE5xPext/qXjR05gMqUBKRrrQiqtT0dfOZud6
6/hEwQ3w/8uT8O+SgkYraSGeZmI8258067II5pKItV2TOAQha3Tp+sYeRH2FhyWPtAyCykVpvfwM
fSK4zJJ5IuRTDftYcL+NP+2hKArDSSf44RGlZKrLTua8vnej3ybPNWM+0ZMCV4ICKF4nHclhgpOo
GgS2piTU0Ue5brFwBZz038U/VGhT3P/k3/7uUEu0B0fXZqU1/P5N3yhbFgqkpiPj1x7Ac/2gbTF/
PaZAn8GW6j/Vh8Lryd5jvJguGW11BkVe1j7wAOy1wV+QoYp3trt397B1PTYNs9MHQXLa1JrewS2u
4/V2a9Pdn1FOendLJKf6xqHP8/DCYYSQOwh/FoNvI+wT72d4NS7DoUp2VTj6+zBxEQy4VvFs9Y55
z+KKCgmc3PSJMFGLTctBoYxQZmM+NuTj7Y4nogiR9SX/h2oHIa7S6n5CcyYhzD8CvHeSW4iWq96o
FyN7XFf8aYV9FChpgtdlk8wY+6ZWCaqiVM+1kuSQDdudiqNDlkB2WKgh8VowSvtKXHNjpyfQDDZD
kJzYjVYrBfZc1clu83TeFtxK4I2vsI3uiR705JEjAUKmkl/uhJBRgR0uQOXPW12ru5EA7SvCp3UE
9j6nvb+O4KR8ojV/Ad6PuXLO7Yjpk/YcvRQ++p3SfcPFZ5l9obZUBVMlvTDqPEYp+jvUL7QxADM2
oKDWTRHxD2VSD5HoUiCAOfDh6TqhZlq45K5kqXFBqjngcNbMqVFQwETHHorK+ND7AvYLQsAsx8lL
alFl51f2xTYh56w78BLBin8XaMXPRjTieOIWfQZ6Q5X5MrksRrk/Fc3p29N8eDcovcDhRseZuvta
chOqhQGJQp2ALOX2ZExrq/DamBVtvC6+u0LaSXnSI9HRH098rG25TwTPhK51Gvbpf1EHL6dYyHpk
BxaCFp3jQz8HYQDoiPHFYD0TEta8dGlx56l9F8hTLXO8nb9PV/hEloaZP4ujXcHHN6uZiENCK5k4
8+SEUeGLIWFuoNjbeRMp8hLm0va9FjhYVeE4ZodAUUt/jtC4/h631ND2OIFgsJ6cG0pz1ZMpUUKJ
3Y+N9XqpQa6PzOnbAYclQRncs3vnEoekwJZEibnQIDzWWkKFAG0KswZGMsK8i8kZ7SQQmVv5JL/S
M+drwnZGjUUd0ig5zgzKcPiRjPfX+bjXgN3dOQ/JIasAGq0oTQ3C5UJICBXN2r1cP1KLh4uAGHFF
VhI8YU17iZqtdyYk4jPVgFkd4fm37+V8jJkfTZ4+WmCR3sOTOo4EDcN+fYHdgPIEM/2lDLuxt2wb
MDaqdFsutVJTjqUg3x4iqeOwCEsrgbFHZsBR8Z1jl8mujXMLlQ12n5P7u4WDQ1UxQIs/db7w2/rU
4JkZwD2F224+5MZxolDIfbe5VkzOJQYWnlesL2N/+XBVo6T3j81TTktmnw01yOlaPyrO01tBs8AG
ikjupriBsjb66RvBpi51/7GgAFzGmUzs7uMua52xss/lAj34cNI8qTyORMu2gAqsKEPpEAUckVNU
ShLueSUrNCCmrgdV8aT+Jl7yuH/yq+YyqY22eTivuXeORcda4xAIfpWT16Yqx0mfcyFpHxo4Ixhw
Gi1ygV7Y8aU4+63XnMEXffO3j5nits3RLgf8eBBVZJyWS4wK5UUgs6akpfZkDsEw+ocQ2ZDtTN7b
qRaM23WK8n2LR2rNnhmKjxyYodiuWGyeDf/qPuFvPyHWkQSuJVTFNUD8A0lUe+yfXxgcLNkYCas9
fmCAxgaWfMZbymqdYDrJKHSezscQCuKCHxKNavCTRKyak9RpmCKpAAQ62+J3yw7vTMTd2WVuOd1s
iCiMh6qHd7bvP5VJpUY/HQ/L/9nDeypF9lxRKHvm8Mbgk5+d6vfl1RZS6QACdmJ8tERixnTLufxQ
owhmHFxs8kNE3N/Z/FnOJss3r8IRvOmtgQmujLo7jLKvNNnoMj+s6srI6Fohc2m3obKXfZunfg95
NWYWC2O3WLxwGq3DTw1dpcZh3yhKPBAubRMCu3Gi0adRK41SsuIUrr3beAoYcExgJIZD4SE0h0UU
0ZcJS01dhXDlQQJxf1g2DS0w5RZQsFwqIQApVcviyYMwaX4TyBfZu7SgfTF/yyf5lIzVQYy0pVJH
Yjx46BdQ8yTFmFLm+lqJ6M35GjJlMz8MAJhTxL9qBgkrlVL1vH9l4IHOI/pfbfd6ytfm2fG4g7qD
3WGqzDfcqG8aeu/QAGtpS+8Hjd1N+0h7wPMA1guz2xf5hTEeQhzaDFwUEbCRQz2q/YnSZ8ydOznb
XRxOncCPBTHCQn7W96B5nxKzYFXHJWnN47r1AaiYwT/RMnHjmdTCWhvwX/A4viOZbCW5ZtUWw6yg
2ClDaDLghGAetMU3/IgRKhEZhY7ZlGwYdL965e1vcQfXbapZpmGX6TtDkpA6M1s6PcRjTu60HEP1
tiwXcPzUq6XVWaInIDvmQ9M0kjcsCpOj8WDe76stc+wOU0OQcS1IV4MJtACads5gudalc4FMSMIh
48U7xRWs6yQ6jaCmQrFxF5reYnsndZb5KmpsI9log2VRdS5cghe3hXnBiKUVqus3MkO/YYLoSeXk
QSE/ob8hJESTSLUwPvXaFO7KpIJbooTuZizvNVzoP6/3cp1ZeINmuvoZGH7CgJBUD2u54JSq37s3
jcPOndJdZ/lyL0aMFj3UK+JbT/GvnMUY9gF/7tC9K9YXpxSuZmREAr6VJ8eY/A4N/VhXWedoxmtA
/77g4XPxTnRIYVoEaTYvJaQ8RegOgRVAqSDkSFDGQacX/Mq0jjE0AX75dgdN3TkW/SxdwUb+eNNd
iAUY24lF84l0OS+2uNTxS0I7YjKSE3dQO1cxEVdfCrnWmR8yAYrYwbnqDG4FKgNemRCJVheqtoKW
Bx2MbZ8irF8eOfPtJwnOuKS603gXrqA3PG6SqKYA+tr6Naly3DdBO1DOALLL3QzW/YOCbPWC1fdI
ym465u1sqBzvPQOD9LoTOTLIJa9QBbColzrCinoHpDJJhggHRQFxHPgUVOruGWK4cuDh6KUqlhgn
Gt/yRnN0ofDMD+S7nFNLXtFUWnvmAGNohqwEeaJlxY8hlE7/PU+Pjt/VpKHG+erur6zr1S7qmHSr
aFaYKeIf8CdYuyEkqJf39Y0XDK3qtD5Y3jtXcqEJlEJXFCoeUKU/HlAxkSBZjUXYICK66wNpawi1
RoK6WDWEIu0GY3Wc7etaVaKr2O7541DQTvvEKkKEchG3Wf4CMRoyq5FGJDyhatRKUs8VquANb9Nm
XZj0mDtkvSSQ8l8Kd35KFrU5eqKEqr93BvFiaxnTe+3wuQhyiYu8/5dPkpIETnbyMsZTVHazrKyO
ou0L9unZrF1BDjO/gCYYZ/D4FfRtLe8V52h8ajz+V7czPZEdwNnseSYnbDpCSNIQPiip0eLk/t7E
gNPEVPiGuqJwAAbvGVIPSPx2Aai7xhB7FqIWC6dPhEHsN/zzqyp4wTx06DOaMIqWaMPV2FQchEoz
VFp3pyDkd4a0Yo12BL6ygEJ2eAwZY5HF4xbIN13+BNQ2y0n9AkLZ88UJz+upIovC3IEwR7phle6M
qh2dYfsZX/nC0A/X5KEyxW2d7IAppXl5v31SmwouZIKrMQz5wmRCbhAc+D4tJLAoK3cxblijstx7
CMIPRF/asFkRyYXrTMA7mH67lO0xqXGo0dIpycH/qnWJSiVk79/tO2S8UTpl26XPVaw93Sf9j5J1
eviVPsXdzOFSvzsEDfh/f5dktivxeWz07TVGlK2thjrHq2cc+glax3721JQO8Eqa3a6sAcq3FABz
uBw1noYeyF8LTV9ZqRV2xMg35bZ+PF3wfqkD8HkUwjOl8DijUhsAOkV+W7PNAcn9tn1Wy8b6aSZF
IGN+ov/i9H0x05QPsFCUfKFlwHuUXcyMqb0V0YTTSVJgpcq5XPjVeENyeaSGrjud+wM7yg88Zmtd
YjOgo62QU1SOtKgN1CDC2Br/nvKnF8JJ9SrjP0h7dFe0Bs9LuQ/qGWbUZqB6GO9QDved6ItGb6+j
1vW3jvjwuYKYTCExg4EzsbEPKVRPImkZkVgT+8DhARGx7eE7MbH5WbwV6668EqEDE0D8e1gX+Pmw
GPIk+7EpKdwv7cIxbdANxgHI7CrlOfg2KdLqPmm79VmNihl819Oiq9/D+nKWUExxQrvQK7F5pFOI
2hk62mkOrICi3mo8nONzSh4kSvhh6zPwD/LUzoCzSKcdXL5RT83nyV6herAARBpEGhJl6JCYL5ll
c+HBg4XXfmvZBGyWMVYKBuCYfdDmp/SK0o3PpdU7QI1c8+1ERj7+Km+zbyTfN6YlUhS0xDFp7RSv
TCWsU0sRftcXQOnxvDMPFe5VK4qVYoIOxciPDn7uSWL32K9r3HffpWkzEBBQUx+iAk99MMhi+JW3
+nXFiyWFYagjj6Nin4Q6i39Btr/M4kdXYmEfXJGeE5irujNmpwXJZk08IefzJcPfmDgnWm0yhezu
yLQ8NeDitWGUkhBnx76cYiVAOzG+XMF9bA8yDE4igl2tuxPAcENtFjk6+dFWh6f5a8IVYqiIJnW5
bbq3pSQaw52OqeV2lT0MqoXhILL67WPbHBQreP2jEDVva7cMygxl6qrDDrDxfilJm/7exhGrJ2uO
yZpXYNDgkyMsnScjbVGCGolYa0rvIfrMLKELwBnlUa+maRDyHT/7d6LlnnO2sb1z2slWKzH+djTI
/mnbbSwiDiOeMI1hlt9nsbFuanf/nesIQlOyKAtK0mqlNp5T45WszYBdlB5ay9Mr5Tfda0yGa4aE
s6VjSNKg0eIeLOxf/O+JwI27SmEKq5xAFHS84vTfkOWxKsYCnpZ7tEtOJLFpaXD3GycwhQi3Om6K
GB0MqWhvGPn68EQDbPL8PmR444D1qfQZ9U48wx3hGhliImACadXyPStJpyCBw4qLqAKuU6EguXpJ
9N1Iv3PQP7c3xstRnOG9mHQKQTbNFCtjC/YME+cB2DwqBdrq4BPMgo3WVmZIrqWDOk0nQcwZSbu8
3RthLKYv+g8k4v+hg7JmbQGpvZq0OR62723E3UHtpohy4CknSz4JpLuMHI/531NOEO7h/BgQNbg7
EVS2kusj0KsFxBvDARwN3D4wEfoQrkKrefO4m9qZP+1i7MBWvN7XlyJxYMyQJrbWMKl8stVTG1q/
Excfnc+dE1/BuGPcvE7FP7cpjkn6l8A71Z+1KEzA2tM9nD3iRrF/gE5oyngPf2uFBvQWigHu9AIT
MdykePCKGAp9HhhwdbeG78RU8JePqxYo6QrFyGrfXX5DVHsxFSUQ85naiv/T4m6n5PjI3O0nYyn9
QLtVAWoSTV3Fs2Qk8tjkoxPBKuI/eIibt0fF38hwg70wqO54KjFAdTjVS1b4tX3ihgA99sIMgeiA
rOinBAcSaQyFCbvm95BVo4c7UC7athQGe7vA4uWLLVKeK1LWuTXCPZUvj8tl2bCaHjuprt6Y+ilw
W5qfw53ScnQyQGAZXU+YpqY3GkgUubt7VX2cGyG4w+ATtXHEe7Y+Rbqp5HGYjb4sW5nrSugcBUz6
gkQIhZNyQqofcjM/urPSgH8++xrMi3UOu5PjZkRaYtbZiAicsIklnfzzb8yTsY1Us+Z+BepRMiGv
adog35tcfuBVNSw/Pwy550DO79B99bitpraeHN/7EtoUshcdH8fga+Jwn4LHCwHWox/cmK28QbA/
3w9Qsqo8KtLdPwKG4N1YD0Y87Cww8X/5xdJ2wVSk99M80u4mBXjQgvHK9VKClQff/0A1gTdcO2hK
tVSY6jjREfD6Of4NKV5VpqW33C4SW1Ys3wZuBVgEufEjqiN0m1Cs1KpPsZTQ8VbOcZEI9fLC8kxW
7VmPPhmBBt8c9tgDYRyvTe8oV00/eg5sy8zGQjGb/qLtm8paklOsIHikVZ1lS/E+fBn1ns3FVmXZ
RBIfv8cVfHAdWfswu8qUON/5/GXgpP9aeLeCAWpmpa8MLD6xEmJka66pf3MigfeCpAtuM1RTjIUb
Fc5sPXPiU3C9tYRkoOc1ZufafP1whqLRhEmMcW9WmB3Qq8oUnURABRSYnAnhU3VKOXsjDBBPhZui
/quO6U+RWXC6CS7gZw5+CzdRaulpZraoDaAM4rVOYLHxxglacxvd3ra/3hNS6+VVfMLSXxffg+m0
vIaxT/Q3kXWM9z2JuIK8x2XqMzIp29Bodx6NHcDKvMvDt0DQKzc5YrZi5gVR96GT+AEnF8PQI/f0
fb01/ca/fmgoQaZqDv3Zm7BgamhMd4LRm2UXuhUmuV16ktNKpCmRYzZwjp50vWp4BNk9qC9fbB15
mW70Mx0zOB1g0PReGx/emm3GlA6NK/+r5p5NvC+3h2LJcdMhIhzl6BpQRxp2iUkM7GdkChf32vFY
OlcNg7c4BkTHJzSRW7GQnMl8hkhkggM9EQoDKynR/DJXIAZkqeUQ+/jT/SKuh0j4AqKxTaQ9M79x
aXBmVFBzg5QzeGV0FwLRVth49fhrRYTFesmIaypMNjhH1nfJPDH/LJCPlqeslnQovXfKQpdXjalc
1SxuLbOWnKw0y8E3pwj8PtDutVb+30Gl58Im/8ZS6B3Inwst6LDsvacOwZESxL4giearIsuOkaXb
NpiVuHwL19JsaQtSRbKZNL3LHBUVo2SjRFrAnJO+8euImVGqOJXC39mydarwuG70FOKRYfsa4tBS
L//KB5HUTKXFwayb79wBGZLFRI7UXOjQUFbr6CNF0SXZ/rAqFyg9AerOU8rZN2olcqF1jvarS4dE
cimjJNzTiT7OCl4zbdauybSs1bLg44o3vIHdlynOKdIn1UTgyqeaNmdtP802wDtzAZnGBXKhTdjf
//rpJIA3m13A7OFBbU4xulSHdKKbyDmHIkGfS1/EbhN0dGk+M7dzdoXjRfg1s749hyVkqpgOWza8
PYcp6QSEPG/iOCWI7x+SM0yIkI8Qnl82leojSpreL3qYBiwQ5lH2QPFwDL1ComiYkN3WyWLAhmXU
vBwSq3f32XjJDLaBZq320l1jWuteCAPXBdzc6yls52bpxktui2JNuxrNnroJvgdxdZQPfadN/VPv
a8YYyldPcAv71GnWboITcon7vYBi3p83hDE6j4pyMOXJ2oi5mXTIKJf1Bf+IYumlvPk5ySHsMdiF
9E9b/qLiSyDheu7uLiho853XrxgD2HRznSjg8Oq4Rl3lkfKosuXD72cdxtchFrZPfMmmNA/lLQNB
XJSHGtspEViubOv6RAkOtSxf7pzNVrWCQsCBQZBkYiP7C0+kqHTacH3D4ZnCJy24RLqqa9yxVXen
zUeUuhB5XouTbNYXtCojdzadnORbD0ejjuUuQFNoxJE72BhBkj9lCWNMPQiCFyGFMv6AcKrkbmlF
yQ1CDHZT4/LhoPww55lFvJ45QnaLJEH3gw61yJDASNXXxRIIx77iFhiwfjW2k9m6I5lcUs0CWLgr
VXBnL52GGhp1wgnu/3Psc+PXtVofuvMXdjRuBH9IJP5xhEPrWYRaUBMJieTnQpNFj4P03dMKwZ6v
rBFc/k5qczNDP6wOaOCeXjaMNXv2ILwUFLZ0NoyZWcdRJodaCJg5S0EpNa7ynHF3o+0009dTV9Dq
WwXFzfMMEEvTdNl++XXMS0vwrydPbUl+zc94au+ihQEc6xFDYuI2u28G19SoBGIb/qmaTiUYiTMr
7m/TnGNf5gncjxBfiAkR6dNcBXbp26/md1OL/qLA6VRGSrrtau/cNrgkJOZgJ+kkKEtG7+J7mV8w
z2/matdqBKWDTttvfGyMBUwdQdQ4Rf3EjtRcI9oUFqz/z9iC1SLg9BVWzDN6UdJA+MMeqURYm5CJ
tBWM/VrnA6aTQPDzc6C1Cx/E/xgFyj56CJDegT+YvNkK7T1Bomtk9Rg2CJH3PBpQlyifYUFtFzAP
yzEk5hq1/8i4aL61hT4rMaCDjZ3+tXejGTUx8ROuXwulZOgugT0CD9PXomMf4hyhBfWa9AdeU02e
lrQflc6JBJOVi32wwEqpCs6BHDwnY2n1GUrZvENLVGifb6FnoPje0Z0xiOAAgAWBe1Px3hWhniyl
MhLZ8Z9fFCsKf5++1u6ysQTL6zg4mdXtx0THmFlzYUrzKAhL2CdacWecOH9ORgxFA15WVc0X/6JM
zH8MSv8sLemnewors9KE1EEyjERhjdMSzgr96I3OvErm9zk/TG5t7Y7ZDNWHz8rylV9L/UkLbpHZ
XAN9SvPV7aJOFvlodbCYyd61fnDZZPjs2eQKTZ3KmmKiodi9nHjcgc1At0FtJ7+fGDN84kIE+KT5
EAZ8l9OC6ZMT3ddJlYdpIXffzMnEF1HVpZpKVTLw5+1NgPan3vfQS6jLGPnmqcXPLVu7wI7t3NgP
sCIUOYhY8MEmBPJvrkm1sStMOnyIrO9bKaoloA8e4oLkhrHZMNKdLVo3ABuwqfjTpY3f7HppPpiu
stWjLSVP8Z9Rg1yz1qPTAnP1AAlyypNm1DqAuFgZuwaZAMt+FD5VIK0OmRqrwila9seLgrOLCsqd
ZseFzrrJ/1Pw6qaIW6ghR7i2WigSIGRwKsCeQTFhZ0hN08CWWXVbX+i63a+1tPqv6nY97lkgi4e1
mUt8iYSvk7Lf42g5dJabixBJma2Am5G5uRBOg+nm9CorbETbucN+ArGC1w9UDHFgRguqKuEs8DAX
+46+qyGGEnVCl3ncT4p/UzfxpNBiHhMTwLfKbYgE7eYMvyu1nPjvnVWdl8rupwOuontsJi/QDiRS
tn6KjADpK1ZlhWONX+f10EQrxZg8CQqQ61FcoyYhH/LlUwZAiEjNTw9XcJcXs/5LKkNUs4iDwZOc
Tj8kPZ4aYaQ5cfgqY0PtRgZ6VJI9QtBfwGXc1ZEMoj5eTnvoOEPhzW75aDZixnx6dqZlQDzDHMtM
KGsowmH3dX9TdvNBWwciSI/44UqDhLArUv/RcI1jvZTpt6W8q8O9zeqN761TEJP/x5WZ8kAS91Oi
2kbdZRA8LTTHx4pqJUKdVk1CxfZ7PQLUsCs7B4UwEdwL2PnGd8XGhow6/JDN/b1+X6x3pri4Iv7s
xn/opY825qFPaDF9KQfuCEES3USw26QEDrAGLN2OQPfjGOKAiKIJatdcyypWPJ1+sf7QzdkS43dS
MF6hWg2rxbKeaSArHYEK0247E/v4q/iLtVld2JrSIfgGXETNIg4wRosa+puL8ie/t5F6YpfJ11B9
NuNWdImzP1/3FxIo1p6J17hFqadWuKSTnw/dcTtml/+ukG2W5sEKBh1f+2Cz4KXmDPYhpwckv57G
wlzAOriSL8HYJC+yah/sc0k5VJ7m4w6dydE8hDK0pnJfso61c9RWGKscdDwBJH/fuJxMqr1qFZ7P
LUWUx8Pqwwj8YECd0C3aGIpxuCckidqsr6VOxA7SoiulHiKRhqByeWbwidq8J0evWs/7VKzkDPDx
fgiVdwr83FrBTaiS1hXvbDQl28Xv+LsqyloNgdPqmdMFOB07a7OfF6qqLDKsmpSG0GdnIqDhvGG/
yhnxSB59NdF5vcQLnj3dGut2CLTYgRbVO5rdx5FC5MINIWRcGA+iDAvmAN1FnIhK9UVWkTCfiKqZ
AfApCvlUlsc4CeF2thaCJuBiTr2/zN8SKn49t1KiGHrIiYBUYA5oss0rUrEJ9VNcotkaUBt7zpmh
U22K2u4glMrxhAREYVgEfFv1wsInX6hQYq/fQKeY3841OK+itCI0nF8VisRdyUK1VidcpowwqYN7
wjS4mAay7Az/Vgi7ygEtpAmEA42N1j+APCPtMIJMFvbyfSTb/IY34UiDoVGMjECYrQ4jdctHwhOm
GF2vLwolMj0xc/Fdujf2czcoqb+ETp4h3ohBIDjiefTI3iBF+PAYoSaa+eoAERyN2pXNCLqb92R6
zcs9VyGnhYb2c5nsan0Hq6jKeb5N4+nTqH+jJIN2U7RUTJ+pwCjgl2MUat+cv4WeTeg2crVMwG4m
L1riOmVi8lfcrc1+ivsrVIYz97uzHbK7S4D3gGQUhkCt8trbVUHVAX6b/4sYvBvZVnBcZH9J4zSn
jJuxaTtw6RGqlQNzQlwMlksABWQjaKWLqpoKggNavTienFvZZPAYM26+aGD6SNaMz8k2Iu0mETcI
KUpMzDeo4z+OAVlnkLFSAVlO1Kgs6XA0WK9ugj2nX0gag93yr9oJoydBZHJFJEd5O3Vc/iOW01WH
HNTzbJ2NCJ32quw7Dp+MPRgkMJLJMkid/Qgx2WwoKRh7gR5lEkvSP/B0ydwYsdiJZpZopXfKzw6R
bmq7mnDa/LBWUhUY5fjwK5SEHpkGBNitMRWhPZkEKT9ovdHa6dSc4WGZOa3Orm7AeoRzGH4Ca7VA
UgSBS13VVvihogHzgd+SrAkCSZNMnlKvLPWDmXH6JAkbrQLQosKFx8f3Qa7ZMV3F66xjppoOY6Ym
V5ZaG6FblgMiA6swM44zo9Ma+8QVi1t8X+iX83gFWQ/QAM4Ti3Mcak0K2dMapuX5fcCq7XVZ6ng1
KsyXSn41jS+Cf3rnnG4NCxNkytn8+TXc+8ckeC3UXz7/vLVrMSxRQGnCHlP3/9TIJLV5QXzNV9IE
3H3n3Yp+i1dz2wJmEdWy2fyTuNYTEw7brr7JP1DpgaK80ldUXaWzFB9vS1DS2Qg9kV3W2Qhsp3wB
1OnHCP2WzA3U4GAkAXgYx8vK1FpUSM+jirArNZ3/m1FFZEgu2W3PCrLE6VFJ/ETA+EzTSTtcAif3
2gLGH9cB2q3yOaXKuvWHJZhZYpfbZs/PF8MBE7lcEBoyawxUdCR3Nfmy7tZNNsS9TS89L1xPyhmB
8IazlO2oqtTItY1UzO7LU9vcOxZVU7GmSNrskzE7ccGJZtSGpridgjhzH21kxPFmUquVmuFx60FI
ZoWoaEgLRv4Tm1E/FJ/8+gPzqa6z5TvPY1akqNE4WQPi/uSfjvCw8SSfWmRbN+L/Qr91A1QIXC+t
zrlceeehjZfBJZfDviZ8foRy00LP8/2egBbMd9gjF8UdS1CDmEJO7WlSiovjntZeWSKwcAS9oUyx
WSsZuDlhKTCDCyV6pFnJ8TsH7awrXhKUomA6HQPrEOMksxT6NnR2o0JGa6iaTz1ZXykxpBMyMVtv
6qW9C0+AmBfzX3OcAzaAmonYfh3Fme6E4GWtcQegS8iyNGNZRYAWydGbnU0OnFhVvNgkb7gXI3k+
z7rgnPZp9B2sLsHyBHPqmbYQe1YACkgzsMTCJMQJmocFdKOOqOTO500IaHQ8pP9FldhA0e8v4K/4
N7D5QW+bCFvh8t5Lq6HEHUu94t2CEyWPubtLMeUBCYQunMCMrD77bHMpgoPqWDLrNH3Zmrl37cUz
KwbEoo4576wvKNd1j5leFz0xk2D3rmfwAHdpGEu2d8CEkqIQgIjoRhOkAiZLaYIg12FFxOPaJGJg
1LuN0mXX+w9ltn3GBFukDxHTXmktgluYD+W+34tYmEKKYy5jQRHLzZn4SbEVDthphyQIhB7vkie2
x1cv/9bSJ/9qv46VTI+9W1a1wofHOHqLky4sWhuQ1tIDM9VmmegtQJn3ImMOb3el58o6m/0SOs/3
yZIbsfkJaBgUr8S0Wh9LTYVEunaMfRMP374K3WfiXiCB8+3N3/IBgjzJylFVKcMQENPxTdG53I95
iyoEqwQ01fZ4py3ohDHrQUXI1enUSi0cJ9QDiDYrPqq3Liw/TaYcC/Pr4LPv8A32xCIoMv44prKK
Ti4P5b6P45zYaVkANNcYphjZ10CKB1H2OdCrYRaE1rBqwTFFctnFVbNLyHQJcTmpb0GLuuCNPSy5
WRF7SY5bWfSzsPKN5A6v1+nEyiOcwzkUEfeqZViOyxIh1+d1j+8FdKdvDYYZRaflHTypUPh/c37O
NdsUXIPD3DWPdVobOS+ig5ehZHYce8avnuGZEHxmf4pdfjzToClnJhhaPsBhF2tUzdM4/xiFR424
JLrAiGzwBF75dbIOUaI2W1v6EvrEeTPpwLNynvw4shpIJehES/Ep7uOr897k9egqfNy//zEALzLS
wnExhUBwDPVLMazmIpSJ0DSEJO1T8/88J/t9ovvddsq2goYN998nH2IxeFHujTssSYArM7q3/KzQ
PROVot+HqndBB6HJfNv7ixdMz6UHmfgfy5yMhGVFUnx1P7dYIWeeod/LDvadzNXTWmyJaK3ITcXm
SEwsDsuWJwqrMwuzHE6vLXPm/szIvyEM5tOew7oCnekWL/OGz/0oavoI2LPWAUFkjvPcxLi2Dh+L
wx0xAuEeC6bSAeFl79DiRHdg94DtGfmOXIlTFS0hDCHigkeJIT9w9iuCEm+8dY/JYxqUm7Tk2wXR
Zzo1/vEbTITuVhoq/+V09cFHmubxqso32pwB76xmvl1kofY7UfKMIDm/3C7/kra1mqAJl6h2RELz
XpyAyeUfkNaMqvUmyOEYfnUvxgXSWWD/GMKV/bwTsc3wCnO+PfL87OdL6G4DxK/yoY/l3ocSskH5
/fT+Uqggcrj6lZl8m0tgyVLrg1ZG5zk2uQu6IYxNrWzziS0ddR+S8vZ8yOwOyK6jC9OtjceA/mmC
xZyL1CcvRQ7DKmQt4qixJCSU65iJbUXy7f6bQmf2QYhH29mKIfckU578dWw2ZDinkUu4kmYiDDRG
aq+wXzKGW01ivmLPvTzjFf098RefWbeiog7sCIC59ycPgfz42wJlB4l/MF5xhsPNzyClmCHeDvlp
AJl9q5EVQGZaljl1vfr03NyRmkw/bfBvtiwvDXN2GVSkzCxlMFBgcoVvmYsOjgAxIiVGq+iQS0QF
I9eAgOL4HUk9esiCFWMoQpM/2lqjWyNsrLFG0vzTnNlIP+RO8dw+1189ES2eRivx/pgc/N/LqTlD
yRiu9S43QW2mNGD9+Tg4zo/KUKnpV9+iYlCcCsFX3ZeGR0RN2/9oQFyWCSAzGTNPujINPh2nUyB7
SKE17sjQmsWaAGtXXqUjdK0fB9R6zKmnkXrFOsjHG7QRsZF+371BsvMs0M5Z4iHYfhHtCH8xoIMv
TnmQcFmH6Bic3r2gnrjelusQxJ9x7x3W4Y8wxBUccAjgl8+ZfW+xi8rU+mmZ+YnoOpVN0VHkqcRq
on/9fX6mvPq8lizEqQRRxuEiRWBCI6ljUbygTZ0yqtal2Nt0+1Bp7NtKOlEB2TIrD4xDT6waz50V
3lyfj5kq6AmxEqae1EUXF2id5Dct/ousoKQ85gZDNQZu4sqEwX5ZeaLBpdD0+jkqoTuIlf6qKeYS
hfA/HqnBBe7eYD5iwnESAEwvwUEvoISOyqwFI0NXY1RJRh8W0YqhZuOGu976jj17ruqHlTnxyYjL
VGNW0vVST7BFu9msO3AQqk8m/htJ0JdtJwIKQ0gMZXdx2ZHtHZA/LmU4gonAszsS/3Y1yXGi9ZBo
VoUo2St2iW80/l7qedFDRo6bb2ds7pD57TQWRtLxA/lP3QI6wRkRqb8Y5ygTZAfDNR/pLOeS2jwy
235QRWxMfH07S7ZKq4sXaPdt40cWIvGpFjL5lsZOsKNzQEEWLa3DCPQ1+4nrEEyYygogZ/E8BHr5
76tbWT8e6948YUttw1othpbmzAiRbsQnZnqfwtsfW53CDKFs+5ZJx6tdvGQh7KTjfIQQB1B6Q0Mi
y7eqWN2skoRmap8VQh3JFt2Yult/dfyZlbxTVZWmt7rHcB/7CjEPAF3YJTuLI5ukElK0k5PxZro/
BPyDFQDmweU+E6CJ0R3T5GspZHRvj1Vn2oCUVRSQ8O6LF11CztlZqa9mTHGI5HcZNviWfsSEIptP
+275lmdAsCHcB6Kq0TzUt1JPQtyg7Tt5hVEk7spQXLZ6hkEQZygdpIav9Z0JZtQ8kV4aACAtKiCU
3bzqImPicjxm+dHgFZYsf0UUzNjhnlh26Ac554i071+vNl1fVYrb6vxQqDrUIBrmr14Nv5Gwgyb5
aE8ZULnvOHan8k6X6+x1O7pAN5+l5jMkHk3Ai843zEYVfTOUW0TLsyO1sg762StTPsiZExTZNdPB
sTEMsAT8tJ2Rx4DJKWHVjnYo1cazRbEBgRVO0S1M5fkleLxEW9jyatQb7rfK6b5kMUco6dit4Lf0
UjVjpEjGrpDCWVtX16hgKU8PlO61MEZJMY4xlLGjHLyHtnfgvfiKLNAYqJ1s6pinxnRwxMG7mzAF
y++ytQMmMZYMDsHU2px/ETpBMryTuKgDchMlIZXbTNhUKiNDS/6qkT222yrNNKAWtPhb+JkntDrM
fYNcOFibL6gJo62L5EX5iIrx13WWBvBbGs+ev5ieqllp+CEtgG2Ml8vhn9Zc0FDxCnPbKBdVVWX3
FlHoj+pHmOKjg+vKxWC3ffBlXotkLlDQ0t8PEtRKrJE2p9CgzBCyKtkFe3RdHFCIGT2N8UWvuEO0
X/ZCIOpQda/nTivHaBMehhKZxL9dABXE38/G2QkyTSUDWIRjs1hlwHR8m1QaQU0f8+bfCZKwh7Wa
GUkW6xzOdaSlQnx0sYFY3NtEWFKmFmxBrx0KLYN6YF8dz1Wjg4TFEs8ZxPz4SyRHwbfpc5UzYxMs
Ncy92ycrgDNgR6y4WODiRkoPsc0Oc5JkJO8VyNPvDN4P8GMGTOiycl8sq1FMxCpRzWC+jqrr8NjD
7ApnQn0o8SYh8R2TVhivxWGPFO2ZW/EolD/6RYlK6FaUxjtmg66gcvRAEg7sAnsOJrvpGZnD03/y
OytQIkFkMsqMas2OYCEDQVfEepSXI3aGIxeKLzUfv0o8ip7Zw6gEXJs+etzp2rRY/DM+B8LreAvy
MYCJdwjhhxQPGd7ctFqwyIDbjNuRZ/sNUg42qokd6hbOfFjar+RAlQBSPtsz/LXIX8vHUnvw99Eb
C5mrxnjqVUGQsGsHrAZKgCKce8ANumt/F5AOsz3Gir2GMJfnuyQfK1z3Q7jMjCLaPyPje+swiWeJ
328uNhSG6T3JcInPsGAf2OmI4EN6wc+BjVPrXbAyzQwRm/ED8afCTCmqjYTbE7YaZVzNnifU0Nch
cfNQsZP2CVV+xpN1hPWJu6GHor8dMTZL7vpTMFPOzZcickLkm0eEIwlYtp4KuD3q/ylAgO/xXSta
LqWoGxf5zzYcfE+2a4nfr+xsHKBdXG+5D4fBG3lFC+A2yBwuH6Z82MxkU6jVBF7+12E5FziesnkU
rHr3/M0GD8ixRD65tEGbOhRqD1PSnj8nNyIJMn8QfNSzARVUBUsFr7gtv7hxhYmzV1xht0Ru1Of8
4L2xF6F2QcHRDoSDSFF/IsGIKvRRDubVN34ZzP7rMomyd+7/aZGzgoMHdUhcxj6+stySimr3pGfI
tlUtQpmFsEYDJXUsdWTvq7zHl0oujIBRll1Fct2OghZu+rrbbE2JzxkfZhjgisEf8jVYc6jnbjA0
XxYyOQV7FFZH2EPiBD1WE0v03QgaIQyNE1zai9GMfnVNxvXQVEFDuXiZlWRVEpxj736QCLf42u1d
8VP/29q/3F7yzVn/yKhvaRk0QfpSX3xns+BP/SfhoMfKUHhXEH84x2UPVHD+5KLzun0+8nSOiOd+
8xVedrfxAu4ZK71q0rhCUEPwMsvmQ+Bw7KUYYcT6F7i79tROdUJpk6VIaX6o1FAQ+Tsoa87XQkDU
zUeGBz44i0ewZcMrvqSFhuwKgkx6CjF4WlWFGOn3CY3VeKHKktxcfFdX0atBMvG+9Mm5I6KtE5Eb
+XSlVdYdpatXwXDJI1oRo2RmxSsi3XTr2MHLkvL3LTYLiwDKu7y5237ZjKfAkTXT6MphbwYv+cPj
mUvextq/MVOSfnZP1t36RTDdsHL3WworgZidferTT0apulncFc92uWUzBfZ8LvYQj0Vh6GbrKRqI
E94zb+2DSnKkmGNoCAY7tkitPktfYjVGFX0knNZOLmU8R/ES3E3QMFzbgRuAsN6jghRz8UFDGyhU
pArv81xkWJCj1+rY9k6kaHqvvEs84Amq/Z3LbpfE1kBheBYxyt0ISVBqaiOelEdYAEYxzSMwMq7R
56o9NR8zgjgL/FlpCfao8T7XShcA6iZvGuanrOw562MhLXnsHPQMtv/CoZvXgLw3KXnraFaACsYH
hWUIsR4X8qk+OcyfWSVY8SitbK1TvX5fGEkGAN0aT3PvpcitvtHhOG83CaO3ACIj3LiT4gz/IGCf
FXv7kQb917b2fcTrS2j2kaBPtbHM98aWOJ3MC5fIzRvwY9H9LR5Zj7rMrQpIRd1UCL9Folw1vPaq
OdK3/RYmQ6ASN2EaMpuUP7X+kE3Gh89X5fEWthADhsd86Ydr9vSDC37/tZzP7UnWWFXTRi3NxvSU
1c0io/LufVbQml/MJPYeejjjYqNRYmAqMuaFL2jJvyaYFUnGt/1g/OUsiOXMy714q4DIPiiDo9AM
1WGUzBMyJSzRlhPtn4622lN1kZ3y1okXOThNnbRx3glfpfRErXTdZxT+bboiwg7IdlEcClShHXpV
J5y09/gCfwV1oA90ily2x2Hg/8GfTFRPVlA/AjjA6HCU/tMyVpTUPgdShnPN2bopWENBsbXREI5N
8pYCyKEALeqWIhJFD8BiIoPVEmC2Pb2/66aj1IxirqsLaKmR/CgdYiObEwpf3kYn3II5bh1wsMJ4
iCvxdkkHdUKzep9Jxe/py8IasKd68YRTrAfIadQun75VroEEP3NQyx47KO3ZBvOuN0N33xdFHVVy
+Rt0RE8+9uBnxG0hdg88+7M0wA1zImy2UB5G1H5z0BGf3ZVWhqaYwEiCIB8imZSe/iA6TDoYvATr
K/C/DkQWweO22WMdyV82lGYd2iLuEZXDhVOaySjrGgLvetvpq3e0nVZRzqqe1iBWBF6DcWB7hPt3
nFe/iKYL6tYLzfLoYGdbFBinnmaZJM9C9To0opchFcdMdSye1L82Su6ePuNh4cHuf2dLTfUGrHyg
aa3g3ZFSrx2kQHWIGUByi/4w+tWcboinIRNg6OH02UQ6EWcyqZ1LkyttmEoGNQxrcyAEEGprDYTA
dEFoutvI9VwRvdRa2keIXlvath5RODU3zTUKj5QXsAE/usspnimUVM5VRoJ92jkIqYA9ohAFU6/h
roPbh9e/VahgMOMhhoCXQam27lgkcKDHc2oYJVf8WWpgg4GVYCa8Y2B0L5pGUtnSsP6abRDtSKFL
DZZoFeOSCSJj31O5twYl0dOOyMsJ07LySdoWk4vP/vmpX/yDZop0g7qlDXmzQjfMwFNVdZQiadP/
smAuHbtntB6pTAqfih62WT+pHvJV9WUaRGZVzQDzomfo1Mj2w1vIt/zwgydeZ1YUYnQMh3DtSmO5
obNcqYIf4cdqOSQyKEdFOqsJIqsk/zroUMweMug9Uh6w0H7OPQmsF3C6Xd0TsGFGa+Wk2HHkzQ4l
O/TzE0sveMFkW38/e6/lGq7zxisg5aUbR0BMEmp6UT0Y2YG+yQoFa3a+qgrMtxBVIYI78mTl99cG
+1mIcDpAKK4S8aJmhSgVlpYHXFpDrve/SCwhr0pIVUcE1lMdJ/jK5FnVLIRntJFvMS6d90/1RJFc
opQFT8RDqWOr/pNKLwNlyZXsYDW1NblTZL6hv2ybAc7oE7dI4xsyGQ2EBG5EadcOK+gKjFOSRcak
9Zg/btovNS6/v/UTtxgfnCl+/xYkWbZnal4OCh04ccLNBhr0EFYQSoik6tvA56gT9B2TuqBCCl6B
y1MDizWYlt7htbUJyhqYm4b8wWjrNIjzSYbd5UGmNc9zPS8/I7Y9sOLjbtbRWLsghoHs79LREIaI
VmNHBoTbcSzG2apTHwxWz7rWJXwviuL7cY9P78KX8O6fC/vFhbf9woaALGNirKT46o5S1laY+X68
eDcg/FA22VV4d3snMEp8As0vHUorMnnCzFdyZHec1tNrT9dYBvyHjfe+DoYSXVtOhauwZdBX7hX0
8z12IE+ABYA8G6BJ9/HiLc81F5ZeD0jeI5EGUyjzVe2JmedP3kyP8T99Mvl9Sp3ZNMCfciiamdJz
m0/ONmLRHH0ZhxdfdZTkC1FBCUv5cHqB9F1P0Z7AbnMP2jxJZ/Kn1m+89iXV8pUXAQN6JkXFpYVJ
6LkydfQaA1KNnOe/wUy+zOxqGyxlAkXI0K33KjmEeqFFhaHIEOxVnwZs9hxT0f1YKpcheb7swpjw
Y4FagLlNLdwfY9u7NobtRs2Wk87SHX3wf21pIPc9Ekrv6hu/JtWmczRkPMRfKqnCQGRRCynawfcx
yvCT/GmymVN3Sx1goo8zBKOE3KrVtkdNj0+zl4zIuTKcfIQEr3b0FKNveEnC3VPHaHr6c/EmOk86
3KQndhtD6znNDOxfCTMhyCihGqRv2lKV5Ap/THdtNtcTZ+yM0+C3fIEaSe36kvi/5vpGATDrbc2I
Y2UhU/wI39tRgy/quIkW/Ku3hDPdoifzcDYgDOe4vf0NwBfmCLoaYt7L/E9ZfKV3pc4f5bRLz3xY
KS34zbr6WdjF0/cgyD011I77yOu9xjjOoyTi0qL7fOW2T7dK8ZCI5jOMK7aOa/lQ4F2t5AkmT9tL
35EikBVa+ONwk55vWMxD1c1ei5loaFBUIC8qr93ineTiJeTnEET1TJ9R08PgdcLgta/j2isrFmkW
zNdMtPy6RRo+prxfYMDrVBQ6B3q1xp7mgINpJ0ikAg6PRfCtnL8hgXYIGc5cCa482KorG4JZIoGl
v35m0aynMgBAa5mVqsSdY5twcNrcXVyMu7hckIZ8k4roniuOX7v3Wa2h3sE5J8bkKWxo6CDajJtW
ERIgCOIVPMrxzCn2zmoH95sIvpqZ0b7G0spPyjnwJiuG1Y4su94gAYQOUNHQfZiZZ/5/XoLNz6Xv
yxoQimBRSuKPD3o6WipX5m6d8Bsld6T5gmtVsvmhkwTL+plogUkapItulmIgyX2N09TInAhVOd5o
p7FuAxiS6CGaN8Cb+yHq3f77SFQuethUQxFkQjhGQLSob2lWVujY2FOfps4NAlfBWHVC9YDyZBzE
alU0Px3n27U4TQny5J9tmdTp4OIXD1ic0VWl70gU0jVpUt00SQL5iiVLxzjK67I5cz702T3l2Uwl
mDw384/zKdQfQTWpwoFymiiqlR1jJrwsUhNV4Xic8JFkr6muPEzlbWlrxn5l6Ki6wCIb6VNwttK0
3513IzOKuyn3VdHaTg6qKdILegzGGflbPyLMTVk+1oWDKsO+oPxFZK2AYRaEmSrXjxCa4vPevq+s
0rRTQ+LlwBsOu/fK+0Ybc9WJnm1VypJjf5g=
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
NQ+VUcyoS5XGYdik7/sh3bYyfAUd2VjmsIQtuYjVMNH/J0SToRKLLH8V1Y1clZutb3vnsMI7LZvU
wJG3nJNmkEm7TZcSq+QJWjxn8VfSfmzB0U56GyWLznJrgkHZgG55E15MqQ8UPdxtKqe5K/EgUF9C
vMyE/h6adcQffmJqx418wBN5R1BfHaOMxLtlySrCd/7b2m1VS1QZ/eJdcE9P0hZ4D+XKYHbpW1iV
tcW7Mj21cw7csEkn66qGv5sAMWMp9ebuVlbh/jYndZMWuGkjY3HfhirLB4YHaXafw83J5awnklwM
+fSMH3sZuHVFHJrkqj+/RHtZPy11w4iuqBDZiA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 6400)
F4yzW6dFmNtF19366N778YaBEfjlQz5SznXpW9gnQRWYHUDphCbEpcUKyxWTbCTNlkyfpiOydIQA
IB9z1TqsG1jj49Cn4bB7udhY7pn2hXetMHvZZKmzmF9G6itHpcd9RaQc1aJfPXRx4g5HN0Up+Mcp
A7YCQ6nwWnCa6Wnmln3R1a86/qZn4tdxaFTB9uAIYVtQ4KulqhvOD3GGQR/XzNxEUTzScaBW9t8s
Zg461fGcTMHXDlv/ZI70bLy55s7KOF6wpDfeqMG6y3xJjJmPeScKStsGEE6msQW7q/apQX1pIMGh
hA2z0GFpZPoaw3PCiGsciRWJIu45ftTDt6r3OTmP6LJxsnlSWkqPSWBLmOVoufiYzgqPeZel0vjp
52OrtOkgGDvjksHxMH2NYXmOjGf/iAnJI+QQSfJ3819w3DnHbtfqE8kVojGXHy08CXFLIpfcH3n8
AEokkXVoWV0BZ9g9bkrocnrNRP1vzBi+ekPcXJXCbDnM/x27JX7O9no9g+eYu0andRCjfluunFAm
vM+BTIk4bF9LLrk+tk5xhX3RkMG5L/kNd7TFdiHBoJjhZ0l2/QgOdvC2dH6fUjQVQZG+E+U0GmGp
OjQlx31fVvBnqUSgEOqiO4fVvdq/BxW/DCg3O80dhfF11/baoWz+CYtMQHJ6oQatiBCM6Ng+vpwz
SDOAUADe7f16mMziNYVN81vewOjtf8b2CjIVZQF0TQA6Pd5OZSdti24vQGtnc96AqCAk4a3pRAXj
wohwYysQ0V60aETWKNhxSMRiKGvKStfUs5DS8ZcBdzxPfpyXD8YevZYXleEvqkHX2gYh6qkXW8ME
U6rz1tu44hDGscdYcgluZMyp5QjETuY3Sv0nLXjad787qx/FCjPxpDsGDWvamYfMlQ3G1yX4zUFb
NSNxrVBbqaXr6rBQfCxo/EN19TbMuQyCiUhlJlmFlOSNihWUxQfzFMmb+Y5EsHL2KA79yw+VN51X
RGNZ9KfHtCljyQjwoPBqWkaOAZqr5OhPUQ+3ESz5m9qz4whYr/zF+2JcXYHzznNKsT493qyhIcpk
A3fDBYypFeNbfjbBVofEZAYENQ85aY/B84ElpVDF0vB9xIwR/dj1Phgpvj3SbNhECYIhedsn4cLD
/9Sm289R1sChhYNV7pi45zOF4Fzgfn0ZAmcQYryBfIPPz/Gtdtjv64ZEgneoDrOY/SgmKctBoT4s
U82TBUrPwtPqjwsp1NKPjtRZhKsfC6JOwV36XcXnsquPWikD4+kJVp8RgNbwDxRK4Y6RAyPz/Pbs
FIvZ4PwoIAbdgVRNXYPicjjebh9t1NraNa0eg8iNudi24oSHxmi59rFk+JEH7gPHdOKbR3/ZXugl
ZYHKobRNMWmMmdB4xO1EqS5K2rymD5GVD7e+fDtTHMxhsLxLcPgQlTwa2j3/f6kncMTbXr379wQc
WcKhM0VoZnP5arNRC/2EAI080WM/6eNnt5P9NVYK0h4l+0pIdjLwqNe7ccd09C9mLuYg1ygdlwtl
9KEXbkA4b2NsxEzG6BkCK1sKxf2C+P6pelJRaY2/5GjGpcegrhaH769/O8FlT0aDE98uBVAjM6KN
I918n3c7Hd0fx6mWgSpW4Phtx0JaiGqPzRwxVNd6yaGgDkGePqn8ehcMLhlaj7OQVRo13/EnnPlX
WFlfmOZPAja+HJtFgnwQk7O2MaCY4MTqJPlllbiYPchmCYdyfyitO+gzq+wEv615piIX88NSxbUP
71gCuDfwmqP+aQubPcC2V3WVzTyDRA4ckxlaO1QsYlWRSYn4W2kK6vFGgweeAtYWJkGVLGkqFU0/
3g96XuB+VbaQeC7myx+pCQc/Rs10rJXNZ1RoGO+U/LY1x5Rj1sRXvDj7uYrQ1nRbd5FzzmoJkeSp
gzokloAMKXWht2nqf0ADNM274AALTBZChLc2rZrQl1VmYoLFgVjEdyhaBPkGopXp7TyHVc+rVjKa
mZcIvjj1Dk5JuyilL7bH89ekJgxvglhjq/mWVup/Jy52ogYq+cmBl5Lo9t3U/7Fw7Gq0Fv4mDmEl
M8IkxCXsopuk8zMpQix/gvFy85DkcTt84UyuOt8cO1i2kmOB+yQOnj0elQf/ZjIuVaWWLYamo254
sU5Ossaf2i5aJFnETJDtbJV8/hSGRAOMPanlXc73SOMCpu/heTlAQCTv+MMmXkWBzTVtflWhfpQ+
TvDINLoTp8ecTxrkKSsp0DNlEAeZwaRXurvNACfIJI6DIcl3YalNpJb0LMsIozdL7PXJV6Dskeqx
FMehBJfuaR4gA/iqvCcCqPyjeyP9d4FrOXSSL7s+yNBdHjKj+oIgAMRsH+z+qfoipjW7uDup5gcL
Jxtwma8ifWHFZHxWm4MTRQjTIsylEDyjYGmWfRFffVERZ/kbgDFRycqDnz/gEyNRPArVlT36DVJD
oUC0yl8qJHiPhitfUBk2WKiP/7Si+rjTPbqrapZiUygwJzj8qYRdBVcZ5i6WyyP5lKj6vNegv6/l
TYpmXb2i009BfPpS2uzTlFRXk1Sszy4jnytBOwvBYaoQL5FjZYGXYS956oqrhmhbZATdttCyzjUp
SRhINtD/QCJqZxdpyj3TCntR8eIgi8bYpwij6cGFM7IlTkF54UCdDdk7HcUgWENk7ztuApMMsoUe
8C2QHuWfyYTn3C3qXZShncagEFXoQfPxXMqKD9Cr4zLG9DXQtSoBUN8sO6Qb7bOLYzoIPTko7mMw
HYVcZQE69rGU3hPbpGwGWDOiA3JSBsxr0scmzz6eyxz817+a2SCybmDDDtoBKp230hgGOBIeIC7F
rXQm6lt9W3SWQ/UOu1tNz4Hf1ycwAhoYV1niXGQDLwcnDEro1T+CluJNc/N0LSUZwDACq7qNza1e
SX6G8+8nmIK+I9V+FcqgK8X4XWH9QcsaLY2skj7qaDB4HJV1zb33Jq80aWs6pGXD+IybbRL9ZQMt
BIvfy7zpz70yf7eh36EtZINad3oHvQGs8nrn5Te3QHZ/rQ2G5D52F6/o/qq+LkXEK5xGkz8Zw8mM
5CB9zQ8emL/XMB1xz0n1CEsN0zMOdWILBLJSsPQDA4pQoGbf68EOuTNmy7K8lVqNHUB+6WPcb6qn
F2JmrO3QGBL2glCrhYj+bzAqHTjsRtd8c866pCnlS9Jol6KZ12TzsynKGpaiexLMSmFsFUAYN3BD
5KvehnMgfVTTxqwUDGFfc5Sf6z9LfaVpDM16hYl/l+/qQbvD11QxxZQq67SIoaaTmmqh/VbKceID
HUTOwEfwUIeETDO6Mu/6pgFjS0TifJJQeNekuAnHHb5QV8zfwUPsbMisCdw/xd6Y1zHh4Xy5uRdb
EdPbp7aKl2p8EIW/7OPzzrt1oJi++iS+gcXMJua4cinkuGfQRF7FGXpAjB0Wt6WVFtT0GXdkw+oH
wbWpBQ91vieBonZ2oBMd9hIDIQ06h52g/wQW2BwMJYfnh8XwW/Xyk69H9E+Ctv4r3BOEC6+ZgCjL
78nF1CEP+KWxUc/qLL/lq2Ilaww0eLyJa7QuNp3pBUazyZO3j494EC3ryG3oXeLxoCxBbtyQsziu
1H/k1e7wLhzNgiYO5wZgZL9U68JWws2rNBq/8og2XlN9hapAwiogYNJlvYVAggAL1O0OSRHUvV2c
+3kK0PYRJ6nCt+3zwnSy2lUs0YEpo3iMimpbfl5TxES1SBMpKKXao8KqwppTMOmI0eIVU73TZVnx
iprHvflvTo8HTNeVbtOALp3lB1HT/xPtIV1nH853MF/eSkoM6EZxEk5MHXz9uHUegyy6xilfm2v2
jk7RaAf1tcruQ7kkOaHU45svp+SAU1uMXJPhCmERRiN2PjtsMkZpAGgJBmxspHrzQ0RhNKAPhiZd
A+Wc3pMwcdhndxjqz4WdymRCOfwHPtL5DOQaWxEMQzoAaDU+inYhyNXmdGAHhmC6hR1KqvNJ3p+X
mIv/i8VhHAHhrflX1x3Q+jyjdHHaYbNz8ZOu1l7UYyxpkuh1hFUndb5vD2dz8mIT86VGK8MMw1St
5LlamQnZ855Qo9nFztbQq5H/cnWg+sTFH/iyysBwOCl4wP1RoSUSybwc6oOyor8u35p/nMFkCiKY
VpgnfQrCoDFzNXEB7+e7UfMyuM+I7xvFeQ3nIVXaWmya6iD5oYDa23qJSlMDa3ueZbYxrWUD0HY8
roaJ00NLnqpKLn1tzZV22zSthjsBvzbcoYl2jQorr5tX53gBJ0ceUm8CG7FvzP92lITJhX+aMtDI
vdksGytXCG1u5OgXqM2UiTwTdq01jb0SRpgQ9cl53oAjMO7Pxwk1NjQzDYqVD8UAa3RSnKdkMx3l
h+GO7ooCdHhQ5Kp8PCqBarudAfh057nZwiCyXzqt6jos3zHy8rkg9vNSadNvS/Dgej0rZLzgHpTy
jVIMQu9piLrdmSnRYvXMtbKOpW1nz3sIecS2arwFMBk4xohUEm87cpQEKt7f24cOdPtIt1Mvf8wQ
wUp+ilnfWAh4F3OgTXeI+Wvh3n9yxbK5ZZSe3hLQVXSnrhDpgChR0EhZUE1+FZJtftDOChVcNlma
CL95iaHQ1BUMKVlYAjvjjvlJ8YhUeLvfdBWERFYBZgwJB/vX0tRSehArFTfkaaRz4fe09N/fKslP
6h0B6BqoZrYdGIrsvkg5m5s/RovSgv/QhTQwRgvXLOrioXUMGay+esbDRMKAV3uJeGvU4Bm8dUgF
cpdjJa8PyV4D+83qDBlQTSeB0xeRkIkEkmT5O+Pc58xvac5MMIDaTR7dhIrbl2JC7mywSY9uF9WQ
siF2zLbO9F56A1SmfWCLfJH4UpC0OxtYG/FSogmh0/5f9Qivr9YjaKykAA/96uI8Yk/waO7Sf6z2
wZRiGEr6pLAef03kw9fEtp2HIdVFSr71qsKbjtYsaqlguhT/96/hTVFBGQJmPMdxt23Vv5NnhqgV
l/cR6KaC6Ea68+9HRijCkH6kYw8/Q7vwCGS1z8xl+8bKAygmHdpUB45x0/YtlrnhZ1qKY4OpVZ+c
3fv1i+hjE7QR8QBi/GPOO0PhQHPWpuW3s6cq/SyxqCkBFB21axJ4iyDToV3cL4/FLJZD1Oip3zvd
lPOp+hmu7+2c4MO3wAE7H1AIRuCl4UlI7gocEBFGVIYVzY+ufranAygtT6RvhzBHHBiFTaNMdeCr
hgJRRII9qtxWSltFSc141oJByLt3PwCcFaB1avk1qYEacmzL4cOeFkU4zOplxuZlhOBweydV8zKK
z+Y1QfhlFdhJ+gipWKHA6RarSvicMNLEd3rhBoqId9I1AOp37xfhRL2qWRL4kCpH4EL6GnRbFN9o
0zhVOcNa3QRM5tLxSUmgU+Ef3q77yUv3HLzavrUPCqSB81c/Qm6Snob73vKifRtNvjST/+8CkF1O
uC0mb8+cGFD4dUF07icYwC9gVCAjyC+1Teot9i11adoK7Q5U8V4wktoWXgZ9NvkI4yqlaNiCn3PO
Uf0J/HCXWt/tpXUKUgbL62y7w9AdQL/EYLGlc9nvIfmCJqh/0owWO4XNyufLwynzdbS4P3PbsFgh
aLMVlghvaWolNHLOxQwC0LDvjtXeC7bPAVsEUyS+wtZjQSjp8nA5lAnvwIIpOexaAeggpYlLWr0W
AxRva5GZuzjUE5iFHe8FNcL96vT/eA7HjeVQ5YhfYBajDe3gXbOmqals3a0kkcKtlEOr0iKg6lox
dzAq6QGb78WxrT/C2iW9mbFLDJQ3qvuvQ/SrazALY+vPQQ0XMJJFPbJP3lYI+Hicdv7TfbCnplmO
GalMOAknorYR0E1f4bMAon71NUx5dTZYUfqP/WwzMPoyu73j33b4WhBWEPqt2Flj5+ruQM7kWNJl
8piGOg6Ew3yycD/ocJgJBXBiGaEIfi2ve2T5VYc9QqdX759L4EfTFCwpQRQPRLdA8+e27Z1J7qbq
XXRXZRka3MoHTvrrFULpHn98gAcYqRHnWn5SwFTHZzfRnwSgkXA7+3ymhL9BXVcu9dfs7y+fPhw3
V3G+dM6vrFHVRsyyBtq5fE9nvL0IlJrVfxCBXjZlIeis8vIhSZaIRmVrjFrsbxT7W0pJaVSeZjRs
VjXaGCV98GQ+1xgqNKXH1XooaiSPgwFHQgecKMBA9XQdXnHRv1JRsw9Bu2+A84v1/eqnyK0mDkLF
9SDiRIZM5qA9ellnnPePyD23Y7Msf5kdCZCMttftT5B4LY2apWJ3e/IavrTHNgRvtijNdhFTK98K
B9FStTWYk18RtgKCSLCQevCUXokyYxFGBND5PIkWgDcj9R2iWdxku//cwc1BIBCYu1JuPkVfKai1
sNdXP/eEWG+mhGdtSxPZu1lxBcibpMRbRBskyDVn2mDTC55SlF+OxLYElymDolzzlubEW3fUSiUE
4WOu7ogxZlEq6VEjovU8Z5sgyqwwXlVMARNg4hkJFxJ37fY5bcUYqqUczGx3mMs4x0xnuVGgGVyE
TRjNLIaH7EqE0xWM+tFYr1C2Kca3MXYNDTVB6enNH4sjeqdaPHQPjyscK28tEIfXv10anaj1dWjt
0erUz4OZ96mNd+IOs6xJRpXjdBBqIFZa8umndKp15OASTyk3g2wHhEtMXvQZECrSkhjO8G2C1+BK
WE3YEAngp27qRJr9dzdxLYuhGE1nmIPEsM1lbiH0dtV5VysaiBDqgwtPo2BQ18aYSt46VxQ9U+tV
mupvMIwH+2zuaAQ7uAXCYWvU2Qb+Xj9tjAYbqn5X0qA8HCK9TGz5cAJqq320awYtjI6EnhmirUgO
AEXjk9pVlivRG8zJVqJW0gDZfynSPZoJSi3ltJEmLHjAiFbXlLkc/Ve4F/cwp1zXMISanK1FKCF6
erB4Zyna50lXGkJK4ijE6z48EItiJbAWr7nz32zdh8uggkFGYsO/2+mlG3FSp0D+rVsQbQKTg6nw
+rc4wD/T/DJzcWo8LdYh/LJGwORKfp3mAc8T8Hd2NnX/UYnvgXSkEllUec0CAckAxDCHxlTbsPRQ
ie1xTxidEHm7Y6mLWQtQ0ONXmonlZT9PN3sIcbkPVRK4Jbf7WDGkULk065Kss4uS7S7efE0C243K
YJBd/cIv+Yntb9I+Ab0dj3Ol6T9yVYVsuhsO9Lpx6mUhDE5IN40m/0Oe961/k7lbvhlIH9AMNma3
j+dmXqJ4YpuKxkmCh/2bAbuGQ7KLn/bG/62+GnILXLJ08IuygmctVKjxef/ezC3s5JxjWlAjdAE7
0e/KRyOjVQi0NesUyJZ1tmNzoZV9mrILV36ESMZonqh/e1WZfnj82oxYe0wpUTyRMLRIPo/6zUDG
elk2bkALrb2S2VU3QHEPZOkOixitDrqT0Sq4QKz37MBURdCOrPiMNVLcSZkKLsqub93QcMPYpRTT
ZXBTMd29S1lZoOL0oc8dZs7MilLi+MiQAwe5SEKJlhhur3ntG3JlTpyqIaPfKZLS6vnE2DFjdHRz
bDA01WGIRTNGLjr1RCTqXC1dxC6P0W8nDN7rKvSLpjjhJkRNuW0c7ay3C7fRLoeY0eYWrNNj4h9K
vZ1MffoDfiyqjxA9yEmVMi4XNVzPy23HHDpvZfBgNrW9YiDOcqbmy07PXiwIbPCebH68p6QYzM3i
EhvHbgrIvueifc/VZh4qh4LKXPh+br4eUJo+eYq9hfri58XgMpfvnO5YCuGGSB3KVQQAdO1vn8vc
SrunLHAP9e0giMxZ6fGpgEWWL/TTuondAGrojmvwbB4ynjJM9bVbPqf2T6sMcS4TE6LRcuwK2LXN
8mr9pO33+ItpmBzhlif8eluglQeVVrQQSEo7fN/fccIXWlc3ybvFyp+IEtFS3O0Ysl+0hAju1mgZ
tRxc3ZQcIR4zdYei9H/nbatldEQd+XO1Y5NEr0OFUusFv5wJxvSdh/708biVMx+XiZn6f8wjgTGg
9faRl8JqJs/sQt1yvqDoSQoSG7iFtWjlFD6C7OVzoVczCaAC3a1ARR6hLARIjAP6cweRcgT0kFRE
ixiKX7QZUTui1/kM2NHqUMRaja4dsYEJjtIaudqXi2MwEw4uvtgiN90fyDsIDQ6q4pBtTa0FIBmd
cwXpUbu3kQKC5gx8zUUaXa3bH6+syf7NvOnpDuYT//t61yM5wSuCxJ96h3CMSNlovQ7U2ktRPo2N
pIBuSuZZrgFPYPzhSm8LEYf7NO9YgaGaJtKIg1hWUmUgGiCemuNKvKLCC6rxCTL0ixBMXZJaipp5
thmKdEDGWdI6FHz0ZH+y+bdL0dUwwQzUPe0C/PXIiKqYgs8WUhmMqCyb6udUWVfRT4yLPDGgwAY8
hDksGyTFLcN0AbZfXZkTjrX59D7GqNNb4JZYeq1vxGqSDC2LKiQA7dXCTgiCiPiBkokmalH3xicW
mJaSSyD3WkyE2FURl4B0L0uEZeEqeSivtDB5ky6ZWq4sjbuRpJ7VNF2az7ND6398drkbuXvEz43E
DRiykro6ZnnQ2gO+yunidmny3F8aULmiPYXOO7ZfkMqiTJpQqfseNH3kwCikzjHXtebPoPf9shQO
xmzQdQ8mHqoCGEuxrmAlzg==
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
kxrYa5p8vjBPvkiY94wIPl5zfz/TQgWKbcVkf9/VWX/e3IlBUPrjBC6zfmFRwS3+
KmuBmhWlQpAoiu6N5YYIMhW3uLi6yHRaiI3jy5gYfXcv3OnGiQbcNiXI7dqUI+Mt
TQ/ANaP0fNfJK47NaiWVvrHWn1FTCJd30pYgwhh298Tbm3+pFAlGztpCLO/qmelz
AL8W2S7xj21did32ZGXniqbOuyD2ClJ2XFCfZLQ9edJi9nIVHmgRJ/oAggZszpFu
VNp0u3YYYZ1+gjHuAo80IqNgLcrlrXEtJC8b/GYYAB7Z9jZK8D67+OFm2cS3qm+R
tR4kaRG229DOm9TSOkTdGA==
//pragma protect end_key_block
//pragma protect digest_block
5eG4AmB1B1RMdIr0yhDxOlO1T1Y=
//pragma protect end_digest_block
//pragma protect data_block
sy8zufD0gT+YZkjfyjIcWGbutcDET9Cav7lLo5XwXVdsxCMsRVti2/meVoVTBtG4
Ox7xgHsNXaYkE1/hlDlHgU6a6KeTsmJAGRq2ewn+l6s0s4N0LO9FNH2JDFqCP2tP
M302FS9JAGcs7SRf/QD2wvbAIM0mltGDrB89rwge/tBJrwvCYTxux9pqs2u+mp9e
TXUNL5ktDVrh065vlmNlwyLy0VaIsOIhfcY9NJpxgEt/YdQMLnhSzCBjtGXGZ6cx
FOQZ+g0ZT7bDD6Y6ioT9GYjIMLD76Sxo+Vfy7/gQMmxQAWfP15DHGzHrgbOakrIP
Up6wwGJXkQ7lWaBdFHLG9MCVjZwDTuw3I97QL1bA6pVXQ8RrzzVxSfYiZG71rqID
yvERrJzPX/GwtFXsgILmzTgBs6nATPNNkXd2aawXuCptf4g+sm6Dk6sztpKYoMyF
D3z6Z3A4R8XSjYpcdhGGwbr2+RgZVYCPDQLAv8wvOGO6UPlGPI7+36DLBEuPDpy3
pP8hS1gX17JJKsBmyf70dA/MnX18s2wjmVU1tXK6GJRhJT6ffMzepjwIOuU5hB+7
FLoNRV8rsAgJ1pBGpqqQOKoQfXMXEFUAdEFXPtecSlxD/dkTj51nekBk6skrxpPA
dWdC5to4uPtYKghK/1A08EybWpBXrRCzHe8OmzxX3X7VraEtrz05NPbcwt7VfGKe
XwSZdGPcklWVeAopOvwktcmP8WUHMuNICpOdJKHuSROhuE2yBiwMtSg1naEL00ES
qBHqWgWGz0fpeyuGHx42B0XEw18Gp4BXnvmnbCu0kck1++by4Da9GshCJAupZyIc
4r8FDQtUv+VLSPRINTBdpYiDE/CrpVcjdHR69P8MWk4f/elIKQUL8mjhwed3BQhF
tmXXuV8ZnsB7k748r+j+AAVNq+bjC1QQJo+KMjgRHYiIbw3bz7n5+bqkCMWk3C/P
PVTz93E4f2Oml+cN1D0T8Mzj8XhLcbfU/Y7q0NVtWrqhrs06t1gXhhNU9Zh1kJ0w
Nu2A+EEtnkfkEjhrjTq/U2B/X/CUtQXSZuQ4ovF974LSWi/IUdnDvh/zZzb8uGai
hqPCdYWReox9v+1+8o73q42bG/FN/h2Lwbjb5u2ZRQx9TQNlbW8K2syltS7xxEL4
cEmg8iITqSBwhw3ano8U5CRZPmXmY+IJBC5sm/oHyraH5tlgGtpHduE9lsG/V8uM
h/JPBeapA4FpranVJdQKnpF7GJiF28b5HZlLrATUSeImAyLwuHuOi7zk/jrV5biu
ksQ4EDNfOu30TKHziLIQsG2l+PHB/VAgJ7wpkBJHyZ9djWHbEZAaAwHnhhytYiN8
by2W8taNd/1/9zdvGxVHMo06mCCgSjSa1DOu6D8qI4HtHnLNDt4ZkkVsel/nScby
grIb5NX9BrAn7e2wY9uxCjCItDayDZG2CwVKwblwPLN1MWtUPHnxx96VcSNomExX
HPn5EPNH3xsusb6PMYVxUIU/SSJTCitr5n/V6OFdml0jJgXVmrIWP9BWsyKS1mtV
9lWAovRhN71fJ05kbQElSCqxUT4QR+7iKtCJ9epOZSBTy/HDETNq2r+50PKOL/Ed
2p46tfIP2Gi4MFg8HaaV/GowqvY3UBVxhkkH51nsr9Y6epHoIthXE6k9JRVlJcVg
yO7JCNLgHhhX0W/KmC4b8ex0mHzH/4G9K6vwFiLM2i5rn/Ee3OHCmpBZWoDYsYAC
WmAcKSk1SAVvvS3DCfZFzIgM7tCr780RU4bVXe9JLz2xcwy6x0ONK+8sHum4LXjS
zkCoIStj+ugoYoMpa/ZqC8nCoR+ogGD43U/nShVg6Spftuz2/fNB8XHITRxSR9fW
kxQjMG63+yL241J7ntT8mCJOBTtYK5rlS1T3TwxtnnmcClI1gA8Vf0ER8xyRwfnv
MudG/Uk+PWKuTvQy1Pugxr34jow6hU/MS/8FBn9LeYXaqBPYpIdnmJgYqyVj/9tE
9FUFmhuUBKvB+jMNtIc9UmoWyuC+JlhWErC7qd+s1K5P0Y3xi4Te1SKhWg/h1GZt
RtpYCZWj1050BqWvA7cWTefAq5nqWZIdMeiaY2p0g40bjxlI7zR5MMLH0t6CTRFc
DWAkbf3f+Y47MIuXOq/mceHU2aKmmd/Xcx95PhJGBVis9ZII3v1jtsK6/oE4BCy7
m/MPN1wP21MaZ6/BixaKA6WGrT4971BLteN128/Hi9tybHrQTCZW7LA1FefpV1u7
wE5F/obCdwK0qoPlQhBPb6bs2WVzwLTxAnjf9fmc4uKJ7KDSPnRUNz/rj0/BsdV/
VArNnHvH1dnFPuKCd9t+LflQvVxN8gju10FbUQO6NgduyPi5DORO7GQDWCPhN387
doElJAmWcyYWmxUrVlyfm2MstDLjbmjYzs2wNg4y53sU6rQsJdyq62oM7c8q/i2s
3OTAYu+kr7CBv+15/PMSmFQuffXybPzmbIarJTC1iei3H208jeTuSFHT3oBGcGVt
vn+oTZHstLVgYyvLsrYu9pVedcCQglaMg6g5BiO5kF5t4x3PeQrDxG3Ee8e5zc8Y
zkKp7paFeYYbFTmbcGxu+EpRm5LF6qzsa3IOkqgxz3RsMN3JWxNSmkfgFlw24N4s
nf22IEjt7coCzYc85rcI/3KJZBRejqUrvNSTy+VAEoj4O6sB2TVNt4Qy7pmS1wzf
PCZYNyfs8wHYHLDagZFwURmwDepChc4wPlA8u9IcWk06GIcoYrOrN16EiEmn9F00
i5QZ76Pwjn7UxNu4ygftLYKlFpzvCcDBU5o+j46JusxlxD7lSO+txYW8oOUUaIAo
h8nH90898D/13F5do8ObKl2ejpi8MUP2cJigxjo5sX2RythV2KZXCdk+EQEH0PgI
NJ/sMf9+FVBL8aT5WGwbypyZxrwY/gD7rxgMgRluHiX5RNiFAJOFEMsP0MwMESni
Ewq8HiXA0TWWUQG3znE0r7/2V3S+fXKBavSig+xRecZFq4QBgSUbiWf0/9iImKWZ
mw412uSGsrxsE2/7FiI/Hj395I2jLy5WBo9GEysA4hI2tzGZtxtVpswJqH5/qvuC
mKaYCmkQ9c/vGwLgIOcXYqkX5kk6wpQmyY52hxofH0FVGIiKvkEiYjQcM302/6ol
eGrqL99dvjbrbEgCKnsnSU0Fq0q9L90XdntEo68Y4JCbvySt8MHNTLB+Rcpg7z8g
Wh+On7V7/Rvv0m5xkr3MVvsGR3JobbGnlv+uIUvBOqA8OrrFA/ZVZ5cIzUiDKbFs
gJUPzF8s97STSYwQfesPisg1wYCxJek1Xx5wteBcGD7skCFAFWtZSNnsSbvJZ/zf
RBUYPKkfec9V/TRN1IlEIreH9a/FNYlFwpcvNqixDv+TM93MryovpcFVMXOsUgJF
DcyiOwpw8AORbUQuT1BcXdCpP98PJh/oh8h05Xqa5gZcn4tB7yrj4hEsuJIROpnR
9g3q5sodRNTXWS73EHgb+I0ACiPEqJp56GhNPKejUvkjamOLREMMgmiE8SBSBcbE
y6X92zBEXjHkLTC2XqWw63ZIrPbOoQolA/r7PSMfrRHjcbw2Wo0NClcV+u6UeP/T
+TBOrhhVVfASVm3e8TCPj+ZaIHzRbo+qem7cuDAKHHS/aOw/1D0mqKRdO+MGEIKf
gymSrCX0VWc+HwIcpZCsAVsz78cukXMfMUP92w8GcyVAo1CJJyRhKCP1Hm9fz5Jc
yqDlqrpefdkOzj7JyvSqsVVsZ7hcltgGzc9dNyxrmnL5Vs4FuwxqVW397QxAHkk0
8QfKL+kDKwrjOjXLIL4eCp1ty5hE9L4ZBCErQDJ5LFGaH1ieLMp5gwTCMvekDHtw
HwGa2O37nMfK8bbI+ljpm42oVHkJApaUgnH2FpZ9vOoF7GuUTysz+V7BAjFhDySW
w4V95OrNA3XJ5u0n4grrd+v+X072Tl8XfRiFnXOj6JrQizq8jdnoEaBuPVNurjpp
w0dq/I2d3zUjHuXivv8v7+kJJSrdWQjWk3c9m4rvoLdHx9jjRNyBwAMKHWrLYnRx
pT4M2T7Y6iLkfJKqGOfhybWqiPkNXFl54SHM/sgZ3xa8Bxbo5QKfEURaHmq8mXYh
ANlUtFYe9uTPT/jJycf+htVSL5+Cyxv+Yd24gMZmmrp0FxGb8q00VuFowI88E6vS
edvlWeBO+qepQH6rH1MPieEDdZKEALCxUVL7euk6/aJCd304a38IrY+jeSz9ShCM
pH/mGrVTocULFlwuPy2bMmQZM9S9fDuQs8QQs9YkdbIMT8uduHfAL+O0o5T/pX6S
8NN9XygucccBPbuFchG+IZ9C/Ui/hQCurSVnFcqruGjIgqACVK8m9cip3s+zyILn
G5aQTk58wbROWUVwz5LVg4SMMBsrHg/E3y9K4lYdsycSfHLCN8MzOMa1Vet7R7rz
w9ZioBhY9Xd8Pr5RhOZ7fK+6lR/FjZ5GrQ1F3qIw8Fid06/Jau+ckvZ2C9gw1rSZ
4+8KkB5gwrh4XroaXqzibGyYhHJfO+GYUvCl6ikQcCITPN4UxvWg+j2PUwodH9w/
Ds1ZY7XVFp7rTaUBurN69CmEY1ed/cWldFNpyx06txe5SR69B8VAZAxGPhPXtrd2
eh/o8/NClggXm/tv87w27m/MIuj2AgBGAUWuUnq986aX7zrG5nSlbWYhab70yMQc
eGsS5KOenvKoqMgku1JH59vVhJTsWu7lcBwoOaAloSNcnDW5QBVtbf+lmqWXBqc6
FMp89tX7PJI4I7l7SKSnG4Ch1doNBdGW6fPccIWJSk8FXtC+X31+d2l/Z7LPMVqI
14yqv16p9e9T+xObPKAvJvHizeQpt4J5/tDoWHH4WfsMRfFCIi4R4TTRaXlH76IF
sNj6zppEgNlbcrE8o2TEkPq457Zjves7TfFKsF6CH+QS2q1aptLLDjNleWdZCzWL
3V7j6a+6SdtGywjPHcmf00WkL85my5HJSPdbZr0Zd0m5HZaRjicTR2e5pUalKGKe
hSDIjx+fZjFjBOl+HAT/o1Ax4AuehbiMbiiXzwNi1F1Uz2l5EYZBfrjMZcAxqI5F
pwL00xy2JS0Y4aKwwEbOSIVkYeks5elORcFmMMEeEt7ds59whCLn3NsxdUweSPQm
dpfu8Svq7O8TGiXH5zxOcSZJPBTehiMUMSvr/oxXsAjycDW6dCzDhonoNBiIeok0
NfxLaO8ZIEMNmdTEHaRPGocWrij54EmgzJMaAM5vWWhk/8dbe6zkU14IREhFJXdY
UevPpmgA1eZbeF6eFgaUp1+7STSbzEKkTsJXuWqO/WPCb/GsCSsOND6hu6Shwv87
LnycXSnLOoZNzOFfggEnNpwRkdxwaK8vLrLcnPQqNWJOcT5B0CjeDRUmoqOWNSYh
zBOIfYi4R1NJYNN26tPU3kLgWRPMF1TqeLg92awkVR3wt7gtkeSeuw5Ab0LLLnEd
UXD3M3xQUN7kYpSyQhXWzYhdojGBSh81BRXymkTFDlJbk5RYI84qAZhtKr9W+P3j
s5lqNqSX7SHBW8acPo9MI7afrPN8YO5DsLegvtcXk2wAOptPzX/qgeZkTU3jlHbM
Iu+MFsMFSSoJT9yqQvL+fsI7wlodRm9KUENNXxA0U/ua5V+XNf2kRnrYQn1VON6d
33QGAPvlVfj+nGBlMUcHnGRsF4lPnWqe4QJb//zh3aALOx1OjkQ2D3Rc++QzzW8w
pDlZ/jGD+L9+cCQTdOWk1znRZvZmz1EeYKpcx90EsdOQ8CXCtInoOWu3KPQznSnQ
dzO+kgXs5+rMpDG/rM/R7rK4qCbJ60hgyTjzJ72KKHXgYQ1E+KymF11wB0ANhGS9
s0qKpbuSlOw9oMJWSIEOLofwaOi010Kc4we3l8Q4OfVqdkVhkYN4j/JmInRGxeu+
jiozbbyH8l4B1J1g+nanYWd3i/ipB2J8KDFEnQ2n3PXA77yD/w8in/I0w+B++Ug3
ywkkNXagsyVp4cJv/SkPipIlSpNRs0XUIMeZ95/qpQx91TXqTJggFY1nmK0UOICA
0x6yw84IB0tFPRV5hpyRpr2TfvkVIglfoq3WL98rYz6lO4saLQZUrF5pPMbZkn7J
porjPMhIDaI5ht7BLQaOeFRixmJUgBQXrV85gnUqCbh3K7pb6meBXYoZMjVIXFul
dcT9ATQwzIg4NXjlzJaaNF2h6pkdKx3bt/KgF13Av6XdejLhAQBa0FNB11EJDw8c
jIkF0G326fIWdlr/YhyRRBp7Dt2CK9h7/9SmDcSyKrclIZU+j9ytqHLSyil7JS6w
g0DmCYmKxdeKi24CMYnWI9ec4xrrpr2y7AOGI4yAvgdLufcbslfPXxtD7mSPwxsm
uZ9TXug8N2pVPrevOpHVyGnsO6MV7jQ/XrjyKXN60Jbs2EhHnOhkCGy1ijOZLkoe
xRLfr/Eajxl0H+Dcz7WEwo7VynC2VasMUr6G8FBuTdyy34HQQRJHrEb+uOsxm91y
LD9ilYwIROFbell5Efot+NQQmzciaFAXrN1DBD8zehJTSWuWc4ZmhH1xeXngAYgm
VcxWmoVWtaGY9ayH95jXlZMbr2ARKyBw4j2eIzqUer5z4zVYLlmeroQ983q7nHx+
pKsSuGoHavtepdNLz+rV1Rr3KpWxQRapya4wOPeKwOmaY+U+jj0J+Z4uJ6fl6f4F
bX+bwh8khav7HyPaZ5GCHF0zTzZEVPf/DKiDvcUhFMdvgX3MTqXKdjvFjgXrhmqc
j7WzPHCPH5v1gPfiIsATp0/SmxUdaxx+CMSqgPIyUrmKF/OcemqNrKDpQWtpvi5H
HhhKmLPsts94mZiwgGqIKIYdBy9FWE9T4JG+hjmyAIYoDfNio/qigHP6Wt+3Pu8/
41IGJ92ZRdUfSOR/BpU3pGN6ny9TDBTm2oz+YkKMORayAg3m3t0vY5bNRLHOmyWv
6JrTjJ4OVi2erbigoRU7gM8iFSAi1c1tnnA5Q8waAG2Qlq9NB+OFq3lftb4Y9W4N
MFBVRb9uJbzp2TdqYlS8Bd/1NVU/NK4mkRauT4U6iPHfQX+ArljImA99N4BSMmZb
rfR68px6l40SCOEkFJgrZZhnoANMYB0OOo90dK0HkE6Ron4MsV4vg4XSJKcLJ3iE
+tfF3exqHqkUhNab2oqpCpNfCskmUXh3TE4y5NursTxi0uEo2aPKVDtRNhXMMiS+
BsARBLdxbKKCLrO9VZ0SGmQh6qxYGcBqCC4mRgAYc9zRvZzDUeSN5vOzL+upLmZ6
5rYsLOBSi1CSdfMrHu0BPw5Nr5X0hbzcPhw3CXmOVC16CqWlv2UhdxYaPgMQEhhc
zVBclDYKmgoi40o8TJ6EiOVi/kTk/guTRFUvCDfhDm+haEHqsK7F9PQ4440yEsbW
HlPUH5iMBGlvpgLLegI5l36rEBV7RrEeSkEkrRraqn+hO5j15VMPEguSa3uX0gm4
NY0KDTzE44YqD5BnQWmLcuedqRP2wIW0YgHlmHDI1LeeWcuQmaJVkjtGysjJIfdB
5HVU4AM0ocOdTrn0V3e+Yai3VIJmZeQiGNNH0ClS6vHgQbXKQWW3IrcwjWAPBHsF
SgyKs0zlJaINDAOuDApro95gfzk8HU/bKS0+Ez318IVBY99lDW+OSjIOMQvVrbDk
Sd+JW9WKgmHPKKrMebQBw+zRxTw7wG7YuQfs/0Etp9oMPbMcXUk1kISr3wQa0TSe
t+2SqbHxE6EASqSpUTm2fIFJK3Egzp0BGA2hzPgmMkaAR1v6Wk1hvGgEnwM7YSDl
F4g4XN/0SfX3P9+n3p9PNbHqjbQN2lgEfJNmQAtJF4nhX9Sedfi1TWMgKPbzGz13
z2IRixDYqhmKdm7HPia2YFt5XzIzyrCKRiL79CHU1DsYaMgOouK4FTSDFX3KkcYu
A3ZAmaaBVZUu2VMaqnJ+tKOlsXsf84u2xDBOBbhJbNGZRyyneawraxsfWJSVcxQ5
9fzxcMLlwr41Vt28mVxZVQF53/9u1uRJM6SX0M4L4sZewCITYU06jDIrZcuz7Fz9
aZULVIM0VzuIhqeVrsmCkCz2DKqj0xON/7ryPInXoSdKgF6pZ2SH1LY76btshoUe
R1nRgtnzZDexBSUosZlY5kpAHVQP3g7jARwWHPRWIxckiAaAVRl1l18tUrs0xeX2
1l+Gl9bAogLjWZuBDz4F2HynaubaAiRQ6aq88e05OJCFM3yyByrd7h1iEVdRHOmr
myq90vKZDAYPX47c38g/CrlsydN0L/ONiGBPCjKuEPQejLdF3yF3pIBafLknUP4c
MVkvt2/9oP0HKax6TF2XlXLyzp0YdFdrisK0+SrtwllQVT52rIoL+Jxd16A0RVfX
+sPUDFVG8xu0Spet3pbUXDpkAEJpv6XgekhTIhU66JaQYF9Fa6WWmCDQT9xySz7h
2OqjTN5Ym5NEJXQcSkTMnoLIZUPV7vWOEjaULTKw+VqdJPabMrCy+kXuBjRaFffH
bd+V+8o/+2mOOWwU3IsvIA==
//pragma protect end_data_block
//pragma protect digest_block
zF0UWiJg7/i756UIpQPng2YOdWQ=
//pragma protect end_digest_block
//pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
QcPhabDKh8ancXgksfgFAI8nvgmJeaf2HCJAdNTpx9VeHNcT6gKq+p0f4P+dzQxD
nCL0maZ/ep8KQg7kjJfVoMoDGVDm926DwuoUvC4NPjJieVOaxs9WOcuMxtUHLt6W
evQldRZ9Thm7UUTcCiDfU0GRG4ijUO3mE2MjuXDXOtk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7664)
IKN1AOdCicE+FHlaorqBrNQeDpUxg5kQ42rDorau+ULHlazAamvtz0ixtAoyfxAF
Cv0labke9YKa0iWosVAhZ28wayW1Ez3fomfdKQ37NoCP5mf4WxwABEjBZa1/63Vq
oNYisny3hDw1RgMWZErRgVtc5u3Ut2o0swkUCVpxXvd3AHkk3aAFoe1GMs3w48Sg
yT7WCTm1IIKh2XxNPNpecX+kCF6eGcyOT4Fj+gnimDleSmR4ZDTn5ojbZ6IIBExr
TkuLyrvAIMCdVsSFa0eUyu7qpuzH4R9yA1KRXBp6No2LXjRlnzQ5ODB8W9vXwDf1
8aAwtnRscv593zATM1gRuerNpEMsB4avIcjAgHxU+PYTIknqY/rRTsXcAWqZXSPB
igYKXKcHmoRgSZMCeIU0aFrt4SFK9vgupTWsXo5J3F0fE1goUrXzlP3NhEdPrIjK
NFIOnDHMiRP7BnyUAp1uDZ4eMnbXlvwbSrGcZzG/jRfXGqBlua3ntpO2sJFzy7z7
qtC/NpL0rGaszmkdSXDUm4yDJGmlK947vF4z5dnXpd4100cS+m1t3grwp2jP8OWk
Y+DCB4n8DZXeqThoMZ8G6MlVhCo0wTeqATRB58r8VaeGrm9hM0M/eeXmAuzmLIJt
zMeK/ap2uF8qNOUZaqxZCbqK0Fu2FbrKDBxFQJGjLxf/U1a43YZt8IyK9z11vSJC
/jI3coHPl/qqbtjUQ/fcB1s5bgnuvfsfC88cuW84EewCP7qecM+Yyu4W7/wDcoas
RE8hetWe+zicoB53RXAZsrKSzffvPbKcoBDjKnAjrktGoPFfR2mLwZuNEOI/3I+D
FeWVHW+pOIbxkP5hE02i3TOoK3l2+QyK1Zy4W+2cc+LKYtIAXvA709ECWADlfdT3
PyYUnF3qnoEz7mERIQUaHdZPyJHYRYEk9Besi/ULmNDSmPE646z+N3VCtdBdigCJ
7/n6lNZxP6A+pfzX1zge29R/2P/GNodD17mJv3O24URs1p1nySJyA9GG2o/BeS49
iY49dePhWes3YtC+OH+EGHs3sQKmiBFmbUQFu3suQmdWWrd75IPe+Ssrl3nzWgzx
MKiLjh4TTiSIfdYDFqJtgZZ//4A7smnuPnImPkYIF6fJR6V+QICaDTchngYsZc9s
X8raa3w9xpMpH3I9xVFURe3I6t2gC4NITas60YvDlKq47wtLW38x6bVvh+1dHb4w
WyuUgyTv3PXa4ozNWIS4YfC7zYJVgJkHARbYDvoH1b9aFOgL14ApO6VIkVq+ufh2
bpTpJdlNDIrIic2yD66kgxMWz4E/R676gV/yd3KYC1p/8QcIzEz3vyAHGTguGa1M
vJJnI/ybsJHfhvSCdNndY5+2NoLwaJwmv1MiROjLetpnnNhGtqCvvf8MgLraEg9/
MN2DDA3pM9F7bJJoF3qynkYQWMdBvBQBoAe1Qk8PyCREPSmn1wfUBhF6hcMbKVRO
NYINZcgkEvjrxYbqXaEu0bDA1w/7cB65GrSsvtHw2bnEZW0Mv+r5rx+fhd7k9Ldy
a6l6gWUrH+0VNKAoYLZpSRsEcw3zc36CSlIW4bMuJbepo0nfbTsoZP2OLfk0X7Bi
qCnfe+j/EXFAQsu4JeIAY2FTQhxb1hUg3ZyLry92ts45/mH0lEDrbkUnQmq66YKK
NuYA3/sbjX9NKRtHOE4r2hh29/4MkkikEBxuDgKDMJGXolCNTWyih2MVuJoGBgXN
Gomz65PpqwifwnNrMJXAOm2hgokv2p79VmmxD5+VMJrnMTCgkUWGvQrK+QsMcjVs
I3mRhLRIKO5hSBrYohNUBwqzR19C0jgXoY8aBN5tt7R3OIoQ8FKpnJHHr4lI1isq
/44pbxd8n2DTLYgOUsOd7rCG3bMRx4Un7CFwo9X1AUSoONhMyGl57Qnv2Ab9oowZ
q8Loh0Pm+YbFurb+YjaiPzeYolcZwjEO0pMS1/72Trlmw4NjaWNXmqoAgBpFoH33
VBMnQxcOUZgn1TY5FZCLbLGTe0XYTKJ3EwLWCHGjU9zNYKzD5Wue0m8u3Z1flFpB
EsN429YmbfHRFpB8p651FIAelYKWZ9LpTwqNfQbtaOk0KmBEdzSQuWvjeXkjuZwm
KI0OxTWqJ0RjZDTbKCPtzhClt5+jf4YpQJh8xzNb8oWpb639rnUyGZU1d/N5BLES
SWi7/sv01nTH4o1TqlsRpvshWX+nGHZaZZZ5MhfXEeDlBZ5wi9uKUpOYmnx1r7fW
k9TSniQFGLv0NH02ezn4f3KZuguERdes8YLt/1CsFqkH0VCxvpkceArlq60tLdX0
En6/5JSYFh29cXmGmSuFfQgqqRaF2e9qneDOZWnk3+3q4Dbhqs1SDCI8DlPGjd9E
ET+B1Ia9Ef7XwKKymE7BizJ84OQWin/BlO0VCcP0CLhS8xcUfHNpAU38RRCWObiS
I9fBninqaTv5wfEX96blxDI/MvEx2pspau0+rKoFbQ+TtfK9D4xu/xWE2BF7mCVk
gLDLaKX/JSfutp9mmjDsL9bhmB03hJBkSLgJuRqJ+45bEIXeSi8B9dZYa4Y0HXNc
oBAdYIduMaW2H7A6+AttrA6CfvofUtTIV6YXhTixhCLQtpJQMxVXwdb6Ilm4gcBj
uXhRhIJ1ogUGc/JzQvmOXbUDMeXfT0qneGp0orRPpqeDanVvjbK29m5mUPNheceb
I7M7iLs/fPi9VTo78jcqU2Ve+GiA+duSDHy+QEu99Fy9K8kU61y1AcylVYDQriuG
KZndOwRvsyCr6Jxufu+OtzGRq/a2w5+aoD1ZeCmYDJjGYcFm5m+cge5Kn474qndp
9AfB8xZdmCRxt24Pn45oFYs+dKNwuLWreS27Xf3msr/I1DiWoCVyU6AKLOhpuEJI
esosm0e0AB9hR+/urVaM1khEdkiDiz9opt16uoL63EXJ1hUZUH3KTq/YO0YUoAcw
D/0MVvA78tA7VoJmNGRkHC7E/VzkyLbQ22uzw9SWa2Jo2oNtJi1fa4TVSygUO2Fw
iSw4rmSeojRGE1wkGnoCXT22UGA4hEnSnt+KJjjL3RsqQC2hgx4f4d7BS36isfME
XdvVQAFjfrYw1M0e+VQdwq6wMlGKUDnPt2k4ZkWcZLu5giXrUWlHLm2ztoAdglfU
yjCwClcOwGG2ZJ71eTDzngCB+okKwIt5+rlIEOJz1XcC/HnTWquEIvOIQK2WKr7M
V5F2vzQ+WVWjGUq0RjpXJcup6tdiW7xmQrSu35TGodyCreahe9eXUwWdiyeHx9L9
PmftjPDJY3kUIqNGGAb5xj1r3XmeyuLDFNR/dMxmj7xhw3SLTRBde2+760RMozLK
b8WaL5FYXjGl+y7OrA4z0izlU86Vfn1viti5UNp4EjF03tg6kh+o/100vSvVm/W0
nsBnYjh74qP9Vr5j9l9+30HxUkfFjZgTPFLFXLHrPyLRiKCyrYxpoZshZNhew2u8
852vGITu7XVBWShtsSB4cwzRxZh17/lQNVNJaoroHE7g9QFuxpuU9VLDJObXFZWj
6SV7dn5wso6zSI3b8+1lITAiwukxccX9JrC+FZdTQMAVBI7kjnLxqBjiR2Ng8fbn
/8/9dzj6GBj5o6va881g9Ul45vKuuqZurg9xeK3Y8OjG67yQz3Pp9y6pPqCX4TSf
c9kx7mJxkZjpXTBzgnk6EXaYPseCqJ/w7CYURz/6lbCBtrJik4UVUptpUFlmOHCy
yvN1CK4KmwAf+ON/Weh6+PfPBGk0ay+hIE7n7XlS9jjChCZb9ZcFrHdOcNYbaos9
WFhhKVHmc0EMHOY5nQx3wX7Q40FNZ3wxYfscEXdo/r87h8oMDLDZ1580TfzkD2uz
ziyXNI25OPoOtK93D41dJm3DesOc+Jud2FZ7uqsmLEF5oD3SXPLz41KT9BYeVMbs
fFCW0lujV6Obqquqwz78uNCPN/774MOpM4LJIb8T06a8VGfpqrSPYBA9bRPnpGZf
kouHHcf93TjKL5ar/F8/DkVNy9sx9S0q+bdtDlnoelC5XLFY1dkHTG6sukepa4po
0+yslRVVuzuc98p7FmYO3edL3AQ3hyOhDSGTJiZNgDGoifjB/AYq/rlrlrH7dRmc
3QChofgn0qYstEH/Ok+Jk9Ff4VDi+b35mSCSXAU4LNYFaa6J1yDsC3hiT/rxygsH
Ha3fa+QkUFrh9GG0n8f0W/z5etQdsba8Xdoqo/NQTXHSE1YlgrmgEfb/BBTDzRiu
jaBDgxxIebPMBB20HzyMSwKsPmPctaayWsAvKBxE0mWXbhLzIsreLucP5CBQWHMF
i28GdvN8pum08IwYE7Ed7DtDxfIEcfJnZ8iFLkTDvZvGCq0JaMmz1fiHQI7q65Xc
ag1wqcQGKRGND+CR4Y9zbLPG3/WhlQ94rcsfBerOt1rZHRLEdEJv+ChGqrj4CO0G
C7f0LmvRQBahSD33TIjs8g9M+x1F4rg8wZyP5DxZrbeK/PV05YCJN3wISVTfgG6s
/InZICD6W+5Nyv4kBmWe07YAHt4bC3iipludxwUcgePIPZuHPoUjV+/g9tDj4f4V
YCMPBritauB1oJhtq0VIsablmeovvlbLB92RPJi0L8T2MPHFLjqFDWhpihRNCES+
OTLAJpRxHvmWurCR9+FOU9e1C9NAFAqH+FmO0NNRWG8ks6BTdaWZfKmx7lm/T9gj
2wMs4p7PIrspK62YYLjTJMwoIJqp8/j+Jz8nKJAajbYoGfoW3kZlaFad902M+w3X
V7pPEsQwrwwXFhKo4fzkbKhkwaWWCEpHjPSaSul82WpsJMpSprR9xJxa2CO6eDKh
sLnU5ZCESMRiK3q/onqR64G4xzkSrSJwG1pQc/85ouX5H5/upuubtKmdlJ0KbAvo
Ys0wiMIsNnCFwjGr+V2wGhkKz4J6nyIfXQduTnlopcK62W2eAV78n1WXAkoCaVek
MUICgRM1Z+5XEeP2MoCIxmJbU3HAA9/+8JuV6Ig3zkqwGRY0BFrnhfWBXEHu3m1a
APFxA/IPSTqI1wEOvHOTPamsPXpmuKgaKhk2xIWUBpLKwGf7C4hPeM8Hgp41ZN5/
lMFgaq+RkFBuKSGLKZeKmy+gF/hOJS9N7uX3Fw9PdlyvnmapxEuRL12dNB7tFSUb
nxcqZA4dj47XMfMe+6f3XfAJL7hLbC9I/kZqkrYEBEv0NsqIMIy5HWFDRAeXxjVm
H6UnnMW6adRBMSIJvKmArssncoFodfwSHV8+Nm5L5BraSIsiNfKJWmQ7k6pF+nUk
mAgIhf74bIVhMFCcWoXC7DbVwWJxOrVOXci8lIJdkz5Dvw1uaV0ysf0uW623JNis
NabToFtPEfQVnMuq2fihgtdyxPuWbzLFJ4sytRQExaXtxSex0qA3qNKATKNv9urG
cL+5bkMR+Uw9XSzmX6smXN3JDVxh1SvoAvFf2U6EQgNRoiH6z/CIFejgTAoQatLx
W9vmXYSw6njvC/FSWuLm1luRCSAQbiWGna/wTilOeumNHCnDWgb6KqUzEBDgpYfa
9xgHHZxGrKIhobCHJ/I0IMmNTqHcyFiUOx0YOHVHVQ7AiqjJlOvc8GeOpJzUUITZ
pwcHQIMZdZTIhDWxjzr49cCZOBOF/wWJdzxzO8bQSouHBcxNlxWw0QHxf5DvbZpE
pRyXT7tW+8OgZNkIvujz+lwcYmmwbCC+DJxW7otlaE1Ah7x9z5+D4l8qZU+tzzpE
Dzmkz7KF6UH/LtS/IG7THX9WRipljJju94Ugwnb5b9g54mAXr8oyVvBz/saWivq/
rj6y/QIBNddaeFZR4CWep2QSBW5Naa94CrJGQKXjXUCLldEt0kx6Ws2ERO3WbOpK
x1NZxUfLE0VbXzsva2LWjsBt0me6mQbwmHXtBXuLZJ5GNddi2VnCo1hZhcXNNSRc
KTs9vDbvfw5hZgC/cz54mfayQUZl/IqYNrAG5JLkXZLBvYKLGFms4gfKZCXYduw9
terA+aShUJw9c2F9jPwK7jkuV7PIqnLwNLw7embhjHXXEiX6r4kUQeO642enu/es
YFJN8C5GxtOYmZdO/YPbZoLtYYr8ugn5EbC0Y/zPqm+3kH+TNTcBU5dk2IiwrZoA
miHa9eUmURFuocSJkVGqPKcmjFOwdBGWilEx6aOn/YowqJXbLjAF2qMfc7g0uytL
r9K8mb7RBeGqHjJyLJ8lG4jHKxbm0ako2Vb5t6Ws+KQwlIUlyBr6aJ166Z2+rerw
BWuhSC47dJFAZlJy+8Y/zooz0R6sR4GFnXTGY7T19i/OJ6GNNdjoJb4i+8kGO3ux
SQu+Alzbl9bCjKaullj5NZr0OZce14Be3QeywyslLVwwJIsFAw1ZbawTsiWl7FGk
qRnq/O0fdZ5UDHpf8EO3LDpvS277nONmSNk3zmpOZ2t4IoD4KC2P0YwsrYfjbJEZ
ucnX3yVzSueG0otFsAVCytm3oinRWqO6TvvfXzZDqrjDhtABZmWoIQrOF3lvaEJO
7uwrSj92NJ0JVhwUbBop2qsKqSjP5t9KFe3qIVdASVeoe0/bqnp1Gw53yvugR8Yb
t8Oh4eevbS66QEVDzgD9Y2erGkyIZiWwxOY8l8MpBrwunM63gBg8SMnkhZNsxRvh
zWG+BWZBScJ54r1bhRbG0xND2rC5YgjnKO3duCIYGG87Au63S3SK3d5KlBEVDEiu
nT1Y9bW2VR3sYXdmclkdoPkD/lmeXlFtu9rB7pITXsUjhijP5jSCJ7xkF6liQpDc
ufNH4nwY5gufHVtVHxkhVogSSUi+UWaLK2EemWJVJhQD7EfYF90fHgUZiohesYrD
43CoHOg4urM2g00cuH+f3v0hBM9/VajTXp7N7vL36lzuMatVkow98QoH1zIyQzjt
6HR33E1zit/tb1wr2jHxVydkjm40s4tlidgF+RXFo0Kz3X76pTHxkGek1Ci/QKUJ
7Zii0CnkbBTlL4GTS5vJ7UhxINUsZHnVH09Di1p+UgiLAddKnXz4ZUgPm14vntO9
4E5K+PDGXLiIw8pAOi5cQvj7xBaJHe+2G7wJfo5GL9AKCKU5+nNQzO4fo64SKK+c
X9jmtyewjyxKlEcQ79YnTke5i+LafLM2OszP+l/pPBe8u8qx5XvL1RK1qk3zX8B8
aXF5z/q478n0QIouLIOoOZ9Z4hqtKzqz3iL5fP51ZK6IHXnH1vvHxcek/uNHdkld
1dGvhqbAufJPG60yGyF3Hj6lajdERaUWds8g/8p7M40vZB5zor+3U6hCBxzTqhPc
5j4XtmAPi46ud3JJE41kCjAWzz+bZc5WIHGHPeir/3ex6z+F1P6BjJPfC40Ok6M+
l5HH92Z6dPl7DLB9L/IhKW2HimJo7z3xTCY1Z5695a0u8sd0tCiD2ebChl0KdVAZ
boxTLRdqeNPHpbru+8g95SlY5cACf+6ZyPoGqEvXIUQW73ET73ndD0sy4xo0ayZi
T55FtHKRIjEvkfXaKsCmmnB69XpRozsLto9nld3HqRMeUAUU8CqsV2NEMbpcMzKR
X/wHIDx96qKgdEBP1ut7lfQtnxusjHuqpvW5wcePsQqBSv9iFCBVIxlE1oRbyYCI
5tKUaV/boI0UIvrQB2EGt4z8XWu5p0Nqi1ELeh61o8G5J3vwwbHhL6nlJE1GH1t/
Yio2YPmS+uYplwRP4XpqRLzyQOTgvyhVV4H7Y4UZw6RwLeGBjiCJdreUrKONvFf3
i6yhwxxWaM1fx+WcwzMUnHApd/heAZV79zJEoK/5SoJZydpZuWBwfbWNLTjx7BTs
Tr6IsfUdWhQ/S4Fymiwh6TD7B/iya8magkI+Nc7JP/fCTAkYqfU0KHAfVGmvecZg
/lG0RCmplw2nrJXN7dgsxj19Ef65iobdjOvpXI7lYzcdnJ5H8hbLW2Wzxu9NDOtv
3cFIs8CNiZGNNRZ8riUpCyqs6lFrL3i8B9B/0KKeuLmVt90+vbKN0pL+08hX56a5
qluqBgBTOesJiuwTcTRzOPp0P1vG37vQk8TKuwgakTVsnMV5OJ6oIWS4ZMjTZedS
48Vhb5wIlBy8jCBuHyUM2UdUVztCE/NrbR8bzWi8zEBTVjXnyTOKNE5kLZ0Ie7i0
OHe+peimUHbtWkE/93olxUAUN1U6aQ3ejloMe5e0zEkYcAYZW0BGdTxpDgLRXMqp
26JniNOxZpJZiu2U98Pps933a9Fx++FzZrN3bW2cjf1ng/RDpX0CdQnJEkpbsF7G
w1L+4sZCW6qmmo+c5Z3Ha9qEBGxm0LSfKj6Gb/0RdmPmYF/f0GFKjdS37F7Jj6KZ
jklX/M2lu6Us/jGiVp/h9QotbUTjWRtFECXQEMpQFDpLId4UgzN0aBYyJd54jBgc
76Mw1yJT2gJzCBp25lf9lTapjv0DwZiLaw8C9zXLJN7V6kGax+78ZzVR+d2DQZrb
fI9DYoBh9TmmBNA1eSGRV84EgXfN5tQ2ENdERLuhkRXIFnVUb6IcCq4SIk6etuOg
q0VVts91ae344ieWxxCqABdgaU6X07E+0P0DC2qcGXPa4BLPVr/Yr/ZxCwCyDOvK
2o4XItrxjqUlHnanGMTQGeqOLQjN1nowFvbhRjbKiOfGXBSdc5zHr2X/yHMTXDzy
uwJMY92NlXzHx5GMT1+66aJp2DNLB2JFEDESjCNbyf2t7dfAYScaix+mS1NJeJh9
1eKokUui1cWQJuqew3fHnQWeCNAjKyVSJ7c6YwfYsotKN6Ojpu+PrLrhMMBMJjWd
p5Qsd/h9Nd+qseB8176bQmtfIWXQOJLdqq4ZupmwIIH66bepyN/uMMPQf8k0WIQe
j/9UcQ0UQrJW4IaTUXi9ZL3nS1pBZfa4z0EHh/h3UBtJnwvR6QODSUzEAtJM8DTy
01zog1YGS2agC8yke2su2o5KW9miL02M9HtjPj/p825xmSPkOA2OsNpKFz6/HXf9
Y5nRPFzPmZdHdHciOkprTwZp/3dRZGaJ9oFGx4WqxvMhr4wzHFEykTgojuPCbjAZ
zrCn775wGgPO/V7fKvu7GzmnUh2xlcgaBPVS8W8KSOstnsq7hVDzEjs4w02TgZtg
LzLGzLu8bdSl9br/E3och8B+2wJ04rRrVF9fxQvS9UQFwDMGCqxHJwfzHAw6mXYk
gcZc4dMpz6lUmk0nQidEnc/0LNKz9UeJ/Z606AHNCGIqu5clBHwlfKCn/IKwZLak
ybFHmlzrdIh/eqAMG/mXO9GoBCb9c3Uq4mOC21KVEXgHwjukVujUqvdlr8sfCzOo
7xNSl9ivcRl+XaEyndA+GQ+b9sHCcdjAP5l6SVsvLSkiz39ifd89gI2Dq4cCRoeH
Ad5lvktXKZBRiGqr4YHHkKSelPTMHcXxmz2k3GpxxX/68HblBVgwQwlX7OIjDN5f
JO14moxOCoH/6Uysry0K8JDHSfEPk8Mp6KOOuP3cn5dyIi95nT4MKh64gB84/5BD
uDk1qG6bcHUcWUxg0191QWC3yTdb3Od60KntCd8TfpYO5fi4x9RujEM47eDQ673T
F+SGbKMN/Mqdo0zhhEyXohk5s6tOc1Rf+uUgCwCb04KiJlpR7kKskOgDQHROrevf
iqXrF9lJiB/PyobIbymR87b5fCKFxa/NnmKYt5d0lgGTIhHHaRb6Neu77JV+Isl6
lrb2YfsTyM+Zb+cgeB6Cl/APtlOMx8FAAxznu2YYOyQICbykcwKXVgzSLVF22dyy
BQ5sdsZRsD7ZyZPR6r+NZ0+TBOo7vVpk0XpyMJ+DjHng1Gi9fevbRapBGSOcrRqJ
Djr8oG709Q/rThNeUBW8YNngNJeNLjGQMWnIxs/x6pIAXWvotqgRWT9vK+z4kY58
w1P5kZWxGaAk9CB83NfBrZgfefPkNBxmO5Qf+wKVG6BH0l3ib0MX95l3/sEMbVHL
XMzuyKmvfY/y5NZ/fg7uisANLW0bnc0X3PC4iHag+deqVmjMpOze2aKSldggZaET
/yYhVcnB03J/Tun3R9PCGLalpxxNtKNNj4cK5dqjJN8brUGUm0IBegjy3YT7Qcwd
we0Vm2ivHVBYERBFzdsPGAMOb54723n9bWLjG6gsuzqOZxReSfTfW6TofZhBa3UU
skvSUolkiyAhXupKZl8kbYg9YAh0CYMM0dk3V10+bBbeMx8SzvazbJQooWZnQFSE
fR7twkStoGuxm56ce0dv0xCLR7Y8QeQlvThGjYFDJHPMQj7cVRQWxXzyNHu/r+YM
Y1N4Y1minQvsX6WKpWZTAzD1hKY2aRajvyguMyTJ6bk=
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
3d19eZFc34O3J1NmZYMciwn2NekFluNLguULyIeNrSWihnGff1LUE7Q8GzghkHfl
TtqSn5tHufaYPb/8CJ5R6dkiECe/WS1eaSR3/U8JBrf4wVKN4+Gm1CE7vdM7Symw
o9ekBfss/HXgTLEqsghMzTFPNIU2NEBYN9+7dDwU7iU=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 9216 )
`pragma protect data_block
AimUMKitDNG0UYnCDrINmUiuUym4y4I2qaHdWGUVsm7J8Qt3tFg67LxDe5Y4qVZN
z53d1ay3csQL1IsBE3x+UIABc+vlm3VSNSxv56WlwfJXkx9bs4KEiRWyZ+04BgP7
S9dzO6VRwNO6n3jjx3CzsR6vzwbrvjCiQrAK2N4sgcnlDKL6ePQHrjts+WM+8yLc
h+t0wt0VuVxrSHMHXtyq3bWmZhmoqDmiqlmnsOUAHdLFF/VVXyDR3PbjqzuuzgeT
FCn3VoHjt2xZA+Qr4rQmR6wor2Vd68dUyT9jlQVLBserR7QmEyNEbDYrE16tA0o4
7twIGI7yhyRXibDo7OubjyP9oI8q3xh+PAxM5l6ImxepI6s2Akqx+9TtrL536wMa
DVcZrXTsqWukWNmQx2Ka1rV1rJnlkYOvUwV2GJ3UWGs56Ss/pD6C4wlJg8K16Og0
Z4T99W02/7y4Krj4ouhD3oui4sZXShTmWzp7Y0UsZNTYMzDVGxeFWiTWSu+FvPjS
5y5dbV7iOymU7OoMcoGtyoMlAnzbvFjiP0zKJ4JNiBJp4OR7myKIWwZoC3rtuXWg
H0v8xDOfLO/MSrxeIJb+tU0XvcVHiGv6XKPNljvm0qovpVUom4V0KtOzUrKXl9RF
pIVxqKzTHIYx5k3/uBKesYL3hewa6tqjGJmNiJKMiScoe//O4whsWrqKKfwBXluy
9NY7ZE6GFce3hLLx5fIaWuBEyOwHF/byfEV0OXy4HV96DHS13Cj5gz2qgKJs9nbJ
/BwPcvUAZOZ9kYNqh3mipcoMCscjJ01LDPsI3RX51Rx22jeT2CKExATZXx8C+OEN
ibKt1bNUztQBVn3f+1UTSu2799vMZx/1RNJUgLUIFIMkKgi01ekYlWw8NPazBc+A
ucHfH3LhyV1Fhml68hEu5stO0jKM10vsiHK9rYqiJpIX2MqXsI6rO0WNhE8ah9Jm
TQOPzZM15jqyuLU0ALhwNAlqOmwmunWXVCNV5Pfubq/OuGUCVomBaoRgfyg3s01G
t/ToCsB0eTDEhpNftGT5cECgA2v3POUBOEiQhKg+AwNxstuyh3xzUqJ3FRyOr34m
SpNZGZ0ZiGBvUquJtdVqVIBmK5GuJlGc8G9inwTqrJp6CBp3gWiqJUzxRshXpCMx
v1O6tnOUN5ytE3LFxSnjnWVz2Skd9SckunxXxAiW1YMx2HzBVJed3gjIOY8nbI2K
76xT5RtBWSCb6E3Ueg2Xm+yWmut/FgBsaSis/NWK1ZdokkS3XnCcYTz9zC/TSxSM
FruioN+qlqh9i2rCtqE3jzvoUKZ97aXGi8UvAl1f8j5vbAt/FJ1rHBXOpR/C6GLu
RauAHUWV4WpM2b6FpJHlLwMPv5ectz2Lk6YodVU8z63K8oLi5i2AqOnFl+fm+jdn
6CeFAk5eqofBfND0+ej2rz6tjUEBMxT3zkEmsT40XWZteW03XXaBUhoPiK3KK15z
Mr50wRat3RQZwoTr0aFK+GrwBNaxjw01pwXjXqBGFcxMmWlVoakInrV7H2i0EuIO
tDZlycGqnZJXpSKiGYZflP80/e/+C92ux1cKz7OOT2fH1BDtzG9/eMVRnJUXQ58/
KW7/fqJ/qIX5xbg6c9RA/THP8Xhl5uLpLlwi5t/OIEor1jHIm4uKVvBu3EjDK1dw
t3H+dZ2Ehl5oMcxgPgmwBpLeeBOgm+zpxL3ZhRPYnAy65U6UR6Sbyax+ZPh15w4t
UnF77o5L4fgFTG7iJT0076eOkV4F4/IqYFK2LKePFMQ9Gd1Ly7TZKnotbnO7t1+0
WGiJ0W7pNUyr6r1xcIMvpm/y+9TyF1duZ2LWVsIn/F0xraMl7W1rut6u5QNgYb2b
oKiuvl2KlA9D5TpxXeqd6mzjzBXQAU8WnxQc/i+HvXF9gskaSuib7W+ndeiC0B7R
nYPHvDyctwgt/NfTwLn7OT819f1LISUZNFNA2HEZclmq3POZPoOqmrj/eickYkGr
1ZkDnFYBB5fxHdepwdx8gLLw3z/2wcPAieuw/pi7rIiNVKAtJTnn85d86FDjSSK6
ZblUJ441kGstKOc5sPSixPJHa6bHvfbXNJXmTCyKH4MpVSJbLtJUHcaMGCwj3XtM
rOKnCds6PZLz0TF2gGsQhFVt2WKp/5T8Oe8NypNLgwrAdEV6W0mWmWg5tqTV+/b3
WwYN13+Iv3sp40bYtiEc+7iSuTSTl3qENf5KBTc2F1YFmenQwjWiqeBGPcEd7DeE
7lpGnWgeet1ffr08n1oS/MA6OeOVFABLPArW/ROjo60wH5XZY9GKGfKnnYrcVn0o
Hy4gptIm3JHZbwyI2ih26BCLsmHkwSrtvg8eTYgdZA9YhTSn6bB+YyenomSrJqmk
L5dQeUQ7jxJYu8n6E9gUCC6PzUAzFw7m/dEWSUF5ZFIWtedbgjJ+SSNu+sox8nRi
5JxbN/GDnnLdG2+/6p/6eTjTRXBsfgbFO5ikj/HydHbNOHzCCetCoBCguhU0Sod3
UCBQBwoGIJPyvNz8XiGddmkezZEExRuAgLbu3qFW9LT09J7YK1p3dphE5c7lcIQ2
zNiN8IyX3Xyui62WcbLwSjUeier8QupSy+/27zT5b+n+ocjyhDSdVLBNn0Xulno8
arJmgitB6IT2OzV6V/ufte481tkXUTcL35AuSVmok0SNEjEMzHJZO4DdJuq+fbpH
5pszTGODJ+tHSD46Wm7q4XYm/4+na1a9rIwvp0kjjyRm116vQOCOCh5rTcERq1MJ
JFxfrd0wY6QNdAOR9l6vOgrtglTnSYFpROb1JhN0fKpFScIKF6+HihgrtICHt9DE
WXKJg2L0zD4hPeJX7VUQe7lhtzN88wYFQA7jPYN6PBUcRCZaXqBvAyFWhwU/XEDz
FvoCBjx5NBe0nSZyZ1bJDaVBhvMLHxhwCTvM7EfFb4KWTipiS+PzRgnit9DnH+Q1
Lo6H6RtFvnZM2g9/ZhfRaGVcNt7yd029CUJjWkGOvtnJ+NPcm30sYUJUb2tGjJOD
juBO+oCnYm8XzMMv3PfTVJB1+yIjKD8a+t4vWpozJtPWlkEQ3ritbR37B2ipImqx
blVqhFxdelpVDw6QGZSVDbZw163mXQ7H6EPcQ6m1fFIR5DzN20UPvm3KtNlOkao0
j/TxIyJCCe9a9YljI1n5jS2spl3m7CMcep2eZ3BDs4a6E0TUsObYcyGDluqghSmk
uqHousHAPNOsSoTUx+JRUhyyRIy+lREx3HJzyBwFKere5Xhbiq39lb1tSQvb6vSu
Nhyf6fltIY+5ToipbrXq9B9xSHBx369OM6CqGrBo27cEXnYMRneLasPznJ6ky2jm
fvRvKKE3oYrtV5T9YPxu736MGWLheQKwdBxtwkVl0wQGcyypkaPqxeVmu2RajB49
oQTSxQ82rY+5EBMRoy0hcTEI395u3+k6ZpnIkVL4p2rhz7AyWt1hkGvY/bzt+coZ
KoPmbUY0Ufi3TqnsTHIn+wwn7i9fJXKQ6gxzjfzyGsPBiwtVsfB7+fWMuuaKY1Pd
OZnCpjOvCuM/JNaFGfHg2sK3D7VBWUI9s6O64VijaRyNjleAfooR1beAoyntAUVC
6GRDoeDKHJMANdmLI9snFly9EM18dODn/QwqC/5c0r4i48G/r8Ur3wsk8knL8cDl
TBMAfQQpbRi34KVsJJXLkDfS3lHQVgHWX4kiwZ1+nEZ+RX5feZ+3fGn5VeiqV4Ty
LDbl+mdPTU1aalLSUr/3Ak5O0vNy/Yjn6pdL41thhjLa7Kpc/9CDVDakExk9cbdj
vIBXoVxgct2Q+I+U7VdRk2y1x24QmXC91w/jL2oBBYZ9djo16BnN/VGQGgf6kUgK
Vm3HHOJaLH2NmNNWzo1ipdxoGXk7QQiaTryDL9qtc2Djp4q12QBjAxW7J0G4b0qP
We/8Q9muPV0bM0T1ryvVPISQXlhPqnHyeJ/fOZAxIS/kmTv3b61EBrPiFyS+53QF
NCVI37NPlZikufHUPw3qqM6adYvELmbua5EqJQ6nOrP436aDadKUCeXN+V23lcip
XzxTKiQrylJXNcoM0oxK1nVnlKC+lkK6dwkhy17C3oVhh/ItkepRxIQ3AFdDzJfY
OEP7dR0+NbknI3ZyzKopPB9UoHpaBFLhOUbpkBzbvNW7OTZPtCFtgq68HbJl9C1V
o/drsYwJdMk0pWYzjtermZFcXZBubb0MNyBIqazf5BKpZs3YRbNEpoAEhm/1H8EK
mV9ZiGgYlaER45M15YcubXupVFwQVDS58TFI+Z//7lgANFUi91aWHR1HKPG7ckko
JVw4sqH3IV9BJyFgU7Rczg7rWP9ZGurWQTYmen5N/mVc8c2A2fu/bu6e0T5AQ+bj
ru49mkHAvOAd4VFDsQlr4P+0JV/p+JSMvoi6Qly7/hyaQJ18OOZSkILTXub3jv7n
HfvQz7uQGoZmJXYOnsiJCPS9hpXkba7Y7JDBrdIzh1ABk8nouiRFpveSMiCV9K1P
CcNEm+5gSrVzl9r6p/0ArxfKvoPxZ6WjJBotDzCz7UZ+Im9Pq2rR9URukajq3JC9
MbO/6BisignyMSZb08Ac7Ebx4CwTxFvnlhuXIbB+LNHrkzll3csYhnxKs6XQ89eQ
ZWIar5//BQPgAPPpVvgo6a26wJs8MA/+GKJSgdq5qpG9gW6UFOOsuAm26fBlujuA
+w+cNUXI4y6ZjwIxbzya90qzTz2fZPHq4Li1FzdUXcLXkszFL9kQUziw2pFJhWgC
6D5T+4WB0SvoHVwEGZwPyKEPAXnkKxjqMEOJhnh0gAc0CQ9F1h41Rj0bTg07Xiuc
unNVhH51398C5NbtfrWtIus10Jy/nSNWo7O1m3ReLGqhw984YETlJnmOS2e0vtoL
qBzhJfkzUyUh7vTnk3em+W0eK2nYNG0Wj0L70GdO1F1YR3y1nrIJ+NlCObWpjnx0
UUvE1ihm71MuzXPT/fcOMGxvQsnpGLsu45zWvykbmTxyHknJFXFL4qAu6ht70A3/
+zdz9KRObBz8KWk5iwiwuJenUz6kaCphGTALXDmLwOWN36FCwA4Ld0cDdXyKMBxP
GOUxuNc0nargllXU8o9BCDeNvNHoIs2COvfPB0IrFMcYIHFQdwTKZM1ejtP9wVqz
Vdc2xcLVGuPOH7OiS8l73qjQ0/YxhZdd3fNVcK6URu7YMKNbiUXp6a+IllwVGidD
AcyaQj5Qeub5S9cQ5ZDW2CTMsWvP1Aami4Z37tBczTA+luf6p3YfvvZ2BpEOSabQ
sLK6c3rh6XFtfee93uCTJqROaddbbS2OZ+NkReG/aGYhA6+VvzNcdJVnSjw9Be1x
vcQZhWHlMrzP8pYYCSj9jEoAXjZmZ7CsUx81mEnjg6kv6Gef0oFOT4mDlUoRIxXB
d75k0kr/zFQixI0+DULdw4jM05E/inaj11K1bPK9auSoxVSxVRtHd3xDEqz8oE54
pBMaUCtEIjSCUaUFL8FBE5Q1jAUYEvLkpiHHHad7WFzmEPBDeBGN50TmUSAhE47+
O1k5qh35XfCM3zzxS/RgqJujfcJKjnB0ND1mcIGeqiXLQ3+2H68DxhSsSLIUM+N5
d1/BfJ0NhMDI4VUmuWQvgEbAiAxpM7rkx7wzQiKuOPpAkNTkJmA0p5jbMvI51Gjk
k0PBsxRD8ibgdPQ2f5gJAalpZybPu+anFMkSU7azMfFP4lmIpAHXhRCcntPR9nBE
QSTL6kLGMOjItFocE0INMiZKNQk1zVKVDkOYLvtXad60KE8BVXwQ1T29bcKkLIz/
T2WfkyGTmrblwbggKmXtrUsBgGN6c2ODq8WE12CGJu7e0t4kNqjdzJ2wN34tN07c
YQBUUnXIr812SPNudEDySGucDJ1isHFppe18VpCbQS0e5zY66frAFueRPK/Oox+/
CCPCGw6wPKnr0qQ77LKQlJaRJ4MCfY4hQUSTYgijsegHKgDmd8liydO3cpiXrtnP
M0y5gvp9879JVV/In7qFgbaAb5ZMRYcj/mMwCfwbBCbJVZmQD6IVmQMeVdw0A80v
IGhrAivkQBQas6JuZ8MsYRAwsF8M0V8KfH2v+l7xokHw9ABqLCpIvh33CqvJdkMP
Mq1Vwoa63fJmzUUWbhGN8JXqktCgWeTLrgMG1onfzp5yA2yr7Y2Gt9NVGbcLIS/j
eblROLpggWY7AvIshBNY0Br3YLgPYpDNGECtBCxYPUIrHN1v+25hjS1OCCo0H3St
rZxcpTok859JB0X4g0Odvsh7Pvy+YPSEBd1lijImg9Y529XhzxgxGhSnvB5RTBfq
mpJC8O6w9DTMwmKRBcRHqSUnGiHA07uQSfszZpjRAKLwcUk7gf+tP/+4d7ahFJhQ
XC9W7cx2LiZcP1xGQPN1GH6z4NNd0ZzLW1RT6vavKlHAINMaSCvrqCd1mNpFcz9w
3C+wThgOxVrIO6GUujE71m4OjUyGaXq6NnK8eTeqMsmuYGpmY6gBYquPL80XzPdJ
wUFf6C6Ik8zlcuofF+fII0QZ8UF+qEpXF+3Y+F0/TsuLrxNK0/E45OnY8R9xRNSD
vglwIrEHsJJjxQcmE+mcnWfg6FD+YkiCXNhhsQewtPdRtrznmanaMfN08h15M1/H
pBRrp6tvy361MzpT9hCAqVIdWPfgBqFUlkozKAMAEuZ6JDX9upA8O1GOtwnfx4S2
eYjXarkJKpwHHSYyAlIH3AH4ingWO/71wRDoDn2Xn4PL8ejvsBq9BdVOO7Z3vEAY
/1GY+WhCwot8rKesavzUumEM6fIzO8jRGRtEC4BQrQoZHeLc0wMhYloMsPdCuuph
cXTZQUxjwb4unuSY8R2IpWa0swhlVsnSuFM12onDd2ci55mGeblbJBZGeQIJeIjk
ohESWRzWZt/7kZedJbGnCxNeGegN4RI3XRsNy32gDwrD2Mffbc/ePxLpRhSLP07c
6a2uo//xtY9pcfjTgOwQ7X2OYtMSt4U8xUrCFcX1iodhCqPQVqVRxbK5CyzAeRFF
FH4PUKhknckFksERA//c8aVC0sRc2OU2sMw2EOZdS9ai4UOkmEQ+xcPuqoSQ/+D2
TkytmwVk8qX3bvQygPVFRhAqFQZLPeqn7PyF49CGBd4rXQDLAWXLjym+qAoQWQAX
zqHFIIREdKGSQDeQEsdBShtiKjinqYVlYGc88T5lZgqtIowcAgC6qrlICLl3J+cz
ayTnavXqE176aPzJPDTsAV7SWWvv55DUnYZQOc73D+Bx9D6uUkMbS7VB5+vw19rT
+0kxV+b6X1E7E2duxXs88rHbP1Gt7Gy8Xg9UeAoymN0FDf/1AEvtJ6GVK/162jMq
EbwRaVErSBgBHw5FQGqL8e+oABqPZ+hxSOWLJl8mfWlBmknQ9VmPk/Hn/ISyNhkx
4Ken4QjXjVMdVraXz3nS8JMWX/+7KGfl35luTzVrsyLxkwHleLyUP/DuRjQ20oMT
DNwl3LSTFJYsXHhdPg6PB7IdzAzWNIBzyt0kVwt2f9yAGAVHxLyW3cXd56KiPTIe
5sl98Xtq7TowhDaWqe9C9BdMGcOgxDt0SIhwtxp2lO0WzRWiNBR87TrB0ZcguSlQ
0vVU/2RtSpHRwP2/L5dq5kEN+N5VMbLmnsvt23S1Fo74kxrNXDukbK//SIitWYcW
bKfuaFR3J/fWn9nXMsm/nMFKK6AXdqP21iImZFASQtIErwYQbzxQSZCqKnvHI+PB
kFMAPqWtyKzdBLxJMyPyg68TXrnDBOXZa83G97CvZXRH3hLcFxc4dubpq/fnsRaU
UMp3DjvcH6jyoaIYms3ynU4FQWjpyKbhBVp7CkPti3SsPRpcywDpV1fQGl/lHy1H
TA3m2T3cArO6LUEtiKOp8SKHJkXBvKUF1nbA5qkEmlsBTFo7ydeRhih8WZT3ky0s
1XRGkg8slHIzPji7TXuX/jG6qvLbOe5Z5O4Gs/3svt/mpmG+XRNBrUrtYdreD4ZW
2aosSovKga80aRta3yQcpI+Hdy9JSkhlmV58b7re9Ib3XlnmWN78p8VZ6iXTZ18v
bqogLaI/dgG1iD13g+0eQRjSEBbWpzZWrQBUzZzi9r+ln1K0Je2fJC0AepV2vOYw
X7VSjOuFPCylntlNqG6VXQAD9o/47Li2VrOwDG/H6XLnEaxefTbgY1GUeYlbvKIY
w7HaI0KY5QornV1rZNte+xdjNaFFG7lsuIKx2MxA02GSEXmTFTXk1WHb5JKKqpld
4FiZ+goS48tbJz3L7X+jQlbIryrsCOLSBemneDELfR+XhG6LbgR+zFWTAoVgbVQ4
MIZQFTtNJ9pNsSd8n2oFQ4Dmkfi0UZrCiqhNRQ74ezuJFSJwmeG6yQqfqQ+0beIq
V6eFnh/cTgx+WYl/nZ0PCWXwO97mhL3pj/5JXa8O72MigFftzUVJIZMxWh7wLXgH
KmezD8YRstWEir0XrOKU/Kl7c/HqgGtyKLLPxEEeaAWKONdWeA4gpFUs5ya3ohFt
Viovf4nmDCcm5Rt8Y/oZqTG3yoGtZgoWQnwAFeKGQJe/TxRLTBoj46hNS1CpLPA4
hhg/r1HmCtawi83yUdSNJcFBHhBnNQOqrHYjfBCHN+/4bs2WU2drkkQK06Whxgwa
g3piuuAsNvQh63QK7UBD5hvjvyffmipt7/C12o18xKS8EI45YV6igixt9Jigxl3Z
rO52Jj/zw8/TiRhWaQrZ7Vvh/GAlzdueBv+Vv9IlDS2K0OWOMsNLuqIlfDDkXn7T
HzFmxX/y6FdGSJzRk7kGlexLvRo1VaOe0Z6M3j2M13hZpKUsqbFYtGcbXYmizEu+
JEJIA7kk4s5P/7SdI1CCUK0jptVlJnc+BXXffS9UBPNkfA5Yvpf5Or1/Pq4i2877
rAHsSfT6Wz4STtxM1I++6PN6RCikZujr2EhN7JtIchPcBET5vZaIonvvGZ8ZulHW
acI76X548Lx/nR9oo0vVzUdTyLxZtt6ttG265fODQRao8eousFukHNu1SrzmN+4N
2KYEqimC2THQInCA4obAxQsAiMw8x+xdg7fnWoMxFa0XLGpjkhQ46DYWhE7fMIGR
HpSoErLYPyuhxDl4GMe5NdHbPOnuQjvUeeAUpjCzCnxL5FRL4IzOb6FABfIMH++n
AYi+WaOCu6AZwoo5cur+zAXokJlskwdKzzOm/AGF1ttILwTqP7iKuzQF7oRG6Dd5
AjswryIJSpGcaT9fZhFSLLMOsNmHWGxJc8iJwyg9DlN9vojfItbQADwchs2AE2JH
QzxABk5Uy10DaK4V0PQVQnOFvP4zJ9dbORBU6jPvuTkN/X6PJtETmFQRUObcnDco
O8ywcWZUBAMEnWhIjwE5L+LwzF77D1v9I1T+sIEDW+D0+L2hGHHny2gT0ONNc38B
5qioYQ+A+NuEtZMGD11SSbWMHW0iOZWNY8+sYf13X301rXgLDoYB4uaOTbZw0AEb
jJAgwc52R4Wdk9sz38HzH4NsN6XobpjwObnPwaIpBtJXoS/8motBGVk31sjY9tK6
ZLd2swPrH24Ll6MvukeBvBGkhlyM6W1gg9SO1MKsqoyWf1vQ1CpPxiHlPfMbRStm
HlwrpVWdCHvrKoc54vpXJgAUbZQRhyuC0EhB/dk/hHBbshlI/LmWMe8gMr1jbUJH
N/3DfyndbloHpZW3y648GIuUTi6Fhxkyq5TFDDcBWiL7qbtsm5G+u/dGQRXENfS0
2CaRK/ioY366RKwjfTIPfxWwDmnDMdSurUjiryh5uu68Gszk9Iov3sPe1GLX8xYq
TzbpKqyf4zLU9Wo4FDWzdvzSaFslPfBVffCvHw+YyxKBuEfMDRlGZ3g150qeUi4E
X+NvayE+ceM3jkLW65+ynOVRiMN/WM7oUMV0mvhL6AQC77o5Cp+F8IwW4qKSK61S
RDU6VES1Rr7q3fnHlLe90JdDR1rJaxtKCkDSbcKs5Tku0kk4f/DytN9AHoiqz5Rq
xAC6wxcaXJLCqfCUNWhqhqVrTeVcYwuPyEryQXBaaTnM5beKkuW3Ji4oiJ/uFAKI
s5gKnQQzG6lT3HFIN1SEAp6TKhIyAGndT/HEBON8s5YFy7WViVPaF1Rc1lVNHage
TP4E5E4yk0jtEYWDJxhOjjX1Uqy6xPnO/fjwC8MDoPomg1Yxs2U98aqaRchLgHzx
9JmDIlAWAkM3AEyqEffjNSAnjjjnPogNk9sWwWWrt3B6a8fImCFOHxxHMrkYzQBb
oEX/fo4/Zhb/XWAorUuslsX+/7u8q8So2Qxux7NLvX+wtaUiyAtsbFnaeuTMhL3D
DxIKtD8XH66DvhRz2cHp0b315eQybS/kZwc6QGWk42IqiE8X2M+1QqpG4R/IOwML
g02c2TRqIVmVon2I639phyM41ve2IyztzzIncb3bObcRFD5ib4lUyJB5cIvF1CtO
3rF7qxZWdivzrneerCvIBDmiInJI3D/ApIPhY6zNvgGdgdjYry+SRN+ONTXjuCXS
CDkgswJAFM+ne6+R34GeaL0PQoGch+0w+rthTez1Enfl/BhvN8xvJt7jdW+o0mX5
84zEGCMWzm/tXiL0IoorntRXXY0RE3DjbgWnEDiHNM1XZzdu/YL9BoKglhuI0iS8
Pp+jsbQvoTKts7Y2fpxTWsBkBske4X7i94KSWB8IeuyQZJNSUfZvhRwm2TsNtKgY
6QZMUm1EOkd6rHs2Rb5by1GtcrtDs9uuQPoasHtg/29UyswEdBrDUgja1YyUbEA6
fP0N/46Pf03yH4lt1HeB6Eo4nWYzbu+7n/f0T5FL51CQy2MXE79ZirXRCe+w7w6b
M+cJHH2Dk4A7e36Ft2hiGRBNviyP90mbcBt8RKHB8jYjCIn5ueU9RmCVGUxL/VmI
WqDjoJekYp2g1Bh8tKH6Dl6+NkPmYoUdxyfw3e8ufxanyhCvSZEfJaB4sCJXfb/3
MxbVvWXUzLIIrVS747+vrLpcxhvNHcIzGkz4mWTmvWKtQYuKKGvx0KZQyq4sSbVU
NYYQUsfa7dhahQofBKMCeUhtPixYV8PMDXxCUwhoQstPhQZsF2WVpUz+dhZIRKwy
9L5fkTS/Nh2vVmBS8+XXPvriStrTUnTrWpRFdLGN0Ff35KYJyHRBqCw7YGBkpZy4
bW+y0s6JQtCPucidtxJYsVXMM1whu0j6RZ6wolCVbfgq+HdLaBRVtPcQsXaa2TMa
y5AaPLsaaQSSqyJ8N2SJc8TomdWGoOcpEKgw5QGgyM34GaC21/Za4xetuWvEliAS
Jwb+U1sIboHRahIYcEB0sm18hV6mH+hdsNAdHE2C3oJHqmyl3LcQd+jXrvFsAr7d
o2QGUxlMQIgoaTQo1jpvjJWgzxqTvSJCYFsVhicQ+b8IMm2K3mELUxE6uWVVToow
egaNPpyFgS9NqzQ+MSFHfBT5d/T/m9VRd41Pgkmcj+HugWPtFHGSbdBkRMcHgokt
WZQ4XvNnxrpXkE7ICtcxdv2xpe1OOUU64JTjhU2MPDMkrt+Jjsx7FT4wRePpvMu9
esHYegXmbkaGbbU79laPxeUIbiMCgaEAmK1OgfqkaHqGc0XHslspu3KfLwoFhY30
XJHPPYAc4ktektM7a1BreSIHUPYL3rr3+qm0qARHOJ43W6pOiYzjSsrNDxI9K1hl
mJ+1cczke3qY5U4QLRDXKTC6qOhqVULq06aak3r1d5btx3jE7RlIaGTw7KJwrrNP
1LP+vWky+uJ6fn1lBX9xnwvvHIf/N3KOpJ47XUp30RfDkZkfygFDKjoffsfZSMFq
TCYrQoGIoRh3TOvvWgJleqR8s7I5QO1OSQSRQwRcWc7CJRNKQ2lUTGep4LEfBUUT
5FNH1JzXexUln9Jrzs3/gU/um6jzi+rZbXZLb2S7spsO+ajthMZ4mSRdmSHI2bcg
zfVceR1697dHT2TtsHIrTdhI0dnxlArRCdQu/G7yQD4ft+vKS7iWWuHAJoyi7ctH
NctwF2sRSrWbct+hxcYml09Cp+zobozvhAQ5R2q4y1LMj1WCQSxOUHAmwlOFwm+Y
BEapQBiRwmS7Vou1F6HGbqO+O79pY/45VEQ2l8gaEhtWl23BzLGZoILYoRdtjVZY
lAEE5IdCa4OPKUK4iQx+aOfYjcRJ2hV0No2rcnkX+NEzL/TMqfmzZDXZL8cupBxi
tPicHD4iKgP92LzbFlLgAMh9mFCdMr6pZBZ0V+st5PvMn7Ni31+44eD7Sd1u9C1I
0NdueRtKwa8X0iEVx6hOBTGybv7td9bZ5gWlmfsgfIBYkqBHIbcTe7QwI7asLb1V
KfZoyZ8Yf+f0XMFGBj7tnF3QPARY1WTpoNilrspl85Vdd2y2eYUFazDUrW5aaJxp

`pragma protect end_protected

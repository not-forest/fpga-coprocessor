// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
WhFcAWLW1GO3y5VOWlfJPHIRWXHFbPI9AY2Elk5BIbMFeaMo9FtX5ykULzhixGyMRwsTJGK7JnY7
gFa2bHzryiYGz5jiGbAK4VaLEM5/GLhFnHJF7z3Uc5hWD/tnlK/Q7tss6oAI1xjqiWxApl86Ys3l
WYpNxfOC1Z8+nz8LBlvbMgF0dBDzNG2PMbgu/3AGQJRolGd6cWx2YFfGxesKbTk3XS9wYWI/xWuC
Gkpoi3RM8I/nInGCbphSV/PldYukr7jnv18cuoeKVtXST3eSwGUzgvQFWiscFveYl5p402x7SMld
vQ8wQpI66aIElIR6tRU2IMxFJePfnmdCYl3O1g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8736)
VnJiHih7DMy/srVBUpQPKeVWvTr0vbjP60VscuRfi0s0b/4EoGTp9QdIYuDBu+zw4DgmEalulMpU
ZfvjtJmq66oA60yd65eO5U0p7O0qqLjz8AkkW1NWY5LEQiMcuWYNyL8FTSnuEUUt4i0dpQYGekkJ
ALEgQs3jPl0zlp58yKcxVVLKsVeKXBaS1d600XOBbyCEJ1TdIMQBr4vQRXbtXZzgk152zUaK3cWI
Y5hJdSCO4GZrtYH5RB0zbmr7/dR3G/yoZJR9yLzE3mtkNTB1GpPOVoLUCMsW4KzDrVvKvBNxSOJ9
Wjv44OZEZJR4fMT4qlcJvJvsu4XUgwOFy7tC6s72IDombU/buM5o8U+dddcHtb1d+nktQwQ9hPqx
CosgqVq6uSobiyAq7FNMyYL+DsrusK/Jb8L/xsGW3PGtxqp8mqhgmJtHjlRmFoOs4ga3AIV4KnzB
8iJoPYhPB/LI/tBMV3hNohkf/vx9PpRsXmELHzyRJx4FLqDNr8Nv+b100V7F3TQtQCPPxDbJAv+5
DTqKAFagpJGLrnJzt5v44WPuyYN7kWHulxMPJ0GhD0ZAe3BYqGk4BCgpI0JktGM7cbuV2fLIATOz
4akvQDuW9gVangaqkrZKKA+o5hT8mQ340VJ8TA2CGWnubFQ5u1282SNCzvrK1XxR1lrJU7d6zgkf
2voPTyOZnq0C58H7R1bTN0pRA2+CUvC9+HT/dLMtTlhUnxHHDrgfBpXk3TVLnABUHf3Y+smdL0p7
oHAjaHivtY0zJfOohzBtemtRJZ9sxGghvM29VaNcesP/+v7OzYCvBzmjcjdrLTzn9ha8nmQaihX5
Gqj/lba+po/yZD5RKD834jWm6/YIk8vFUnBVD1ko4MiS19rGhrADbWiSVafGt96fCUNPLhAFM2Ho
NQQWABugn2osZZcV8sXBB1rGw0Vlv+nbt8BxQpMuOp5D9JmUgQDaRDzQLrCzOpHN+Ith2bbElH+k
18gOk5IA7RymBmtggfubj8GMtmudQw+fXWmRx5yGPWse9eiri9wiOE5aTbhH41GJpq1Sdtt3XjRG
EHYwJ6j6Tf1LoytMdteH5+09lTnxJiqX8daQG+tPcr6UNyEplRPrhsiSCih5S3Sho5MWPArb6mtB
QrQ8pHUanoc20cxsTsSWOte6QqAXTWVcSmTSg2G6VqbxANtPWWzmB8CPbZEue9969jAQ+iwM7HOW
7uAMiJBmhvzr/3JfeIJyfdgHLoPpDNbUeIjmAsmqHD4vjNCfMsqsxLkE49uYdYE3RyiU37KA3vNh
FesfFNvbM/ltek9tMNuOimwBRtRdjlx0T+aY5uFQ2oPa01gane/qOI2u2ZL3sYfFZRc1qPkUjzTl
16m+HzuQ9luixEYNm2ATUrGODYrP+SefXj7SvDIvN5yL2Vo4jbXU20xfWtnSdkTYyiB4wisgiOn2
Y6Js13E7A5f/BGlK7kMIEjXXM//cW6K9BPUygQUrusPr1i3g+aWfWFQPT+B4hdyN+ZZlpcw1DrLp
/YqVatvbaSk9ABM/KUy0u74At3WiiI0RGs9peTqnYu3n6m/XmU2jVegGHAGfwMfcQj7dUzyErTk/
Hmd+QMnDJWLiZU/qo4J0Up9j2eRBfMQ9c6a+SKRh05mFXkzjVczfVq/jgPJulfAjUaVNuO0zNicU
ZHZH8edhwspd3MdXixQ33NJlWSwBWV8+aLK631kXqmEmFe6gPVoNn13GmBbN+3Tc5HH9/AMZtYuN
TDXrc9mMjFnGrRQSHs6DV3LlexR3qd8PxWxIwRTm1U9ErE94OYnmtCy5C38b4nRxKt6ikBRpZlRe
sDjXg7lrtqcSZll4a9w7fNJXlQWVu8B3sxwkBAU7e3frbcwZGByNXtO7al4mTojA+Z65jq+3tO6R
rG49bVEMfRaIPelqxXj8+6ebR7IdUiVcCiFiN97E+P/BZMUgukCcKN2bT/0ijKAmTW7n+9COa6DH
v4yhKQSOGSPKb7Ar83SVdbievv3RrCET0J4/qf3N0MrT8WSALGDBoOnDc1ELis3LAdEH6JzYf11a
3FxL51O5uFvelCcXsAKd8SHaQhE8giemnq45S2rxdRJkGwi1/XjdirzTorf+2+A9mpbIiWjDTK3R
Hx4Ky3KUvI0oGegj0YgKsMskZyH5Xf69nI58ELSV6h7xblHId4NO9oBuiwRNgwwl2AyqwgGbOl9R
o3E9N7NNqoVQgM+2VIYBPef9MSnfqz1memnkngpLI7sivIxf6+yQpV3N7FmLYUvagH5DCH9UovGB
xroGwuKqtbKZhj5UqMd9spV+engflzPQlo2pw6njXDBolohQadpvJPerOLleFJ5FGxjkaCbnD2vD
ifsk07ho9b/KSZM+aZDk4jDyNYqjUg8UIhNJtrUdRmM8GKLLiba48A21Uvzssl6n9JnCKHOkgCrJ
PNEgsHjUVorivmFypy0YBpWXlMCM+WnWLPoYkmjNXm24YDdz2JTkv+BQr6XWZeNWvqqMFs95MsNn
9dQn7aCpuutng1mRlXU57im9FKPPYiuOr4UWIlJStMjpSZS+NQYSvuCXrcHSriHEBhSktVCdjA2t
TppPYmtreRTa7dPDrDw9ijvZRI6N8Tl5acc4QWhBTxBBxSm02DPVDey88wXqyIYH38LoN3Hs7xj6
vOqICTyEzQupZWulBaQrzo3YzCoGXe6fe+fFMARtYBgXjsDmHzI9vfCXwvohcPY6cKWC6M84RL9L
bxAjYP8zyfa3Hxrgdp7B2/HSPwod6QlH4LpQJERukhyhOUKm2BI9yOpa0/Smitu0DcY2aTaWDLpp
4G/A83F0fJAB28HXRoLzsX8IzB8VH/Y6R0QGutw1EGQtqoei7zmxs7gOYcNWhIJ9ul3WA2Lc4Oza
aejldyXfQj4xGFkcsnuFW5QGb+NaUFEq1gt3Ba149AlajqVG6vbFf9BroG73uIA5KsJFCE6VhnXr
/7mAfLjFjOTCEvixDrQOHxI6FWBRuM98vS9XkNhbf0XCHzji/xL2gRikLtJXTU1wnBmeXTIVcxbR
BHRjegkKVGgdGs+LXWfgLzCqCp91ZqK3orIuXhyjB79xCZVFcqcT7zZLV9gwO7Zd7REv8vcOWM5m
4PJxvy/WQRC2LQRha4jBF97I4mLzMNXOU9KqD9qG3rhoYQ1TNRNI7H7z2yE1w/xdsR4Ohk2nV/Bo
DZ6VMZqoYROZbT60asCRJaBlQi188HxJEytsIu0Dpxcg5li+WML74y6Qe5gCrdBEytg3iUbMN22F
2pFVLikjpgQsYw1qOTtSd4ieXZrtwTevbrbTT/ke/gTtqwKNAxpD+9lvRcefO0mk06lApSguOE34
Al1iINHildBtTEwun5TQROD0y34k4Cmn4CDy4yUcCxknrLBmn/qusG0TsetrrY1eZlb9VkTED6EC
8nmuarpkp4KndfWdlw/zbFfFOKgwesPVBNqmuRH3GqCTFrcxfEH8Nc312TkcT+CGpBd83cElqGMb
noI6lon7nPe3wf6Wgj3u0x6doAjRAkxLrI1ku5CXl0Hqch2oxM0xt5m9+ivs+JGhFXZcgyFAnC5x
fbunv+F0bgNkqciqSoV/F3sdrHPSWXy/N0m7FzBIrX7YTh5ywhQ4v0rtiK82DcZ8sQfL1QTkWKMF
nOYmeDOSQcJgBdOpGn5V+T+F/fGABLym8TmaYp3ihAGf1IrFUB+Db9GE3vEmoFHtfbeVxNtSKKB/
/c4EQi47TV2RF0CstA/rMgaLB0hyr+lF89F39dW5Rs69jJP08mhvIubBFhUOh/022Ew7NxG+5aTy
siNIjJ8JPBwv2uZywmb4E2usx6w4Lkm51IfoOHLIgANeSiG490iTQWLM8U0erjlKlNaUpNG5aN6y
DAWEcXsyt3Mir6Y4bcXyIPBRGoHxugdXL3HgiuDKr/qPkHOB0Z2ChQ0FX+qAuZ0dQEbiqVEu6HZf
FDqFJ2Fn2RraQXf0bq7dfjhcly6z75u2mtqoZWSv88A4M+ZUYVC/YdJJxLNNCdg/L5DZyudO+34U
X2egtli5r39YmgVzOnIv8W+SHHOZB2+F7ACtiLtrtNM0oFselQnI/3VpEpQwpENvm1l2CjQr73Nm
uks2SDsu88VsBNJDojY5ZcF5XOetMNshE3h6r8gznqa61mHLxRgoy9XVM0ZlEYn/Y3qozJoxAiTm
0560xVuxIsaUolLb6Th5cNP95K+OFw1NT0kUMI8YXGCbqxK1LCtHln3JoTfTJBILW/NjCHPtXv0L
yvfx7CoZOQJfXf7QwHdF9k+ICM/jaxLb3G9n7D5kI63msHBujVxTk9HiJkeK8Wuz0do0fCEWUqCF
4hifA19XWytOOHHB45tuQJKTwC/hcBjc8WsTOzYbSyj9CJwaKh8dGunHDhIXROg5k5nBoJ2RzxJS
g3nK8254mrTJcGjK9REPt5dXb3glGEC8GoZb/mXuaYQYb4gqVPGA+9S3Xp1S/qasOKa6x/DYvSeA
rxEwwfNVDxSm1ZAW/EMbs9jKQqYvAWwYt80s0O+3n9qAyl8ewGmrs3dXaDOvzKz04a20ylPKjCl4
u3p2eChbVnvLbHGr/FLNhPoKduXM9GGOQLdBWgg3ZYRB5J4mTO5uYWxTjdkF4BjK39pUEbFgbXXZ
27MXObyA2aHDTDsbw8oSatAnz1ttfIk26AjFxnDB1PVnPZHy38IXSGzQngWjfqaax1u+++Dy2e9e
fWEoshZPc/X0vjBfEgdUHRUKK+cEA9gc+G1Bsybg6AMu1BzJYgFfieJpNnyDTNGgbBYYlimMxi4z
o7AjjxZ8BbdVOGSnb8Xi5qpbOYxUVWNbf5Q9GYEhdQdND34Uj3T7yOty1fetdyR1/JjalvJ2rRn3
POU02bRz/GnT2+JlvfHv/dpVPftzDe5xuhxhcSKtGNwChfninOX7PJlNKKWH9jpNSFrdLglO0APy
ozcnp3tPr///Kz5BUHMRQPicCcg7XF3LE0YVWLpvKdY2NT7NZDTELJf78uAByUPAtBZSbA+74NI4
fcwXIGAbyg8WaK+OJZmigz/EQwZwbMDoqcChIMmDjfEmI4PhOqXQ2uuiy85ewwia6k/c3hlXPspc
JmKudDYTSRX/Fe5k9RShlR5jF+Eknxy8vf0NVJ5MEayWmfoIwu9gd5b15BvOTyWnOo7CeCjU1KrP
QvBUzXDexMNGYlGoU6FggEY/MmwhOZjk6lV8daayBB83di/a2Hq+VbMWmgHP9IISePwWQe7vpgfh
w93Thoslrd8rjSQaTXLMFVkdbYw7IRM/BV4S7GKGebfYklkUPbVdgUjcGktyRrqXa22VEahhk/Z7
GCfx4CSs8X83pEQ4e1q4n0ckuuCjwgn4gZ/o4IRDKrMtTaKehdOXxJK6fIJyJi9qzMv8EmXg+3sg
FtlWiO2GFjLbFQ+CqqzkzJZvczEXAOVtQAQt9k0hoHWguE9qkKasOBnZBkBjNL7Z1vkK58hVvqR2
LGu27/j6Fq7kUlGxVPo8ZY5abPskenp+7uDFz/McQaeNWzjZU6rYgx94L+Yz3bqaEAjAVQmBIW0/
3T5Jfu/JBxVKS/QdMIa0NWQUsOptB4zbjE8DZec67bldl00TzSb9egvN8jvkDINPfUowj4nn48JQ
Pjucc4rEQaYTCmq+WUgLYwv2+CHwjqkMlqDmJA/dxRITVGwxoTUzYpVWmY/T7qxMO3qYMKHVNYIV
cyM/3mh7pn2ivloxIwF8aBVsTidMBc1ww2e+wUaty7zBH2E5WTgeYfMsDL/5C0b3uif0au//DEKO
lcJJoHNiyT8FODjx/QQb40wj76trawL88v68pxS76EeDmJ+u+oSEK2gbOEGf21OXaB1zV2Ha2P07
dTGUpxcglZT5qvbeP0VqA6ug/PKOiIRmhwETfe/2RiExzSzKrU68pGmLb5DsFYIwFEmbXpGf2NYN
DiJJswndu2GVfvDK3inCfslcrNQ1q42DO2bCQBgYUms52N5MhdpC8e4hbCRAMtS9+81srWP7Ino/
3g4DNHwTO1k96SXVhHTu0sEBJUBj3OBU6f/9fcCqFXwBxJ682t2bvNkVE1hnYbhmbMT5AnG6hLFE
I8mgKZOyei1oyLLVaKQ3Ctb/cZSTHZHV0gfAKFuwi1IxinkN/euEkQAPmDIIW8/Pi6Y7Mc5i3AWM
ycvAC1V/SDY5qm/WgQEcN1KEe0Eyo+6jO2kktV2yjalsg3X66c9YRNhUehJC5fTSoemGteMzStax
MFH7Uq9AzRvJaV+6HRwq9dFhH0YlfKx8TE+I2QaCNvlpLFAPDnOedBpCozriEwsrgB78+qbr+qZu
Kq0R0wwBcNq+KRbyPuiJnL+riMQvmAprB0BJLCOD4k++Du5VfwFjl5VFxGYyyWUfpOmN08Zgfrak
f9/3g2sNpJZ20cnp63p7/jS/PLsCL58Sc3JGLJv82Y1hMH36d9OfbmRoGZW8R1P1hisRBh20PRQx
bH2eQiOmR4RSVqdX0jqI190yJgs+CCgtCS7ichKfMeahe7icaxgZz/waSd51ggyz2oEDwAy22FSc
WBUBLWvaplr7yQXyCbVenAqb9NM5kqMbXOQSKTJiNRbFSUPj8GtbpS4i7IXeWvOifccaTSxnlW4b
6O5BwbLX5raMK69fl+JKgbQxTW//6DIg3qQ3+8oK6BZ1SQlTA+rGur+FzZ2CTRgUIarrcn1mDK0m
U5guzqsNscwIMAgAB/kz+EM+j3/d3QIzfriyQul8v+loghFfjn/uzFOJ0rNTbAAqAhmYIYHE9fTd
v+vItb6m2wzuFmVDZ3hTFiYjb9ylD5ySfFGQUyNF3LEwYaHE3yAjRy1tr+H1W2scV7OdPNmrjKn3
IHlUC3I0ZzGrV5anKA3gJCL2uK0Yj0G+039UAMyA3eW/O1yFhVTPbC16d4L/apvHgFbmOeypl/Fe
Q63xRXmXKfFjF2xhdjUQpj5khCQ8671J6luk8YgZR2wlqIMIRJN/cRau1grUtsR3bJzttgNw1i2z
DwUO4Kq7yIWCQ+t4BZ08flAYvkJhEjOvySxNZabaPEyiSbX8mYb2pf8FgKfgkCdRHQaSHtwIlWUl
6p6A0wbSUYg7GpnxQp8k1LXpnfedSI+PoPp3BTCJ8QKfwUV7jARHDU/OkfPkBvv0scBo5jGcRN8t
PKfY1tOl5AuGM33Ls8ExjYMTSgSca4Uj1xK0VtWyWiEQL9IfC2YOqssDR+PwUm8FUiywB3Wt4MVL
xaHT+Q0Jx1Nz0gucuDHwMsONGjNAj9LDQKX+tTbDRHkNIfnpANmOmoslKglqPnyLIeDdV84xe5Wl
37QTNU2ifPO0DZ/pJFNGovRI8Wu65bZ9xGneoC7XUMkuKZ7x7AcIlLx8a6eZ+SxOfotc98NxkOrK
fQ+Whix1iB54mIhlua85jmGqrOYrRMLZpdUHy2EmNBOdfZ3GqPGh6JVeto4jRsQ4VoVIQoVcdMOJ
kn2GCFt6qGJRy2lub2TUtfQAc7ucQsecb1v4PKeG30uu8IgAH/8Hl8Q69i/obraspxgQOjveq/+V
e5uajN82EPDv9r2ALR3bGulqgQ/CXC6OKd40NkwJrPiaHYMdiSQQdV4i3Z4l/VfRxGKIxp/VxQ7G
zbBJbvm0ede6l8aEJyCOLDG2GOnMDMNmrexRSKNU3JEHJWsrNyy0uga4kevOxh6eDW0Nw0Ihh1oK
Ebtfvvx/pjExXxW83xWbe+cC4PAiwvHz+aUwH/xnRvrJg03SRzmIXotr2FrbuLaV6DcLt1JSlwH7
zuJjZJkWpLd8xKZBHtQaBxa7KQdw33Oxc+XJIZUbBaRFYNmIkMDNga9OLDOJS3K4uACeZ3+VL1Cv
5Dc3tm9d8yFmRkHlhRyNkadKwpuCCZk8lOZCPHTxQb211fxYLdUyuGEhW8mMcTSWh5y+46v+5jmM
nn1jQi8ERg7HtNWDLQWfUaD4zC2Qv0jeazumy6elQe5C1Zz6JQNjwtTE235oJFYJJJJYGKD/L818
Z8R56MbxwDr1DJO7wfj1PtZ5Mg79NV9j879M5+Vzl1tap3SNXv/hIolNbLLJPFSR+l04IKfNI2eu
DvynPDA+Rn0o/At34FOA5yu4wM5U7Y4kOPrbfgCb7MOE9WeX3kp0vAsfJ8BiHUoRtur7/0aDrdQ/
XLnKbiFdZn4zWDcw7itGSwEH7EW6yiMX5CI3tUwAnmyJPUg1qgnXxx0DB3r1euvl7cQwxtxlVKdW
uocv0jKzyc4BeWDn5aqsf0uhHS75VQv26FQdZeNad4fIXLziW3RMZDExV4lQniFKaa6OVJf1Fvge
pqO4YhXvod8UUHhmP2Jlw+VONw+/BSPGNNygcrk96JRcavOlaLjN9zfhldhbPvU6f7KCV8qQ2n4X
aLoJmxcZQqH0XSoeeAu1Sfjju6NHCWunqrdN42nKjHDKcFVegHuLItjaQ4URuKRWaUiZxxGcnI2v
3EzS3NIuhBO1ezlT8SrY5WF48Z5HIVmmhuPQ4lAzYTTPqmYCJ3NJeOv+knkQcGNtUPiiNFznUdYZ
fNm7Pd3xbLiP+vaqNw+EcgSJ5ZqhSGl5erVCBevLFRAw04Uc8K/YRjcYKcm1ob0WzL/oePTkSFBj
1NgOfyqPg9Ybjq6fXeypn8iQGnR0A2ipWJY/qDAk56fX1wUHPHnl8nIGJ/1cXVk0IhNxCcTBtosY
KhUVn0/qbsHj6NIVCpiMrPwJGbEAuViwQmAQHhgFRY18aRk5+ZpLhcZo++OrIxe8/yRbM+CW/aEK
XoHtpAQEHXD2YC23umPDktMIUE/ra6abTIFdwwUBP+qgKDMIZguIUEHdNJrUuI2zDATLIfZ2VwGV
oX1C85v0k8ai9s8VxxSWSkwMPueA7Tl+MM7aLo7vhMq5czQiryRPwI6lE2hYhLBLdUB7qiaJJdjj
1CFnfScrpjHcgG65/X0aHuswC4Q+3E3nZSSOyqaLppvE3esS41l1hmDl1fw+7kVutrQJd43zqKeo
OW3ZhZy922mQxIiwIkhzE2bitNUZy8PJ+5VttBbDS6lX+Z1N5+tanw0oeT71h8M3//1g2ZH5bB4E
nWXSe8TIBFUKev/ydz+6dYTvxPyPJrOvJWrE7TTjTWd9lHbkFqrd2nsJW2XqX31QknF1wglyZlCU
7+YxD214NvvA2ORXGLl1DQw4XCXfY2Rcujgn5l2ve0KiPRC0LlFa8qF1sS6CjNP2IbThuUrCLap0
gooK2qeg1llEfQLjh5T+aPMWaJgOToRV7NZU4ZTQKIlnM0lQvO2kN0QryfcBj2SVQtKKefjpPhSR
cTZKeNQOuGj/Z7oO4iNRQA1m9P7QHwLjuE+kDqx/A8tCGTQaihobTz2xU/BMMOol5j9ljD1Xaw3U
Bd6X2eOWzsoZ2HTtauprJjRXqSwFZ0YSiQKrBwsU6erL3LY9rOTYUx2JPLsbL3qkeW4M9kWpg1cT
Q1EMKRPnKkdKRpKeY5AKBbgsu/T41Yzz3W96Dq77O8q2O1Kfto0n4vQVgk41FAYBVaE65fXB08Fd
J8SaJ+KdB6LA6zZleUsfA4Dv1y4bftUU8GAVHFZ7LL2MnLpRmsv08D1QxuEIMdYwz5lWeyW1MPKx
4mtI06aGHMMor6/YgKWAEWBcXGXEMNWuY/SCcdwlOyzesXAe9RaH2LZez21m8zWEDUvIqtHKFMk0
pSIitx/cuZH4/br/87oRTxJlQEiGZ6RHaQnWXrzsfbzg8hCPNqxJNj4EQbbxsIUDj07TtEV4AJtH
huccKfAHklsT7GlHqewg41zbSTo6AQWps3+hsUMg2o+ctJ9eqKOATGAdxVbvKQ9zNRbLIIqYnxGe
Pll4aA3qki7oyGSVA8WAYEFo+Vp63z71RL/Qh2mejfmc9OT260AjlXPZxy2dbfsqwMuSX6cvLLXc
j/kJPsysiHFXljlfHm698wNMlQ9lP6/LDn6nfaUr+4pA65WlhOwkM3IXDTmEU5S2xrtk8p+c46rw
fjpjHQKQgZP9b+9XkCDy5FmU8gssArOUOUJBSFdn8vpZ0uAi8ecUL616VJ8MhG5iWPoQjNA8sz4K
OcJRdxkgE+VAUKM33Ls/7VLstxC7FQAAlfT4ZgJ0ZwgVjO7Lx+17+bmkyIdfmLFpIkVjwxYci4wY
wnj6fjgdT8KHKdY937HF5aSdK1Rt7JQIICEbDmP6njcg5q2JK9jqQs7+jew9OK4BoIYJo3kBfuvt
6llTId6QDFDo/t3s6FhowuNOt5VRERw1sW9pUqdZEa8UFitNQCG/qpfApjbUmkFDOsvWcKMqVtbt
B5DDlS28bRlsN4eFDxDOyiXptGWSmIduzFLolJWq9t/yW8lqF6iZGMcHY6Us6ruQsPlU11HTO4dt
4PKEqA4oFZfMI7tv5HHX46VY7TmJskRSJUNvqgEMoy+g47KxocnjZkxpalKJa9w0HcsUQTiymJ48
prBEhsJQiAfnPsFaPqrI5WFi6nLrCtsK550J22+uIQhifXyqzQe/FjBoqaYkMKYJMG+5GSbB3u/0
Sartlv4GVCjbQQggsm330O4+GAt29bpHm5mlr8D/XAfkyiNcAmEnUjL/268KCy5llJ+bbUQ9/w33
fHTTuNxmHQhazRhdRsoHHhSdlH5dmUNOjy4zmph7uOR1BPnNdi5phxvqTU801a/3fuhukG71IJ2K
ZpSl+oFefLhCfWOtGLrslGBB11Hp29RYKt5/wvRYVDtLd81j24uKUkn86pwNP3W0I9KumWCtbgBp
+UzkTqNVVrzbK6uWmkcpl04kgefgCjsxMbfqOaURbH982xoocZ4DIkZ5bunDni8EH4CE9Ys4skn9
d2wHDJ67kQ7+WdEmcoPmq1kw/EZTfvDTHDiMZYmvBjEcpQ9BuLHNUGa/F6VGiFSckGTg3a338XWs
KPRs2woEU8Rs4DIEmKrwbKXo055r70cFYfLbxr/oekR3hDf6ohBQii3L/n9tTVRPYn+M+Jb19qEU
q/IKAXj0KM+oIhOvmx5nQaZEq6p0Z7cA+3egUo1hrE3zX/DYH3KcTN765YLik+oB+OrxaC5EFpY+
B1/LrPJkjuHczrVSb9jOJvj7ZQfWRtPyOtvf6xypdtqnB63MsA43OmHmlrQLv5YtCZKEa+GOrH3d
zarUYOmfzuu1AtMIMjFfGvzfjK2/e97RsN34kQrf85N9fBpXJzDO9YWFNILfhB1ufMS22pwgpUOO
v5Cuw2haHue71Qg3VcGI7OV2h3RaA6aoskNyHp28O+J8bEQxYRB9PAtZcNMrPZoaQdevWtiWM/f3
tqQ3rhkkH5xRBI3K9ULfHxacM+axsLC/Vh0WEn+UbjvUwFRx7RVncfAW0NaT+fkNqh093OCUIxWM
8/2s1ELD7yfDeTV5sFoczhnEPYTiRaBSAuOBofD0XjcvgPbo2Dx7iE5eHBXF1jbsJ+S7KXv7DV44
kw51C4EVIP8U/oBW9+8a0HlXIXHpmxnCS62G0qaiaFVV3p70Xfb4sFbqv80IP/F4bbFU/0f2QhTo
76A5hFT6FYtxE5BsDeseqYRzZRPmjO/Y3PBqkFRy1P+XoDZ97kfKznK/YbaEROqFDV9ilJ62FRWC
lwIbmgNObviCCCEqm3di7GGuhLKK3+RqqAdWKdrY+XrAXoDJZDouvse87kUwz4v+X0nYISr6/YcE
PBUTRr3rv+XqcYrbCNaP
`pragma protect end_protected

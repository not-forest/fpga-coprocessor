`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DAjaYT4WJogQ4Y1vVH5jTaf1EV4pQ9hPfQZxzhNJSUJbTmELlNrKzI0vRSM8RPa7
CAiGwLgtx/mcmbxibg6rbhc5IgUXHCbWefdYVwULkDYVir6xc9f2Jaj+5i+VgOBu
xqAVeGX3Bo/K2aFcwgXVBGPpa7ZmIPQZwPMqo/+9E8U=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2400)
btkucLfZTWWf5GZFPzYH3UqJQ0fohQCnZR3GJgReaNgJ+K2/t75E4IpVu5AYfJXE
Lp2O+AoxTfuPzATqkCPF64FXJbK9iBs1e1EIZfMkRUr+PDPB1wHXnFtg+suKxCS6
bEGxj+WOjrWgrmApv8G0NO8f9dLwfIx+DTK3Oz83ZJb+lwYTJ/JBM5suhF0YRwa5
tirVXVk0SHvAdAKsbLnrWTucn8YryaiBCSn7wtiH4OuDB/3FYslzyiTSkB4y+/o1
sUBnUUgIA5Q3TsaqN+LSY+kQbJrw/LW/Y1UaQjYONi7r6BlAkDRBmmmFmAGbC+Rl
6cNBuj4FGdedZAoMc3eVs+kOkqKHqqGw0RV6JgxX1ZBFBQLPcCLLAtVRS0Gn/jJE
UpWsySeQXRtkAUbMa4YCKKqKO/qB+uDGShOQxa2vT/MYfiz7CcCTmOXDsNLwnlbC
NHe5yXNs8nWHfscFe8wm3NX2kUcdwlC+FYF8BIX4i1c7G1brngf+NqI1iOJgGrki
A+PuaBUJrSFEpi3UhNbyBq8mksHA66e0dFhsTYCbm+NG6qKU1vhzEP5RO+Q1wqSq
oEh7vXS1760L7GKlNhWESTX/xqLaXGxUN6owkGWXK8EkNRuqswb1eJ7ZAMbVQQPm
FZk2QLAFmxEvf5Op/e0Y39ZmDrIb15xCXLA2hzc97haeXwE1IiYNhjEDgOVZ2pvX
q6Nobv+eQUL3q7Jh2lmUlCLTM2U4H9SUlda6+HQ9btPbm09znWroLUy2g9upoXRq
th6cg5Qn1V2glJRH4N0iyK5ULilfU2P+89VOP+vBOzufAduQvlJU7lxNCKcBumb+
SXTmigaD3ejyy4WfMYOLFBa71MEVBRSmlRpw3TU+ZxUYKKrZawuE9FYLkP0YNaL+
Ak2IPCXTsia72Ld1AELp2lcVe/F3M0L0X+3xMg9JDzcJXlSYwrGPs51qUen2xK/J
Vw2mgKVj2sM/qpW7D0jCzxriDiQjU6H6mN6pd0Jxg6od9pgi5UUUZLrEev8fAQ3C
ER97uaproWkfCcbF2bLZu8gotlKiyYSp22BYEcv1EXlkdtURbOgG1uroBrGYp8bd
foAm3wnXvzvmi5Hu7ofVdpuzq2/M29S7vWMxfxtyLu0IvOjh5iMMPsvS+ChzXYgV
Wy74kYypSPkR2wz6gwKn9Hj1gBHsuTYKF7YvyERv7NklrY1Oe/B/iyLjCOAwlZSc
VvQug2ns/ZZuC6bKDEBtKx26ciQHgObuSQAMK+A9W6X0rM2ljcAN/FUR14dA3tsG
30qQhfV569CSx4kAQmeYMJYhGBUAI7eiSsVo3l/SAXaYNNlPg3CtU5HQnabPoFmE
xDpZjw0HggB+F5HyAU5njZN4T0jhTFombcXrWzlsxWzu3nQ4VAQVTOlg8snPd2+V
AJMC9OuGTfH8HT0WpKokmVkYDjZkQhN1/+hLcY7ca7c7sey8wPsLEZtzwB7Bsmaf
G0Lfg1edZZSckbUuacGeBwS+6DyD8KPJTd+6CExYZGqrA/ZBAatgVKN3sxnJKFAZ
HMAIpOJIltGLyLgn8Kav5NCMwecTX9JLylEPph7VOZU2bm+RtR2t98NLW462CYuA
BmrpO8IL1/mFMriirazqg4brkdc7s6FQ9m2stQvMtLqH8Et6EQuKiASYIRXaYLDf
JYSmPA45+jvf/FfNJ35U6t/V71WLghI3DBkx9TmNgTGncn3B12O7KmxAE56TuCUp
At71VNJPxfbsHSGwuuJs4A/N9bV+FV2Ha+Ny1n6QPOz32YXnsvUxU2RGLENnvZKK
LM3wCtAjv0bN80MhhKSUcPohNufCclL2c2ptqNRb3qGxox7mTMerupwiNYarhXGF
BzPcQA3KGXq1dsmj+GuXbGAhjFBPwFiBgB5fs3o+0W8l9gsur9KE0i5hvwdJiS6C
eHs6s05h2n42IpFsmG4os+wN1qwfQ2Wnfr4NmY65F/tsZ0Ty2QbbwZQtH3qTW+Hl
tO4aiJC1oB5Wcz7ZvFGijCUZqwKhCDFcABLpXE05nG6PlVaWQQbE0A5P4SVHTFSK
ZDNB3YO0kBb1PsUAqSvskJMb2Xh2+/1HkxXx0NGuIALR/2aObdQjhQWjrWzwL6GN
gRvi+bmIzFPkySl15UfFMfRcOV7l9VXuZs7521EymnCEsKHQ2bvGFINspqa6zVyY
MgvvZaqjuaxIx4zYwyXgUsQ3ssDnQWmFM98edK6qHFo5bi5JiQGK+cMBWXd4RbIG
vQJFuWQWWH5LFzXXMb0Rp9uIRtmBKltSbwIoSWgva/XHS3KTEqW0dn2rTKuad0VT
sPnDKxb50cYU+kbYiRTUyjrPTFrAmtJDA4uPOlbqz2hgS2m1s1LDHzcdxjHM/mGM
BOQbtEPp4kctMmnTzd6JpjbUkhCOEaQs5/2LpPQnQ1FC5yuKQlmpdX8EK46dXRnG
ZPZ1DGImhZaoSxfFoxEfxjFZpoLKdOPySVz5Qnymy8Da4zNIFXCB9YlQJntavow8
H7qmS/zQaZLMzwZ/ikR0XaMNSJs1aH7GeYI9HoaEmbNCrIri5p1yo8H6zExCWpAb
CcfVMLJb1FPy4VOh7LPiivpWljia35MpQbfsIT1LYPjKLQV5MgI2yu2Y07VJZzps
j9ezcDdV8J8yxpIQ8D6YWnLExqmSE7E6Qt0lIi0C1GUIghma5fx7XT3McrDjfXiS
z8zEKFviBlTaUsSnbLcjFe8iL7F6sq62TUiboz8SkBl8JpzqGLmYip8s4d9IJ6SI
vh5QF30oKyjG6V2bypcJ9elp+3YbwJWsoIz6+Rqh2D862pwJI7fTXMcfYzBRVdlt
us9p/AaQt1IkN051cNADcsAvc1I1ouIWI0EVr3ynBIWxQTOEzFqPrmaAApDlDqGl
HkEHoJ5xaD9eJP6LWZ7pTzJBNRX4RxurwZLnuHxEStsTWsTJNHd90HYtjf8GktMO
98G+POvRtCc4XR79Vqe00yUFLM8wQnM5PVVxDPX1IIpXtKPJURVgC1Q3FLhFLuRO
eMU4fjNRrwTD437y7BDFDiBauYOm+uCiwfjRKxbxAUpBhTdm6CfZcNsJFBCQboxj
ZEmInzK5J7ElXTgh3KNYIYR/ceRXMRwZaU+OQFdZCpu2e8d4eXiZ1V6ilhCSsmR8
uW9UYdpF6aIQmCasL82IGThUai2rWBgSdvw8bShArMNi4AdwM7sy3zYv80Z/458a
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
Tlyw/wnJflBZZvQAh74XhIWLWxdk/s7IB0HfTNJPOodejSANy4s1UXyLrm2M0nNT
YJ3GUcuE/NXPP1j/UVhtfrMBfFto7a88f+R2I8UaxEK57qXEcdc5JWFVPuvxmTI5
F8f+6DkOBftyBXkksWu4GyyTT4vf1PKi0/6a6IJxgCQ=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 6128 )
`pragma protect data_block
aV04MV64jHotUBeN+YqlV1S/Utap3UoatfS4EO+M0/5Zsip+0VBomAmIrHOiKVbV
QDHLvqwTGrxluci2Tntc9iUx/R2azwRxMaBDc39YkXdZJFWD6qrSlzc2zVScqh5u
lKiyTzn2BnQuvcmxsLbt/67k96cGgGjyI7IaLPQAUhR36Vub3mmcwu+nT3mZ5/VN
sLqZvLu8KcCNyaY7JvicPht6eD1bVN2/rHjGOZyex0GeqxPmJdlaKsl2JFXFFPpi
cQW8oSdjUvrgLaLrDEdYLj+NX6UJEzxlblHGI6E9+s9HHtvg2onDSyJr25vNgnsH
yxYG7Dphsi9FoCo9K5zVHiQLT+QV4r7ehT2IVl/LtQU6lAR7YOJnAivxAmFe8W0O
Nx47V9gD19yxBHrIk54P6EwRMnNq41JDub02cwFmdvDp4xkOXG8Gp1hl5jR3SORv
YQDPE0YVpjzx1LjL5jde4K4XWDFBCxdoTUmKG0xhBUyz7n1QHEyqqHmwJNlnfyGR
7QRJh0td5ufgepC0UP6oH/raAD/iffFpCtHxVY8bTogqfKybPDaejPAVPiITbG+0
NosNHum9Xjz8Z/cTryQLHAhZfc2KyrQFRqBSAA+vDMJeruzVmPlm+glnhZh5qOEJ
Qwd0wV37BNITEJfB2mq+cAAXJNx466TSg8h7oH/hfcjnIIKa8pyyP7td0g3lKHeM
uy76CD65s494zATnlOu8/6CLayy8lksw9zDTelkICVRR6xg2zzc084244/vAQsR7
Ekaieb6ZsSIuRXocJBMJQVw98EiwTCaUhdTlOnSAWjtiOqFiAznd83hGGEgh6Nk7
azYdIdimvyum/5cpypH0HEljNSAopeXoqlxgqYXM0dzVkON6pA7N8cNERRYxg85x
kBIexSsD1ZuzCQW396BZM4Ri6GQg9lK7TqKk7VYoB9xf0pfjVU5LHouX0GQaWJ9o
804VH+cQzthSoeZ/D888zyyYCbk0rRuK6gV2csyWp12kNTrl3YLHpiYocQ4hxc7g
S0h1E1f/EkM7wH042n2KqQ4AqLQici063aGI+N8vakL6GaFml/AJjhzMtglzko7r
Z6K/aDRgOtAQADaQ0HwoMAEIBAf8/PI1j6k+5TUfJMplOl7qxV0+lAj/U9cYLQ8+
IxjthaY+c1MdmaH+XR0JBG6uUawu93HEDrJN1SE+CjC1H2Tr01uybxjphOZKEzz8
44royb8+BXoCNK8MFwim1X/UO/bkaTILYC/yczXJMvM+A4EZX7BP36HDfhTin9IG
WPDPvknTUviQL6HJcJGQoNS2SO1HThDiBpPQEYcvmugCAY8dI/nDPaNngrg5AE3B
+SZf4BmRa1PH8BHEs3+rZs+poJ412EDEbGgdlmOAIaTUccgkcMuMdpubi4aMtt6s
wGv4tLQYRQWPFZvmd0dEVxqjoIphRy+qhflzvqht45528TM6lDMEwlCRhNAGlzrl
y+rbxamqe4AGCtBKRFYnK31lUmiZcJ7Q14GWM00Ht22GiHoaqLydlVH4w9x7xp2Y
av6FUa1pN1gPanM8Wau5wpw2U4o+CT3S2Zk3SQugbO9cZUJW85T4JDK1vz2p2Rfe
AsViHs2kLpAWtzoq6XJLiMnRP9VOzm5qC7NhFBHxnxcvqiMa+Um5e6jLwQ6zjO2m
rKC1Hvpb870e0XJVx6GFrhVDQZoNphvdgWD30/ch8USMPALvv9+VMpWC/TM+x8vv
wMlkr8kZn9OvEOF8dSDpbpxK1a2VDaOw+9znf5GEKxjVBwCQysnlMhsFf6eoh7z4
IQt2PuOXsGP4kZRxNFjMehcx29visibLVOa2BcFSZSAgNgAnDJt5e/AVtNCLyxrd
E6LNxE2l5SeLjFfkjzhUehpi9SDkvqMs9eww9UdBy7srDa2LA/IFg9p8vglytmIq
udKSbMDJ9c0mCcrDa0K6J/e4FrJLg/LbWtJ+soMWgU2dkYwplBmZre8Xc9NxsJKH
PnVB7DfIMEIR+TJN7S0f4ujS43Xl/JSkPYzdOyYgmSWlMr+3RD/X6VTjPp112nL7
MEGLG67fl+GNO5zBwLseK2VmVgJWr+R0OxNrY3GlZuMWT/l8/YHsDAxpw1MV+SCM
l1Wj2w5lUC8pHpI1yQJrXmedW/UL42jZ5zBUgGge4II89c0tTJD/9Yeuf7OeNlMN
hl18n1TebxIL+hBHrwKGU1r+vjFHFPjSxsBFxnxYVcDuPeYkZlb93PNPu4p1jYHk
UwWhrrLYre5lJSM9nMY/YGJHBieyUADWldvLWuF14eHKJu7Qm37et2SZW6RKTD72
EiPzfAS5ts2d1Xg2HEyuECVehjgfCl3bwdbFhSvl0UCD4eYMynlg7lMYImvy6K4N
aXjP/7YpwE/VPcQJHq1EnYzc45Z/k8zL6Z6NB4gD9BpDnNe+xj8myKA3QQnWRznT
jYBRbSr9SNzw8tFK3T/uT+OXI5s2GdjiloTgj5qyisvqWg12bIKb9ihdpFCf4X6z
rkSRXRzzSBC69RRcchpr/jIejocVAOLqrjaCABm8JPQ6uGFQAIMS11vrN6CktEHS
qCXLrVdRLhmgqH6Y/jTJELjSM+Dw+Va4fFkQqQPgeJu/iwZ6I28GC2LcXtvb1emF
oTJ5RcfY8Vbo6KtNIJndRXxvF61Yw7nLu/dxE8oTTkOV6syC1oyPpCVFeqMy3v74
XbvOUocZ+o6he3h325fN/LrOcEsOahc/mY2uUh33cn/ke0d+uJsA6tf7xFF3bO1T
0Mq5oHjEo94F7v9kKIdWGAWTPZo2tInRIc4DyG+PoQqjI00rPpRpMMvWQINLaubZ
nSqeENoFykWwAk5+icS/e6kSwsLN5+hQ1/EL3bgDIyNwK0+gYVokyStaFUtelYL2
bc8T9VysBkKKd316XIZJQV1FO+rHhDO1llYwSt8gHHHfXx2/OnTSDJLttpz0lxIj
uT5mPutYBQoXEX4j0emqCRUTmFXSgQgcu9lTf0vJj7MBRcayJnzkMWdSW3ByMZ56
6ZFxUhV5vNQKCSiWCI+DOK1ZSOTDXh8QeSR/LF3t+vtPWdXsOh2NCjQd4R284Qs4
cUleEvnFTKRbM+Tx10jO5m84Ayaj8WqAu7er9KKdQc1ojvuWiYSt0OdAg34HOIsQ
Rm1m+eRFMU4yR425AWTZQToITVdoOx8KRtoRFVweto01toYfGY2LDZJ7S1uBjHl/
JltX0ZfuflkzmDApeX8MKZbkkAbNA7flBP5WG1pWnU0RbPMFaA/3fO7mMMNC/bw5
GGJj/HTGTful++z/43zvR5qAUX3BQr93QdUbPN4r/rmCIV1HiNeMs3wiRvQai7JD
WY+/fl+hTTzV6Bx7MGGXnEh7heyOT01bnDhpOQQ+vCyBcDb6vpjAA7hKT4FBJdPH
5EWcuxDkr01urI4hzig62VInAv4LrliQEntsGuTiDwHuWnQGMQRfkRWjyBiSbLpt
nSOmmNOf4oia3613S8dl0f+d8ZApFbVSg6NNo9+ZzY0bXkzz1C8Ql/lOXbYlL1/P
UI4iAZ1idlTS+M3XSfOB6ahktZEdbdmqaXPwVmwGnSCAaaBIL9iOxfSCGfu3bRwQ
TSD7zCeh7Y4u7IPW++6IZRzwsS042JF62B3exTIiSxqJfyhWX1gwGizkpLi/K9B9
LsjpIX+nJP0w35UlgSgK4gCnUKJrWKI2e+pjbL2xg8cJ5kajhx1bcSrtNPkdQrs8
zGGqTmVIGhTf+NNZRvFb4c2wLjwghQBA8d8M3ltdWD1r5tgQSuh9kyb9uTqTryuB
99VpWPn5GZycGYF80yEaJj1GOtCfELSQ9W7z+VORnyRwuxN1uS1uOsPspRTfwnO3
13y0Mkc7F1eMXlhzcFO5iddNrtnQwpfKITfV8ryhFriXYBe+3Lw8QgcyViUpCC2y
DX0TGpHjbQXahtmg+JSxBmzLM2f7Zkt0DcrrJs4C4XRnWK4dEeFyepkQmAnlO5Bq
dxqtkDxW9SnIwbYCzin5yVpBlPuQYO8/rdmY/L1IwXI9+sNmoPVQuDKd/lFF1n2s
P5iXhud8vb5/WA1zeEfyamdfX8vQS+8aQhd4ICbfE+veZ8P7oav7Ufk2ziKPLeGn
yp90B1U/37ylSWGEp48i9MJf72TkAGOtYtVmR8PD2RGOM1tCC15aeVvRgJU70Kcw
9UhT9QAVyvJoICWuzwaLKmea8yEEpvprX0/yYUPbW824YxAGJRBr9xwXcXgQr8h/
ty4VmtEo6sqXWaMGHmOgcS12qLO/dPSJ50JJlgv6pbn9adnvrW14q3EIABx2MOYh
y2tNXblN6+t1U2zPPAoKcnBbMo7DOscuDvEVc/lC+fRpbWv8rOnsScy20okjmKMn
KXhoVJCO2D+117rQe0POOlugIe++E+cyffpqO4K36b7r3yAZ1i8TeyVc0e5xPYSo
cazcVZPhG39wj8pCcSLvKSmDFZisrsNLKOK+FFSNsaRNrWSQ9xFEgN5bi0uRQiDr
8f1LlnuDSy766NfR+og3S7Q67xAhjbTZNKCWpScLj0SskqN8k5LhrMR3j2CmM4lA
B5lvjZ17RyIBNhMqYxPmmOBlc5sK1QxF6A6cd8NRZJ5rrPN31DpCoTFKMFCu5bE4
dTSmehDA2awm3i1tqZpf/IwsTXoOJx6d+/wpPhO/7e7y8zxAP0XQH1Kdgmk5xC2N
mlcvKUh9sauhwOvXScLdi3n3wGa2/HGc3ZBHz55cQie8nSZfgFiTuMVy860htop/
VaoLO1cwEIKZ2z6JlsZRRUeHQuP3Ka927dAYYwNfuZEJdRX5XPadPszDjLMlOCfm
E5l3ykI6c99TaPIicy4Wpm7E4Jo8j/Wdqe8paxPeN5u4W6lX3hyWQgyIsnmB02DZ
UiptT/dAL4b4XbMoL3ydF4fshAOs4H0Ma8sFO7oRoSaZYFkcUrS1E3n3AWr2UsoU
clg7hyorc0fFL++8KOLT6kZ4a87lAlMcVVt4DStYDvWdMb4ly64p/1cl8dY3CMYs
tzvX0/Rbst2SavM0F7B3MY7io70FVbDgq1wR02YM/YNNNIMB5DssT1yTd81YJcZD
dFGFfSuG+3h7sE1ss/JeZpgihdSfeJm8nlDs5GMbSyvuqLHzc5AWRA7zuke7EypQ
zBxsigXI8NEAcVv01qzciF4H/hQ/plQKuGJOf1cTcJzimZJpsS1PoICdvvNh0Xoh
DHbQe2ECb/cqzdzzGSGqCr7XBMFfeErhZdGaI9BoJUzyCjWbsPH7W+Uh4cT+YhXp
KO/ebC8VApPTK4lFfVI7MNnVyWMWl+eQUgndyAfKdQ2/3jWFcEKPUTryMBrzBA39
trWm58KXLBwKTaB95HSSL7whU4tUXbliV2al4/3SvH3LOqEDS5WkU3L2BtqR/p4/
ho7ibPP5D/3JCJeHv4Ult6EMWiXeDFDaxVeAceesiwDjLIgZnq5tQzvpYx6rTkK2
7YV/bb2jqHh7SdohOF115F5y4fme6q9R7PrbSoI8m0PErhRsejv3Z2+GNYXJ5DG2
PgfWsJU35vjUdmzWiXGZ+myQdmcBuRwQbyZRz8tblHmvnWB8hJZQ4KdlhgVEP+4T
WP8H//hurkFeO32NvWpvfqZGWb8pIxKQY3oQfNQPViYuh0M6zCgARurZ50QQGkbH
z3DVB48Ixfr41W+A8wIx/dPPGfkVEmxd4qpwvREQOf03zuLOmQ1bJ0+U48/gpW67
tCqSl4XwtVJXeBnjAGeJiNZ+gVJa2dFGPh3qIHfZHkWFkHy+N/nP5I2FHYOT/Ubt
pO6b8hJPdNxsr3ifV83QTo6HrVBBpmeCJxQRQ9CIC1IgNiQvEtjFbhImxWI7qB7t
GLdzv9U1IfFknWHES1KAsxki1YdI1zvlKJjAvVPvG9SRqsd91OXsU4ulzyWhjWg+
VoIhFhk3vzZQDhk7mzPZhDa+2v0cngqKFn4kZMf5QNdP876kT5EjLHKpVcHLVfrt
kX2w+0S58vMDU5smaFGE6IraVYxQNNXs/KolqaudoLEXdnNJ8zU97SZPaoHSQTBJ
sEmnVvSNVUcMF50wdo8tJkkH224blIQcn9DMl7daVnSUiTKxUA0Quy3lZL/nlltQ
uVKFP4r57sxlqXBYzXtuzzU07sojHSjx4NWWIgW3+9nUPZqJdm9lEUgAQ85HzS44
xkoWbiwQlvUEvcCXrecjQex6+qXpSMQu644CsAHcydURMjF9319ARAu5lRXOX7Cl
31bXwV8/jqmEq1MxcYkFlcpeqtsBAi0ZsNCgey4nWKh8FhE1NSo/b7b4ffmcOx5E
0ry1idQyEnXD54vWtA5AxviPCDYqdFBt44zmcen27xry4cvM1bliNOs/7J1/bT1N
LUSK5UFsebyNWGeP2bKoBZ8ARmKTCCXB4IvwTTsyYJDGhh5z4z6zPZrhEhRj4JIF
KnONg8oxUy0FWifeLwq36UfelrMWW+wQozoyNRpo4B4ev+vxKj/3WjwQYeetu1zP
4e5E8n3uIDsOWt74ZS7HWxn6E03Rlw3uemwDBjblwFrzvq1DttF/LBjSfy85JjWm
AyLpqoK7KPAt8Ekw+VoCKjtAo+8c1aoc/CTQdNcB9TedA+/ckPU7DFxv+OGP2UHL
7rLk2leGPQ5TqcA5OsttSxun29bnqSHjqhy3j2teht6cAWV+O7WhYbCB8fzl3xt+
NIL3iTHxkVuGWuFQkZi0Wwh8HVBh4BAKwgTnRmGEtxmwVwMd0Hgxpi+hd4DqcSHw
0OH0VMlnsUDTTpNTV9qM/I+8Bx1VCO/GzW+AaKtQE9uaRw7IfI8I4Dao3CYmSk7J
TeNRHLFYcJDAbv3jlPHYAtHELKqbmqP89FhQMzOZFm05qp2fV1GGS9UxsbR7SfnV
MWfakNgQ48QjdULS2X8/RGVIhsSWi/5Xy4sTgtclCWnywDcdDgBT1Bn8WWYPRgKk
//34UdsahsqHqXuzOHImx5DXskgOsyG0owka/Kmo6D6JnamJj68uUMvwglLTZQir
Ye7AkcFh9LqGiDPzd78p1PuMOMbVdSwjkyC7/uJM/XxNdJcCQAwAZICb6HaXtaTC
PNfEKuguo7Xr7k0maZQxn9A3e42sfcwLSkaZTlGX09ZF/SzQAC+xcxHs++14HMcQ
4JLaL1b9s2YuEmjE1IIY7RimLwazua74bJj9GVN+lxwOOfB2g1nYWACl7AT0kZyn
0dkx+kZeSrIdLN0Gu+BUN5SJRWSppHnkvJitOClrBAkl45W9Y+HM9JfebudEVFAr
wtdxZqWgAyU4izi61jUT2o8gkT7sxKp83sda8GeQs1973wegXxf2xrsgPPsl6RQW
C+bEcPv6fAIYEkXLj9+uOypkKGa0Glj5IEmU9pUwfLThRFub+zlWXqs0holI11Co
uY7P/YT7P4iU4OV1qw2tLEGbPZuAZksYUAVX5FyjFLjRUA3Uiy3RgXh9jHmFkwVX
m5fin/UseDaGeJp/ionN9DUcClMTsjk3jQIMDucUlhcG3Qi6aRe9IEQ5avP8abPX
7MqQEXeRwE3zwTgDBGG2rw9Uu0O0EXxO074E+omstXOxDLeucbkJefAqKWuAaESn
wbaFOnt2uo1y3Xri04qbPrL+SOYB4hrHoLrG6Vv1SGQ/FF/wvNxFQ4ERnp8PtI5J
tk/ogm2QWezEKbjJukO/nqPDQTFVbL0eUD/G/ns92l0Fr6fVFIt9xBJmA+jzZ393
JggxsXnl6Rsm+7G0c+hYKcJmcnw3LrxdPVdsA58ALS1KTvNqkWZE/9gdOPKYbx34
kSxy7mMok1SKlaVd3Q5LbYSAyvXXKirEC3vNOc54BmhTMJ5GgEvu8PAnWIAXeKVN
untiJdT6lnfaTZmrGk/LQd+SNUgZ8oOcSyJ9+YgftmWvwdwJwLZ8hFRC8jsvuslQ
JaO3bKgQrf7V5dzKgA8xURHwDwTzljdp2hZJ62K66joC707Czv6QlO39aWEaCAaE
DqhWyzDlSfrh+nZPUwoGdG03WZG0OsAlwZ2/Zsjtk2lsKk2VEBrHs9XfTiuHJxi3
Evd/dCIfc/6AYTqZlye8ZJqZAccl/BcYRp4sgmRJo/xBucqi8fR3Nq425FmSdpo/
diNQ0T2AAcDFjArJ663jiU+l+0DFbF5TmzFs0JE6Fevj/dBcKFXhd2IITa4CU9FZ
ak3wRtlPjNKz1ac3JJXG5F6jXdDDcGmTSJygL3SaNk4=

`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
KzclxTJho/l6frpU2+hmFfiOcLwkLbU0w5GpznNEbhJV9JnWscwyA16TjGREJXbQ
5tJDJtVB+LJlJwO+YK6hEwsDXubnnjGCtosmyRKBM2HnIpLdZ0NaPK3zH7LYmrJ1
t2ONYwps0DCV2dABd7c4Vv1vF01XnxMBP9iCXFCOW1zFZB+AIflMA+5lc1bCGasD
YTgQGKQ5r70ys8utFFIBkY10dTZBnUacIcU+O3Ro3iZX3YI+rChnBDqzwse9xeAA
h8YFFl5mSQkzHyTG2JPheeF/JXnBJMX2Ljs6Vem4unMbkFu7FFi6uh+Se7xzZcOA
SowMg4+XdAj3Mv2n7/rRZw==
//pragma protect end_key_block
//pragma protect digest_block
vOTUQtIaMZuA+o6lAmOL+uhFqy8=
//pragma protect end_digest_block
//pragma protect data_block
wZJ8vW7uvL0ghs5fthQbngizvc2MfdMErAv1Wx7MBY1ECGkzM/j8YIhHW8tX/f99
jiLIPp88R7ObiX3n6I9LGWN1W6N54k6NNzY7TVnl7219kEsUaPXGvkIX+Zbfx/z2
oSNwxuLQYW9OB5NJVC3HS4LgxALX5ZyoycNniCxsPMV+o0v+zBifcgdL21hI0wQ3
OSQiKdYcathlqy32dRrFeHq39HofCCfglHyZEn+57YG7vR+OCC7+Z5M+naHnQNNV
GF9dF5ZuRt6e5yHhiwK3qhpZW0jGoE2B+4ThDjxiazpyfEjYBOuuv5AcTRJZG6kx
YIXgCCt9u9Xz89SVmpifpMwo6niWIAqagbrck4+oRIJLzEMujKY5gdQf2pqIhM01
326BTJvbhTUTwVggKyuRu71O5RpEwD0m45zFdTvp6XQ6fyZ66/PlKhXmkL8BPzhH
fk45NhOekxQZy+1dj9YEf4MTrgslrYw9Jq6NvhX+QPHO86/oxnLtwaobNtHkByz0
G1tU/KuhHeagVeE82hsGokzQTFYNdKqjae/FfiypNOiIza1c8qbIl8JtQmMm6A0e
C7n3+/uS8PIxx6xRFTKrP80SolikWd+Z28b98xPlqx+UfNuLKkHzSEsiXv1E9ore
qXZTwnIpgv22lobDxbxRq+8TI/KPHa8n+CQePRpq8iI/S6DesAFfH+R5ZDhlTtrx
V1tFIlXtw06nqUJQSfjkP9uwWbhNCCnM97Snu8nlSszR8h32CZ40jkoV75WVdRZR
8sAV4ELxWyipBtjEsOZCEuPepIPApmWUyOZLDz3R+GUXsCD4sY53jlA05zoWnc7o
+EC/931hr7wLN7ufdHeDVIg/2ij04ijF8xUQnFlgsQLhn8gtNYF90EHQ1O1dYHN9
ZrvnXUoXy0iQ7OgRPgT+ELEkkTOxJJJiJLlcwWM63tDWerGvFUq+GiL4DVZZpUir
S6upz62oSqZ7WAYOrSLINNNRvYXyB0/2FNYrjDCt1VjF3BklJcfhHPf5rxRN2Hsp
AFOwRIAdd/HpI0Uw8bRVx4zZZrQmk5Rl02oEw1eknWfWJ/d90mAoyvVeeCSw8Nap
AYWY9DqWXv2WX0B3ZE/EKdyCi8fIRqSipOHeQg8W/IQldPGjhqc/dZm1T3prvr7k
B62rW0F6PZYz0t/IQuFEEVXEnYsJO53mmxmLwMXdRGsZXG/qixiEPzmrT79aVRx+
n0df6JB8+Pe/9FWp5jNgEQRcVYJnG5m94BHHgsBNH/4JwY6U3EZ55iNX8cQxjzPt
RwkFe5Qlk5t4V6hUjblyCe36ImbFi/twRQpt7xxMgTvKXEnYDTKHwwXsjjAHuu6m
Y5v8Uirv4GvTMRT161d00KuxM2QrVxpygysVc2KMi2WjrbSDUBMFd4c0hNXyA7On
+wNSJ9prm0YDLEcdRePLvy4tg+Jeg1GxXlyXyGOizaDdDLHML5d1Pq1J/CFT4BxA
OVFJRqGtjXNiGu2mx3NIfERB9bfiSz7IRyvIonFU0B7ER6s4RNop8bRwZ8d9XEbc
3GD3LdMoZwUQILaoloIei5GE15tAZUp3P0p8wonwUF+8JNma4aU7Q/3Eq9l4QOdh
HfMaDweLc0ho8Ei7GBp1fjmmooOchIgZ4JAEiOSvvrdQ+nnBqudes456+Ur9g5SZ
NgH6BpZilwAnOEoLHzFLagPV+pDb/sFBmZA2is7aXiu2f/rFsxcZDTeltKIWrPGo
JNRRniQ0FN04dEbqAdemWvrq8S+2dQx3yj8f+mRDoV5wDg4zNKHBaWQwzzFlhMeo
cWJ0PWf5Po+Aq/HB09NYr0lZdETOFxqGtzVu2zJZ/UXn1u8azN9sPJ79GyAP0Qir
nKYKWFsbb7AXGstQnYe5/EF9Ck0jEhmUiRHopdycJ0wVfTCUwpLZwlGofwDu7vck
6LzeznbFdyQcbsfJqBisVAYmkdYHlQ9rYqzVij+7L6DimpRxSoxPqCR6ZML31hz0
AqYI997iPTqmB4fhmaMrvuN4bEIgG6OZUU5VL3a7EPxioGo52EjZFgl7pWSidDkO
WG8MiWmcj3lFEToG6y2ialC3mZNLuOM3LVPbTcdmFZHSfXhyniXUvDhU9g+l2SHY
JBKlZUWwtP/n+fsLZLzXkB0S9Gc2EmT9vrz60HnnRmu3yhE6HXg+TVD3fv9grQII
juRVQ7Ld3mHExvatyk6U4Z3biCvVj624Ju2HKFtv951meiTfz6CmhsOS4XPV5yWz
Wt+asSkp5zxUNr1tjQhkBp/SyYury2w5zxnlICb8CB+dBF0/6sBtxBkNRXULeOit
ZUOBnzazvf6UrL9u4IiBzFscjeAQoelbR2hMtJ2EG03dif/hs8bOw3HrPFqzbPJE
RFdImMVTlSnxTo3yeitszN8BhcQ3CfcQE9fFhTeyeHO5B/LatukMzHXOdKQty8Uf
a7WEVlpsyBRDiDoZGvPUd7wtCK/dxUExkGyoShWD+eWTquEzrJDLZbt8r6q4RCli
Kyv2grahzE9wuO+iVInUS0uxI7QVgfQ54kT6b/yVJEJW/vkKaBe3HpugxeT+dke5
2I0uzALEoV6/Ib5epheyZp57QBeacyZOM4buXGTalCAjF+NS29gHkYRhLqfGrRaQ
gySe82/vOAz/7KPuFvDirmd7aBDfqMmEc3WorVgpTmADNPeX6/nmTeemg8W/ubqO
Io1ltcyo7l9oKdZhxwHp8CsM4Y1XQxEPpc81vMG8eF0lVgLuu2q5Of4NMwe3c90C
RLmguRnbW1mTg3J2k+5CRHIvITAqJKlT1HFZYk12ZlxikliCChWStfcE1EjhaRnV
pWYGDXG1brX14FtrGy11vVpTxLybLRXCZhoMpr25rkNEhdw0w7YVr7OmNFD8epUB
CgYoWQ6FKO9YG0YA4wLqcimhSjRoT4CDWpKAkyJ6LxPa0rDx5I/S8sBGsaNxHsHV
yD2BYAMiB+xGZrmduESYDea9sh37JisreqDmHdtRlzLvtWxle6DP89qwCRI9Bhsb
IMg2LiLUA5odb4s0wBWSDVVuMZVSm8Bf882QycBNza4Ce8ZRfg3i/3YK40cSKUq8
mEeC/xS6SFdmgh45yfselLFAxZ1mDuN8LoD3CWsOlt5LPhvn3Ss6ZNYK/r8ddnW5
DNaqgwbFINGPz9bMbVCkvlH+vPgUtsKuu1PI3gk9TqdfUkXWVFNvvb2elCS5yPbm
k9anDArWS8B1oZll7hgnhvQ746Kvcp0dSh9vE5Ic+7HkHHRoTBs6IR6buwuq7KX6
QF3Hk7PRVKAaaYiZn222X/rJlVJGKR+r90l+7DHfJuHLUuZSt/dDwQQmqKcAIetY
+x3/aIhSOr2o0c4OTtihBIHf39r9F9K09TVmZIafEwQX7KdJT0bxIb5dYHj8qVo5
HOFZZCREI1NuIwvdOQE1BfyCLuXMQ4Ujnzaw9XT2csO33CyYzMQE12mu1JkkbivV
rxUJxvFgZsl1xbkS1DvnjOoCeGMr5oY8BiGy9E3saHmnkGj5+cQTCFlduzea4afh
AbgYgkp7Sal7cwebgMEkHahdLofAHSk5tzlE6Zr0cWV0BWU43B0N2Mo7B1gyDHOE
yZud4fNgFg1Y04hTExERULrDe0nDrJwcQ+mOcd38LKW8Vb9EI3VI+6H1c0I+SM/u
L0K0kIRL7HDu5TPbx/u95zD91r6Y05KGYEDyivWHK0p8rCK9oz1rGswq9c3O6Hdn
JlvD+1+1XW6ejxFsOlSkJR2rT89RL8+JOqUKNBxNMDChj9BslwEslpU1p9Ut8TNe
TyQeEscvCfCqtPWD0c3cPgcYY++Z7rUto5/1+gyroD6/8EYl5ogiXxx45rLVd4TI
nLYjmQ1aqh2VoYpeB7iJekqNIb+21UCx8jFedXVubEaptxhg9oQ/LGPMa7EcKbl0
MNAYmt4FZvv7BXLW/ZoIj0tBcJR6vfBHHU0IY3Vivt8OMaCYHLIRFHry2CVXO6Kv
SxYJ9uhKIOvAebxvF/pCj6GDKwpnMVIajItNa5VKTNB0vSSVEOco+gSFYZuTFRi4
MWnMPNy04RCR4SYVRveRm85rN1lonOle79g91wR7VS5CNt0HRAAbeys9QODR9PJn
BVJ5zd0N69O7QgRd2Kr8fhqx8R3f0LJUOssRyG0cmD5t3umg1N+5POzv3ZLdwKPb
tBMdEKYxhMS7Ic1OfbP/c7QpTRf7WMrHdh52cnYjv88WCaDilVgtbwhuh85FPl2t
C3HVqg+Mb8+6CwgifNJwvJx4gbBQP3ZJ5KxGcvTECn0140hX1yDwrMpgwX13W13R
wSaK8cC+ZfqhDo2FIxjpoNEqpo/hm84pD6keKATUxhOe/OyH8HI+LkizSXCsD2uf
JaSHlIDSnskn8HJ3UsdAsxkPa7k4NVerchuBcxP7IEZ7OMX4IQQKKq7BXWBmBsin
untpATr0kDyIYhfWGCarw3jfGsqNuaMNGlHMr6aRIvIHhI8eqAbKQbyV1r4vFaR8
tqFnIGafbGdsmzwFB8cfp1QuQcqAP+A6y/rl2L9U3el/GnpzGLh5QQZ8Pv4fi2te
JqUz38LIPvWxDd3sArjPWz92TSGAGVD9g8SnFetrFSjsAikBjMcI0osFbqa/CUj+
ZA07NtMWx0IcU+Y9vZqfnqGUMWpfUEE1eJCQ5x5g6T03SZqKmMjXBpO6jzZGxJxJ
u6XNkS4W3E+hfDkn3XBZ/BxW1U0ifxFphTTs0A3kKPq57jZljUYjoUtrXjjXMYWA
IW8KRfOlPKemO3EudEmCI8RnK2ymGAzQjJtClWy+gOPIrgj0Ow7pp4R53RxYR67d
skixrKxdTmULk7Knjy24n+8U6brg/eJwUSrIgvRhBpz0hMqpYV2NJTNwZv1lmvgk
T8iqsk95xVlIjOpN10EShpH51EkMJcZaLG1z+OWxRGwrY0meUYzJVFHTwxm6uAJ7
pEYhFFMUf64BKxSFQahLIZsXTvVO7ZOk1vA5IZ/+JgLE7rsml+R1CVllZwKBWLDA
8tq5tSglmzH+UoByAN/C815ebCwpwQT2U1hfY7AMxg1udM3d8eYDPpr3k5UZDHtZ
v7+HbSK5JH4HN+X+BkZYOba5db5YakXp1UAZl6dvVlcvj7cuahl4pLPZckQrrcr2
Pv/m9hTzCkFjkmDMssGu9IyWjzPu7pjhod3NGO6IzrVvqs9pQNKucWQQp2e2w3N5
qGUdL/TPyyN7KCXJ3r7QBhxWhErKU5gyGWR6VIDJwBOEV3jlC0FTksky6eKG6X9a
jBU6Ui9+sIc6LEz4bDndM82aw1bECnwDeSXY1OCUiLFaVt4+0uWMjeBdcngSGpsL
G67+XlxGdtKc+ptGyne6UVdHvbRJqwMI0dYGXUeGdbXW0jKqLUn+VUZouCISMnRP
ypJ6Kswq2+ndgzqwki0pI9Jsc5Hl/blmIqp+11mpXxqF+539Vwjzhq29YOcWpGuJ
CxYgFoe9vq+Ld2SvJgrjYAjwIcl9WO3O7afmULk0m9CKvoS5ImUTWED9mgNlcsPC
V5kDmRMQCESpWBP0pyRpMxTE2ogopdnbsSJJYO5dmj8fd2fDh7lwrq4t/q7VbpZp
2YmyBCD65K1nD4pbMFC4SaWazRE5QUvVpZhQO9PTVWak3GeXhAQQ6VzVa9lZH7xO
9tu/NYIZUc0vvxkF11CT3QzTs7vo37MR0V4Y4VDSiyf3q9PHiSEDmJp5RrGKteHs
qDy82Lc4zr4TSbPdLZt0op9L9N1mzRbBKeCAL3RQhK4egq+pg8z5APaIu6+4Qvwh
id/WKR9rc4DPpAAYACX25EDzcl+V+ZPVTQSiV5VuycjNacXvxgYcoKaSig7m/YCg
6Q7x+vA/CdIfh3Ika1fbOR63e90smWPoA3lt8tm4X+MdHg6/wgR662Q9aY4W0wPT
k/XMlMpUdP9rdru7tLvxCJhbDhOPMPMHVOtzYFQvAxOamVWZCDxNdrqrVngsUeXI
q2sLwatq294LoSPTF2QklaLnEt4493aKt0tHsQ5jyzXSCpXut5Y62Hx4qkETCNO/
zekfaZV+Se9GBCpbQ4zc0QhWb+mKF8N8UUsndxrNHkoRzNRNjpkNxIPV1/TVLRm+
Rdp9uZPO9HvZE5l9Rz+G+2F576AUjxh3rWtP44QU2CYPor8zG0gFTtBc3pxZjWUa
kRnr1PIafIGmzgDjF9CnJNfLbqxQJTHvsDoMqYi3IOY6odfXS0iQ8LI9Rhh8FGwN
IQkzGtVrvt6NF+Ax1LQB1yAY+LYhhNvJEoC9tL8m5Pa86/9FLntGXN6OrDHhmCYl
VUwQSCmdZ1kavN0VUBwWSmbcrVmK0e4dWhrdqTqfc7W/CEfKOmsBcU4eYijdE8Gz
X4co1gFfOZHVgaHL1SygTyjyke9g3g8H61lsSejzzf67zEpas/AmiEqTIWzpnyYm
JkM7dNSJV71dFnRyhHN8dYrQbH5VcJi7DH0Kn9pwvIm6P/ZFvZoho0+VRC52EUju
fMtZQIBeFop2xRy0mmoDNvFJelShl1pIkPTjFz2ApYdAUvgQa6Dq1OgJTbTJolr9
fJpFuo/mD9v/f7mtGnJaXJdfeLyeVYs3kjPsjN+D+M5iDIQEIY6GYTtRggw3B99P
4/tb3jv9kTBUoFnwp9WG6ZXMIBvlIXc8obj/hOjq+1tYd803qJb8CMy+NX2YTn1m
8ALo3yJ6Wy5jg/usEG6GtDWb1yfLUeBDMWcEJGDCYVPgm7A3OhIudR6fTFdSc6kH
84xAcDNx5iv29C0CG+8srBQ5VZedgvbmu1+hoBqZkz8/jMsb9VbzCxp3cEvMU7tA
Xz7LnXib8beaaCaMnolgHrzupv8zoa+Ti+KaqM3Yf6Zt63liqjbwnsBfdpuGotI0
Bhi0JeXO16ED+Na2zhb02JYsm2phOjRyjEjWubUa1TBsoI2NymPhbHkVosa5+pHE
4QMbk4krBYaZhxseM2ekXfcrzBq4ZbSejC7JXUJHrjDf5r5Y3u1MN+qhxyWez1un
Hkr49mH+AXHes2GaPERKZM3RaNFpaxpC+41ULh6LUCSfM0JltS98aTJTVzIwDplS
ckAK8LZel+OlslqD9+4+CKedtP8DNZAPTbjJ5+q/8ecXO/+W/A0KfQbGiMlzarvU
wnRkBkefbmBjW+pfqJwkSq3G2hFj1LSbkD+gYUDfIFdvKZf8Z8BCrmpKhtq7eEIU
QUHzpyeaBJc+D9hJ0rCxzs5o22RyowNgJDBSlUVxcNTQvZMIRM1M8800jnUqKerl
rWw4FuDl6uDoKKQ2eQMtZVIqw2RTzsa2kXg7MmOxN6jILiO5mEvqyHIBCzot3aFU
+0b9p/a+6YlCoIH+qNC/tGbeNpdHfsA5A/Ji02yPLfHpTShF3SMpNW9ZZLKKcHh3
4JW7LDEIacbVjQ61EngHmCwJTe+mVeV3OJF+ciBeRvySIaYHEHw8rMmJFZJOpEb+
kEZCX0wnQWgfi7LW/cvQE8gMiWQUmjZZnTXM07zsiqudPoGVRghSiesFcbPkiwxN
Mp6aVk2KXjSz/5hSWgUTchtkdbeoD4R2ipx9cPsLRljtHMIbC0vDqJ9BGKFAjqxT
VAk0LXDvc/UBiHT8fbCrHKL/cHVX19Sh0t5tmaRVYpSXDyKUNcceBWL3ISElgxtu
CmWqoeNX5PJi2LT9CmAfgKxwYw+iYXmbHQOQxbqVWNyuy0auQhf0ZQV8vWmK+kt1
NeqHCiKvygti4+IotYgd/mazYVZvh8iDxiYsThyPYa+uF2ozz/+ER5nCX5ZWjYDE
Ey48tRFm1Mef+KnRLMMZmpC4P/AdNYdO+QGQh2oxaAeYb6uCzKBO/MLIypfriYkG
gQ8/s/gxRfoVCyufLa3rQSyZ4TViBlnRZ+8EF/sU2aGrwf1O5V7htJSi5FqRmBTN
/U1Au65H7IQNyNCkDXxomt6EwSl6ZHcUGVGiU9uCQLJJ64ONR1Rk4zTqKP6pvLuK
5Nph8vXrx2L2gUhSbLO4THc46pZAYKt8GUtrdyBizCymyOrLS7D3AM3/jGFq+lQP
KHO2UST+CVUSrN9L5hW+DY65ndByXClh7+wkmlqywNY1n+OPMqq+iEyuFML08VcW
RAfGmsgEoaBW6FiFRIqcoOZAKfJF6er2MC6afGJSN7Oc+uGvlbJUD40mHlnHT7sC
vS6BVTB/0aXvcC6FnMCNuNEmJtrCo1WmkdiXURYnv5f2lX+KdYrUNB6/odJPNk3A
xak0+hV2ht9KRxckm0PqpR0/EKM1RrRLKbxKdY4TJnIQepGVrF7GCvX1OkRTiigG
FlqwhuGvpclCKgPCKwTElCfqtxFNadlgyLsXRsZUYMzhBtZzchKvoHT+qlB82nXR
koAXnmiH4R1MCNQIOFYQyxvWi8eGO0QKmZPErXMcEHf1KvB4ulq/G9aQKhfWvg4f
6uotNyuWkx3fcwulRQ1gWfWK2wLAlGSz9jsM3QcBrw3I2c7rOLhco8G8Iom1F2kc
FGa165mkvPmM9ytpWN44Hv3L+gTjEeKE1lzYvN3Oj6WwsxUhbXzhoAH9/woiORxo
ko7OkumzMkizS1sqR3AKdZ2cCDqVEKHPqDBOdBCR0TgO9Odp9WyDEfcl0IoBziws
MIorkMh70f095lxBXtryOVq+yvBKMxmrvoD4RYTCNAtS16UDcct1tOh0bD6AYFcS
HJXAoCA+LWNokMA0x7FswtGAyTX5MGEkG+RqwProdeuLN8g7MF9cnal3DgzUubHZ
3sel2GWX69K3ksAVyQSHSwhnUbOgAo+BKRqVRdiv5huIopMewjNBY0Je/kTzbWNy
2rs0+TDSiPgwmeYK2xCzL5P5Fpbn6EELKRM+vBaXd/Js4AdNf0CMfOCTjK+zK0x+
vWcIuPxXPaNOImaFGMmGmLVTWrDBvooltD0rmKLzPOBlI0ATMsw2MiNAQpPjL1Z4
9x6FEBxJKkEBeF0rI9/U0vAMFNp5S4yI4RRE/fLutmmumfwMTL7432Z3Aw4Yzezh
b0FGV0N9Y+m8B0TnwZTvQbxVSepbnA2l80KToVoqeRQ1yW89ctVABZlJliLzxGx3
8ghSU+hLgZ0ouKj0bHcPuMBzyVWB8Ikj/Xtti1i4ssjtUga/kwDEcFGwa9Bu3JKY
jXi3dOuJkW4HpMXjRwuCuHpOpVV64HFkz5+dsV5uhDahtQo/7kQolb/SD2xk1mVd
qJ5Ec6DjWwjZMl6SAD+pJNWzMKClL2r+dSrCQPfC7EGfdj2uJuIawV8OXKyONC8c
N9zVgB3Q/MtCv1JhS10OvkeIeL7HA6tuabtl3TofPICZu8iSBwP0I6RI02WbaSY0
l4/VlUIEETopxqFRCmXs5ivbBYc+9TmCaqbrO3O7/ywIDcWsbe8FyEPg9iUlv+x0
mczrvGtu9Qj0EqiM/50E15fCoiPLEhY3FHdRD7EIjmExeZqJqaDKt/2n6s63o4Hx
wdIBBN1TC20jZDDrC/CX3Ua47bg4GaGJlpggTigdDNgiBVTDQTLGWhcGIqC7YasY
V9XI7GTQasqYR126QHyH22wFeUuuBgXXxbHiLQDZTNMgNeatw4Ru2XOYokHjKVJ6
Qk5kU3P2bgKrxJjQEF8b8KSh3anOJla/g9iQwPrA93mpgKYU/JcqpwJda2/WFqlI
Hag7bf8E4YJm5ddvUGBpv2BUp525RNeQqdsZB2z9133f25HpUDrTcZKEXk64xa2n
5I47wiWGcijFiOffA/+SSunJk46lgbLhjUPGtR6kI0MHE3m/0V2pII7OrLaUSJqh
xUZf7Vx8KKZerk6HbvPS4e0RMsq7GJsxfsHeSwsPebX8Bw4EGkeGCi3FoNCh6A58
2fXqUsCTHxGo83vOZGwYn4BGWkgjXwwjH85Lu6TIznnVR31NVzMLKImUTdqR5LUs
RW8z/A7yIsQBzTP+eSN6LgPIdwEz1shMMH6NvB2UXtNMYqKTY9n6zGC3qjttGvbO
LRXtPd0o5oNbfxenVtqqioYjNNtcPC1Doa4/tCreM1Fm2cyKBP9NNzLBNpVtk1hH
O16veOED90oDW13VHSwM0Nj8gyrZMkeZu6OcJExr6Pm0awJu5T6nhqJR8Ld5bbAW
U4l4WbLIfa9JBxMMF5CWjQ/8BvONmSs4iA/JILlYf1NFrqi8E5rj16bFm8AQapqa
GzgmTUv50fMUVn1LbcpfskGe6il/zajx9V3tpwqvBiTmZQrxEn7loAMHGauoDSPw
8bUwT1rHo3keXqVVM91Nqz055SE8hi6Eb/9QwOCudgOqQksAvtdr0sm/fctBHOpP
cUiZTz5LQW1y1PYsDNcgpLVXUqhR3dua6xHY+5DLnC9leWnF6uWdvDeB8gR9TcZu
xX3HVVf1Dqcy8gIYKXolunnV91Q30yDpkAFv8ysPGSKIJwIuFiLHI4yaxfnNJt6K
wzJdo+Ias+C+l6EKhEQJ60sOJC3KLNWl4ILVjy8Ai9BGi1N/AC/c/gZNPZtf147C
CYz2NeZZ4QIXIf6spACeh23LuL8HoZd8xA3CsCqwCQucPYIKOxFRj7vVWXHE+OZB
Zyc1h5rjNwOAjcPPsh1SmAbco4rP+h27hgaWEtZv59FCmJn8+BY4IX5e6MCgk89M
/hr2zaHMzJXYpNDvYLbn4JlOkGVpXJBIEsX2dn6wBWqXVpMu++5EtgcoECY4nLxc
jAUdtise2jFQ7qIJMxjAbxHCshsybD95WRXvYb6yWCFobuQFwPihW7Z2/EizP2aR
mOKaPqABX+ZMRepFDitimZ04aYIjtWaGyk7tQfuwgO9Hq3vO3YB8KBRQGYhXtUZn
MfinRcCiDtr9XcrusqYB84IXLJzKEAXoml4NmYDnAGrnrl9z/57ySzX8XFYSko6Q
62UP/1YKJ9+ovd88lfm5LmeA1Z5p6c7VvJjmn0bzqjYp+xINK9PZAUXazvxZSBD6
0aqowRH+tyV9OcYs2tevt0JUsc300Ip/6P1XsYy70SYZ1I4GNep/KGK9CfJ9lSiO
KuwJ9y0K5f0klopOdxBce098JXovgzix+zplAWYCWYeYbuYK+r8y7uP8qVb4zBbz
gLqRNA3jYmzeLjSw260+z8wyqcf82DrN115b9lg8z5gK+rM37v7ymyMcxO5s9se6
4i1O2A9+QrkL3WyErlYkygDxmCt8cW6SmPbsrvRqLeBsbFqZmKmZ6t1ei4Lj9KSY
9ZE52WbrHXALfLawBuTgKzCwRZDupcZhis+Dss7cX8Fp4mzVMQYRoqf6Kyyq67Hz
BmX7sxB+I4OVuCELWiXQ1d2QXE7kSwTVsO4mDqz8bJEIe8Ng57Lm4fjergdfgxRn
c+ahKMwyEU0/7EqmfJhZaCLMCQfTWwBtbyMbQO+AWsZhQNY1RibOV0iUdVgVkbuT
3pR++i1Hfl5q0HMfkmIZ+P6c9ahdxukFuLevQfLWmIdR2b3kf6uHHE4ocqRbIC4U
NbOrIBYyG0F1A8fpLWPykLvjHSTxPsLj9XxfEC4/U8H9YddB65TgDavRLrMxVPrI
Mx6XE8p1un1w0YjtZBjzEFQc5sJ6mZELpmqrkSOTTTGgAzHXz3or2ca3qE/vNtLp
aZLn+KbGFNYXB0eOnoJJxiYcbzrW/fBNkUjbNCMdubr5KzjlCR9E9t2jO48pEvPr
7xX2Da2G2pR+MCmW5JUQzENCQ/tHFetSBT3OfZkBkVBeN8G9fOisaf32e/A4daxd
k+l08Nk8bdrLdqMHKiks+FNtTK0XklbXW7QZo1y4w1Tc3M0ExOZiVXu9xllQ1oXQ
yU939V2UWQcQK0mr8NOc+G83uMhJWmu+Rb9YMRpaGNIRwkz5YdwqtwAo8Lnf4AAj
iydNdICrJm4auqRvUkJhiyn0zFvu3kuzZ39iJg0+wc/ca+abugKhHQBLmjeQwnEc
g3yP/ayzjw4YK+/YMUZXm3RfFW3umQwWsAnxZHK9wj1HOD9t2sD72jjITRg9WERe
82G68vE+K+eMAdk4VEz2Iqm4f1EFQOW2bMpXK8Tq6+FGNOkKFEStq/u1fkIRTQhe
8hSkv9YTlTPzUuXT5+MSUczS+IbtQVhCAQL6PTFZGNgxD3tQGWMwPAC34jme9YYM
KLDs2pJhGiTkYrqmVAISRHWzCid6SQMcwnCzUAYOqpn/kow+9xRJqLYFlazhm3mP
JfkDSSxrynr779D42Mjx08gWGwVplFIB/L85qX0p+DSd8HOhu+iAb/y0UzYDakhu
pNNCjlM0c5h35AHcNZiR+CRtpeABSwh2tkDFWmMAB/qVcvrWHf2FneFtzQdlmYbD
SKeOvLc5MDZBVxvgAE0sL0fPADAjBXHPtJ1oNE8xYpO2C8aC8xSbaXp9ECYX1gT/
JmM54duRJE4Txp+lr6jAyBYRBfSavtgOqnUd0skyf3GTL/YR6ytXzIzVzdHofH9w
fOLJn4AXFBBwia8uKSEju8tPdOMZlHcHMvB8AhU2TR01Qjl0fFvLKGMqLg2h84qc
sb21hbXif9xcoABI+ySIyH8WuRevxPHGl7NE4FsAIeNtEmuoMGYHsnZJt1zWryod
2lxfheuaWbKz5LUeEfaudDp7kROJ3H6ciLzisuzeAvf8Uo/QprxUh2eAYPHo0xXK
3q1Q8LMDjDCmbWRDMmILg6n9kYjoN2hsesBXMKl86mIvOXG0goGi3PU4A914poG2
3NmMgiIwVhwS3H5/DLO5klS7oSXnvf5EQ89IR5KqonFi5yGmbQmxiIgbLqkh5J8b
p0dmHJL2Y5kJzdVBmYfCUAgDJ3jVvoHvjl1NAlTgz/BBK8qH/3XY2l1MjPlsd7f4
rMMg9tnNYoOY2VU82Ei74wxeNMaiixn38oUeMOpQR8coATRZ2FWrtVHiMofkkIKp
HDEtLqhZhehlvKNC4SAwGD0p0lV1XkC7krcEDy70DYahgPo3yMETbWCxftDI0BFw
CG3py4WtlVcMmXwmTom5a/nBPI0teGTwvzeGte2qSULCFhN2Hr9/YJhOSy+Z9waH
b2H9bm9IdUdWTS3xHROk58zBAHZ0JBLWLJj+8uTkXZs7m3uiXUtbMgGjXiVZAx8i
pouKyf+V3zlJuaE4l6RN5qwLfWkfgzFBXg5vVZ7ye0LvPmOhZ7qLig05QWZ5StYu
fuPsDgIqHT7ZRMr0fzpDoIdXYSnLCBCRAdXglQ2SJn7Mwlfl53OdpZwI9iff2Ao1
qRz7YTpB5MVgFGOp1lsI/4BJ5xsisCtuD5ig4s8nGwJTaQE8OAq5zgPv6KxtFQOL
Nd+h5fdGoCTDWkhFKzX06QBh1jif+crjjqGn33y3zoO4Ho87Unj7QbRRgRWLXAmD
//pragma protect end_data_block
//pragma protect digest_block
5EDe9JjZHX/yULUiOyeR0m1Rg7g=
//pragma protect end_digest_block
//pragma protect end_protected

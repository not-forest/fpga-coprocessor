// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
zOdlHaqXCfsFQpgA0wSz02QN4J08AOhC43UNZzkK5PnUTLEJyzkXnK5aet9cBGTq
IItiP3sm0A4b/o7/KfJFx94axst37clU3IiK1egGBTsF4QnBYU2ezmlIDIHeT8sP
aRkef9Tu4mvbkgeVpsJEsNIeow/okXn7wCy1h34o8gM=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 15456 )
`pragma protect data_block
cejxEznDRGK3p7EDAClDhYoJ9FRNiUdi7V/LJQ+372Fze8PqWF1udioL+m5kssLL
CRzVhIz3S5lHWNJPMk+SsjdTvzrZntm4mPdGXsRFAL6m6MYCQZ7dL9Lp23GqUslQ
sNUVOMkd0uQ5lfWplgRXd43RgAIo+ftLLbShzW0Iwd8vxjUMpoKhP1MMQVbnt7J1
Siede8flzJORQQSOOtEwu1/jrD+mID8OZUupz8RJdz8RHiPcqHJumbPf/wXKRZwg
fPJi6JEfJkp3D748/oCpf363V7SlZXpAQULD1gitNyVNQdy6hRp9v58+f+vHhD+s
3Dj/5JJ1gzJbucgIm32eCdUxqFgn+m4s9iEB0y7GcKI333J7AxpDPSuIzer3uqK7
PVw/3GqSftWLlQ/S0uiF2QktvuV7RtXiat+CuSqHXDpLfVNXz3uW/O8eTiCFjSZy
nKphiRm4F0+3EkQNguMTrnRFzOaaVqybJdyfbt0bgqx4w/KagIWJ98JVPeZ6j8dC
hbPyuaQ+5T8Ybyt+LRW14X6n3Pt4dymzya4/QP5QctRpjAnOcAkuJr7d6H+1Pph9
Gs4zFK+oPPjENjTA94R0DVI4qX8Yxd1dYHYBbFlIS3NIk/JlL5sCnXzfuREV9c95
QuKepr093U2ywCMYgl0FBmaAF+0QJ7uWTyTcXZqeOz4BOga3arrwu9xVjmmqUw6V
erC9trb2ClRa21f/ziFw3rGWPWtNoPDk5B+1bg2vO16+2v65UC2KFKYcDkxYe+JG
i7z2Qamk40zJjTRPRPnrBE/fB85/GpehLF3tRp5BWPCDex9qIXU3JKNsoXmUYe0A
LQl5edOU5NCmdZJdWP/BRbMy6LVwaF4dywSrDbwEUA6Ub0h3rLeAsd1+OFo2DGW6
JJPnV9e4NJBrS5dnVNIr8JF+uflDUiMpJQFe1QieHCDV5+TQUn+muyNEnIjog8OR
EfnZokAja29WeYbV29DUdThryPpeiZLe/hI5HqxtdcCxmv+G1b06MGPdtTfH5swp
/Zbr4Hg9bdw/AJZ/BBRvt9qb3mh/Cg4LIvJf/4Qf2xZ/+nUPabaaAa9OjbSf/5Xf
kLSotDEpfTV6mhZMVojsOasO97H2R5L2Zv/yovJJXa7oqa6HdMhMNG2PSjfvArcb
os94EKCSdRNZWOAjrmn283w5xW3C4c9OT9d48j9moSDNZUt2EZEk4l4rlISEcYeb
mFNKT0sqZvrcvLbEOvwvnjLnDVoc+oHIW4lN4qL60xdIttvPXmTHtOQtZl1/PKZX
f0TiZlDpwn/EkumUvgFFqNVrn4gdmsEnVzD+U78xhVhikmcaIYQaPXKWUHkU2wmq
SST1hWK9HYyetrkghzUzgg9gn7U8xByj6zkgu5TB2BXzOaih1/ccaZko0IpuTB12
vbp4zU9K2DU/QNcTtsBoxYOZk8O/EIEVImChEbuEvMKa2XDvV/Q0W6wIElV4xmn2
WXVPNGS1y2+Kmy0BNRJ3bHNtKgd1Iag4+O06jO6CHdNabPA1dF9EprilK2+f52GH
EsXmf3iFuJdrxugp7KYxzIuR9M1JZWjpJhZbntSZBZWQZ9gOUVfpnVNtSyWn7Q8A
CIwLg/Xk1Y/jMwSUyAPuGh3ko6r7Q16lkdjP6Pob7zV2zf9XPuNu4R17ZLB33tGE
zaM62YKW5vrrdwefDpFstSZESABAtahvlCx4yOeNJFgMmoKUkvUDi51lVKTGlcCR
YKrhPnitfYxK89s9ILj5HcFzhrry1GuljF0zUhW2h/A8libt6bAV9PIzQRYIfR4Z
gT4Fbg4Bq2CcOm3pFtk+lPySrQxyLNc06qOWphI9qVOPqrOuNIRoA79syNBMQlDJ
D5UiNg+/K+iBb+a8A6gndiRw5VuyAT2udio0big1oTnIgdLBZVWYmO2I/kxDQqmv
5yaELotZj7S61DRWek6er4Lev9vQ6lSJIcHzDnjzYUiwmxCze0XiFL7fRmo1l8KH
L3vkJUJnQOSOy1F/yYX+RPh/0a+aHJPjAa7leit45obTdw4f9Avyo/3Vlc2x6XDQ
S2hdezzKLI1a71y8anbfES0biaZZRcsfILe02b7y8wYrm0dPeJCglEjyPl2rT/B7
QFBXXW5z91kJc9JHdx2ecQBBCGdBiDMOVMp/pH14XPv4gdKQcqnElkI/fsu0WdWx
3W5LPRR+BJPLwBYOjNTlHbn4R9IkHPvGZAUHcneC+4nrfO5iF6aUzGClNlDO6SYG
k9kfq32jzS+fh//ButTvtYSgXPTq2A6udvkaIlwvraxwXKnDjf7wb3Mgrs8PSgMe
QN980F2g9RqSqojnyv7zCPhGQ0iMXKtzjp/V4ut0r82WbMGCX9yOeC6G1tPEu6jY
1AUpAN9TlZrbCbIzYjN9so5qEEJQpOSV83VcAwrJd+uc7y0tKCMGKZtct5cPyYAM
yh97U+BhnJMRyuNNrk3GDjvwz0thjVlFR8QLgRPwiyFQDVzfGI296oGBWtxVpSPH
BNli7oKsjDcfSMwY7v9qmFMhdZ3PbTo1K/7454C1P/rv/8aJMR+/ngDtNS3LxIuS
4XRMCvrr28ZVxhntt7qGdUElasgB/q/lB2MxyK/pfEJ6RbWAizkA+Lr7bbE8USCn
Hgaey1YIRlaTxezUpns2uIekf6rIxs/EA8HPntwYyKk/YPFQvuCtP53MjBjQsyN7
X5VT3EEfUPktBMWZQSJEVpmoYOSbKu6IuWbBGaoJUshXpTdHKx1gtH9JycxO/r9R
KALGBeiN2XTuR/fqIBsVONfD3n6TN7oUBjNpwS5DyBV1EG09+EZdp8OEgyrA2FRB
nh2FJpdsKT1h4z6RzoKtd2edV3p+p24T4BVSOxyEIRhjLF0rm+yFqavm/8wClMTS
wiqwCPH70D3EsVOVQh3aLp7ljQlQK15FcuVmqLwnfjCthpyHw5NmprZMwHjncIB1
LV135LKPkyErX0eNOMOYu1uUYOi/Idiz44Mz+PtFNusxC5mO9+YznbEPGe5PinCE
m5tZcRnaRP1oL3EUAnK92mW/QmFzPxrD+JS6K+Mlktc/P+kYCwvxH4h0ZzcjXBfp
e9PDPck4sUOCMOOKQauZBBvfi/rVdLRTw8tEhxp6Z80CDwCJrkiOWQ4SxKGPLyr4
kGfrS/fpAasgNaV1pg0YHayUawQUwpsv+MMjKP30/lxCQPEqQWo3LJ7dNLxZXGhD
N2+PMTm27FXQm6Ab+mmpTuzP3uhQELMDDhmnY19tkpTUYQrzRxpD3Fk3GLCiD5tb
47et2pArz9Iy5xcokKrPGHhCe1uM/MZANntpf3/nhTAds5jVDq9XTIhU07ANLJTi
9y+I9Hj6+Qm/cerq2giNGw703MhFBRss/dNlkNcHYYHprnMauQvYXNwxWu2Mz6Po
C7yP0sVXzxdV7p1WGivrRyeXMILJAkCoYf71ZXEV8rq4tovmnvaECeQQXnjDA1gS
UBmjRjtEuIuc8VvdrfCcV1fG619RdKFWih5gEE6gYJWc2npoBXUv928Mkl3cbFeI
gaWUoshHQHJSozSqfFg4h48MK1a9WSwg/kNLvKbXDyfaaDCfnAjDZvMkIlidX4zE
uyR3YsO2BzAKMs8OfaP6fcc/3z6n0g72VDS8DsORWLLWWO/G5kG6N//OFscvANfb
MakylwvcnDrmmyjKsL7T5kHOJNDaJ43f9+qfy/0uqnUr6q61OAIhWKqrHMtNjQRB
yf93GT8Q/N/nWpv0sAIqxYa8cL+9xlSPOz6b9GrBRpF27ZXIvW70EL1DfruWJQ7u
e3trOWHRAw9WQuVNEqnlmlAzzM7IaZk93JOR4/OGNeLUl5pCyiHfAlDsu6trS+Kw
f0JF81pm9KRBeplol4DDTR9YLFEY2XvciO//RCpXVYIwy3zbuYb1U1y4ws6lby1Y
ikKUNKQ8ej0LMLapBgHY9kwl1rY8+72uwqLACOWmcrRULTNM9tw8SRT1jJzTiU2u
ffhubXR56h//kRrqrHG9XlQEBatTIsK0+ZytaXnxZSkJJzaNrR+OK7y4/8slGxUX
xZPJoWr75KgfhVQ6LWL8PDAHZZKoCNdv0np6OFvamg+98VkTzIA5sBEAzhJF0KdC
SaghmSNjyf3mYEFcFa287omJtPo28wxQygJv1jmxf3/mhq2Q51TiyAa0kRQ+OIDt
aw9u8HG+EkPbFBcY97H+2HrNPDnjJQlKtp6OpGErOKvSWqQlqYkdLGaepFwtZbQ7
k/4/Cq36fi0Nuh0CUvvRhuNzXX582okk5UO6t/1J1MED6j9wpTsVPsTan7Rhjw65
Z+LRqEW6Hzet7n8/RtbTEFOWSeNL7isD+fajhe2NBFy4nEjnHozQzuVHueK5obfL
ppTyUfGTiIQ1c/5udHuxBdhv5hFq6Vtca7hc/HKozmX466DNdS2m9baqGraXHmef
1zegnoIKMwKN52T4A+iUT9w1X9zI4p90F1HUkX2uxS+wXtRjnI/2dPV68+g6/saM
xJB/jhtG3TtYqQCFa1WBfiA5E2Vx34iuqRQHbloLOmfNRHknU+DmgNCLeaUiAPo5
TXI7Kz3N4lL3YWdG0ndEzjoR2huHNVAD/dE/ucy69tI8cHiisvnzfi4b9+BW+nhx
0HaEqCQI0Pk4CxvNUqzDxtI3pqjATfsIqTrD9oDtHFfm3yimnXMLtCUpuwBr1i3Y
xZRCZTDqldZSNySKMIoqgeOil0X6RhXtWzQSLkXZDfzC1ol09F7EHISv6pmIlvPw
3oWkxZDIZl0Ln2yjh500jQqaysvv77mUlVzfEkn9uDo/91kqM9TfayToQ4c1cBSz
XoTO5OSLquXWh0JBMvZ3A9WUzzVfDioJWK/1S12BD6rbRyyIHs/2VdHxYE/FiudX
tsrLRpiAKp08vPiFmxyjrqi7vtOJ2zPkREVzL3nNfP3yHCQR0C5NGlEFPDoR1egy
7xf7F+7t32dgq41TnabGF7FInYxPhjXX+7jX4BzoRieGTaiS+0ufI6FTC4yIskNi
EiTHXwHV9M1x65pqGFFCWNC/HN/ri+SJrgImWGgVSkvZwCS/pGZIyYr6DhVkPzDF
yiQs7t+caepbQ0mJMb4CI/5VzGdt4MMy6Y50fAAhIfGnlUuW9jzErRkzIDEM3how
2DRyj8OKcZ7vAOwd2myoyoEuQXPPDKCG4wUVBrrYuJxmIF5wN5QTlLKMtouhWbnJ
1K3rY+F+DzeMgCrea8ItJtEQbQj0sRK15c1n4Jij+kS2k7v2tOl1QEJr4Tc6a8Ts
cIY78UoZo3MmFJG1UOj45itVrVDZRKNQDYUMf5psPJsao0JNCfds5dzglI4vIpto
I+AJO9s+9DyKOyzHd3/x4cKGtjC5dfqEjCrIrn7YqwTgMKnkjlxse5itL1kSAVVv
7h5Czl4yfY0jIGj5VSllgihcFWuca9RucFs4UAgbhtjAgoymBoDoxlO1uGywi3nL
Bqhz9sjqQfHaBJXhGO9EwxXwKI6mOafgbnWNQKLARfGI/wneSyE133qSJTEUnA8U
g9S9mKbaYVLBGU5cpi06WnD/itCCQ1NT3DyrctRq0IxU8EMaRcPbkDioEryuDwh+
iPCls9W5B6yY1X/TlO1XBYNqGp8Bw7PeqpSKy24OYxiFN9wcCcfiINlu5OePDTjd
anE7BKN3LtsFxie4tbFAv6Iy03awFDaL8wQwLC5a21x0rKMT1tz373UNLepDDIK7
wRHLWRVH1eChmbvSx9QiFB90RcqAhMKQzsagplSJr2eDaDkHH0IOruLiV+jpRkLc
gA9jZvFipLkzEyNrXQWaD+k5RYaXbL3g6p74nmhlQVf5J4Zl4SMr61LXmv171iQU
Bjy1PSVvo86hTYqHsm3FZAKvgDSGFNwELaSiE/JPZxKvWpk9HGbo71k317tMD9Vi
5AAzz62X3rKuHoGGMgff1Ep/cbBRvL8a7VaqR+u//u03/S+oYFKPLYi0g/aTajLk
XxclVCKyLytH7b+8ZFrBpVTYCGokRD3EyDjEjDmIHKzerx+PKiU3JX4CGS5o7zYR
vUMqBxyu90X4TlkwQ1mri7eodhVdVWVJqoCKx4nuWIIdux3VMjZWB3zRSd+H21aL
RThfRvUfYAeOwPV3pviPcwRM8iwq5lk9tE/DhaU3l4ywsje0tai3Mr2aK8zU4HPI
Rd6UyEXgRzyEB9VLjrr8sdqmd2x8fQA+lSTa/RG2movbRmUXJcdaRvFrqVP9K5U6
NFhlSYCFNl7u2/uyYHGQLXzktvlmSIaPUPivMc84JHbAYo7hxPOZx6qaNekX4xEU
Gt2EAbmX4H6bLeMxsAqa8UARDhkte8J4obmh2Qr8rX20f2+gTTVeDrbURdW9KHr4
MZ54lY3TsZzFgPCmxe0pHIHvVOSU72HlQRZg7P9daKs5I51qFyMVUZCqdCPSsAay
xVb0m5V7hlZOSv2cdxQDurcA/ccvMgOhfDvnZ2nFB1LSNv9q5d0mJjUzajflbGyB
yedU7lSYUrFXBtri8x/nrWT49wzzjrY6tw2OXSNJZxH0UtHPUpLaoBkWf+4lZ/47
JxXD58tuAVFYtuHfG4UiEPfniH8K2fTEmSHXdOBj15yZOs49qeZSEq8HyAvPKt6R
EaFlSuQqL6W41qXxzCntfPsbKQ1U29OZIU4WpkXwQpfRJKgqf5GRSBq7FXwhUTFp
D7Bp/RM01nRXeMsk+bKIfg+vgJL/utrJs/4DYxYUr1OsF3oQQYFpydZIGEIJIU3G
G4T8++x1jeQ2QFsWknQinyAt7uUhD0Bnl8my1EI0ucoOiB7RvuF3iesIRCtUQoYQ
nJZzsbx11lAg37+sWeAkgQnXPhPkE0pmurZpWUimfuhVKyhWMub0mYZBQAKQO2hC
95wOoM5ZlHFYylBohGVc0hthdZBhTe004lCysmT8658d7FdXimJDiIwymbTv4SGg
8YovuxKnYCmUkNjDnT/GeUnTng4VCHDVSXucuOl1wK5vgSyCUXFcwcGE7smz+eH1
E0CSnNM+1ATyC/TcfDijnXEUQmzCsOvst+OEpVYJm1j1EgLdE+BimnszZaSfxyrU
m1do6sbT5EqHzN/eFkQQnKRP1u1CX5QMX/5ZsasbZICKCOQxhe/azVSlbkvlbe2H
fL6jX7ns70Qg7xKUNOH+3GZRWm34nN89Q54sWIv4mPJuKZzMekq0l/jgeFjlacBS
iWO6OhGlXBLNuNE9iI3KLHyHLzqgnLxWxJ289mgkEDC5UlsMHlcMxgSYAyHXdDwT
kZA/nX/Pqwbd8Yu19ob/kcH3uhqZvYMH6IqagEYaQZuv8nm0BMAAsT/VoP1f1v7M
NN7joscAAMtnyNN44jE879YmZTRBG/53emCA8zwPl3q6qnajMwDD27Zgk4hjWoDr
4reZvQhMhlJTYfaIut4IJC+kn9RyiiJGQhkLOLATzHy3i5Ole7Pu2u2pUd7iKyDS
J3nqrWb2pVv8rYky+apcfLUrpMJC704/LFyKb33gclPp+vjIKW6U6zi/iXQhT0gd
iv0CsCZVxmi+bl/o52dccGN5dNs8VM9alg86Op0om786kkRJfbNPCMxYtH/KHz92
ruiA3F3nSn/MNCh2+nr4cnHOSdIWmUDsYXh0O08JdyjqP5C8m5ozTeoXmZl8jQGS
xi003JYmFtWW9zicl5JqXbBncQ9vrPbEGHxbsNN8Sg6p0aRn3S0uARBHrDl+Uz9K
54T0xUAoFFm68ZiG7qm/XpzD2vkkhvZ+crCyWgOvEXk2G5YDVlycyecRYJ+wBFwq
gRUb/3s9FX7FsbtEE9eNApTi962z9H3BU2B8O141Y1KrtlFYFd9D6P7OeFPiRENq
v1SSfObSqabcfLjihCucYCfYvUwPPWnzZIYhV1vcjpwdLu7CGoTh/O2eIzP76xep
G/JxQYZaBmHR6l0WMN0cHSmfyympJg80qocZjuNB22qaTSEUjp0wpH5NXpDVI7O/
DlVUxZUlJ2xQ2VubSnaIp6+BFDCPH2Vx+haJ39nRLot+Xyxsc2Nk9JZ0HjtjMptF
yMzgeMlrkh3UYEnhZlnH1etmMN0taU1vQgSQmU0it2RI+t4euN4Ut18K8NoarlcD
nzrp5XFi2f2ls8a46g0aCIpKYeuc/DeaOW6IbJJxdv3npqeska1+8y2QK5+8bvTJ
iThi3Sjiff7pi0doU+tGvHy0LZw8HiYzIprufY2NrV+4hu4vpL0TzaWuYRbmoI8a
/dJjXKLFh0r5guISAkcxUIYZK+m5ZOWpV/dGVEPGOhqu35bX7AureX724fkPmXJi
PeN8THbaESpatNjYLlZDV0hul9pbR90vsqzM/KWWFvURyZ44Y7g3dMF4ypKCwqvT
JTjaPwPxKG5vFPnLg6m0Nz2hSuSQLu6Ei5hibQLQHLtgWVRtAqGdLdf9mKu+ePvB
K95gjfkUajslEw8y+YCkL2aOv+Y2+lngQNTK23oVCvMM9zLL73r/QNORNhLzJG8p
e4OMNDaXvVltTQaUn0i1wrdPMd5YV3MQzEz5ftpS0PLZUd4tsuMA4QSxRObypwxe
276guw88NJKjpq6bpY2Z/FgYG/7MrDTujz1UpHO8x4ByzmMLiVYFFPOosUNttE0U
Tn4U5gt2+pGaCSr4cBQDPxq+V2aeRHdqoSAv+nYbJLY8Rwu9J77JlxLTh4G75kfY
brdz0dOwQV9PO42B4PDsIQtxiw+BXQ4N62kmeLNe2EAWmx5MeeLwcjNqOXRzpk0F
YsMG9oZP6eBDZgNy1QN/RkyAJl2U5ddEzsZvuvlpG1iE+lhx4uW3ByWj124AjVMp
0kbAfNCpSj8gvOPnPpnTJhv5W0UpoeLOkIEByrQWpp8JGXnBYDvr/nwSgJwBpvb8
+nWm2830zTUs+qA8cCIg5CPzFEa8a9Zy9Oee9UGzIODTn0VlQZH8omxucaUJEPOD
p2lGUqxtQkOAXiB79uLLmOSB4Zf/PjayLqIoXZEdX55su8ncf2gnJwZIIqmH6LKy
1wjCim8GTdYLcdAQdp/ueMICfg38x7S47kvOIskd9XNUGh6DR7IuC6tbO++QRABp
WdelpiRmW7zLe7CWga1022C1V+2zQw/5PO/tF242oRO/Oyv3P+240hAr9cNRREq5
R0WGPMZW2wr9Ncb0w7jkpuC0crS2WGsDyF0+QGTl1Xw0ZZ7oaBFwp+bmvtezq58T
BhwfWoPaGS3WcyAluVNJaQpQKoHRX6kUDdJJXdimFkcudTCSkr+Ykkf5yAD/Ifew
eToNDl1oCNikG7OEnRznHUZ4xwyXBXzNQg6232G503bp51WzyKMvobySIVT7Ogt+
5Y6RcFymHA+okvFKAftMYj2M+ewZk15RCX2fdh0r9Ognyg+fHC3ewhGyJHcFoDdg
V328OXQfo81guh3+rgrx9kviDTW5eiMfUsCF40pnHPLX+3qIQLQfP2t9AMBpOU+Q
8Q9by5YrDoGBWR5KQPcoyceXPX1mHEjAStGxZb8YSgz7tCtSTTjxQUoDcrFm8KVx
MLDORDnWHlYJ+VehcNmFBmKVYLH9CQszEKPqef2Trc82E1eNEsA/NVMGZoTEAMA6
bpXGKtSmBOVRWtijCAVZ+Y12XuFVl2O2xOG3BxnnQFj8EVoFFTC8H2jXWB6Lqu/E
bpPxcWMCncSaUi+v5nz/aH5n8+Bd5CfIl52CHhjttS2TTfKw/337OG+yL7iU9Rn/
0ZbOGfd5UGhRfVlbydKNUM94VqG0nhBVkvG0CFz5iy4gmfTgKS1lmn1QO2eCAbX0
+wIguZJqlp12aA+EgT6b3O/ypOA/vNRCxdUUJbwKb7JPSFxLD6sWrnizzLz3UWJ5
zaZJ5JouqXf73HJec2m6p0Nzw3qP59574QYIt/HiQS1k35ZaGyKrgh4mX3uQg8Gt
JyYwQslL5g2ACN1X7Q7jy5bxPSzvZg37fQmQyjhHWcpGAN3JvikF1eSzXCxUiFZ/
V/om83asdL3rWe6M7/WERPny0Kqj8AqSyZSvw0BaisQsNGv9F13hkDcKcz72KYKd
nIir+YPfn9kch9iP2sRSn1ji40FyB46/l9iukiGudL9K+CKTkMsH+PkM7VL6vjDK
FpRCfFz8h4/6hZRtuXkDIRmV0k/gpLCJcdEReEgQBr6CsuNlx1GjVdzT/6+jEzxk
mYiWfq21+BR63MvPA4CaPtIlr+8GsRikb4+oEeg+kfbdq4k4FsNlJHnOAEZh0GEN
GDqXQXFmyodZHYWMyXo5yVJ9SJBfZosMH6pzIxt6QrppaC9vXMMOrD26wlaHtArV
dhWm3pOAyB4R/LrkICeAsZLN6ZO49xwsm7EfPEYYG5HCGYbMbMkf1Cbtn1tAecyw
6QdR8CHep5A9yQ4rSfkP//YilzYLVfIW90f1isDVWq04HtsRkr2Q/Yq7KB7QSWXT
+fxEBYCSbNsZWa32u36zy1X4C2UXe25UAIrUvBVtz3gpFzq+pPp9jJb/0CP0Nt8H
+GxWuYpqnL9EHg4gC5iZl9MGyFQGUFFbrWBXXXqrZxugmOxEoHDbzLnKYLKBq68b
tObQfdqFZiuij16B+7H5pPUbIvrePJXfLIKx+ObdDwVx3TvvIX+MaZVB6I25r3Yw
e4KXmY2tRWOJDo1d//TOL8CcmzTHzjuplwz0BHnE6w0eII/hU3w7IaFeAlm8xsBH
OUiGFNT4+1qLeXqcHtGTqvi4xvfF99eqJDgsNY7ELo1PhXWeDR/d0qUzSJ+93nXb
ZFsmoqlbLalPi54J5feu6YEv9aCtz5CMouqE+vLPbr5x7awxhDVM7Lagwlt5vAID
pFzAU/m78E3UFegAXcnpz7XKATBim/M/7kAUoR0Qj4e0eJJUmB+SkAbMp06uOyR3
v5tfd6whPUjvU14tD+T2fby7UU4kljIVPCs+KqD6y4DKtDRoYqH1wC425Wwp1RBh
NaCs8Z4q5p+T28AKs2EoFI33wS7mC2FYV8+yy7SuFpwSTVgYW+p6fSqHCtSEiW6Q
t/jhh+r1SgWrESE9ow0Uvhz97WTV+rcNnqpCCmjuO5OPtq6kgbkqeFciX0QHXch6
clYhNH04Qbn7JNCkxD1gZoXrZJcsGanRY75z+CoDPlqEGV0aZ0Jmahlm1y/OqvkX
PEx9eNhJDvsQ+4jjvzXWUwH+C2Yub+eTmKB8Uw1oKcVXih+v6AeRAxc45eAH8B/Q
ZnWgIvTQXBNK92UqK03xIHCj/9uV1rOay9eHjpsxXH11D1cfkuvicif1L+dMIrjH
7QnbjO2SV7YpZ08PcZe5UrXYT1+dK9xMIzAz2LBud5Fw0hvc1VGBWsjT2JMvJNoe
4bhmhlM+LrTYnU9ijU30yviKQI1j5XQpXRn/Xr2GrMLn4gPFHLNfOkCYVN4CvoZD
hyRgRKrrCfd2f7snL5no5zV1oUcMGuyEleGsYB6yM9HEzCanl+6cXS9GmAa4axjM
2Jh/Z6GO6hM4hfQ69LJuivAyOF4EGEgZaNSA5HZ+9+Zqa/+SFt2lvAr3xYJEtJkQ
R9fKMvAp24BvGnS/VX78S3Nq5xq5u1qrrjf4j4Q3w/RqIf6phpY9J3XjNhYbbD99
pn0pJNLV2nCNvg/9mw6Smh41siPpru0M5Wb0/yW+v5g338q/+XBXZsz6JqpW6nK/
2K8Vq3/531LPsjeRs5ePVVG+bdV/vIZKTsnhM4+QSFdmKXWEvRDlvt5eFdFe/UKR
Ru7dpVgoS0UKNc/XLGKo/tM2zJb3/5/dqFqdtCM6a4pDnO8O9WUVrR6u0wp1/eqB
yZhyMMJ+mmuWRt1tVsoJ+Et+EnhehMsZneOWOz57NLowkvaEwTab5RcKdiE44oHf
qR4fFInI6UC17CenbhtgVPJxxiDR+C3ZK6LBvD6tsgQ3VEMi41S5uS9iKLCVes7W
6qu5zcRlc3SIzecqTLBC1QVVznRfrCOhNEMVzRM8vARGN6zRasB9k9VfJCnGup1o
bvjaB8W4HQeOgSyIziIx1gZ6i5/Oj+0IC3FPIx7OUY0+tW9jGdOSe9dwlcBTf/WV
eJnUIIK9HRudFRdB3afKWi1dR5CSv7+Cax/ATHJFnnB3HNEQowOUQdfr25WkoWEF
OvTskpkU7TvFaFz+tJGXE4IKW5u2YUJAksLOU2w+ezLt5uuBNXaKyoGWqDaIvyR5
Pna7vB3OhVsD7rQ+lkuN1VYVFBNkvR6FmpRlBEYewEh3sfeOEBvOTZ2m6x5oDvAP
lzAEojLCh442Hp2oMPoa/0Yte3aka5Reer+IOSgpSjAcoK2EDS+JuRthuvtHls9d
8SB1L2vMzx5pntPIm+dcyItMtSIV59TslLt7Jlguk6PKvoOSHgEMZpWd2JemE3NH
3IBB6MatPwpk2pAJF6ndgcg33R8CDu8XzcEYo4amLgN8AUFBEpa0b9jl0Y3rn3wM
kkdvtVertHiMhkKuvIYzhaHAxeLpVWGAmvAfLwwNrO0cTmYLakDvr478D7lAny4c
Zb3HS4g5RXHR5exh5gnU2PlFVwh0b5SEVsMMDiMjEluBH7DrhHLNBdH0VPR3RvVd
ih2H00oQd1uld2ZbBfPvadWknl8yL8RS1qHZa7n9axT16z4oGVEfAJBsZhP1ptQR
YZySB88TIT4gMA784NEX0ee0uoCVGpEGpnKO1Ad4Xm7BxkryYHRUEpp9L3wxb89e
OVd8fovAErofXHrmYeUrvwEk7eGR2Q8amgCXtDfRENsIVdJlO1MsIypAPJaqUO3M
0MOSR7X8c+oITvJxyYvtTndLbh/6mMQW000HrfJSA3AdDLg7zIIrid7XQWB3iu36
PiVOr/ySHvDOrVU4cAKxmGFfqwGwGN/XYyU0sGoyywCGSnpgHpceN0A0VCjD2YHL
EXbDQN0nwfswKYTyoDcjFGDGuADeBEZgMM9KKxVwn8lQpEIESiozy5Mbwmh4SWto
0RSdRnT3eIQNuB46J+GrxmJ+uWwG3RK69M+0k1onp5pf2moqhtJq0ZgublPtS4Yp
DdBzhrP53Pv+KkvxUve2KuOQCVqMZzAnu/qe9w1F+3KaAxMZo0wQws8C1tv1tWGa
qCy563iwM+OVm7VpMWVoq2rDeFix6V/n+BudpsA/3Aimiu3jlw6q2UjXUpatCsdE
9KHpyfKkdK8k5OHcWXc621+Iq6jK30bg25Z7hRoJsFFqPM3I0J9WVQ0Fn5uM4axg
lEK4dZq0oe33zTotqu/IDsmAoFo5iV2G8Vg6SZyZ5cfgJxP4I+lyIuHxC+bUwcSc
79GJ7MhDHz8uBmBec4jtq9Ir6Bp0VrL3pONiHRMSHiI0aToGQmJlLn978b6vkCgg
3yGoBVXR0JGvPE5NyFs6m5EURzdTmR3gzd6v3JXCgJXI/Sm8y1somTJXrifi1kFL
k0qjhADA5VBsQssn4/lBNbTsBIR3+6o0YikJyE2JrYwHdB9A30J/augCnr5FDs2b
1Uz6Y+EujV+wgVZVtdKSL3MkW6KwDQWAw1acLKBKTdwBx3Diind4tsyp/6/jJjWH
M9eHPDfFnd5WyAiHQwOq7EGJtFm4fImNvPUiBpWjJSoEDAftYnTRwLk5scCEWNNe
hAPnNK/KogYIgOm8az8hLPQ21MonWPccugibJRDddSzfxbuz9bUaQO0CPOk4+Q3K
IEyhZZhc+QEngtkDYzoqxUaWLnLDyghzsFfEMb7umzFX95cGV4wgD/mNOWefP7gM
EICEzdVJfNPnGrI+VdOJa+ajHhwwGcDo5w9jGJeFNe/UR3W6gAzppEwdYslU0B/t
fmasEuPzMwDzbSiL4ncAJP9Ig/qck4n3DRM+aFoLRcC+1rHw5xjLvAWM+oU3C6ZJ
JekXT86ALY++wglAIX+U+oqgOuYHZv19larxMKolJKSU21ODRjcw5SDvU0xxAIYW
NgaqwLwnEnHGIvzwLQPdltIXmPtBnCJTzSgRgOEDN0H8ombsQ+JnFG3i4gIwTV+n
IGwwpOUmW5lYVAZNf8JNW8O8EvEWKv+3gkTYpMsY7zClNs83sJsCYaQvznZ2I4jN
z5E6v7gEvYb0eR3P7ghIduRIuotpIWivuDHIWvlYiKVVlC8oClvwqAWb3NZLYh2A
M5ZVOQQ8cfUEkU0QtGutkbKOr5m819p8dfHvY4hPY4qSsiw5l26QUWqGp0yshl45
3u93+3rPnxbhVBiP1941BSiqMAHDgjLZtBv8oYHtr0yBMITetPCVPQamMUY9znIQ
3whMgfRXGa23pGf3w9C+2NnQrJmJBMC4tuFGik9AetA6Wevc7p7Mj//OaPjff4gm
SAFV+PmsHuYLi+t5QaDVV3SZGnlMy1iYThB4VS7z/16aJpfrunKQ+drUpdE0tm6p
8+zk8Dqvuj21kgLPXe0QJCDeL51z9Gnamigpr87CP4GGZ0Kj+QftsgXjQmN4GFj2
Na5Kws0UzQl3xDHldW7VOeSd+c2X6Dp55XXkdqHLxrp6u90BiNSk3DzEDKBwVeBu
WLZMw1xvx/QYVMnuAwySag7EmiKEfKafu8ben9VykyHALMUmjGEFy7Hhe+4UlH/2
i9h5FvXq4Y+wTug5ZuyayPTjnHuGgFrcR/mNSCABD3XA6D7uu/jSl3fogL2OnHgp
x5LirRAgqFk8i9t8ll2nxvwAW+VnktIWA9Td4NFimVPgxoO3INPKLJCbhMhkRD7b
bkxFHC08FF2e7iVdiIo7dG11jTI2adAPcXGVrxGQoSGBES91o+Pd10/E53oHCANQ
LbPDfNEDsjw7TTef3wRlkWJyzTTlLx+fQ/7H6vXxADQ6EBp3mwhEPtvHdtzzF4Pw
rxenxMpytDxFAqmRj9uz6elAMhsYKGO9Oztzj+NRf51A6HgdEdkNui7BYdCX71Gf
z2z7a/siPetVmSYL/GyHB/3acje3MsJZg22D+e4eckCkUqHx5edcfQm2rGVVn/dz
G/+05eJTOQxjKTA44rLXOFAzqjed0aUNwizUfhqd4kdJ6gu0DtnVLzvT+Gz0P2OK
zZwuVNXnH9CX+7wCPpW+FKV25FEUEggccJjLPtrJ+MF8xN7rpUa4d1b0UsqsKAMk
Q9gu9JD7OitNocbFKw0B+NsOWRiO91PRtsDH0slh7Ms55+cysyyiyrkJgkGd6vTg
VweYMXIeddAjQQf6PzHNUyUE+x8O9vtl5PmhSREN3p8Eql7ejrE/InFL3JZBq/Zv
LwjkN0TyrhocsNDd9Zz95KEssOYl7oE1B1I249g1ImIu1RHAFHTGSU7awRq9/Q9Y
gJewiIKLay+8tYx+pHRnLS9oR5xPWET9LFaMjbI4hNIW08h28XMznRWq5ZUagnPh
idU4R5hGUo50cJvYYuviFhpq7KnePKEVGJZmkVIvHQ1cMUsdLWS+GlXxfcJ5dUD0
jYRMjWzotsLYvKEHmMOX8aSlzYWC7UPJ8He3Oq9NXCOFM5StXSDLGNOyySIE3Ukr
73bYHBMDR6GYphSvgbqgJFGpz9OIjbCs399o5oNxaa/IfIxOPcmOdEkvIhB7iR+K
X8I45uokcjOA39k8FOFd3o9DjB5bFsI8gzr3vRWqsURNbjgFMdmOXPJ/rCJO+dmS
pMsXrfY9aG4KhFO4EcZwfNSNCgvreUZ2gxL09yA+kWmWLxlDKLLCYQgjL+ZP/Fi2
zS7JZCVvN4B979H5JbDfyMf8TqwcRAuiqGO5z64SpAIVascrabSvkesjS+TWesaV
68hfLruOdZ2qo6sRWH7eIYufvWMXQ36F8x5SX3idHKMPQa9HyhTJJiSdJu8mmHCd
cMN8YKozAAz/DcseSSo2pc+63HvDQSWz1/86Ms8IWYPjLgG7tLmBrzp6dqmTAa4o
Nm2stbsHCnoFECQefIbMEaIK60jCSc6XxOR4FRVyAFy/7z7x86s25a2gKvDMHO4K
qqcdNqZCRDUtt4Vrd6mipfp14EaWQMUJicRjOaCH1ktrb8AAOykQPkQdaOVfcJvr
1VK727m5P5V5aOCSJhZUC2yhCWseaT3YMkANdvE59erczCHOQa+wJ1pzAweXQrNo
4+IjiTHtlsWliM/Hn0ox0Hbw2EV70QZ19FIM0uYBAWRtOLPlldi6LnxzmZISd+Q6
VS8Tb5cloZ2aPGxT1ON0+XVxSfc0CS9XGDQMSo0WhhFXpAf8ox1KRB6trjZlgp5n
VMhb8gvyOCovTfTSYom2guH2zOBAjtu+yHrCW1wxDAeGl6N9NvUenejQNvkqqaB5
+CautPxmiOj5umU4sFz5TQHC6zMgP+Am78/orZXpbU/Kn3/bKcVPP2Oe5xvIQ6FG
WC0yYrd9zcTQIki8/myFrb/KIiJwT9RR89Z5x+amEfCFsU/QapJ3705Cs0WzdY7w
5P87x2rqN59Y+TRWa+5JrXgihZDixrmxSGa7WOGfeYyWcWD5q8ObC7kb0p/Fy/jl
TSmZMWnR0LcaO/h/84JRX535od3BiqP4ADRYYiRyRvXMRCSK0JNq6F5UxMUXfreH
gH5ay4FUQP62IoBuqeZz3Jy9lTpm6lVtaqJsJmUCMgNd7tiMGE/ZoTrXaO2/qA5M
685uRB2r08LeRzXHJlpr6AlvNed8eUrwUxmAplSpGaj6D0dViLsNok0jzOecbq28
HsjAd2Ay+2Tpt7VjApdiSomTOcBWLfAiNQPYxzQvb/J2HlkmFe/aTK2ZTly3gCsI
hkjvJW6n7f1oR90DczXT0YZFBHgxrcSsyCVdN6I0ibSCk2R3ykbR1Gt3mfVe7Qq4
OTr8x8H1UHi0dcHwl5skmD9qcVQOU3RN0R40kCHY/22pkxV1WGywAyuaKLYvO6ye
43hbW5ZxNPvgfrYpjFfK9RCQ718JwzKUz4DEP6uz8BdqBcJPB7RtTQWfsmmeoZJt
1OyjC2u3aTYtQrd/vxZ96zK9j8IL2EdL5B0Tj3iS9l2TsMNsWlmSrOMKLbVX5yqM
Vsssi4sWD3uCOLSI/aDFHIKbaEHy/oPScUDo9ID6sT52k8sWRXIcM+xYMJegKkin
BpB6//WqCblPtMJm0QNuDEzcCFOY+UdAonhgHtwndIL1CM+5XP0oRNFEtFcPcVnr
/JJMIdN8r70FrWUASRmRn+b3UAY3BAHeoqw7Ua1jq764gn7AsGWpklJekaLqxL5e
yrLQoMB6zLdhfQwKxHfQses9zcJMUOGgo+k1IeqG4ddIKDHTkKFNk+UVol6XF0gq
+12qHZX/xpnmKggeT9rn83OpRtc8hLxmI2Msmg5lrlESf2g6YRIty0gGroX6sd0/
xGVCt9JpIe+qhE/sosizSsEEJC/aTcJaXEONvAWBUe2+li6lD5NXbsDOm5uC/PEt
6kvcSuM8H3owvrXOapGzJFOs01kO9TnyQ74+0itFm2wYV8UP9rFSdWKX+NlNZqNE
p0POBeKVOSjrNBjwrGfE92vBdA+Dw8v9ZlPoC5NGOOeK+KgPhv2IqHQGolVqEA3i
3yWE1U0x/p1l91JYLz2+w42up7e0h3igpFgkm2kqz6zpfdp8XdlQao40gouwFzsg
NgfAUDfr6kNIuAJ+SmzUzerwKq5ppSopheilizq4jEspFu3MxXgyQrsJlWTvuKif
DOEb9CPfBlwVtX4/6Y8tj+HdtC2b2G1TcZNb2pVTG/ZmPgOBLVwig6IKTlX4UXRb
gBiQ/VckQLO2eM3yTAVusUgLpCMD/w08z8aNdrVCPglH9zXibHNl/DFcp/4SXKon
sq0WMvaiFiQoOV9kcryXTqt//madDmDOBHS2iQafUSoLNhCOwePx2HnnahpSmG91
gPX3bOiT7kJi5QP0F8SxufilRZ64Trn3W2HCVFRl/UvBKEAfxdTlowwR96AR6ank
fX765x6wlmb8GFbHZjjk2Wp5TUpFZQ+KTxBe3DzXgDLF61SUQEyZtsUj3hDAlXh/
0ZyCa8dL1W3ztTHVkqDP8Zcntz45kUjZgjhxZkJfyM87UmtbNcTGl/N5YQ+/7Y/e
4RoQC9j1aYFMLNVVu2+28TTfyXbW3swk2BBFW2TjI8uvRuGtbv42KlUoIopgFytH
wTi8zpf21G7UA/pJihme8JNRbn/SWtkx5E6U9XvRRlfzzFEEhpKJ27/NmTE80P7s
U2fUk3gysV6hyXnzJkb6M5hAkY/gbgzriQiKE0spbIYJPr08JSWGHw94DzbGApsm
GvWcLWTvs+y3ibyLRnETIxhXvrQwsI6xarZ8swx8RZNFcjNIKzOXmtr4vscFDKmk
av9MyowkLkQf8lLgIdgenn/oDeBgVB0c0FMEp2rWVN2sbJiFRdqYKmewxk1V8vNK
HiGTxSLji5/XzJpRYONaJegL7GoE8zwJhbnxwYx2BXtl9ZzJiygOQDHXwN9iYaIa
n7OX3C37sjtuin04c5DvwxJ4QotNWlVJ/XMl3HVWphegRLwK8e1veNWemTAPKMV2
wkpcSw+2mDm5UDyBiRiSMUGfz/4aZpzBEirRqqP5XE8bXOagruD+qGQwNSDi7yDw
8PqThOVT8kefUTJYgQIXGeeo2DTNm24Wga0dLsbGWBgTnx9iuVKbHpMjUmW0uSuj
91hYK54rrQEfsZRFRsMzUHybPBBuBlimz869tKQOjbVsBXYfEmF+W4vYXbWnMDK9
b8F0nUBtRgxoYcpFNshO93/S3PqoYUTOHNuAh5emy97ONxZgqH+PlqKNwk7CjGxs
JhvM8PQas4vj1GxRqKAK3r4TQjhqUebX+feT2OZv1Y0RsLkrbRwc2DqUevHkk+sE
OS52douLAym35FQjo3NlNeQiIHFTnMG/h88Ufp1QcZCi4oInu83ROIdPxKU7r4mb
hV7UMzIbCcjXXY7d38ow+z7SwQBVGn9d8RygQtBa402htvB2/mOfmLZ2Ixuz3KJ/
kW+Nnq0/yUcNsqUuL5lCSQPhU/lALI+ywOHKhanZn/GgcWpOVnc3ntYLaanr4VJH
qNBS0l1T85sjYAngHFvBIV/+bWW4aLxvum0pEHt46BXEyRNU9So1ikYGUaE+8bE6
NtMYUrdchP0gCCHQrtRi3tbmUJDlzEx9XGYMfUNRe2lTqMFMyiwAs1j8VyEdW3ba
PVUYweLyLgyRZXBKqgIiZy1npAWX3MXzFeignD+4h5uOz92IuK8tDDVXw4oG7LAm
dm+Tb8DAKj35Q4q19hOrd1qi51UFH/Iei6UwXjc1UmOTgQ/V8D0yKhZN/GPuVmhY
J6yEBdAt/AsbFVAGbYUEiweTUuTNqbJHP2MBNdQHEKQdOspUm0pQc/Ye45C4bonz
gXYn39RvL7uOAni6Hal8GAHI0vKuFOTjkk4RrkTLyBkXgvNAxdfkJn+IDl/mGyFl
srNWCMDFt+XxvkSb1xe57zpX+z6jtIYxGed9UGvmjT0yzak3SJkHuadOE/0HLmN/
Q2g/sZSam7qxOGdZAfZs75ztDYQ1SCwpupde+84561x6kW+qirLTO08E5sXRfqTp
HodQyHH9nJQ19EKLn6yRIkSfRYdMok2JuPzrdf+YYQPycxjHoKTb4VqHgWz9vXH2
GcS3dMgvHK8VyqXHR52vaen79vlnnr/TzFqytpZQWgxbZVjMijcAvUD0frubGD4/
HenAkX2agEOvqa8ojfJRbx0iIcg+SpgHb3lIl3+wu/7cE3NIPTpuJvRhfRzum/Ew
R5Yq03caAe5amvtYMJVSq52cHSohP58NX1oe3vJhl9fqUmFtiFXLbpcWA50DWbux
Yg06Sbkh5zIOj+YZq7FOnf8sY8N7oNejJOXFPEZBfNTDaFzIaQolJlW8qygR3ar0
ccoZTRZ+DnowCb9yQX4pGid4+kK/fsHS1Q2TCI03zltUv7y89u+PGhBE7q36pyjR
oL33UkuD5bWW1cZGGoGuFSp7XCl1C+v211hh3UOxk0SxbzDeN6H+tZ2/RZ24Muv6
YJYKIHSXxoDYDkJYnQFJNSsLNBzrSwzbIc7uPIwSwvEasfS+zObIfH/EQMD3BvtY
whRn/yJMuARknFMzxJwq7cW8XprkVlPlZTpNIe/2Xc9UktW/11WxUXwRlt7aIpP8
7rxyYE6ABh21yAF4+pxBW7cSl3k9/JNizXEgj7QPI4mfRoErPhnbsNA0+RdHGh2M
Ie33dDuEYg++I03OEO3iqxZCH889z6qrhONWdKc9LZGqsBFUU0xQRtkS+E+jDlRn
9kdiwhKkZWmick5Oo68gvkYQMbQKiFuBltMA0c0LdjwHApXw5arFaBCbDxMZ5sTc
3ws4tWcGQ/jF+datPR2vItX9uzeMpI6NlFe52sdKRnIYVPppjAfsFwk3YNkWL0zO
MvYYy+JrvVBM3S0Oz7CRrh39Pg/jDnYjUYQy8JzPccmymc+YbN6wSfAWH/gSbekM
UTf3yB7ttYI1CcoliCFqHIumpWeVY96e3DQQkcjpIU1k6xHKQV5UP8MCve/DvCFP
a8nV7ywQbPt1j5FqZKEOVH1Ad9Zi6eGOMUcItaHbLW78zSusZcaYor+KwiYISlnM
xlD14iF+t8tDSvll3HyhOkH7vG4r2bvrlI9g0MQdB3Qa8+qPc18f8s3KTHnDDC5t
TrbTvdHKT8tAJiGx+oboqn38GwP4/pgv/iFjvu6P0xeBVLsvr23152VOerHBGjWB
dt9zNfUItbIvjRg/g7L2+FN63r4d8oT/AZSRFLwBT6RAPbLUZwPRCPK247Oca2eb
tPYwc+7PBoGpNtIOb7+DI6n7WSk/8CiWKPG+32fh3d9i530SayC48LEtNbmsrplQ

`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
UfAomkwJ2cY4zl6i/trA6GZiSpxcBBOAtzXxsNcXJMiX6st9co/bB02AywfLd44JIYLbF7n2N+Mg
sttGpB4Kr8qA6uJK/hi7636LLzltArX9YprJfyx/GHGV77+eY5JOx9dobPqeUE0APShi3G9LwHEj
44fAO3YoP44nuxNDtZQ15VP6W2exo/W00vx9ejusOOGfYSgZ/FL1wZm6DE1q5cgNIaTsCeRsdfZe
18tQONyp8x3klus/77BfopCpZ6StRRkUcqz7gn3fZIPnRgd8NsxKVxk4VnF0zuNyUpaQMPY1Vkuv
AHx5dGL0y2wvu1PgJJT/mRtHk0edmuxfw0gCUA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 11616)
Wsm9yFBdfWfw1CRUuLoVvnbtJejTLqHNZCYkZSlZN673FlnGC77NBEt1mmpJh9bdwwMjl6eoyE+a
oiUdKcRyJB6qumsFdrP47LkZgMUlBaNJt9RS7JbRP0u2ofbAkpwAMF6SLBRsHe103qFM6Fx5pS55
bBI0ZfyZCMhoID8g4SgZKVErNy3GchQk9N3ONkCtA89JKb3OLgo5DxAWSGG6sbyPX5F5CA2iLien
Rgt+1izofKtB0L5LEtMaDSSfQzx9QxyBPY6aYwRJGQi5AVGEvgdhWhitYX9MnU/9Dy1/XI8gtC9x
LFv7Ex2PvEISK2YtL1tzGG+TJ1vJnk1Ou/bnc8JClOFf4AOhArOXX4bq2SJbXu62pYglelCrn56+
OeypWAZT+Hsz+RbgkNU1Uw78x2ZDydV3bwqA39naW99Ullk4I4z7fIxsyhy9PH5Crc4WLRuKWVJl
aHbKLyNxjZJrWD41rSInFlt9cyJFomT6UsbR5dYL/S6eVP+bQF9vW5c/PWNXA/vwaW56OEgIMoaP
VvbPrHCW0crG+BmPOD4PMlxq2Da1bAx5WWtvKhL1Ws0RO350jP5izmKsJjbro632eioDUFfbsW/Y
jk1VfetM7zUoI+X/QnugQ2SA2oQ892I+5uWo+bu363EDPHrRWAVeWPxY8lnC9nZp7ajymzFbS0I0
VWulTfVyYZwYyo9S1FPrg4S5qN0rFA3UEvW7kRnqjAsbQYPBUc9nklJDY/mFEIyRohTShDF1q812
RTDUVM41BkBK0cTLfcJmdAVPdFHDBtISuIqb+3V9l4EQdTBNxsTuYY/6SjlM0d0IFWA8zcaNumxK
BMVqCBrlodPPzbdUrtcn8BmZawoH2YIggIVp0Hvqp91Pi8us3Jprwb4Zb9T3Euj3cFp/q2/6cpoT
Vs3IXEnb6q1hL1+jT84nPgGGZyOlbSJSDL6K7+RxXSaL148QNnVe0d540BbZHgFj92/uXa3sIhNo
/KUegGVDZ8LmsKSDa8y+eg2rhdIAWMuQ2sNU5AZ+y7wQL3ULOa3kx2qTqpGHRrLbEJRYJFejd6sJ
hY+u4jTPfnJ72K6/Xa0moIQfMf+tLCxqW4Q/Egb0AgScThQ2zgUetxPzyfoC9o/JagXhshX4klfs
owOlZ0SlATLytrZ70IiQXHOW466XcxIftb1kPYU4J4QNipG7CD8WUvzzf0Ux3xNnDBlIGW/cq38B
hc1foxh1T8evtKfwXhyG/D696iyBjgaSfNVI0u+/+pgIOhDtocC+Kd56X/EG3fF6xC1ELjVN8iJn
GRC0ldwb/QA9ZktWD5bBROroJJ6oFdAYIXIhppz14BF4jNDr4HEuqROpqCAcsqCl+MnD6uIlYwxw
OLlmatnCbb3wfoqWsIkN8FYTxD9mRW0FYUpARneMzw3Njy/xN+7+7Z7ss+biapO8ZFLBeNQsSa6D
VdzqOdt4xf881xkfKHyPCLDWoi1lb89SHzgB41MXroqX9aQaRr9TrlVAm2pcDIA/FZ/ZGAsrcflp
LVDMk9tP/udF1fF7KMmboXmHEGv7kEXUEfAvKiq/naAkUkSM0EjtVv85x2qVu3g42slyLgOAy0Aq
N0nyVP2UeNmvmHInBrnBl6AxTf+TZ9YP+JW563wNRucIr9jNnwvRLGUrF+7FF04u838hokXFZDCa
bF+ntjqjKDbewzCYWCNGaN+9680NdZE70fHWgOvOwrxZMHsdOxvApw6t4odaojyNQ+MGeMg5Da08
7yQ2OvcVx5G/vtBtusWxOyROpQ9+2wqk4PRm0lLlNxyx4H2nhdqHNBsY8xhVgrbwmCfMCD/0a5j4
819YqbwTydbmw8cuQr6wNeN+YLe16Ire++P49Mf6hGuLVhzJas75ZhzDCSzr/N9JuqdBGH66HYWA
dLTpgNJTqqKX9JdUouxVxKG3IS6KJ7W8F8XH95zT1vcKWvm2wf+ITU7NaWjGgVngZPMk5ZIDMRKW
SE3iT2cjUUsM3KLZvu95HQbsXjFMKGI2VOqKzlnr2VaIAfAAPc5HSmaeLGW+QJdVqczd3JaQ3iSR
imq0GmNu6j6jOgsrFzTO75dtVJtCbrtPrjfmbMhbmqZGPQZWzN0V7xTMKmWrBh3RcAYRuQ7bUKBg
GK2CSeSSk03HwiadedVu4rLimqSoNEkSygrhwqH1B+6Nv8KWiY9IJf6a+gvLFBzz+hMOWquVCu1r
jeOV2/MvEC/3bhuAZh2Y5C80AX7aPzw/IcwLNp6k0UaZb0pbmYoPqDlthj8eKyZJIGFOqiLpHasi
ejwBQoflztYFNJM4iNqkarQXPZfgft52779OmGSQ4iWuF2ORn99qTT4hW+iJkVpdPUsDZKTTraAl
Tqt6/7RJcFcnb5RYL1EQQcputeVRIrGZoeprTE9iuU4yW0wUjXEmhSExmQ6+Kt7YqztmOOapmBRY
iPCGCOEesAHjOMl2XW2jYcABZMJZGHfVnEXhUU+XVJH1FBp1Bf1hKstr/p2OCSxYaIZ5negqk4+y
B6e4ZzxSB2jGhTqJjMrl7WDn4XtOoOKc4171vDJo5oShMpBhOY99EmvIt+nLdvPLeAaIbP7OLUWW
oiMC5e1qLtGtMX38BS5H5h67FH0KO1InidDv9UrJ6n82kjqMFL1PWcA+AiNcPT0jZjQCbyWBCAY6
Eq516W6R/xLJFbMNU3HnqKM6xv9B7F7Y+R74FWj6QH2PnrkvAaC443E2YiW25qr6rgOyV1CsUhEv
RlvpLzkMc27uonJ1zz6knTafMRvNup0uEBCmX8G9B4/aTeo9MLDLpgCMcYLm3zwtALbwOMCMWH0o
YMTYBQ+wDP9sanLjmyZRzYCL3k+q/N1nZxVgMNV9uxEQVZSMNRVyzmjJsMaYx+WPpt6MGk0L3fox
hxnOMg/tmaWUwqWX7IKB5QId26zOHA9aBHVrOgXHOECF4w5A+6D0BQghmTbR+CdR2b5t1eTe6yps
OWmbf9i+W16irHjg1/PlBoV0FQ08jocEX9QQS1W/fCKAKSAHaPFapA00V0VM5VwZ9cJmepDIApLF
tUhjLrBX/mx+lC7Xz0CWBLe1BGwqr4D5vXh5rrCOye24QSTozrZCTM22XRjI0kJfqaAXov10s7l9
k3kh8FTJZcIkWk46+ohNZZ0nsGvuonsnaYwCcNiQQc3BhEaZ1Fi/lD1Oky9beV+qUbViv8T2GBK5
6qd39TFXUjfH5j0wgDnunDDFpYVW7C06xjpzIxT2DnF7czCaNA0pqErLTSqj1watwawnauA710rJ
kBpqmqG/U01kggEkf/TbfjJVsKZg88RYA6v0NTuzYqCq6rxEEhPgiDNQyUsHnr5tWgTYbg7hO5nV
9UVd0YvmH4v9pEFn0MagJNFYPErOAQSMk2GnTKn9ekc1VRc32Y0+TgpjfHWMkRkcbXab5rwW+4az
egPm+k80vOFjbbIFm5YSMlvZ9/dzCn2kRmpKgtjuStz4qv+pFwZh+qCKu36/lvG5bPLGO9SuAL+f
NoEmSxxrfysCtihoUAd+W7d0bLT8qvAJcVEWoLV7hgojB6VBy/rkUYFae9VpddNsoYa1EWdUiTZ+
sIJq6XpP2imhpRAFLpCsCsNkJyfvxgi8W2SElAx0GzaSPhKVbOTksZG9orxuipJdA/IRXidR7IR1
vXUoKVliKMTDG8CsVA4XuVf7G3DhC+V/qW67/XOUb4vtZYeSCqdKYekOcM0QKBP48an9Xc5YAsQc
Eg68X4FFmXIFJ2VHK5jptXNovthApjrkKmldY2HypnrJtEBAXxHjhrII3Hy5yOGTiA/lMKmEbUgZ
mnXSByvMyxMPQkYm5BaaYC2+22wiZhP9fvynSrSNdi8HNj6SNxT/n3prTwkX0Dpilx1YG8BD+KY0
JFIKo19gFfl20HLaARCqBfBdu0GvaANPvvvRb0gg7jMb+FbBsCngURb/pGO/iQXpk/SK6w1DZBlP
rldpQD0LZ2QBr/4aV7QkMJK/D8i2a5+Wy+Lkdq8ThhMu6sCZztj38XFdqrfWT+Rc+KwkUlJiqQWH
+Cw7Y3WTQxJxjtR4imo6J5tUkFPxbC3SHXnsUjoTyZg4Ok/8UOm/ic1KPdzMu58l36mlBHRoUfL4
CU2GXxT+epoZ0udhuwXqajRIIkBI61K/Uzkxth3GkIzXiFzMjs2pzUzfg4Tej9ZBRGcWWM1XKn0T
FrgEcR3X64ri84NsQa24aOuoKVMqQqycNUQbO1CP4jeGHtyOu8F8JiPFt36Ea9m+M+mcLTgnQv9z
wcuBtuzaQM46wrm6CVTsTcHbVmtF55Jzrpu18ox0jax+2A9Mq4Ndl1QfGFYXp+7LN3uCf8jB6XGV
EXsCxnaCRjg5989powfCmripmg/cBiqXfDyAYx6yXwMPjRewId9N0T4S0Z1tVNu5cicVOMDqhwKr
KkB8dWVm51G+RaqXnEAob17A8+1B6d3Fk4DsF9BvlEmIZoa+RJDmDcVfHgxt8RghaihImiYfIFqW
AXs05YrodbkvSEp9rg105heUuRZR1reCfqglrY/oR/plp1pvZ8dMFxmHcdEjbpwto58mglKMc5YC
5AX57Aa0794H09RPFa89ALRKVoiS3hYiwzH4gqc2cUjfm0ljnD1ROvu5EdosooOORsqr0HYZLRsf
7mvSO0H1w18NtbQhJ7+tOs6yPtH8axsYjmDzS6JkWVv1LnKcTBOZ/8hlmVkskkxgVCNGsueDo9Ba
ebCRFyNlx2kZqDWnAbGvAYoexpcQwPU/LvOmPkDNF4s4hK/pa8Ed/zjGdzROeJZGMbWgz8zrunNG
TXvPHUs1zCNqMjbZ2J4PBwRwolUYYGbk87VSHscpRBVqoWgiPiPOwGNqhJfRVCMVQDiHVmaj4RVX
o2Q1/bebJBWFiAj/v4aOWkjeRQxx52NEAKoXgAISODaGub/zWrTNAqrzV2pKyzp6O18D/Pyi6NBN
YIra8C8zKjK87RKlaqMTgaIMb5OJ0Sq4n0xv8KGhXRhaOfSW3re4guHFtTH/d63RS1Yrqz+B+OD7
bfZh8KOJ1CaHU32uchLwSG6VFQNGSDFq13xTRUdGZRGAtoUJrGLdplNV4O+YS5YF2r6n1UTPpjF7
hY2wfpqmx9yKeDuDYiZklwIRP5re9WndfKU3r72iOjwqCL+dWnIj+s226raSUh9H8jHjv01fJ2hl
alXEbNl1kAomqjH1dkCwVil0B1budc04mcAqd7xjV5bn+l2lpZ7O5S8yW6aXeWku94ag6W81hs1t
EE/cRMaTsOhFDYkicoWa2lzDtURLuisIDplteDF0c/BBv2hTwQbi7vqM/ZFPDnLxOvoGdZfPiSHY
+W1sxlePlIA67NR88VlC5Z4j3pvsQCstIL0IAJ278aFgsJh1zo9G7FFmn0IONWx1z+8uspn1YaCS
l5TtjfTiWnjQfi1q/gUrTWBoG3duhcfT5rwEjbinW+nf9z2rs4UIOs5iIq51HrBHorGzAnTTvFC6
Y+KErHr5gD3TzdZcDGS6fOTcA+2Jp9IJajR6N/JMk2pyHHq0OdLh83xtAJI8LqEd4jdZ8biwWL2s
baHLm3oEd/R++wt30HtiM4SuUMwrcxRmMH9Vlp7gRwzx+6s+GnAFO4ovEM8M+Q1gFHytNUUZGiuM
32EMvDSp2rq6FdQwDb7MCgb5qR/OQU7HmdyDfuYgOVbyJvQbqh0V/Viqs4X6mcWOz+les+V1gv8D
tl/xAGVNVBpinC8oNxUahG4R8hVSm+XEuII0/lgpeudH/gCpVkQ1RwlS6WJ5lf3WYxhtZN7eMxpS
N9hL4cDwz8YdIEIDHB1iHo1odIqAn4bybRERVo9D9FvvS+EzkBV6YfKmTzAa260JC/uw9LzdTyl9
O+YXdJ38x+4v6JXCU0RsficwtEnY17bh+2z6K1jrd4jdvWdK53LqWsS3OoOzNij6507XJdt4hvkC
tfrQeoRSxp4s+alnRHoN4nsDoQ74GyWDj0X4HBA4rZLXlFg2e9SBGI8OWS0W/pYJ/ItpW8QlQFIY
4aufuxPMH4eUeDZu7QlVyKmECmPjxAUsHfJ8M2Aj6CWaZGHh+6VKNvvUDWsUH5i/1xsdq2XpRqX9
vCpqSBZp0mfUNj/SLy+MLEppB48BIn3IiGNhRg6Er/8BfwdWgKS25a3EX95WRna/qBfClf96khB6
NTFJIEOSf4Ln+x68xzOaai1nCHKAdsMiplDCVyicyvtIJbDYXiM78+K30zj8UVPYZKfnxEplpLoB
UtUTSm4Sd0uEIjJxPkPJOR10IkOpT8A1wri3YsI8Yix40+DaKbloozLj5Kb4OlcBzEQ7IxvxiXwd
P1GYNZ0XjVuifJViHOm+i/PtkXQP2mNmex6Hfd8gd7xkpPuGPXb47IugIVu5hYqXj1BWZU7M05Hz
iiRIsWoomoo0sKhXGETFJHmhafG4wvkzvFHwf5GotbkFJXpcUSGJSp/IuTxqax25bJD2aJxJ7lSX
ImG2+PHFcsYPcHqrvHuy7lNYW/QLnW0L37PZMMuoP9H+bNFBGCRfscs8VfP+Ni31FXa/9jmaDH3D
FjXc5/L9kRKkoGHVmwuPLTDFiWLoc+2xYAJQ1I/YPA7+2oRQvMFVSCR8mNh8KoMHgDMxnqxC1Vg7
QzcVLHV+1Hm3OO+nnVELIWqET7mjLVMu5tTZPKVwpyf5JZwcrCp/mtuK3TmiggBvKDoy7BUKjptq
y/O4k5k6wy4MFW8BdFCcgGu5+AJOtqN8tqNkkgH8LtmXFII7AJxtPdU8hViLkhQmuZnItRw2n4m5
97ciP3qkXGSneaFK1qcO5ommDqroLwwn2CX1pI6AwtQEbtqUPw6vYOf/psz3AZ95rXhVSUVSYRZ2
R0TylXMnFY5jkI14w/FIy0Itl7f0Ij34HGi7qhug9e7JMqxc8AIrhq6IO36UhaHrMpLooB1JuTnq
nAkIQzH5lSwNcRfErH4u4L8+CwG/5fnqkjNV2AWwlXS2p/9i1ROmVskhDqt+louWh3G2O7N6GDnr
IR2oZaWkIqV1nrIoneMgFFp49en1y2vEb5NPnYEaVJvRmWRnKxIOiP9Akmm4bLnLRVpIeMFmNY0J
O7AIvh3dwjTw8dcdk8y/wbP8on//24So1Rwm5gLOCVetzVkoxWQkKdJ3+Pl26RUSC/9dDxcYm3E1
OBGDxrO9QZhOX6FwxnRr3wpMciX3S9WDSjXI1fiSL8zHtWwaGsp9LrT6mhq+t6uyFh70pvWFcjL0
QHd2AWmXRxk3jpEs0miZwP4ealYKWjSLiOBDI/ILgWCwxhXmGNDSTin0pc2AIOmST882DVz1DWpG
BqkE4o2HbBzL+/YWS5JUoK3mU0OLIUN4g7g+9C9d4tRobhkR12BbKQSi2Lnd+Em1NbK5QfU4u8kX
ficvmC9LFzqQrbbqj4RHAQ5jjU4VLKRAIIeStO09fu0PCatqnweWI/91+J1FBFe2sjhVrjInz5nC
r9v8WEfn+LbDL204B0XaIncemxdydf46l57YevVCUUO0sVXDQQWTsVrZH31IiSYRT6j0F5Mxqzg4
9dTcMTfiah+XTsNCgReBNb086ey4r+Ex9i5EoWTtXCHVMO6DAy50KeBODdNQpnAXZjL5QoxwfKeT
ljnEdt8mpvztLNRZg2GZJIjdI+24f2CCtXukFx2NKMq8Hpfrika3ZYFVwT8ezcl9TMut1SLwCqX0
CukYBUaZd833eiZ4aCOuMuIgj5Bwigsu5HGhebDPr6K6jy9ayZJrSPmpIj3pZy0JfW99WME5s3ex
uDPl9sF0nP5pnntuqUd50B0b9bU7GvmqpEI6UgJnkbwgfzon71l6cOnoRXY5eR3DDQuAp6TF7FG/
YBmMs18tqa0wHprzOuxPtyBNYr/VyEN85XPATQNyaLUggIw6IPF/kuqAhfS1bXb6aeP0qY8dae/B
ul6v/ys0CoX1oCXj6fb0uBkbMfjfj0FngCvlqfUx98RCFZ8EnpvTK15bSNuoFrz2PGxuTMcCMS9+
mQlJMsSMo1HJEMuDi/xYf3HvD+ogSqXmPMLHRPlFp6XRySrRbP7CQ9QtgiFfLYijNR2EWNq7b1mL
dgCRdxDKBVBUectSymgBMCD9ehmmI+AvPqVPrQY5E43ExAEtb3SgDsjGg9Lb133G/bb6xW54WBNb
ooe75pwUfPKsv+AhnQdvRNBmzSY4y1aCIou+5q0koIt+IHTjHs2Qnl6UpOqu43voBi2CaEd33AqE
rWRMHmUNWgbmRgCseRiGl57oEm8dobwpkzy35l46lYEkLPax7CALknaK7bZUHMt6njyHcVGa6EeH
IqcpfvpI23ZFm2roO7mXshOOBPlAamVBjgt1yzo8tuhq3JA46nBuIkqqGpFpw18SaV00ZVCiyDMH
Wn8vv0DW5yyGN9qni0OVWOKbYliF4l+g7+z5oXCa2QCkudKhTM0uRleLPyrcM/mG1DGlAq9x2KFG
F9rApnZpIdBnTR+hMQwx1jYYTNWp5oSeoJQk+oJZ0aWujq9W83dJ3f9/cCNYMBxys7kLPy/yl6xc
U2hANt41UfxgsPU6ynJRraRbjcJ1qPTb8Q95ct+PO9wQ0VnKHVbupzT5rA0y5BKEvj9Woj78XIwF
/Tr1X+txVce6yDTy0g5bUFkL10CdWys3lc3VTdSMVKuu0fwdx61etoSGG/1WRHunGVLCFT8G4/uJ
uIMgAOHwJLZ2vU+95GZ1yUKCQUDgeWdX2NxjgWPJALMxqggl61xUWoqLDL42WJZdeLXjkw0hzoiB
1a82ZCEAk/pAyQ1JXWaaPho+uLJDtIaYg9bx+ITIAtTmLxGaXmlCwhjpk1/CaEJ2E/WYygWKYUEJ
BOpwdQ9f9VsZB3A8J6qGmFOHcs62ydglXrHzTlQ18Fm2aeKN3BPz7wuHOqriu8FsywD0BMeBtHi0
dFzhHY3Crfvq7h1jXZSpNeSyqUDf61K0CddIlHejnCuWPsqqBbMQhWyvBjSrlRP3+wSEu5GyEf+O
gOpZXcuWUYuKjrXn2EyEaNOQ52X54Xiobnwv3Bk3O1Gbj8EZITkasanmieDeUYCGkmFJVsLLcnmG
3osXkOxxh60z9psm+BdVJfiu2F5ZuaQu6Nxmdlr5dqqJouuIbt3jll8jkWp30MEArEEmYJW8neZB
YZjOcxXDzaOIZ6QffGfVBwOiNJdnf2vCMf1fKZuZDOquc5iNfkBJRMQuMTaljNhP5gKuutJS18MP
l+TVTaznMW7Ja3ZaiDk/QsO+nWrMJZIWgxuHyE3705/3dExL0pT/5b0UOfdGgYJfcaimk8qUTuxJ
atxuupo9J1jNOtw42gqwhsqE5OTfr+9JH+F9kOxxl4vDQjKvIFmika8QhfpBtAiGdcu7CsTC0m2+
+KCqZwbNQX4/3WzrLLmrDinDbP9EMzaIr2QdJcYcUDjenNVAP+jYObtMOcgE05rSvgKs9upyBqG/
XHRSfjLiZlMiVasfoi/oQM+YJPu1e5vIdTqnPPt4c1cqx1Gla3nq4m+1swMqzx1z3eqHFqijfHs7
wxmmXAm0QZ2scVX10pHWWhA0GISqOLahrSJOyJEV8T26LeI3ATSL2MAkgE7BL9YFY10QstEW1KY6
UcsIHF6vpO8eL2w4Wf5BT5MJcNmtMya4lKvrcIxwh+6aTwuokXFLGJTL1UDIWgu1aqV4tGQnwoN2
HcidWILonmc1bW1oIPQmiOSzZlvdQ0qSpuip2CksdOjHrTOewKiou4ihwVwZK+UuvQwqLV2K9U0v
6Uv/99tt7aKZD9d3+p/km2P/UhnhqXPddk2tKGSZJWT0iROylVj6yIPwUDRFAGUqDi5FdgGi+ptf
dlz2CRVP94YX8K+XqjcApaAwrzXguRJR4aCs5ozPO0DDCoZ3wBL7pkC96mRt0V6isqX8CPAXLdH2
nW216A3UfPzjRb4lPJbdlea2XzK/UG12NigPlINKQmel9+B5tNANLjld93QnFIAY6/LBGE9eEt+k
FwrNfOCriBf2HkqqqA/MKy42V/XGsfm17aT6C6NAa5cbpDnMR2vujzFXqH6XFfeGNp0bMUIT6y7O
5eg1MZ2QCAXkPZhuSyxPHXmqGUCqNj8wqxDIAmw1f7LXTkrYxfmLCFO0wANywyL/SDRQlNIFuwbp
qywMgiHyvZXUVAEi8dNM3tN3bpCiepbhwCTnfIFIstRkTX5APEjJQxpes20FWsI25368y3hDS6q4
HHXkyf0fRFKRNqJT3y1mj19uRuX7NLRITEA25uhpJa0CJi89Fj1iqsJUSvRhllv4rq8zbyYyDekA
03HuV5BRguLdvoIwJmiqANc8GGVn+U53u8qv2MFgMzzNZC+mTNcHN0/nxlvzBTncQduXOIBuG0Mt
XYQVapYgRyD69Ju0lt7PHUxgLSarVUz+CtW34en2zSqWXkxsZdFGJV3lt3feDO2GALv7qe20FQwq
mwwStb3R+dXduOMESvADt41hPYnwnirngnLsdlUjFYhEz4eTiDyp2n+I6uhWBl5CIcvaeCOdukOt
Qm+jizKhXix7YI4dnW4NGlSDPNUfTnDJ7z05O9fUScIuiwuqecnCtoSMrNcyfwkDIeG73qI3sLPE
mu0j0WrPzInSuGC1TcXFrDRa36Q+cVDf5nD4se7GRTjSNPs86sRqlDxNfqFDFTOvB9X56mQzZszy
WjhT+4zbshwywJBkBid/agcqeVlFvD7JKGGcaG8OGiKzhYBI7C05MiQOU1ahznoGnhUDAg1fCn8S
Z8j0reMJ/RbKRFS8X+wZmSSmaJ0it8CuWxpDYKtjd7bC0WZO9cNmuKNtO7xBFcr5duAvJC6vG5WS
dq3YYcTnsb7CJM1iwIr6DiM77h4sR8g/IccF4iltlYid/0vq+Bm6lhgZDRyAE0NU7ESGel9LX3aO
fLtNbWuL7Q+cIxQyr9c9kMhDbbAXNh2XKB2aJfVc8661HmtFHKcdho44XrIG25E4SRm2cCbk27Ji
PLfHOtGXPC0AcKyIAy02TboI9oWT6sYDFH9iU8q6WcAFpkpKrJAWzNHN6yqCf5zkY+vIDcLYmFnl
q2AgXYU9HxnfjoMDqjrmBibSCBoFY3j6rYaPI5TAvkk5DYCwwdraH1sK5dYta3f1+z9PUVaSWB/o
aOklTLEf03OTkRrS49evSvgpO1vur5DghxycloPxiL7xqARQlS5c52t0PfvhzB+P+CUz5XrBrFwt
AIJbUtWTFCX5HUbqsEZph06bcJyD8dRTnA/BFmGQX/PyYR/SRlA8cw6OgjDuMrEK+iM1YR1eeV0w
7me+QFe16ApNB5FA8ZUjzCWqS9LCWG97Cwj2roSN8llfewkieFxT60J9Fx9g5Vbl2ADrgXA+h+Fa
qZuFkm7SSCXCe+jWb+4OBln4t8czptzvYkLZoJrOkeAsnxCOV/rd0HneZpC022nHKgwgdcQFDRcc
AAn+4Cs8pSoXRtpKlLBXZp2ptY3JgX7VMlTj13CwJUD+JWIrAs3ZfY8YUr4UYHfIUu9O1Rcp+C64
d5ZBCFrxsDA5mdR4/fI+GvM5M7S1SigQF/WwSyMcPcHn51QvfxtpgZFPVJEhhrgydsyI5vaD8Aq8
1R7AD0juBmGOB3EdJLXO0FU0yrNj8MKPBSDLB98l7lMHZY6MIc7Se5F7sJa60wpbgfJZlPork6cW
jbffx1yzvxL76/wwZ/7Y3ftaJuvYTsJWUSMCCML6W7ngm0bduEMyd0TWWrxMowrTS5YTje8TmqLH
6FHrwQGZX9G6OPxPI//zz5P/u4DFBOLgaPDhyiKrTi5oqpkChN5WNa04yAyN2GVJdmtCG2JJpn/9
uUFBbOKIEraHb6NBE2SANYTESk9wIzHlkU2WqjGYl+FLjOSsSuOtiw0+tIyLng+HrnK4A9/eDeo/
EgfESHNfsen19OjgNLANINnIqCr1oX2tWdE3VmUrmLn5Vi6am0IadPAtheC71BLxYlJKHuoFFKNd
3d4a119+AGd3fiVEvkjg6MHQXlyk8g7bXXcS0+8ha5aV2vqiGsPZNA4GpnrgSvu2xfLmGHyFdrmi
hzRz2k9apDE+SyKF8vQjdz4rEQjvVxFoTDXZnAdAScj6QMIqN/kaM3nssgsrchLZFtSiX4bvXrVg
MkcnyC6oQHnJBz+Fg0cJsAXNWmjdRV0TDDUOjHvJCyrfpoT3445TrT/ugsb2KKsgdlHg4VSTKRyt
CJMmMRrt1MaJwfgt0eLSq5w5Q1VCIhZIxfogu7wIkDnKHh3MohNhlyWIjoB40rlV+Uv6POQGm88A
/UrcyKS8Vn43TuoTOS5NThUp5iaIjLPaDX0oWgve1oUZ6rDCJCkpD85xPbcmvhCrKdzhzQBqtBm6
uGDk+Gx0YRkxQEDn/ijjpMgsYwMsErbEwZouZi5/ChHMk4l1AWK+1PC/c/Sl1fpeBJu+uFKps7bk
Td9Y4Qnpi0m7sVgBFikDMF4sNtPc+HsMJDbVbPJ0VADtMCtGesSH4us6PHbX5K7A0z4bXsOME0hG
JRPwronRwSv8YHYDYCcAOnx+PzkTk78e7d+HZwK7BUl7fbKICH0QRxOXIauT7zkmLw4PmAKneZBh
JiGjj/8PrEVu4YpIYAdeJUhDmR+EHeI2nqY4hJYXD28JXeXB3hBSpa4brXO2cOSbMvriXEuBVs98
tD9F6EntBhYm9bb7LKcuivod61WW23GjgDmNoV/sNQRYbX8tfxfo1M5ACLCP7R+BeiUQ8qT9kVv9
5v0sSt3LuQqwoPRJiBNOMLLk4jEsXa7ajE3FFM8bIHcopyWK2D26b2GS7zi77ZgyXD3fF4IyXtL8
QuQMI2AuAsjfDpNd65krxx/irVymsAKIajr5q4CmXna5N6uV0bHqUzfVHjCGMaPu6OxCXDmMGdOk
qUX+nIUdF3HcVJ92fkZfa8AfyEOvKSV5PmMcRINXFqT5Sw4R59zjquztk7Y3h9jUlbHbrj7tMSbh
pk7bPvyp/YxTKNH5eIuEsfTT0r7fYdGR6B0Gs4eoWiO+moyhMIKJHEsAPNZtBjYN9UjiDdhabIge
fZ1XQzPpsEDzsH0+GDmhsN5DegdIg+QJVNstovG3Lhndr9bHhuk0Y13v+fYaRHSkjDkjFMTGSYQc
uFkpuZjI0Q4OyC/6s++hwygABNIU2YElCM5YoLOOvh4KvbYDgllDwwaFlYG8X2fzksNTln/nlLwv
fdUvR3t+TYn3aLNtobIOZgsPC6itZ0O1/u+aiY8iqaCq9jp53XQqbwG1ntR6Roh7TaH78b/p4AiW
gdq3cSLEbFNhY6bzU8JV4LZfdpvi+iP8oi0UK5h7LrtBMCqUcbnPWhD9T3OMjkyKTKJxo8i9osgn
C+2yk1SqGI2WFF1zF4VMPpSuIudVk0Cbov+SYg+cylVk6GXkpBtJTJfvHxozSxH/zKWnqAPfpQVQ
999YB5zIe5WuzT+2L3pMd8iEso2hWXuu+NHhMPBbdi1sfjFARZLji3fZqe1eNR3gDb9ey0cs7egv
kBHmBQWg6jzSl4ENfnFlP3BpWdqQSOepapqvUOuIYgi9KN+2ty/LRG+w7nANapHxtkbPXwhkN7LX
olzKlMtsWYevn9aQ4nvx8XJVFAX1d7galzBnoUVZxz+HA8vOS5adpJCVwmdM5RloxmJw9AHC9vww
to9DhTDx4kc4ELBwYj3xuPaqyQJZXPqgp9xPWNyztSCIRaEXCQbiXQ/WM+kpHoPmS39Snz23Iyic
UCpC1MAgPd6Ru9FWPuAIcbYqwoo8vNWxddwk9uqzMiMZkMCTkwgMiNBAkY/DKEMbqjzlw4rol/yQ
yfbhB15PMNWorOCekq7SdWuwUlqw5K5uxVbyMpw6HXEIHw3r90A/e7oODUYj9xQpNbu/Hlx0iKkJ
ff5qcWUitPzk7h3eIkRmjwvAkTn2+D9FiAFy9Kryk+NYNBN2/ZYxM/Y5EXcbPISRNIdPmhjYHEZP
L5OLQyvI2GwyTrf89tN52Tf0VwEs1LMF3aHbLHji3Y9ezRFu2PwXw/TIfHdAzNyh+a3lWAbxEvH1
YkLowOJ4ZE6Bp4P7lH5LgZW6GTElXqs50+M2uAifWe9adBx74G3RsRqGOwUoYFJL63tj0WKaECAa
DRd5GAzz/8jjcQjK8aItz0Axwhx+G+U60Rfs/fjN/Y1UCZMCG3ISAeg5JX1xE2cEFt/lqhQFCOwS
qTzFPMoEe1vRSJFMpt7128BS3kVW/uZCpYw4K66a1lhHndAAdxVNKIy/IUhYQG5eMi9qzdlWI60p
qq7jB/nQheYMHAAvOTvawlfnZ1M71Bi1YLQNF46BdrezEzSThQkZ8lnAvvfvSu2rpqiW5BEmZNzO
JQayj2nnl/L8FX+rk6HKShTtrkCW73j0x/+46vep5g6+6Puze4R4KPVFkFUNtA0feNukyR2kshLs
B5L6lFkde2F47E4NaIDPnRh84wMfQEcIzZQHqhTAWMprLfAXDWGxzN73/n6FqFWO2Y2m2eYTjYRi
hYZczqHDuouxGuY34mQgsBxyGYRB2xg44k1SY6wsgiKxZPLuABI0RpDcrLyQ1tfwS92YX7v5mgCG
TgjrnwsOzgz4kwOfCOjnW7ruhyEKrEKcLy/KzOL2S/a88+eU0EgYGEgNYSKe21DyPLB+YghrZwza
ktNJE5xHd2/yAEEsCLmVMtNHF+jdjQrad1bYgjzBJP31KElYUYJ3zK6W/lNx8y0G8GlzR2hbaHev
n2htmpxymS0bxMuC4J7KDzvbmj/0546ObF9hgrQrY7WnIGPqO6u81oWmwYXk7V1sFchcHcfFJV41
mJMpCNmrN4x4Pr3RvNOQvOlbtEDbyiBXI6AL8rQBwCOI4JcMk3V/pvyYQSs3pCDBthc3vmGEU6u9
v10FOKgl+wEhMYI6wErNTtrpT0uf+ir/DWySnfkiFfi9bnzz+FwBGRrfQDo4sZnh9nKmHoHFq5OV
E2dlnbdgK1rtnJbGeIMf4pahfJv0QgriDOYAwge9dpAea73W643f0HQ7AORAGojHvLbt3JpsyLB6
eNlFuYh6bv2tMMN/Q7kyznb/2AW+JvPI9i81g+LoyCiJC0wmlcmys7IwBCGlu0arQmLR6HSUWOQ/
Ex8A4gMRF+geM7FrUJ/i5AX5VZ8l7+C+hpMIYCxCgbTh6OuxXzWQlBGkhwuUZzWbh5x7Vpn+u1Nf
Ln9guHRE/M5ccG4AlwGvYUk2QkP1d+mh3Uhhh4lS5KjNXohgzyBMXkKhzajj0lFprNOQD9uxxDeN
j0pZNb8J9z4BlkofI6TYpCjoE0b9Oqi9C89fpJ7CY6cMIRCBPQ5+z0GWcv4i3zp6l5sHK6K8BdNY
Pi+dB7qvqN8cD+TLq9XmrgL5iDUC+1hOfx5A45n4wa5n2MFDza6V50aBXyfYC6VTMxGhnJEKeNQD
IikpJg2T4F8hV6HNQpEYc/2hJ1C3z74ifNbw3+Y/SxPIY4X3o2pgsiCmFEzMQqGLNgeMfmOHGhC4
WZmIx73HvbYNTc/o3WsfAAIX1fPTrFDp7v9FxgL9quuXZWIoVLbLHwfJl3Jr
`pragma protect end_protected

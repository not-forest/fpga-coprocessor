// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
lPaPagurAF1kuecFTuWvMgCOIGDI5VHmrzY1eiHXEMqdzQsVh224LYs0HVDr5zU8
8IBJBH/pMjNserAz20hZPe3VaPSzR1gtHy5U/WUdB4mB36nqjZ0msikSntaTHS5O
0Gcz+2wPWg77OMB/SClIDV+8sUS4XVwoXRZuHNBa+H3LeR5H+bJgAleQ6amuopoa
Q7Ym7/EegZEmDVS9FJFSS6j6QJKx1y/yE+H25OMyIVfvKjZOoQxPzOP+KrOSDQul
cv0YkEUdRzqWNlklKcLjWMFJIAvsoHojN/m0fztiYgwR6Lh7kk+zYwaldYsZusvQ
aNoKzATepwTANQ22GisTxg==
//pragma protect end_key_block
//pragma protect digest_block
PncG5GdNj9jqpWA1HP+N1P+LrJs=
//pragma protect end_digest_block
//pragma protect data_block
w9u3HFxRse53hYGGwcPpRG3po4jMZLM0TjW+g5sN03Q8W21kCLOhTHFQIa19ki9j
zMTnSbsiHmBjosHYOeDoGRrBwqL/OjZ1ju76jY4/sLJ3dosUfyAMCC3hTpMzkuYh
0BO/rysKSF7kfS9Lixhu046sU8fltPGzTXC5RpYat8BANARCvuPcO2lV/D3FNmyh
Z72nioOyMyCvafy/QGYSpvEzC4f5eLsTg3f8Qk5vQKzRLdcmxuGRo/EkbKxtSUWW
+XIw5lk+8Et+bXE+sNJ4cJQkCiyJzdQgN/N3FcCwehq6BcWJq4kAY05ni/s/GwoQ
hsiIROXDmaMlpiDnHHdrF7whI7cJeh8XLTClQ3YfC85tCSwTnBsYZwdHlHjx8c91
cjRqNjmsIKIwSgm5X1V7aDHJIfhCNk2MPJun4NGNfXfyZfpd1N9JanHa86VYn2Wc
ds9y5TzFMhTqRBBmul+I2ggu1RlMKtkImR0dM0m3ZOrkIx/mC/64Sht/a5TMkmDI
3/5R9GjSfh3ewTtTXDI4pSYAkkQ00o/537UhrvvEJQCLa4hU0ak4lFZLhfjgMmUm
vJoSviRS+8CXoyNohyA/TTz0reDzkMAOZbSnvcZwenxtgbcJS0MB041QsdOqLniP
iVlt+yoWqMJHy1xMYy37hvMxInq79bjyEy/Qih5wFrsGJWX+yrR5oxkvwiWnjun0
yduc0aSG7BvWBP5TE67wsIlvWDXJbUUaNFT4XL4hLafWfKJcyfG2DMkAJtaFRyCJ
SNp5HRdikd+WzZA080VH2ol8HiE3y4012pRo3ANRJZxA988aNwa429I9v6hc+BNy
xed+lytGCTPL9ibzJ8OfhKkELvbqKfcEulEFxzBxho4QeBBdqQ5s1UHPQlYobgiO
x7n/77X1KsL/QXFNvcTKyan5kZ+QKObV4p+cCx1u+sdpZJOBpaB3MdpKc/WS8C3x
s8ez4Deat3lopGPLU8SyqOELkW3IyQRlZU2+TwyAvglUGRN6ufZHdt2bQYa1vZDB
/udEVdcdvTIQuF/XtrHJbQ3ynmtSBBzFkctpiWm/rJEnefyCDq0pBlebbCtAUHNv
e7Ijdt3G+WOOLfnjzZwtNU6rqx4VDONxbFcekSImVKoku5UYJUGWfKAuMHQifUVl
9RlgDL2VocnOkidxK2lpxrj7TmRiLms32zd1gHGdTIWGkNGIrp82veLtOKUCu2MF
C7Ncffyh8FqLScwhreXaCL9z7TqnJ6aJ7opgoZMaLf/7NL+tRA0D+4b6tqrGmS9U
/aLCcfzEJsHtjn0CBppsE705mO4/IY2furHFpd/tdxSXioI6K6ztb0yD4O1sBrGW
bWP2Im0LpqgvFeKAGOKQJMYQYNEulh8BdXERYOBGNaRT+D0RcBTXnmZWWO3stqFh
Mva1pY1ltvo/sUTMRSVMXp5hCgTflZhsm6uP9X0XVFGRBJ4TN7vdJGZFYbMaB2x5
YUcbjPdlHvZjqMqPCTdY7eCOBlWQvD8nQmj58LGA1OiLUBqBaM8hrc4NPe/S0eQR
gd37Y39nIO2fwdhyGWzNxqvD3WpoBckXR3yo3uGpQw1wJx7UUQlAFD+GgZSfs3Wu
8Eu54nAv1RCXO243Q4GcmvEmH9ypS/yLT4Wlz+qoCuPltdJ6+3289iiO1kRwoJBh
LHptImXAauV6YYaihxcuvQLqWd/Vp/qsZWdIohf9H2JoxbwJWOoNWIliTRSe4JHg
uQ/2lluUv/kS8f+At6UYRAv07j4G4qTujpnbCOx60NAXMPqM3gYdivlw00rvSuaD
gL8mF4bwBcYtQFhE3g2SqEaEcA1RizgrVlK29/1yGtWIPas1KVIz+/EYnlXOQZoe
UklXcghmGRB3EQTgIhWFHCvdbLAnNt3b4uPz3jYXFX/tdECbv3/OyBM+vQ1Tx8ob
z9ysNgOAOqGuiMSMbJicuRDt4YH23AAz1E7FVZzd9HxIZ7or7aBvVeWkiOOlAmn8
qP/cmd34UfoC5IFIiPk4l2HzTk1eezLCsScHnQVPML1DA/3ytBv7Q7D8AX3gBBiD
wZDRU1sBXe2+qERwKvXDgwbA3OwfIpY1eGp3goJ1GhZV7qjR1dbyDJXCiPkz7wkw
WJfhEkhKbgJxPuo+CpJyZ+LQ0EyikG1LdcRKyzq/1b7OxPpoJ8Nt6FIDVjNYi8Rh
JrtLRkjHtgRT+s+6EIdO7tbZ3oTCSLVC1HeVkW1Cn5hiH/a0eKFSbd+hJjUbEwHP
j6YYq8YAdb3imzO1CAET3NIxZBLuI1dmE1koNdDHWR4/uMdDyBwaMzNCJzGKTVpW
oEamFMzqVtm+ZbhNAnO3KHqOGCEJGwGm+yZq2xj/AQZt6Xuf9E8S0bG7w/HSqoR1
NTVaRl/ipde7VB44Hdo87CY+WgPMWm2X/byIpVtq2TNA2gyE7VYlWFSnndqeMS8/
08CWqFRZkptCZT6HibhvCweXEJEapWltIVMuBTau+yRd+GojQwomy/nz+xJgO+m4
Aj2d5NyP831GMNyf4ScPp1Z+p1Qax3jZiIOP8R+tgEm/WsmtRPq2yHN/APXfE7BJ
Ebccy7H8plBxaZuHsfiW2gL5zH5mGHmYjgAPttZrHVpTrn/bHKpQbuy30VS5qMRC
o1gdeDi+TA7IPKlkJvawmzpKNbJLWXCyANZIbvcBqGD4vDQCc0asKVCH9zztyjlU
lsv71f7sQBy616MKXvwK28+3Kl80x7v0cV4h1BvfNLa86WRe1fLrNd6CKANOEdlS
HU6m69gRUxtLZiChGnMapXAQWmz117klm/o67eGrL/PdOTbxmkG3JvkHoW+E7qxp
ConCrRW2XjJ3MXBVdE8GRW0f+2FAYTaefol1d+1ZuhEcfR7EcGpij9kmd/KKB2Tz
kNIDwWZ9I6fwbv783gB1zub6O+QkwTjmzy85sMbRLtyLyuBv58rjehmMKKa5yO/e
xjIO4zOxjmyFc0E/wGC1Atf7i1L2n/BrTvj7GuwLcUHn8EGydQkzxNRizPssG3d8
gcBBpXvk0zY2+gTRKq3kdiTciWTOgjKmTyTN6b4fRgatscmiH6+PXvr5a1a99eQf
GNoq73XdnBDVr8vVnODJ84roRjoXhTaWc9T3yrtWJaYj5j7q1Fu3m9rDkCQW6OVM
a5O+RbXZruO44uVgPENRdhIOomH5DVZBwOxcNaS8h5nKkzML4grCu6PVnSbXiZOi
S0/bMQAtbXeJBndUrRKA8k3eMTrcsaoSI+RVUPLzQJfmi/20kmQWjikCUYo7AlZD
yzdPLU06+qEL2YCXylijcsztOR/VwJ9njfQryXL5+2/+h4UBARewWZiz7PSsIluN
U+MP6wczoxWkgP+nOJvPtxx25Zczw9VnVvKbcDgqdrU3gHFVNU0mfanCFM4eIfJa
TCDTuivVY4CHqfOeRWFJi5WDlK4/MDaEHmu7mdJj6IIPbTh9RSYy6nWckpPhq0PH
KoOq1ydyFHK08q/x7Be4jJ/od9GHpzxiMdupwBxfN2UeK9WmbZJ6DF6pvR7QRsBb
FlOZ/gQszMp6YHcfmhvHExBqygT88KisPaSGyC5nXVFUG0bJV0HWqJyYjPqhdLME
IJPSOWI5JE9lyd+hCb0nJVj1dfkzmSzOGlZWK21SMBOHICXRc75n7Rs9M5Q2qXk6
mRHeubSHz7JR9Pv1U95gSEoWBEcnXke1r42Gsyfg8yCqQw6gdSfqk48P7urojibn
vGQwCS4LkZg6l6LDHXyW+9Jx3JdDJHIy/07YsW5V0VYSxBgCZkYEdcpt3C5Esgar
GxdOamV4MNMNFGplV9QvJX3rLUbJDgkFxzGRVcH7y4Pvo83AfJ9hBQo0q0z87h7t
/KOCvmMeDSnmbo5aZ4vCKeLp7BBFMrps4QooCr8AUaadMv50dK2jLDxs8LrxP3YC
Fj+jHh0jR8cqSFJG3v6v+Sx5aa1TdkNclbnMQn/P02otryF+y22ougDAyVqiQLdf
Gczae1PAW3DFELU2hOxwuairdjGiLC3kgTVh2iVXS21J3o5fy/9GpFn6pM/Pwz4C
CnfGkqEkzDr6SqnJTiyZSVnVwh0S7oBxB/lAbf571C03qDBkDudChDPNvzBSRYmU
GibKAASnt8COWgktAeKZxNPcCycoYou7XstBpu3s1JFIOU/LQgceAhqS1BuOzJAy
29LeqKFfs7x264GKWJFI9IdN8WcPFtY+3NQgH94WCNS7DzbIeMpu/trNW1ZVyK3F
Ck12+QDI2d6MzvEvj3UPwjQ2xUOGHj9D6g9JhZW5vVdBYsOF/9jFySVROjdMXeir
aYboN40MSoNREMC6jFul5sJXIUW1A/iQeNWP4AiX3bXkzBkuxjq64gV7mQuKhM48
hJQLEmDjn0vQSokM8FCjdhpbij02SyCGO7Qtt9oNi2SYsm2Uzwq28EddjC6MCY/G
xjzbFUfj0bWSfaaSBlXITOqkYokwv4jRT5l97BENyQ/Z90gpJpbq19tBcJxiC2+V
rndzgJ3JxisRpnHJqELJB+MGOPx6KNfNjI49UrAJ1LPr3POjLpjja5UN5eyCmI4q
Oa57kz3Z5/N8zhOEnjUxQnYNwSep20oUjs/8CuQDBkix3JyIBAuAtqwp3T6Q0J/9
4gfX81rxXXuF2QqcBZAoOHS2Tf6V6V5nAWJ+JKeBXGRGv41v97gXncOKWYS8Oy50
Lid7H4cP0i5BPP6Lsg/sdC5os9zpRuYx65m/ksQQPwWyjgS6fAZ7ZnUDyBHl+3Hk
kwhxnQBcJ9EYaEpMRCTvz6dOCiC/xELeiZwzX6IEy6Y/1I4FBdjzP/6vhcTwFlwD
1p0hTNJWc0sb0T8OLaSHVP28WF96cJrXX4Qk3I1wnV43aV5wxYR4B5hsNXZoSlFK
ABf30rDO+spENcY38lFyxs45yVthNgBLp4ZttCoZTRSYxCAGbs8cl3Vc9oO+4vf1
NQCanveRZ+orYkAjcL5/P8/aOrz8t9ol7McVaxzmY+FbFKVLkyXB0/aJ8tV9+7V+
7nNxxHZuwIaWiFwoG+b7vJBSB7NB2gwOcCT4sc/UDQTXLGJrAHQA62yRUGbrfkp2
mww4jl0TIwwL+F1QBXxohGnjI0eOQNmj0SDFxdcwjfJi46btSy96yjPtN9DEKgY8
Qca1f5XBSXlv8e+hYihHB9i2Rt0puZz1/3NJ+wYIWJ/ZqLB7Ao2dsSPwdKk2ENVo
jTkssmAClAnGeRIsD0ctHHPZB4GiDzfkJKop6Xf4CrxwiB8u9BEzlyBd5bbD+JUr
id7ZhWF0z0Iag4bLE4KnYYlHrQqEw/KX9AHQYi/c5W8r30znaNJ6ZaGsUqkwQB4c
+AfYBZ25vBCf4v8IV0HP2++OZ3fD0fJjKWXx4R9Ki3jianehkGFl4wFguEjFKwQn
Dr6nz97albfZQ566gTKkiu9LHGpRvUZC9lzn3+p0PqHAGzhpHvu9KgfYCsACD6N4
dbK+/ZHg1SGM8CJoNJK78A1r1LmyfSvUQL4obnkPYEaDUDMeIS04YRlcH/GauC4l
eOwWMqsyj7sJrqkVi1jvTK5gINZr0/ZcP1/+9lFYOKrN02CSDm9YBNReDvT4W/WM
HmppzszGX8xjBmbtEqOfbH+YSNJ1YY1kLkBfhOC+XdwyZfKWVORCACuU8Vyiffr/
Zcsz/asCO48zlwo4GWNBgf3z9hGLyjYySqXRIOXDbFLjtEHMOyyKuV9u+7lTgTZO
0bXV4vmTy2VBrMJvfaDBDY19tpfWUA3yRw9VeKmXBFuj6Hx334o5fPWzwUkp8aqh
uaJ4vZ3HA3ePZJjpX0EbcwhfAAPUFfAbb6a2mjqYt2qMJ1ATDmNJQZ7BF+D3Laoe
C/Reir8cTslmUKzzRV8nn1omgEBWEhUeDQgRG3Xf49x0pcHJVWDxjHc9KoZKjvdp
Zoip4CxDApsf5ow7TV4k5eg22xJdKi9ki44WMnl1n7YBmc/d+XPqHF6lkXuwxtCK
N0ajFGgRApuseEsl1tM3+4H9BBCK2HJTRgHAgx0m4TyM7CwT+Ja1814q3gTEE4an
OW6zKv8vACU0xCqy0dwCdM04TlCUSFJEC7yzbQxPi96OqV4iy5Zjd/0kaW9tiHTt
fpLfg9ZaAZOW7Q7n03gftsEgg3BTRMf/QKhwoc5l6qj7sSL7SgmTXB83GAkZAacb
cLZ1vU4oq/lDf+axOTyEpXlDs72QgbDtPa+Caubc1x/IdzfdHuLtA3xZHKEfyH0Q
8AhQXfHLst7p6zY7zY9tRdYITupEiElWidD2cIgo758BxFIgY5SgZwk/PARtER2B
9idZTrwi2UMQ8BM79eLHn231Z1WtIZOy9XLu8ZKydtBvh0jflZPCz0Q33I0ZvIhE
lDecUNtGDjxiHaV5QhSSsqb8YJMl2JjGOInHN9LlDIofXjm9vWrYwFSxh5M44ls7
gukXly8vgGznAk83sHaPgDzsBnprrB8XpDvQ5nM7oVe0ohpM7KEqPo+Ufa006Niw
xL8JToYYU4gIJFLQCZXPxRqjlA2pbJqvWX2tBz4QNRTcNV5K4MIQSRmasEkFDtGC
T4JhbXWLbSd5JPaKtdgUhGvBLT2mydO2/XauRvzv1h2GbzuJFP+k2PwkszwYW9qV
+yFiOC1/4zELmQufB+XZ3C1MChdHZLOMefQImjoDYt/QbMNwmngZ5t7NVNTlhvsf
dDG2Z2Y+htMpm3KDzAM6t5pHSWg4uuIXWdn8t7BHOBR0D1DBuEXM5JLkdf5zFEG0
JxeFWd4VVcCT0aGa27Q310Dp63HLjEZvyBTtHj4UO0ASNtmWjds2zhQJzhoWU3Ge
4pZvNJc1Cp2qP+81yfinHt9UEGjDChfdW3aNVxDjRTXKSQ3SfKw9lsl01OJXDMFh
GNKfsBWHy+tc6mbO9WHRGpA9IlB2yhT6a0p7BMUkMLdV/kUSZ85qVZc6nTtKN5LH
P9dQKdBwdNdpZcIh0w2SdnKm/04EwCc+A62BQJ4tqq52jzJRm4GMuw+4GuBCDH9q
/iTlvwfH4M/7GPVpQcfHaRPuuarMeO4dTXra6FCLQXcPJvFH+ptBQrvnfeapcYHS
+QfvMvWld4A41bYWNXa5NQLJrtGdih+k/fHtk62VSWvQwhmEZvGguWmH8GT6UPiB
VVbvMG1xLvCWjTyVzkEnharOfUWNxZ1ZHmMrLq5jNSluwqAg+ndesK/L/YKsoNds
yX+ZyWnl6jVlEFDNnoKinj04w4aYzimebVCmRnqJSj9DxxD7db5YQlAYBktWO3I3
IJZHh6bnG7i9giKP6G9n4viOybixn4WQ9kLVNq5rexKsz8VKSXTRHUNdzVCQVoZF
7IvFjhFW//lTxsmT/HQXUnq9rwnsY0ra9RgoZVuLAXCcwuZ5BGWMjSBrQH9a4Uoh
FrFOSIBqQw+YcFLgzHJ+Q81L3HgLlT/bHYO90tgtrQSctRd5vUvyHBUXccS9Kt/+
VaQp5EfB0oHioc143RlIlFrQTSVMqQZoX17fDVh4tdhBRdlyaXULqdgOwGzr6mfX
PcqhrXhQSKr11+3gAgce6lbV4Ao9XXI7BA1ncjcq6FlPqTzxstClUgtJOVjlSygf
/eE2h744BTXARTDyOWer6FRpIf4rL8XkT8Ye3p+PgN/t0sFuzR6L4KaErx2OoI9s
E8iDv+sSWi0QS879lCFQDDnEUXJWrcDz3Y02u2tjc70b7pyzJD5cHiVrvhyG3LFe
HYV3Bws32mZM0NDNG2JDmLxoCWHxXfhM5YOGF4WLhiBHyXXHnMfP56FI/v+q6slA
wTdaJ46J+OBDz51taoArJxE8Wq7dt1O714wlyLI/yxxI+ediC0bj2R77TgEX3nmc
znGEuEzk8mKuUWhwhkQ4a0BX4zRhszZoyYGdu8tJtFUk1WkhWm/pHZ4vxXE5f89K
cMJitKmmQ3sLH64y4+wUwr6gcxlZTf5zHhNzCXaUrAKfsNX7Sf/+G/EAa6kPPnmD
aRAyK+U3GPhnlLaD9Sf9VQ2et4PP/4mGe9ZS2v61m+bioObVS4e3jdT9yK0bSZGm
XUt2RmubZE/8Fcqp7ZvVWOx4ciyzx2ktwjFuIthR0fzEfT81x4EzkdSDxhWmyp+w
UDFLOo3WcQrMsgFQfR9zQBWOxocGIuw5dQ2scbOr/No2LD+9buiQGjpwCmWGP3Ih
WzBeS19Qe3Qu4iJuEkic+L8n19PeNsMkCsY7vskGPd/91AaqOVy34GPkunFa6GiT
qvbB/4ILR3vOCvHqgkg4ut+PUHbPy40Ql9D1wkk7HdXtg5LVapIa8IQ9GdU78fjw
jX877NTk8StOy+SUEwwcdsKKBLevJF+qWOKXLsUnAQuVuJ6bxDwzz8Hf9GwIoKK8
KDlDPHbMHnex0mikaJldBbWuVN+5CXOZt/YiRVgFJgWt+G4HyUdWUmc1aZ4mcwmJ
w08Ja/HdJMrUVjl2ciIMyNeu0rnE1lY8e8QO/rDQEoVgbD1xTY94j+tdYOHE9bfi
wMQQUq0iHuwtTA2DEaQpgxL3WEwn0u9lzY03kp+/AX/K45CWdxvJK4kcp1NswLsx
kLvhtBXfc6xBXH2mpFvttYNZthx2Ef4zDFFt8JnH5oVaKr6Tee/xj5mBYQn6igRJ
Vzuue8673PjatC+5VmTKhOs6fB8+0d54PusCbEeZcxzd2L1oWZOGKAoZSu+dbi62
QVd8Onh8wbZd5SPaJtfoedWdY1JKEvg3rIj8K8s9NYIXbmU/UOdsWIzYIaTPaYto
jQgf7EGKTdO+l0VYDUsuw1RwxNLYfLMYQ1A6WH4OW2SZ6rILI6iFax9ub9P4g+yh
o2dF0L8rMIPD0zGENaSdlteUxvTLRHEk95tPlSqUnRfWSB6I7WgOF4GbrV8EDq05
uUOE0FOU3uJX+SXhAkmpTKaKbWpaPgENOMPYEtj51vM8P3vDFmYH/EqRc5rN1xRQ
3fizNSP01OA1aKAoEH7LDRPitPsG3YwqB/ksPEP6dOLRIHcKRKJuirjqcor4qAg3
mCzOUpPFgmWLdWKPEfD1CQ1PZ7baMkcqxhRev6MzWi02i/Pjzr6Y8TDEouoxvBqa
dBD7/vQfZvav8TDRxt6Yom+tAZQXkVkg//X/hiwVCFDnw70QnNSwNR6Dq/IWNrkv
E6WMdm/5Gv4alcBc6vRvqiQqNWkYrMAg4akWvxNl/LtvIeLuj4QxdnpzvXbhFpp3
hrcVJFkfQvEHT36JUKaoaB8FK8IXWcILNOrwObvVBFQyuwYUutZ2fZh+rPt1lKEs
KGFMOhKopxj/8ReqVTwOgFlY8RfIh7lD9assJfYNAwZUv1Y3MDxMVPgnNNPmNaww
c9tTWiaVdV5FEakSfDxE7MXGONrozOYKoT3yv/prSxekki0zK1hFKEuHUENklPN7
A0RMSERQknenZvE+OU6GwDfSlXRuPJf8rBDc32L+pRzcDUDxS9n3fD+l3cVuBQ4l
UQhSgEQGkpY4UVL3Ud/GdbgCBIp75vagaHV+MogwXhR/yqvW6iU3MByILbwbmnke
0iLDp2rkLyi6Wt8E3QOQ4zMxwOF6eMqZp+sFIpc8g86VugXmU9ihHFNXIt58RJP9
ULI3/L2wJx6ThXhr4Be0ijrHkvIoKvqTWA/5+yBpqMufVMAvhET56mylnH3vtIV1
5dcHv+SHdKBp9h4bLh76D22Okx3+kdHl3s025zl/IeEX4RFJg2UaOKtBhD6ZrUN1
EWX0pYeOpPcSOa4P6eXHyL98km/vONX1nRBVR8x5haUVJ0xxZQT96k15CtgHuIIS
ZfAYFcmUKW9ETLxmnBdkaXOXQ6Kskt0pCeLTxUY/Cs9HQ+FoFKeZdWrkcsYE6avU
ZO9VIIRA5PCG5Gf1tmYbyv0eIOaVLcqfvyYrS449C04Yr4QgVO5SaYUVQ9lY3yUq
4w4ua7zzS31YiUyqlsN71/+i8uT9U/SLsnnlkVaWLvlPk6Uu4RLg6pjxMrpQc2qs
Gak6mAsN7Zf89lzttedrqbBV2vHa+xiURxqWtNUvBfZFuwylEpLFA8WoS+D9y4np
JgWSMKXnPNW11gG9lls65BOxcvxFcLgRPH/B+5UQaV2QHcwEDozCHFT3Yb9f0rBL
3PNesWjFKyM6Qj166ty70cW30JpQnSlRxdjKInS4jbqKFjvo7cobiAXxG2gPDAjA
/n9NQCuSwUvlLrMEp2GfhHTeCZF24dL/HmUbbu3SQzxM+PPL6GftVT3y1V8mC9qT
qcWRdwaL81U7h/1Dl4UG5B2qCr7ahS7frJ1f7iZ6D3Sf9AnHJwcQSTya+nSI5u7o
m+qV25M5uQCjIThTvjGGfDT3lEq6I441Cz2P4PvVBjgSrhZVeL7YqjB1000hkEvT
I+MRry63s7K1urGQL5cYO1tgly6wSQ1PB3wJcMMaWe+5sdtvGcb0hY/yagnJQPCb
KDAzgjLPtVYUbrDsUE0U5RedUQEeET//QbQ/BOrP6wc=
//pragma protect end_data_block
//pragma protect digest_block
aSFXigD2yEBuYfHqMVKpG8+XE3o=
//pragma protect end_digest_block
//pragma protect end_protected

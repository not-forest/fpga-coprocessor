`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MvZ7dp/iLmo8UkM3BSWt6b/MCBAlIDxG/vOk8UDoY1tx5ePGWZvxv1nDnk8eFnqc
yhBrxYkyDn8KokRd21c2wnjnTyinDanX2vbNRloRp3y8K7JTOFTVfm9Jb5VFZS8I
aY02sHdpGSHYyrSW3TOdpzoVKCOitG8EtFq5Ta73KRg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 63248)
uk/LZFHFZb2jynxplWImg5o9SYKYvYCGWnNlaq1cm24YJ/3LVYdOq3ZXXj6u5hiN
XIwfmG/WIc3T1K2Wi7EqWsjOu6yvOpEd1ENqtMwM7kKyjjcC/bCVwohdAsnZrdCR
r/OuWb+BeiaKwtnGRNDeXUKaFWN/K1IjkEubFC0FVR3vu2Bm3I4RgvNK0wNEvPsV
UfI+lsn6rMnirPKAVb5A2sfKHvcSKQ3if9H4jL42JsXz4NihPOY1izLEkvY9ROD1
xGY59RBN12+rVL61NfkvFZcLXetGc3m59c9NBaCVsZIf9HcjmDTe6PNRLSq0hvGM
chodDCdZ7BEhFEcwoarSPcXHGkrhISC/mX2mb0ikpi317isBa/TTjsAowo4OfMyT
GOXOSAUxXayotzxeOuNOXwOXX9X5cjBIopN5nu+0mAEwFy6SLKn1gegQ9d9aocju
XyXq6+9QBWdONh4tuKCVyS8DfpsvBjIZyOW8LGecWcdKUrxsDWyjty7xBocxNqbO
jqh8EbFYMoAYWvUamE+ZFDegerMX4JkRt6ugca7BBWuniVRkHxy7CM6wB3ff0ynl
B6MpBvBHGgd7NqLYxmFcMCI2DhLibTMkasg+9w56ostHqYoyATKyFFbskYkWxVi1
46F7EYJWDYbA0opeosFzQQjiL8G/9pDVrNzJgfrMZAIRVXmcM3J2kuTRdwpgZzqA
N4/rWgX0jxguPHM7QF1HPmre5gApKbcak5BYPte6DFNbPn6J2IBCowXZ/z3CVJMa
5YwUY4PS1KQOpd1kf1q169tJcF7eBob3wTyuoQW0uwj0uParfdE4TgGHJ5IvFwDc
Ua/yYgDFEIS0fa+u5R2bjL7NxTRDCydsRBrpBvNkyJT8EbGb96HkGHfO3FNk6fvl
CGmrzDyeJDdFZ+qhF22QstsDMoPKWr3FYyNuneUrTXen8rpL1Br9W3eYjuTjIHIh
3LQRRjHv0IY9/Hctyb468lvlSWfOMWKrUKr/SYXxzi3JBL41cnkR9ZF5CSbe88Xm
clesr7BXLx6v6E2hRGU1gq8kzRWA/JWgSjUtSEzqNK8kCI4pTL7X/pkunBwmMSsM
zj2JKwWR1lhSm0rPMIXtPf1KUlmc+5bvih0kZ0321p0G4eTo1EYLanVR16FTTVde
Bz8FA0zqBVwGfLgaYSlDbJh/nQj6IMGplZ7Jnf9R2hwa5VzsIzoxF5wtDF2QEDsk
uT3xNn08ymy3ARZH0XiCFfoqU3WCIy3fhP3dFZfwHl2lW3SqrQDJnlsnaQGvFfpb
BQNOVIqV/9QoJlCDy8/HlZBd6p5F3hc0N1+DgZt6HjaG7DpbxeUVLHlYuspHMWnC
KunjexQ9CY9iRhchZUgLBnqfdHbDVoWBblWsPMkrypraOVFIjrEVJ0WnDkuBeth3
UYZS5go9CD2jowKTIRqGu0fdBE6DCsyj49XLg0pOMmKygYEvCOPBOGCPs1uHxl11
gLf8UBJPwE7JkT86QJSTYVvNZXRxWGUxbZnO6lEN2efqgdUMgIEW1VUQpDQI3CDq
tCSTmxra7SfPgPYUV9Gyqb42HJ4odIuqt79SxWXetux4p2tjXkTcd/OELC6Nn3Rf
tATdbZFOseVpllBscxLZG9b9clxikadLOAgMrAhVQ2BYmgkrRApH71F5zGATS+NU
FBQVNe+27vo59LtXRr9qMN03YDxq1VdW3eQDB1cmTJvu8p5Fbv56wKzxixNGO0uP
5EeJ8Akrg0trY5RgUhcFtghUUJWf1IrPB1zQKJOZQMlCkVNUDf4G4ax9ygI85B8k
66Q/lgZv4cb18TvWcLRbHz7n9HVO97xbCVWn3hTLg5+X5Dmp4HjkjumSiECW8IlO
GytD2HWZNU1Pjws6dSViqIFH8zl/zbWeheQYPXGty/eVbNq49eGZ11n1mmukm1Q3
WRBNONXYH/ts/S7i5nZ0k3UEgQAduLO9rXKXspOVw5tM8vG/er/jPvweLW9jJdMx
4Apkhsnw/E0KFvu5bsnYGJR5i6VN8k6bt+rd0v4Ky9c/P0X8CFeaK2dN4bz7dIIT
bN4kIFolqPrWB+UVgJsf19gPkl6o+x67SDBpePfFfJ6FEx0zuWOoeMvgQJbmmFc2
JgPuIutCWQobutA5oC1915iab2hvhKxbd62XVQm+if1hcMvMBP4Kt0tLUSEF4VQd
OOvnmxQJ3nrieOeVLUD2a49ve99MfJNPWHLG7joMQZ8zg5XOti9y7EKbJD99/xW+
GCZK9GuMaxAc3HP3cH7dLDnzCqtpPYiL29UiQAwO/lNwHDBoxdekXkvirnCdGYVi
1EHu/TfIrBJzVLrPjlcuw2y5q7QKtcEK3hVrE3dfotz50xTEo+Z4Dv33VXG4G43Q
5DpBmhWJ5S5MLGXdM59hfOoyDeQCTqrTg74zHW8vnO+N69m4BPCx0IdpSHjRTeqi
nkib+2U/l6z6DFwqdA1aN/E9QEP0tH6lkQJP/BzqaMj+5HieIeMgrJxraGuHwU6+
nQ4aqupHJ2058UfGTYMzMzwnYlAe+j6j+5GfNRmavKB2BLrpEhbb7elhOHHHXBvv
dq8hVzg4pvTTy9/gzI/9+vrTXZ4iKtYpimQ6GSugl7OR0BGVfVTsC/tMZdIl2k5m
6sDBWpWnYk9CGKM2VcNyKVupDAMlirB4SVl7DIKm2HnsCUk7H8ejpbsd0+Ww7XIu
nrjqKxLZP5vrFM4TttqhPMC/BH8HhibqleKo+HXMlBJ+rXjkeUYjsMNQjGVQ+Tes
iPxsKhouqsmKfgyBvuYp1ZMFwFBmLNeK4rOpEfbqbl86pv5QkFEVu0rUTvQsOLrw
JSHr449l3io7um06CnrCr2v01dU9wavtEt8+apyMH9zzbWxgbI1L9EmfDEWV4kEK
ww1J8EONA6GiOKe/3Jyw7AZRnpqf0yeqQHmUvHc/j0B9WDmi8t9nK/ib/RXxXON9
Y11qAhoIMXB2Gk27SaqaK2PmetNC5fykQbO9xqgDOM+0SDegK3ZLzuxq14jDbJwK
s2M49rt1tSRLW2Dr9wTgxrld2snzB4Xum8FhzN7o3YVuQ6naEfbaU4PRRyeCS3Fp
RQ6+Ggo6BDLf9qKvW0E/L32eV1dUXzaDbWd3Ey9LBbSSZq7UWB5U/wCcWBq9WW+f
+BoZE/20NW9NeZDtSIkr0CX9D3I6zePXHLoL+G3OYP7uErsEinVGwb0zhyiJINKP
e+q6JOpx/YqOog1aspCCNZYlUxhuUzuRf8CKFDVy7LSPB7NpzY5XPU8D5nqEX1pw
XXcCLj/z2ybWQUG0iNK4XPOgeO8n/qFTuvD/24akybTNk2ll6vdq9Irdsw2Z1lTs
bMdh3ePPDOiUBl0JKirNlYg1Af3OSnqdykON9Ue1yrJDg+x1zdO8OMCuta2LKS+v
tsxxvYuvKnDaUMnUE+xj7VM4IaKNGdc2F2HGb5vaNm+RwJk7ydb5ZigijIVXX1Xt
moxQddBuFnsqeZ4jhVrTYSPq7kkY4rQeZYoeo7SiqIELW0YK1O9AJSUuEmPSeShb
NKGnvORxqyBJkF6LRgryxyrb1HMnBRdcT/eGcBQjsh+IS0dd0ZYQx/MdUe5VYJUe
R0oGUOa5tS8rmUtSj2emSz/GM5FVjfzNrG2Zey60WN93vrz5pjOAX6XQb6R3aTrd
FW8hyqWMpCYhHYKR3NgNaAknlSe+/aasA69cz0AJ8LpAT/pMsXx4F2Z2JzE/Dq+O
SiDRDU9hxrBTra3JPHD1KdDeJgEotyhBdykptzzG/PauzyWTRWtI0u0kCLV1MgpT
hufzRhuZMT9HkpKV9FFyPFQPjI/v5WIS93XlAbW0jCCDmj3QhYL5oZpM6pzlPg2e
D53Ace5Y2Z8wmJ2jvSWP18tvWfRt9A8lBiLLL0ILd7sQ140bgRyxohn68gZbo0CI
vIfs5GrjmD9qNGaNe4nLwCcusV13AKSs4mHGAtl3PsoJla6p4ad80igRn+q1xtK6
1juElpBWqX2mXSZNzOvLJnCr9oEtbZI6xaYef5MJjo208fu3pswzz5dzg+tMjqfp
gnXXLVcEcttM5r+dN6ArK4zr1g9xw+TXS9w50j1zEZHYyM+Lp62amru7U2lpBHRi
2aWPvl7kBn5ve97frQ6JTN+IUtY7qxyGnY5yIpxbmGjRFrbebC7NnP6WaahDMyGA
UpXZZIsXdcNoxKfmq3Bx578efqZj3TdEO1iaX7Wmi7bJz0f9+oBxFNevLR+MBeE0
WJMdc78GBUq+FLv83zScpT+YvFCahPJT9xWG3ycmE4bPwLiOwkE/b+McCaP1YoFX
Aen5cczI2WGl8ZvVaSURYpqOkwAcF/0+RGiQYJcxn0oNn0jAJBY1djU1T/wEPAV4
f4z512KR3OEWJsFohup13MFX9YLIT+aOd9gEBgL+q12Ry26Pj00pyMG3jjoQfS0n
ZeoYSyQczizwos3QSTbFwUISUTdM0QrIJFGGnRCujrEuRbTCE7A1Yqq1jmed5YGU
IIa33/jKiRt+KCBYK2lxXI09iTUMm7Xb+h+fqxY0bs/s9480NuhqE8t7rUxvMeRX
FiwiKkofOASew9I8MdbCyjrkFhR193rJSZJ0R7KfKyg8Lz+ErRsCVMKZTo3aZ6uK
0TlOZ6c8QgjltW2TOjquRMf9iQUg44QcNosHE5geFgzIwHw/92Ar7pd3SJHi87bG
JNJmyjjB351um4tggqp+b1+8ao1LLg+uBmcTO2nfgvhkT+sS7cemwTjGXcN7FT5n
DCX8GCjYoFcqEZZH2YVASCKb7F/xL71UGNu5oh8XNnnaHj68gVhDp/WKtX1YLL3q
L7ylVdIhY+WId+lMk/7g/w0B+R+93y1wodKOFpcIuJ/VtSihgwrxy0qtS2/20XMt
B1gG8FGWSF5sAREaH2eGtUWizN2ReK0YPLr+d9XE1YF6TXvjm2Bq8MYqGlprPIHi
6kYBN7gIjANvDXODNBBpK6wgsW25uaNr+NYnOTVTiG5FkXad1xcfvNpuyUwX84Hz
99h6Cv+KYl9bwdgGw4CmyJrAsY6zWivzH23MzWkPnQ32IVz1g1IDzt7M/3rI5Vk8
yn5CYZdOpTNokbARYhuG5HGaDKlV2raM9I9hmf19bhgjJHnAivtEyFBJf5INmFjG
MW2SOo602kRoyLD1iMHUprlP5jUzjebwEl9Iki05MnlaWc+4/hHKjZVwQpFC1krC
CRoXIn3NFkzumTyhGWuyrFFhJVOIiF5Ef2+O7zvK9CyV+qieoSDKNzhzDq2fCwDt
1p4+Heu+SCojcfrb/G2B2v7WCH/1F+rNJMS6FJp7RZcYHKS5OZIVGBFu7z2F//yP
fK3bWA6MPWDjGKEL3wJ/1osBzvXH8oGLA4UpVyxPqxFsNLNweHAA0MGOIA7zDtIO
Y4HtNE8e3GLAcac5olS/yFyY8dByIS9R2VIOS2TeCgiFGH/GZQRAmV+R/H98SN2p
PMKirZOC7RMKTYZc37SW79NliRfH2/DrnGlN8R17TlZuvzNK2n6cmW2TLBBAxVkG
YFv8mlpXKQfaheA0C3clgaVjIb5BPrHcc1MaewbPaCOo9Fhad9Yq2KV01LFuoJH2
St9qbbjX6FD3ayOYk/sdV5u/MpKmm2H2KVhSlAHoGHvfCTF/32bsSxI8Hw8e3Wt5
o2g6hYYK+LfEC/SLr4E5mL4EyrDjEREPMw81tZl7jBFs5k1mFKlFudW1SsIcUwKi
vrcvMA761uGx6aFQ6L2RpHziu0GPQxFXAZbZoV69WBX7mGTSIJrTsFaze95GGwrE
I+2Rmpj3/A91Mx6h2AQOTkJseZLGJSH/EimBlL/z+xQZV5Zc97Xz8qWt7tD//uSI
0TVzJWh/UoQpSesOUNVJoRcovbw+a8+nQ97dsCgsy/eu2VVeuR+9GDG4i++VOPD3
Eb+/LMdN+wjmS5UNIuGE00/MAbJjaKz6meohiv/eUZXW6jjHkIBzmQlaHiyyroYL
YzMxO0vs9W4I84mmrP0rwgd2PvUR5Kq1KlCuzSNd06URgMUGerHZq/MTUEjermit
DLIAzpOP7NHvpFX5naJbST5WPo/5QfBp/WpP3jiH03LDFg/nYQ9+lH6rxsBUk0gl
vQKXv4g/2Rq7p5ng0rotunslJzWYxCeJqVl0oGP/2gpDrdi+cvIkXeqkcn4S/cvp
CBARh8vTAExWfuUKVix6OPh7EKfmpWgXVPP+KzAYmRzbrHQPPf8uo++iw1Pf4Uk+
tT7rMWnpcvls2dREy+WVq32IrXXL797kvzmQrxQcxkG+AKue5qmvzZOH1Xm+6dx9
sfWw7URCd5Ken7M5tmRpQ4IRj1Zppmyqc4j09Pw+lteJXLCdX90n2SmeF4UeozKy
7BmlZGpP3aE9oZ5U5X4WEBBOY+O3ttiBRNJkQa7ec6A6SHQuHXK+HK5dI/ixaEzP
gGPtNQWPfz97HUV/XqcO461ArqCmbXdsKaVvqHhoPm63/asYiqtRQZiuK9Df4WKg
sOYF591iKZcewkHvDibm2IOueAE7C1hXuXy8TQtM+PClmO6ElSI38n+vOoLCXkoy
R91R3oUZ8Yob1t6/1dS4Gq5aKBjKl9NxbZzycLr3ZnqnAk/JrIQHGUf91YbTiUCa
oSDGar0vhyMe3hW4L6cgeCmJVCmu7rye4gNCpbrntWmylTroAC/xAQppTPNAJHZi
Lzl+eXYnj1d6WCeIazZ3cfIV7qLS1/bvLjGkgeZXRxiy0oVEpZF/VvYDhBmsbzdu
UHdmod98vdCvYtXnvF/s3YoYn5GXkpg0cyA1iEHFxvbkCJFlI4jckY9j+eaimYE3
ov0Et12VxbUyCQjp9nG2sntuj/5ogiVaT1FWWd9HQLY5icH6lGRcjMlyYIYsG4YA
3drBsMcnb8BWQidPl0bignmYwWb14uCoz1/C1GIHzEJCFJK/wAfpXfSmJzmwl3f8
iiX2I/GJ1AvZfMhhleUSMr5BaQXRXZjulcpPsi0HXSzYS177UN/hZqCWw4RObyMx
xSutOF6q7P32R2cR9vHOcVFCGgnh2AtMRxbcK42di0remkKkeQ2Rs621zohDRKZx
BQlH9/Kkix0eruPTpsT5sR9oejKkCCasP3wC9EJv/VDY0i3d+Kv01ewU0y6CgaYP
qDG31g+i2WcspFryqLTH/0Yx+qRej7GxgwoUBs49qyBiwT1N5A6Zli4/ncf4VMOq
KnLA5rZSI9PslgNGcS/kQY9wZ1o1CVk02haYSUdC5VWQVTWeKPMmDyESaSmCMe7j
2X2jnAystNzw0DxQS9dqw4GsC9hVe0O3H18T3qINFyDfgo1pVOECS130J9YONcoW
PRmginb5Rae2ReY1U4WGp5waKJ0gQtFk80GI4Cs39FVp2vQBjk4lqdVdUtQFdDv/
65+b6OCHFWMeEj5InDCsyBAjzWjOOrrzEf5oSy9U+NDegpHIMO4xnWmtlplSOqwU
Xnb5oT2uHqceXVjox25aME0x5p1vCJLJ+1fuBCWsXfqqlFdGKrIcPSsC5JYbWO7N
SvxMECVmeBo0afMNZbKd4yeKlzwl6tA3IFxnDOesVbZKhDiPxNIE9EHJHHksU5FL
1Xwk+xfywXEmFy9KzjXH5MJJk0D+j5EbZVRVbSSk2Jw4qGwtLFFO62OsewaZ+i6y
3CBP5SN2FpA0BzqxAGfQP0P1a6bI36blSEf9k/JEdoiS7+vK1sw/wODDw60SUOIP
fI1mEut1EW15w2yGaiLaTgegsZHGS8z/3H55TeqDMBhR97M0dZPaGx9QvDB1Fcpo
uoJp4+hCi5hVR8Wc5dxhY8Rx4OThpOS+6FIAur10fKh4Fzx6qjHMKlsT7ZU7H/V2
ggcvMrav65FnRjXVYuD6bl/rRsOPxjhoNUsMK5qtvu4GSC7L1mct1eDRY5fTrwS4
ppJjbBoS2XnFj9fPsfI1kffb31hqu3oxKOEvJWX0hLTb+qyu+aioOLmpftemt1b9
WqIqdmP66DksKOfBE1fK7Ch6XWzWXeXnkwT9d6GKOnRbQTXuS4BIbe6RsawbuZ/S
Dw/PNFjG6iwBDK27UtcMnO7xQneGme5qxNNudX1LDQ1DfGAxeumgvpWGk4C+KfZv
ZL6JUR9DWkhRctEX2PlU1XEzLRzfncvsH8nQxgcqgEpOCBdqI++LqAHGS2i3mODf
zpCPQfxRnwYbvVKzyZzh2urnhHgyu3nOdGOK/K1OP3XnfSrCPCvrI+f4q6euBVnx
XqUDDpA5G5Ky5vCLU/k3yNegVjWMFv5BFoXSm8Nty40iKspOoyeKNwBu61m2pJ94
y+braZhvE88NQ+Z3S5VWok0wtVBhm7PyIb/OcCcrHMZVq+g0gfUdJSnHb99613pz
GW4+Za2K3wEmmxk7llG3H4S2mKjmu6NU4bi4XvTwv3NeSRGRl0/4SRHtFI5owwnS
iSxjd4hoSG8326mNopui/jz7OYiZUZgkhAlJU0CNWxmN/wOGZR3qVIlWDqNer3Ya
bvXLygf5HnN0jxQtU+BaoLAUAuNCI0MxOd17WG2cOxG2FJNMirG6sdMyJfGcBLy+
9cPmAkk9rAfm1oj9Bt9HMjL3MTms6E0dYMTaI7R0fjbwBxt/MUur8YnaHw2npcDz
2XubXkibBBQqU3jMjN8XgDCENLaymltevmjRki+/lITcZHKtWpiYn3d2YErKqgZb
FWs9d7hqFOPU7XgHiVTltDP/3ucLwxUsNbunA0PTEH9M+yk9VR61d1h6RU/s+22F
nk7HVNDkp+QyvX6fcW/ErSQvIsTcW6ZZRYDxLGS0lfEJWjOBotOuOhpTu0Rpxu/i
5e1O+wCuN6814QutFS+ln6QoN6JSa3ETiuKFayzxGZF2WitUkYuf7kDrKvzdMkzC
m9BjVUEa63xRu+169+yrim5KN5rTVc2Zd8dABQRelXb/GbxnZ52Gi/z82vr7K1vj
b+pTQLkGzX+V7NP3lENQ59Sikhj8EVkfy4KFxKJtd95CJEttjnfWW94Qhwyoeyj0
iNACf/Jw97EFplfob7z/VCYynfGMm5kamrfIQ2UjBIJWsuQqMdN+PL9DgOKw39hu
8LpE4Src6tuZ9WOABIBE1lmVRYMvU95P01Gqu3W0ZHNxSod01+SR51BFVpAmmh3N
8NHZ2T2ge/H4U3ZvQ0dkaeiuDd35/POz4nDHgraLEMIxv62uJZr9tEtoZDqKAl3A
RPqT6+O3TBZJOCnW1En3FyCj6XCCYGSxsxyztR+mTLp0c/yIysWi7LE+CExZ9Mtu
V2B4iNyVoP4IEoNTUq3Cz6bi44r8AblFunM2fjRnoNsSUNKZEr6GjUD6d5aj5v8+
IRuq3YPM/1Cu0w4r6xC1aUb9+0hf7deL45n1O7IsCKM8Wk+Sbv+7AOmU8xR4MGUI
sO+OoJiZu41OqyPe0a3uSTw6LReBXIBzvpN5YnL4elOByp8L2bzpiRy+Rx7DWG6l
fCc198UPJ5c1rb5OWzTz8E9VMrzQi1H37Q3lW8qTh9bidzYwPPGwiuFAOrZ2hjZV
oKXrdYonLiR4mcXMlThMoDPpdtbnEhAg64KxxzRBWo8+We65QdLAI39Mt0ztI1eH
HmbWfVh3mrb2tXL0eycqmvHHzzJaSzhy4UAKx2t/YEQZgYSUL/eT23MPBRpI8Lse
Xlw2fDFgnAbrqoPc3CSlSCIAzQRo1+yVktglk/pqrnDw7OLsD5ikManBlztNCh8s
lguEcZ3ryzqq2q+Ea+hcgzTK7VQvUGoHn+0r+CCR+k856E3+rA8Cx/lWTMMlG9re
CvkoJfx4vzlbInGEz9i3VoY0NiwcVfeeGkj7dabuHi56mk0tfMuRmHuYjghPoym+
2T39O3YoqxX8vxIj0zr2ojUaiYcch/5kB88qTq6ZacwVomYydPQ9SEJ+U2TyigBz
q7SATC7Oyq/UKgwuUxq8cE2bBnLkuluE5qhSAmcEqPt0N6rTcWB47MJuLaTOIBX8
lkgRw0IzbFvbFUOgJnPw6LQ99Gdabi/F2MJzPtVv7buWGMKzNn19nzc5ANNSON83
ZbrUlP8xcDvU9b1Y9x3NgURXeHFxDtffwo8X62G+x7JpQqfXGccaLqa3BVz0LnXz
R8BtQp32+M/anpvPbgekibyVbI3fJ00a8RbJyOjd/3BAOPh1Da3KhlwM3tX+2IRE
lxx9doe3KCNvTDUhVAcMIB9zfQbGknlszzZp+1UAVq8da9fkm2aG3bk8luRSYq+G
a58czkKVS6Hqh/jCzkh7MYGTVtYjqS7S9pq7J9PPkzcAI3/EwLDAYKzLnAUGVE23
LogNyHCk+Jvf+v7nlLGpg4eIJW9kLYQKzDmWRYH18QEnigUImSNo7ze1K01EguHG
Q6lmODp1LQaZ8HiuYPVpShZ8hPres6u0vAfqrTi9PeMOvAiXtK0B4VYYvEhTiq23
RFjbNEZajIzCCtZX5jYzC1Bp/YL9AiLCgBi0w5BQpDsDkmoJ14a17CIPTADA2FFd
YS1UuJO5j6fOVbpLJOrt/iNynU7SNH9Ispb8g3nZMuTZbtlAONNcqcg2oZYRjAJS
CkqHcagHI6y+zqkki84H299IM3EcDOAp0TvZ/oQAO1YhF8f7iJWLRNwf090ndWzN
qVaDJ3d4pEwxTHQaCaHyoMX/RlQlfn6TsvE3liT+5G9fnQ/ncJ8jtFA6JNipHmgk
b/QHu/JBxFXg6tZr+VsiwaxZ/dblV6nR6VcBUbmOMCZQazA1ZfHp5si11Wm/UMcY
agId0nllehkzZPpfRIglHjadsXBrFJac9PSN6d6RCZvjJx423/EGoHD57X15cm4C
Ez319L08kSMghwtQ7BVTR6qy7OMgcMPo97Fda7Xryt7iPzawqFws6fBVk2yNAhir
NF0rxlOjzGpXiIga/qzL1+lCWEjRQD05/yP7nLMqWsXKV7goX7AoooZxPajcZRc2
1AoCh4/NFCzVAJjSiHJZJwLOhMu0W6SRQKN/peFJePZ80LCtV1gB7DroAIDizcG8
Dev0G/etqdY6n29eaftm1be+M1hW3rGjHEfCFVbSQ3Mx1aFD8hvJkX4Cv4ClT4EO
whWWsiy1JIs1tYx5PuQaTXx60aUlGUW/RPAvHFc1cZlnIzIvLCx3VH+Yp+48Kc6k
f7NLND/iPof/2yYcExlK4h8McmN21poZot91QDYMHydZ8N0J26VVEpsA4W+ermDA
SvZJYgx8PbHTQ/LoRJlasJJqoNPn7SmJaBqzK/1xpRfM4R9xF0JPcZY3W04I4ZyM
G1jPpk64EqcYHv4PsnFlliGPZ1jwZ8/ztwnAjZff3SGGdFnE+5ejitucEI8W10MX
X3O6ISBkJcdGUy3svw3mHte2vwhOK43mYErW4uxshzz6Zo2IMhsRxNb2fhzGTMuy
b/DAo9tCewK5Or+JT8RcngyMFwmyGa+EJAj96sIpcft0A3GwZ2AUcIFdHYzXq6gK
CrtSr3yuxo2kLGkicfFEGC7avYRny5vlCAkh7BhaERxPEJ3nXtNiIqhCRVsN1oPV
etLBi/HhkexwlNugHkDppXhRgmpvL3BbYaexRW4tTvkgB2UrAm0r4e2YI4QTDABZ
PEPK0/3le7xsQIOChdjdFMyJpvWmFar2axGFp5MXLPY9UU1HMUtKoVK+54xf3Gpn
Aqrdz8/OYDY0wVudJYKGjIpNcGNka50DF2+RgLdsdsZce1sMs300TxN46kpWdbHH
txK1rBP5dA/kIMuiAat4QN1gfUHvojVdPoK0qCL1BEqfjqJdg4JufDnSTDWvvqv0
s4Vs9ezF1I1ThHaK+mrFVbOhP/zdPMSiqTw9kLZg+BSCLkKd+/F2vj8twVODE/MQ
5bc1bLNzl91iOGyNbezaQoFV+PK2A134ytpVbolRoadGBEwjxJsr/CMFublc1jOR
6nxnnsCFvhRM9ujS/iUPImqZETK1fjJkHVk5XWcnGUlXz82f2WTc+xN1VLsMT0lx
gi44NoP5Y0bDrrx+UMUOEx7WA+yT2WFX295unmCPVEw4bPtQvusTeedTBY7icai0
+eQBN7b9Jkkjm/IbYFq0SYfr5HYX8FIMn3rtMcs2MYZHt97goeA2XTspsufDllZT
qFV2JhwlA/C+1QWfsLw446eaSvQ9kGuhMG8xs5fXiwTnqIqLS6G/ur7LART+RYoP
GCahds+3lzkAXm+X1wNWYyGfGxjnggunvDPxjsBX2GtOvmI+DCqDoMcsxYzZBPJa
PhT+C5wO/Dyy8vuc5QVArQw4ThM4+gagvKoitfN5ly+5MT5JqHr+GAbJyyL/pGOu
0tNWPJcYMonGTjBPyP9f2YwsEZGpyScXAGCmEgfS1wVvHDFOWrxfgQ48MA3jm0oL
8wX2rTZPp0yqopyzqcK1gTDfmT7vDvG6DOHmComVN5YdN91cQ4/KVCvi0JDL7ajJ
FUbLfcBLKcaQgQEx7RVOLNHOr8Q/NQ1DDRN4vc8DtY2GseR+tCOFkytCtn65aMlC
+Cn6CkNzZ7TskYmLjmxb7j5ddqCg9Ged4Gwjmi0rfKawPNB3ehEiYWuv+YaLH3A3
RyFJFjoFVuqqrT+2rLbDSTc64jtWityttyY3sjVUniQ40ZBJx5yKNGOmLlHNTIT2
fP9UuVBMq3B6l4rNAvF9Qa4RR2sRcCt+87SjB2AaLOHZxQ4G80r4e+2oWeQ+sO+R
PGjQW+3/44PpCXKiGZyrOw11hvpiUTh3i9WwFAwCBvAD/ISLIyW+m9gkw+hCJsez
LhqiW/lpz3ygogiVjkcfv1zEkyLUObq3uncDB5k6u1pxF2x9lVCQlCUJzHaEwszs
gwVqiJf6wzzjEfqqboMDuJ7BbC0iFYVdPyRdUrBtdSfdSqCVNMkV6Kj/7dpawzIw
LQiMRzayiUYY4N1t7iicuDxf2vVCH87EPPQ/vbsRbJH9XqJIYZu/+n5i9KjmFulT
582j4SnjPPfswIXO5hNcPPyqt4GYaKfgogNy+PG3+Kso1PRlIRTs7Zj0XpdW1qIk
3p+nOgfcNJV+eJYeaJmO9gjp1zMnDiImengSsWRHRk6ZG4M7csQU+0QT6OYpsGjx
gNHYuOoBJYwN8fnEWkgSVzvVM/5bW/DNivnZY9IbowtuePbP8yOJe5Fr76/qhVkH
FK+2pzXqp1llwh8GSlwiXB9PdKQIWhR9Ew7eG5e/KQWRu/hcH5J9ATybjFybvG4j
8z1PLvkBkdjMFgtGmrIv4QafU1zbmb4i8cV67GQCZxoIOP12xredHW6MgzFyBeWi
dSvI6T7k/IMvLJqllcIdlcq3vkOoUAjhHGj2wCBK0nu/vCZ8nzILaGPdyB34Jp2R
GP83GZzqsn3P0oak+NSpO6uLWYCfTxXxjbxGVZKVIhlOftwrKn3N7qPYyDMxsZ89
L0eJ1wU8mtozQ3ZwJiB5MF4sL3M9rNVItvmrzBIYT2dqCo2JARbyDEKRrF5yH2ph
aubCle+VCJe/bczDAv+VLP8pcIo3vbrRF8JsCHuphoWHc3KIhJ0pheqZuV1WhKp7
oa3CD7XW7yRGwVmL+u1DZmAPvhNIAOiuezVBPWOjX1fT7iaJ0gC7GvOWVbOis6c0
OIHmLwvcCGumi7qQZSg8b+LGY/G77cEJizHcR4hrpZZMmfkrEUs6POIZpqsumkKE
5o5UYhXuT5OlZPsqGA7KKEBtU3LujdMTuqutKyMHtZ0Gy+n7phOS+uB30gL+eC2F
ucYOel/Onvlrmf8fJnYGelFRw0a0cMTmLVK/8wQQyznqxj9GP2NR/FVMd3dfx1uL
IWf+hFusxxXren3g6h0RvgPbkeQeBoMSePgjL6KtQ3vX+jBOKjbbQaF09zvyhYLp
U+GeCG6R19aT/maUnY6Md42x/UfyldkLtzfUSzo03z620mmtSY/DL3vFPU5gZuPH
e+x5f4RErG7X4vt+ocyhFuWSNmv+nG784RwT9y5a08YLsfDRpOHBVoB99vpdY968
MeaLbffQehgaFq4CLg9Gb+rmtRaWcxiI1BQoF6ljLVdtj3P40PywGoOdpm4FypwU
51hLD4pRZNZN5GcDIRVj/Xy/7kRnpSI5FH9Ij/X3enNXxUZSm+h6bNzlcJqwwE3g
4I3AhwdgXeiaPU1JXwfGYoNqHbznqRRijAKA/hFRmTlxkrm4doBiZzmYs0wu7A+i
LQWlgLJapf8E5cGlFf2vRgD3nuGwSdEAmNds0Kwkb1OjsfDMeukdUALH5YhifjLS
t1cP6yPPCW1oK8D5J6QcoLSbsROCop7B6pM6F5vj8bHL39f2tukKpraMJDh89hjJ
/OL/1wd7s/xWp2o2lCUfMMqN27KyBvdP+Hhzv3cfDXziM0urDMbFW6IZxbXm8nM1
X/DM2afXPq+fS8y58PBz5sPyLltexPfVSO6Krt9hMK5wUX3ZXWxqUMuA3FyC7aiq
Wk+F6LvRRjaPPVwC1fd892G51GgHhrT0UBXTNaeGTYYxtWRd5de3Q+8AyWPho9lN
kB6l1y6RlYqp0ec3SG7v4rfxGUsNlUgqPeyoNAbtMSYYV02xFPkBSIDaxU6ivH1y
+5liqth/E5wA7+z8rY7RIkxWuKgYF60H9iP18GSKDuYVblRRjwSyhzkzvCHxbQZu
jcXPGz2YjtTkaquuyNRiPC3UMTXUXe+gmLe0lc90KNjt9G3qGNSc1QZvPmcBIMDu
iXseLkqrma5EFEFpvbLEF2Mve8ksNvUZ7AwyqXTAfvHAi6JJrHCiA3BCFMrJLjLd
nfl4IY5YzRroOvM4kAyXTIEBBBZynN6atZKoFi4zpILGTXfQJ2nCinnQQP536jXI
h4IgMBKbQN4FBRt2k8uDG4AqkRlUQJC96SeUMnVr8ysmiSFaykhkyzDr0UtSRYyu
YzXQEhuCSRi0JOdjUcP+7zG3jngdDUj+pilxNoyJh3B9xZ3eGSf/a2Lp4Fw4fGsy
ZBfSf9lXsAbvUBSriwCh2bPWnk6yV7H1q2+e/50dthnXhp2BlteSdovWcQk4Lkkl
BRRY5BgwMSJkv4P8yqa3uOrzSQwzMWIBtN6sQ+htDIcsNHrEcSfzQmy2g8VXIHSc
QBSOvSLISPNlpQv4RlI0txtf3iiRmhPoJ9H1IWDCGOj6g4RB1CbzcZDF6P3KtYWb
vMZxUi54vIvGwk+ThJnRdkTjnANdtzScUga7Fw27nZjlyR1sNs90/xOHoJ4Cm9Im
Cv2AuW4ALNDgieqCNLeaNSPUuyOyQUAhVNojjHvmLHGJIWwzWRwD76hzXLJ6cXG1
E0PfKjSvTx/alL7KG00UbL61IGH7Ttqz0ilMEQeycF9yW/A82e29z5UcNFWgGfuN
ce2OuVqg1UHW8sSYQ/oqyt7xs4uqq9ecBCImgXZui/sA83IkSKq6v4dd9z1lMwA4
pvxQDXUDDFaPZSNS3OtZwHRT8gI1sErxCWdnsuiZlsh1xGrLF0FxHJ3oCXpDN0hm
29r0OtFQSTN/DgciULksD4tuCQfrN1spxKEaRBsWtbDJ2q4StSD7ARsssQhSY2Su
Gvwqwt4jeWdKY7/ZnmOyP92LIOzReiWdSP4PlV6l910bIOgWm37uLOWjeP4706JA
WFHvitmoMNSxhRX4bFTv+pKcHyYlX7yAn3PO48aHgUcRM9o5wjdJBc3m7QvXiqFU
KTbT03lirf0xN5lUj85gxRmm293DcnBrpQ+NZ9PqLur9D96o1BIch+eIRrSS4c9X
Rap/L4Z4xJnW3dU29IypFJCjN3XSu4oyvTTEjAdazSI1FGH9pgjavShq2SEtrrHi
2nwerAv3UNbgCOr6qEleE3OchmsFO3/lpff59f3LeD9L60s9lhjfMDb64lJJ7foY
43X4zNx5pLS9iC25yudZiJDyMfrr6salNiUN4VS4Ai+dXQ6eLy3TWmNSS9UfkUdL
g/GWvGKKnvjf8majNf3FQ+r8YjlYnDHDx3ASqUKDFeUn68gYftrmdcAe4q5ZxSnE
gefG2wsUaXIxEw0ttfa6Wy+kFS5Q/tLhCsgXImoluauHweeWZRef5IHL5PJV61xt
B59seJWDTzqbUEglvkjTofZostqpA3QZgIoTDly8o328hWop6SKOe8g6QeKe1yZS
6KWOAd7bKKqqMPWdRpHfGhCsHHE929doLbHkqf3NJMon74KOvfL1Ep1qX/2eVLkY
LT5SvTnyQA/FAzJYYmHYf4HKtZvr9v+kr4pbDOCl7wjX8AnrJO91krjB01JPpp+b
41YVbNacq8NaXLn5famEUrAtq1QC4FTgtHZAU/FEaOMpQA+I4gMaqkJ5VfofoWFg
tFWUZffPIdOfLIneGMoFCWTH5qfCd2LgMZ+DT6tb7EHVFROPOKR5ATArVmghasno
ahAesZgg1+QSGQ4D4groI7r9U2E01qJSvmTEtFd3Gec+zppYiLee4eklWsL2bt9K
7CIYgIyCXbSgw+XaHH3kCevXHXsgBtLcF8kFhexd0l4B05FYFELQel0Tx7F1dPeF
TRNMrhkXua0viHb2hP6tSEUqhqpK6KxWSdH9Sl+pXtolK6msg4Ax9Iut32gUKatI
QwHJisIOwK/mEvwto8YsDIOtgVKONCBCulDInlYdOujkPVIFfUedsosG3L99/CRl
U7guVyGMcTvCNf/Yn/Ner1fypEqA5yqFtl9f3djq8MCATFxFuW9Lt/9humOQAQJs
on6vLQZE2ar3GywPdLbVywXqpnUiczZWCitZbbrcXx3g2bj5XW3pILMdvzNSVy0E
ToYAa6QLE5pKyMzbTuukSSab5DviWh1ouWZFLxGGqpJQ2NJ17KYbdjqmjDeLIJ3c
xarDT3CKkOQd47/RI3vMKVfaJlURqRN2JYa+Vi9iQYi1g0VFY3fv7Gi6tOtWQFc0
ip1t9UW/IrWIgai6y6RtFtNjEXwGVRZFfjSWTpRGON5UopOVECR4O4n/oF5lPFR/
X1Tc9XcdLVaf8nnCdzkEcvBMh0AfMxv4nPYWzqV6hkv93EJVw7/oW6KK8w6ycMeN
0nK7D5rt9C5oGTNeirTRuifF9we4UQ8Agb3os/nXPTB4kboWLazMuN+dcWPTtY31
vwvr5YV2Qm6fyjOC6WisbuEYSb4zcI7TDGOKE0Cxx6y9lE/5eLcr+PtEMEtWxM6s
Bgj9hYQp/KIaDS8t4UeEkjF6hjaFBRAPQjgsDCOc4eVaWhioIqZ6cv03TvhoVxXU
xMcBKcM9xNP3rGOS1LP4WMprUN6Cx8D7J3HfuTB1LDDLOPakjNmhYZ+yX1PSNWRw
xVqcOgTF0dLQFNr8b7eXl1N+lJJ15v1k/J0UnyfClt54bM9S5PqfDO0YGMkBzyQC
mPqSQ7IfkKC2v726OaIlVINBIRWURi6Nc9VnYx7L7lqLzK0O27t9TAzeTwu3kRTz
KNEQr0LhxlJjD4rAkF4OUARHpU+TMFW0JhSGFl7PVR9dnyQyoaS4dD1bJfzL9Gvx
N38o++dk02i/5iB9eY4Mn3/S4bv7tkM0vMTBJfvRPlxnbafrT2NeP369A/QL6kqa
jsH5JvJMro5c5sq4dxtzAVz6DK+PbLDIc4TnhxTIOdgii8Dx/GsSV2GvlQ/ynarj
GEiPevA/kduZdEKzSwC7nhCANOagWhgNfUzOG5azV/OOzHCCSq81acWiMAc2ViFu
EtqtKupwK+hG84vG5PrHQZ7hE2/U+PKt7NJ0YwkEL8eVDOhBoGm7ioPYE48FHDVT
yZM1BNSbwFz/z5C1xOKy5tJbR2rmkedlv7+Woh3M9kjKmEDEmOqZg5Tl0spHIcGU
Uq7JTv2z9Ek0+vayKNn1Oi6WAWBYPwB0huI8ifF/OUcmUYttwQCZNO4xu6mjWLBs
YudymMIiqiFnZGjNA/ibDfJL7KzDSfTvZDsFdE/R5h8jrCNbUdWtpIouchY2enXE
8EGEeC/OVsk4mLdWJUgoYl5lgopNzasEuQUa7WkPJ6dqlb2DvgempYVQUsi8kHhf
aGHmZ0o1C2MAUJxBuzxeFPCzRpDEXGUzb3PPoc2zgqpmiP1m2PibkrKroDqZ0PVb
/pdGJyoQzA6vzoBWYfTa1MEDkuW40EV2gFRENbRwqZfeqT3MyG+D5ahbrweCp9V/
suWIfzKXlNsDx9BAJ8mPlT1WuGfULcWBdSyqJtKlHmI4q0H4KcDAQEzCy2FQTSAs
pQa7T74WzTq//66su+VSovqORcI2aI9jE7JN7L/VjnxwsW9oJIr2TAaNzTo2ZB4n
ah3z+XR//Cp69MeCm26ZLXColTHghSsVgrhvMgO8FSiS8rlnt57LW5yXcc95gGLP
Uw/Z4Dubwq46CyOmWWTYWKECvOE/N1T5FnbMxn+u3uyTQb0PRp6bvZk2AcQnMyDO
bJI3vT/W4L83ag+YkrWTADE0x1/m5muq/tP5w2YMcDDgok7D7NkEXTJ+wUMRo6S2
kzDePjNCQXUUOozDrtHqEEmfD3OOZynnjoXlhDal+TWqxM9vYP7fS3dyikKYBtJe
jZV/tA31+8xEkIBQwwp14A9wfllzV6Ev+GDZy3OmjaEezBLE412ns+WzYRmmcjWj
+lMn2JzAjeVeUHW7U6Yswh+KBZEUle2ukVyvNdaECiD62StS1/rx/2ixDZ+bc2Fj
gvqEtEpb1ZW89H2FsQyKfbnX+XMj2dFJKhUQKJDm2nv+Jxvt5QyuRvLvZ1qmtHyK
xF2xE0uS50vrxAJrUTO8gSxcSPqIf6pXJEvtXMIKUQxunQxV31wqHbhsyAR3NUV8
YFajE+B9I0fTe5lWUgaF1srXyeQrft3Scle6rkH8CtlxOir2tO9iJ1bJa9XYEQAS
C/u27VguF87c5nPn2Dt1/BjEa02Y5C+RT2C4jVkmCTiGjbh48PLZzWYDXLw0KLR/
cOmdbyzP/vo6YH7bf1gwtdLwvZtA30J2Mo7zLZiFo9zQY652NUI5lcg5zWuh74mX
oS+vWPKwZUQMz6NGFRDg+9iiRZV+VBg/72LqbohQbAmYTfyLvuRIU81e+14k6ix+
pWl2IPLtTJgdsg9kYsbaSzHZmcFgFcwMxCTNfR5Li+ZDS5wqoingUGxB9MkecTMI
KKvfq9cE0Tb+STjRFSkE17gLTQupULBMnZSccXE4dAvVGMU6AgF7Y4SflYcTFAjT
L2zH5vU3oCzLFH9dOEGsAymBK7qrCNarF61GltadqrXzlQF2k/JA1cfBsMPcK57Y
4+egbbcJMcTrdC7hH2JFm8uKBK9aCX3/LAk1LBobB2gqDsduezBg8oV4h8ct8kGh
MtiWcbPJb/yPaZTvTbtAwBYkwrQgKqpOcZwGIuDNeJ75hyDmxJvhq+nnMP0a85Un
QJTJEGxYNOn0xtnkB/MsOSWEkcoRHSgOBM7FgA+8aP1jtKHgkf42xmAPdRTVR/X/
vHveGL/wE9lgN3CQx/DaY5i9ODK/mmC18bBXfDdNyusTFGyTjbbpTGUly5dTLbCV
O82Fe87nCqUAkbCpnLdSOhdwLBN/Zf+zDbj9h1HNgrbuBrCyABuNrKJSRsEeclFI
q6k8wWihuSzotxR9ORU8hNhxCVxuagayUEwMSf+wgAw4PdSHKh1WClXY6n6wyM+Y
JsfpV4rivuLKb/5sBhMrK6n0VY+weQJ9bCh0fn2G2gugmUQg+r/aL97wftyzngN2
hNmpBl8O0JcKYfgTz4GcVGE43X+11kCBC13rIQsL2QRtrZdGjWHjqED2JPsvKrOV
f2gw1GN6Cc7abffye3T/tWGYDBK0EPVySZvTjTggGC/OkZoO+xMes4WiwrrTbJdn
413NRWGKV4843r2C0WBvqFENy0d/0U3za8oGQf4u6xc+dD12C3bUvuO+Jnw3P8vX
6sjZru4fB4GYIzqJuDtqZnO0M9m8WxUWXoDBSh95Xpd98lKwj+Fintj5OGiyfnLm
Ff2BvLqbqABgjXmXNm3/wDUtjvWgQEwyYTpjvZmzQIybKvvwYkt+qkPJo7dmhnYP
XzlmajBvZY5rUOTUYTJNK8IpDv7HB/QUxDqmEuxcoo/iDd5SPQCdJ6fe/iw7IcCE
JDyDX04Fz4BVsudydzoDAeB4Ubmfv6zg8RxA5syeGXdCAB+yrS1AgIh6+wYdKYeA
XMtd2gZMH2fH0KRIpdK2FSabHudkpCdrr1m3Pi5tG8NtJnL4m6iW6uZSkzFIpfRd
kZ9p/UhwXd60HogyoDqIHTOM4mAnPyPUbUIaH0r15fPJEJ0VncDEK18qU4YoEfQR
4cZWnK9Ra492+agpZ5TZQfxEB0EMfJQyTD7R/Q29Z9mbpT4znmW+Q0U9cPxc7Eoj
mtzMjN8CJUB4sC32Z+jthWgW994V1uWBIDAy12jJXNDKOI91DeOkAODib0J9pH4r
mWsvkXhT7XMejp8F1Pa+pIQK1VuiFd8K6Jl34w0aNpc5Wn9Sm3dAdA+W7QvkvBLF
AfnhxVBxBnIK+bkp8saGHEBxFZDXWfZMCfO00NvNBFKbXfGodIkvzPa/VWLNjadS
kBS30d9aZHwe92iWScAweevD0cvMhZGjRuvfmBxb4MhI9O4YP08PSGotvs4OTJo6
qxSnQ3GmphaB4IJTO7sQD6WF/UcdfwnJEzXfZLF0dafdRuobh23T8GJZqcOAT3v7
K8MEoasXYNSKLiC9BfEKdqwx2v7qCdiUK9wXipN+sZMObPzRcCBgX42Usl6lQ2Uv
CFDhr0AKVRtCmYCVw6DIc6z4WUFGi7jNJ/wcmdOWwCdDumSBVvj0v5yTJrfzc4BC
seRoEXvYv/ZECHU33zIomxI3knMITBDEr4MeVF5GP6l94m8W+Xvz0oQjqTwSCLdg
NDJ7mUkV0CpviGwziXe8QblYLpnpPQ9lU+QOkNLDhj7qC3ewesrguNBVwA6hpuVq
En+x3OVVXgN+kS0ygEkQ4Ex7GxJAmJVF6xDv87PR0VL1mXt6qosczYuHHoZl++WA
cZIUlyni9qWT18n+sFpPKvwzz4vWarlScilKIhfsPxI4h3aOZRdA1ZZ0xCrm+wuX
uq8vuKXLc7nhh04s/+hFwuyjpXf+HgZ8ZalDCbw0yRS+087c94iMwoj7Kvyqvc4x
RC+tkpvkLJiRHXpVCKMlYiqWbkcb8o+8lsM+4nXlZDAjMml3RJjlHablhVlD8Zkj
YX3rRKpiwLnyksyqdcFpFLNf+jEFxGxjJFQhe0uT7+uvDqtKH4Kcw4woO6SjFB87
rVIQ2l+4ICTs7rbjkeXR//ielVqLV/5SSrinH/+N59RBKlbijccaxlGDNMFOjgPb
jfOhoS2mK492GBwc4OyVLdIgaJzENbUCXoo3FzGtslsYuO7MHS2h0qtOctnuhjD4
ZFfWC7O+FZRKB/Z8QkJ43x1fDNS8UPt0MGuqB25ZbFJcVLJ9cfEr+Rek5pgJ6Ytn
vmAqKoR/6wifg9BaYqW3IlNJcrhUeQgsGUzdggPywLzA47/SSW3/pw7sa+PEFDcQ
jGWXZA3TxlJ35E/lCFnnUdIhxeJGi9+0vgRyz4bs55L0C8LOCJDGdmlSf8Bc1e/T
DR5yHKL9z+8/+TZHrA1+EcFyIcwYSlycVlgVVKzsaH1eydDZrEOBEt0REEm6lVwX
PubyRu0qm9CLQPZJF+dthXKiZKt5TDCfaxQTZxgHF4SvYPwaJaEUgSpy7SJg1AOJ
ev5UL9FWZTkSwCj6hL1tESSON5pzLogwwT8NSI5oFgnWJ9jqR7WnLN0fClfwax9q
GvM6AF0ezTdolRH8bdoHNXTLnnvoTCqGz4cyqN0b7oidQOn2B/XtpeoBUFNsKePy
vYHEDdOs0AARogVQExTNHmVjfdBKiU17mjU9HttXhmv2HMlT7J+KWqLHs4RjSShn
mqck1+cPPHHB6ZymEwicB/f/Y1oQPFvmKGjWn7KPbdRRCgGg3ww1F5ub2q/2D/Qa
zVYXK5TCrS3DqhCAmSLi8hdo8KdX0FnMcg1D8jor6pvqlbqLD/pD1eff68HtU/NL
zjyhsI71r0ydQdUG4PDJnLIT8+Vw+tJoNNbQN98Fs70n/vHcTjxXHFFCTGd2BkIX
PlkffkRKDi+MAMAPhgVjsoFJmLv0S1ovHsLYkjN5aeD3AapH4REmuCGWSyw1BYEF
L+KNq1WC+otFn4SgTZahINEdaA5q14fu2/Pk/wV4gtd8hoJJXIRRDbsp9N7Yhp0k
ZH0cgOR57c74arGX2ujGKX2wmmDexm9GD4JVOPkjGolm6XXphc1S3BPn/2ov+4t0
TLeQ3CGpfoRNFjCZtT+F3A/vsGqGgKSsH4P4JTioG680OaUWb4aZQHm7MeK+aFh7
iBn2A6hoVTywKZ3/8LEYpHwmL8a37uAQX4IOGzUqIrIW9QRHQbtmitDSeqSsInij
JkZk2/SLqWF26MOVfEcNtFoeQp0Xu13NgcMjP+K5HxsVgugB9ZBkFfW1yeAVPzqT
cz2730TID3ea9Rvn1SPdJ+C2CnM0m2PUPI/A1iiEaFBznBMTCHvEpAbn3lHvlQcL
dBjVhy5GZwY5TGJ53zSPGeDDew9kwPxJMCm5pf4MbmLU83/tMiBar44nXODb1w5n
tTc4zZ4uMPPhPsJ2A/o8qaYu7v5dAed5PIWikA9H4pAdd1XBaCESk4C5pAJAjIdu
XjK3ibXJc9WijvU78Jlf08yliGAmQTz3KCgPxJS1OT8lxP6CvUaF9YHhpdgBzwlQ
KEIiG+BcgyGxZEiUypH8Fwg5g6LuqiYmVAhz+Fl5ndzVmWLdBoJhzEyjvrOaMiE0
ZsBOoLI8hUOqf2RTDGroTqtE87zxSOqZTEiaujuCz1tNwE4ZKrSUQm3ErbjILyuo
rFFo2ylxatPEGax5WHnas/Nud1UlKJjcd/KKC5+kH1aoNci/Beybv2UHFpr0654a
YRDoG/XJ0XtKyBRk/mJdxGlktw6D8rI5SGMICE0S6QXVO1eyd3TgU1RE8sh/6XrS
iSNqjTtE0ZnP1VoUIvbODTm1ryaPu++pdiWFKyL4UCEZWqJaeKEQT1zWem0xs5At
0K9hqxvPGwX0u+okxqUHsiDSmxh/Dv+/38a0KeFDj1j46W9w/hcyDjRwtzkZWRs1
rVGVCTos5NEYqTbafvUGGb8u6y8QPKIzpsZkkohMOpniT+/UdSLtsGSemIVHVLHU
MwM5BeKJiUAKAlXtSZrBAglfR6c56byVBc/65fAfB2GJRwnoYC6prM2drfVltiIG
cwMCH5Ya+DGTdwSWy30yJ7KbWM8MPGgt1ISkP9K8JmeWPe46t4VZ/gz/k9XsmLjp
f1ViKqSVhVGqpazwTgiqfGL6/5hnzGtu2ql9wDmKZgUDyMLMTR4lnMTZNNcSXb/W
TbEEr/gFQGYo2uNSpTNzZefyiN0gYOl/pN6HY/bbEAhqT5BHIotIbGs4q241G/KN
wjxj1CKpdRIPzKWrOtR6WjG2cqL1OOdyIURkCfea3fAZaEDfUBb2QKh2HElmtDwZ
9nagpb0DF1L+n+LV8cKvwjxWXzYwDxk6o6bzNiHP80/Q+rAqQYbKYswbklpXlNdl
pKIj9Z8U2fqqzvRn2VulGGJwNhK951v7okwCE4ACagP1x+lWUQcRVwl3faqu/wEG
svER4jtqNW5z44AVQwnB4+4J+NKYaR8utRfnwPZp/5TVjNEF5rtkzjPMYWV4lquF
ijn6Hnrx9HPw1pOfCEmzEAivAemaSS2Uw4mOgfmRTRHiRM3zJTgv+pd6LZNe1eWf
vwT+wSUHIKXYbS7poxPw0pQwfa4VTOsT7hukP6FiUyYnIiuXfjGEDiThQeDdOloV
W3R3/NeCKF8vGVqcIC+ZW9pbgxUoQZszrD68RTNgOftPQo7yysjUW8si0mos58b6
mBKYPPXd5tqFnbtRI4+VY+WLUNlcU7ZlmKYldU4ytOtHkxxelmPpotxpGqiBAnut
BMUziUuQS11MdhOe2e4uKts40S/BRgOc3GIpMLlNZ+NFghPsqLCx3rQfU+5oZdJ6
/rHqAN1FEdWE5GtaWsWyiIyk/MnZtP95dkE7snPMBfRCEzDwEl1a7j+ZUPjPvBAn
z5EUVKK3ZRcjd3gf7eP4lVBAK4vrpeGeunn2/Np0/CV8f6RTxpM4OkjJpbMcoKdd
5zxqoj37WBo1m2j+gDIEifOqE11IV1rz7y9RV3q9VgoVa/+ATkWVyfgurRfL0HE3
URrLZpskoDQMzUjVkNgmrV9dz2ygWwgrioIWE5E/qO1gBpDNhzNCs1cig3oP96nP
wLh6cGnZyuTmxvkIFUysTD1BUsnDfcEJHT1I/tqEqTSDi0Hek8fBaEf3o9RKqggz
pYXuO0wMWRZzP9tcP9r29YpkprXD27WCNr0Ne/magM9FpLrAdLi7Bmql4DjHc6j/
M3mEiMeMQ/y2QPh0zXYkkdvwM1E44mFz1EPtDJn5xMXtmyUIPi5hjWXgDMvzLpRX
+qR0vgYBQe5iNVHjaSCFaAhbTi0a8SSPma2TOhpW73V+UFY4p3lNWa/yXdgS99+2
WL2b98jQJhenzknLVEh82MG/FRrfHBkY+yGiujGXx6m+2TrIJ5YfeW5iubNM7NtD
q7tXfKmIBatpGdSZ8rGejeIvQskalxL1FPu3dSS/4KJFhKocPqy8oTI9GXz+lZrw
7ir36KHKjDOvprxIMGHGW6Od7vdtWt6tT87hZ3QlY4V7FyJN8XaBMg8xGEvKZtqd
911zWmSDBdrT2jJaKxuPQc3sNMBUScVgH6pZkuJogzLhw+Qm8XjZb+P+KMlZzgjV
nWFmeozlZKcXNwFeuEkOcfCcbIln6o8u+7bZ5ZxOubVCeViZsxMDvFrLxGjtoCF7
97CJ/Q/x2XPPK8GcwaoJu5eKaG1VrIGZYwzbCBYlkgEaV4oiDHTF9Lf+YZUm3CMu
PWiSX9359eV2WtZqqKPqb3GuZDzUjSO3THLxqCYPZzvBfWzTpaNJY2r+R4up8DJf
McHHun7WIbLHD8qbMcagU3y43GbXkIhbbIBrZEymD3r5GBeG4VgZ6gUdybb1rmqD
b+iqqhThcIZIVo+q+DcDQZS1NLLV+A24RbqTxWvKpQf3wezTe8DixoSd3oMH7Flj
4UO51CWIojTFUlKuDfGuDXUpDahlkI8l/8+aA7kRRoz6qtsbniqHWwsKpzmb0rTI
nEH6jGe+1lzAnG0CcBWRKUOviyp6tzmsDYpWqNp7CQM/YFJGjVzCwJgfBRUgMgTu
CPJfoU7jRLdHeWlpoAx+XODUJruB+NIJhJV+Wb1EHxdkA1D1orZVRNaEQpVEN3XQ
XAGB/88wY4kN8xF3c5HCKCco2CpmOIIyT5EOuGkts1x74OAR18iQQq8rcOVoX3MK
ulLwMCRksDr/j79N9rQYr619Za/AmqrMsMw7Br4TchRZTiYMlxD3G2ZwBru8+boi
h9Kv3HTmqZhzZycjWWnz3+UxgXCL/N+56wBleerlcnx+HTChwx9KbVt52rkIeqCr
iOGDRwWRoszU75BPjkvt17on3lmyeqdIJ33wXfyGv1QHyEE8zOuJVcmL1fKbbrL1
QZBnMoY8vZcQ9Mxmr6Cs5eP11Tj6r2YT8KfGPEc0VTmZ1xlJgdQR/IolOSySSgQ1
8bAuRCNLD/ckt1r7LuHFgB35N2ura3Dfc2qVueNI5saCUdtVCMC7YhtB66XHRfo9
+JKTapIhuHSaAFrce9FNTgladYpIpltYIi+/78sfPrYxv9kjppT5KUx4Zi0GdHUy
R0H0rr/EKJs3fLC048jKGIzGFuWXQ212hQ8U8yCuXn18/bbwpSLwz6ZW1ppexj8h
k99oglK0cNI5BC07iZs7Qwns+YtCBnqgBjVpA5ZVIym3zji2GbTZ+MyWSxEilWxu
28EPTU4m5hf5IgsA8R1/C0DrA2MQXNJxC82Sw6stP3DtqZJ7Y7otLzezUwhcxRfL
r3j4GP4O41NDiuNd2L06Gdv5IkiPAk6Lj6jOX2qXlHuB4mb+RPPfqysPxmXlHdnL
yoHd1J/siQfBhaiD6LD235xTZvCrTtTXuTMlMYYdr645f0by4YYrDeph/IkwE854
t4qjjQ16ujsEeUnpvu6LDWfGLOP+bKTWvrWLyz32Qgt0VzlBrMh6JqhwauQAnRO6
zFQTFRHLtvmA+WomGjAwk1VHZSoWtF/C9BbkzseKqT2DnoRSqNFZwn+ZJPEeBeNt
Htpa4aSmHrbIj9bnrze0PXNGpV+1tehpAHgO5ph1TCE3DAMXilkBiz89pSEvn9Cp
DL6CxzZMiraQvrYwLei0+BAMlRVz3H8J3ItZc9tlwbSv0RK8DUjgTmhB24dO83vL
pHlU/PwGVqs3s06skdiEYCj8sT0HxKkY7Vi9JqV7xm0inN4X5c+6QBJai26IGIB7
uBU2J0tMViP105W6ZerrAYuH3bKZqfLbHwP51V2Xw/dKglD8wTPxlH3w18aGD+p9
juCY4jxa4QeMHEt3D+frCL5nmMyZwjv28dBOAlmZir3TUA9YamDWMy5jGS1p20RX
t9BzO+0vLi0w0V8iDMjUVN9gxgQLlQGSPIjxalKITnTxwzSr3j6sOlJ4sgJpi9rM
3Z/I17gOrOz8NsBJu8JMNycUYCjMPgafx9U2sUdy2XmB3Gdw/4IzJl2H6yFpNnAo
nH1gkGsapqPKI7V+CRfzAMRlHm8/jxNpa8Jo153SgAvtJgBawBGLTj0/+7HRFKNC
ABXRiDLcMh3QxKy+Xjh9+gaoUXHnmOBelll/e1maY8A7a2MLnu+1XJhNBoy2r515
A55tHpAH1IzjeWEXZMfeihn9Utk6jzACrU6RCiuOHNo+ietd4Ten9DhbQV3mSncw
6n+kIqcUsWjome54ofx8Fd++GUjXGGYyW2k/eWQehgFDd41X341NdQekogKMrwkf
FKMRln37XI4t3XqrkdubDYDAfk216olN55qskyRgO8031j4vOqiKDNb8JFRrt66P
hudmwymqliP+gY52PSHE1cbKxGfLVbbfJEbPapKLTIjxbVjxWVdPENODLpZ/YvMT
2Eotez1PYKUOuUpCGuTYtRi/sOZ5QaUKDjC8dNP166mNLFIeKUgJosW7IStRqbKt
wj01gVQ8yBqJA9Mnnv8AJepBW7o0IxT3K+6vDBL7AlK7Wmv5X5QHlfxLco145QhD
lzAxxTMT2qQXuczf8e1QwWePitgF4G6sAZJxcNYDg3HRjJIV3xB+OYh/ic0zLQvO
J6P4AiNEuJ/2F7noLiRvfekQg/XNjAp+lf6ZtF44u+nGFhG5ZfAiD+oLwBme4uh1
qwZVrG2NiO4A+hlFO2A7HFq7ewRztCK8TKRjVU/U9R+ug9H2WlwenqoQkHutWRvF
nVl+Y5ZnC/ErzHdVTZQSkX55PfjbBhZbmwyMv0uLTuFSLkGcBkfsC4izB33SrvGx
gx2Qcy0SbPqJYPFka1ZlLU9wKVbHwU+LLSNErFfD0sWYMjULCKNASliA16SnaqrT
ED3FQgkRq6PZxX8D+zvVDKXzqjJ3Ex99E6VyfWZYxNVm1FK2LSBwsKubLyGY91n8
AJbqDfnSf0cNnDYMVTVZ63BEXYxfvd3/aM0zHLB4AP8AvT5h3bZzswFKbhYW6RZ1
vkpXmOZ7tcxwsCvLzvXd5EXhWFx8eLckabvyKXV8rLhNPI8PXY2xXjDFsHO6Xx0E
26PSXGTiLE43MQ7Oki+iJisIjOCgayQanoMcAsz2ZOwmMmDWBZCCW0OCakPIFa9M
EcwnPHu7mGyuKzDOZHUhNjG2yr1OTyYzP5jrbn62CIqM1mjF9igz3ayfpF0K19Ti
PdSWbyfr0uGCtZa0/jTXu8IBESXqcx5vJ5BuuePbp5B+UnIXXLMjDpgJ2mAfImdY
bEUv2AxNArYJ0eCHfoTiG4CjHxeGkWxfLwqfqj8zypgpUIB39bcQg1q4HyhV3VQF
0Ll4qJdIccZ8TjPAsGFbIZNCIWqSpETQQi6kwaLVqxo6En6TgL6mgY6eZP9u4/Xg
LysCIs86vwfHuzbsna559E4BRLUcpVJA6EE/ur9ba8ZhtE34A/sWVdhHMYZG+QTJ
jbIET02fF9IRvsgakoMMnKJ9z/og4N81ZPi5t16IhrJJ09SwBdq7aQRaEwl32Pwq
AQdOwOfdEyhaZJetSTU4V1U1QZhTsI1lT/b42+hdJvxurNSyV0I9hZkbEQj9PBIa
WvB6Ptz3u9ZQVT3qEpYRqo+p4mo3/jgPrdvlxHwqiiLvMsnX8JNmb6Zdp6kkbcK1
+z4EFX8wMp0lF4qfQw7A5Ic49dx1YZR0a0nN1LH26JRWyKXnHp4NDDI4GJqI535e
DRN9DD6S9tfGiVjr7p80kmEZVfo9cFtBWZ8GRWWXNVW/qH3DUZhU2B6DqNrCI8Lh
Gu3XrxH8j3HNnAvkeQXpGP5lttFOSPz97ZQ4IW/LXFdp0bH2IpbeWtwFovEhErKq
ZDsOF4O/uGWM1/H3EsrnFO16EOL9scEhjkYTai1V70XUsa7U+Qwt1PIVImsW7Bj3
djtvg1wbUH6cgzbs9fR2e8dfQY3zPzIbt7Fs/i/B+T3b2e7DRE4SVdWqeUkCL/AZ
lhLheUUIMHIMC8+stwCYxXgI7YPm5y6vRDwR/KKcpSx/Htfaju3Y2LE80GYGx7NP
JThf3FFZpnbUzNIuUIWarvDUUN9dmW/3p/hT4ZEHafcR2HINVpbcJpSbFUFe1PP3
7BrxlKzhCCJwZ6cv9XtD+32gfSnRy29UPErW8XQwM3PP1WPbmyHJeHUYkHXmxz4P
sK6sXUsKXLnloCGUm68mL9il/aHVZ09VlA3zSDvLck3C23dvY1woxUnENYiJBpOt
fVMMEge7/AyHZ6oxh35z+1mWsGTh/UUgZMTvypfsGufU+Vdt+8E3Q0CzXMumZ/pX
3TJAAUDEHcQbFfVzvypxs2tXWT1PWVIH88782Z1cn2jj2o0q2ceVOoqHRIOaXX3y
35KxORK3PFf0QQYOqtFGt9J2Yr7mfNi/MpWcq/+e4tNZhmmg/iwwrcXN9wTfhhGD
yW4uhHCwHAXVW1GYXncA1bCzVbMH3gDHBD02cuoIPWHnMPi2iLt0QDvftNgoohgY
Rht+V48K5aXqAttriWj5dQP4j3VncvdUJ7s7VPTkBFmxUdjMVan4J4zFaxRpjVoc
w0/JiNuuaLv7wp3TqQKA7MJmxU/o3exE46ogIS4Qy7At4AAfHBC41+H4rhr4Xabk
MurTXoIr4IStSggmlYTLDRMw/aU/CK0R35lfO+zG3BATDyPsYXgTgftPEb+pYbvd
eKxSXQWBy5PqMiTEPsy72IpHVj83MQsNBA5TDdYduUw3NaGjHWtmkF//EYd/5WD5
T8zbc+XeV5Q/hkSbdHsARpSoOq749QPG3SjSZLk0AucMnlNrvVc1VZJVBEVvFY5/
I+iOSfBgKeFp4F6H2kCWUmB0haOnzEPF+AFddtsSKhR/XAlVyhv3OwI8xA5Kqg4Y
jU/S2GBjSfLAn4gwAX8i1/LmZSvIlLvLuAWf1w21Uyp/EXu1CIgylPt1rWNDE88z
BHT3KKr6JEiTh5az5rmB+fFg3WrJkzx8h1oWcIlwAm1zTt9/JmwM+PqrYift9KEI
r7KkEd7Nbl7msjE8ZpBmXAwqGcO6VsZX74vE7pk93GTuerUcsTYwGCuBovZqtKAN
7bIbsmueR67iIZnL9rg939uq3N0zP3p1oR/KMM1zOs7dvH13vsmMxW2pePtGWH03
pHqs7ohCtFJPbJ2GSegqFv/8c+4Wab8umSQpRNk06BnZc373eakuJYhNm4pnWnfe
NJgPktd/OHuTn6EQrE2FR4dVliL38eXnW9FAbfKExbIPadjS3kT05kad07G7ym7j
ELT5UVQ+gKhlgxAqV27TGSgV770HF1hcO/tuZIInWElwYaZB8cKGvGJwigDZtm51
g2v7Nn+E1b/MKUvEjOPNKyWSL2tKppdY388bL6FsaLZWJGdFzFr1vZ0D58lwHU7+
+8/ibKTcojj2Ffmla8nJY5iF/pqDlNu3LNd7qS6sEJHicJ6/naIxbYsWDPybXOmY
gcSPhnim3Duf7bfnYBTAJOQdikz8h97EGWS61oEzIcXgja22eWJkfGSx5t1+JvPW
Zg0M/GJ8C8GPYnlkPJV77BS/+Gi+VkUAYUMABAqbztctJEq9ahd3Eq0xUOXmlz6A
cxzvmeXreI19Ws2zTpG760nnRbolfPMfAi/NjWlPcV+/R7UlcKvE5P8J+8vXhImP
jh/WUcnB/fJbFKMGMErI7GR/I3Rj6mLWPHWsOqZ+zfMxoTAfUYJ65oe2momd965h
WRukjvywVFw/z7hm87CzoyMGgZKL2j72iU2RDxEniWINR6Xk1jIHHfHXKrhO6G5Q
MwNwh9o9UmJHicSXNF5UzGltrcL35CoEQwGsfX1z4TWB6B797B+51K8FhEt6LSL3
q2wDykYKRzeYx6gyvirB+ZvrmxaFMj5g8UBv93t/gC3YcNkZLRWXVDwzCsiTPRwz
9FWa7sdmHcAumomVKHPhDQUP+R2luPABuiaGkMeiAT8SEQW/3OzjRsF30uB8L9TK
sjlJida21+KlzNtfwMsCuI5TQpm1ceqXS4RB3h9PbztV167azHidJ5Q19YpSgP4F
h+b9Shcu6P8bCUY+T4MQhMJFAJtdjYNGVR5xwyz8uxLZaU7WJJNCbJqIxSUod6G9
h9XfG0LVI5k/q9K/jBlPDCQWmhmrPFxJPmRkfG0MUX32QTHQb+4YD7/SNu2ECuJT
zz5g7+rjQ5RBiEbFOCuFt0G1tVBVOYbhyyS13M4MR6Zqsjhl6pE99bmRchbirtTD
0OtQKAWqQAAOL+NQOZdLNrw4YUIzcFNsyVee/zlVlHs9ADYE8kA0JvtMoSPPmX1L
DzsRMfE/Roz0y2n6q6ithFuzyBIIpTSKVOzMhK0fnzAN6gvMU8OgnyWXcw9AKpjP
DSjv3fzmK8p6EEBVH94VHhjpjdnWffQ5NUqSx+cHfyhiwzpKzMdyKM5Mhn/CIgZ4
JoGes4XTC2eUE4YHMruqmefas/lLAuTxIDsyP/85JoHUUFaPalAkqQbBj7HUSfKE
QCbgjApM89RkpHTk2ae4RAApGgs0umBewzi/8Erkt+zBgoqjKPeb74ROa5Hakv1e
SP1Xc83H0Y0TJ8gh9bcST/YzvpJkCL5S7h7TWnh1Z3DfDIKO93r1GkPPoj9GNYuD
A6XOk2r54nNHLH+gOFmz9k+1n5IOmivXAx5lCiPY54/mZSwZeHPIbnp7AOqFGFAX
0Dl3p4epFb3psa0nRxVZjPx7KsIXRtRQ6Avl9xo7QUyydb+UPDyLndKeTdMW0VeK
lyKU5x/z/oouqYnanaF+Ggnp4S5LNMZG7Bf7yaVPhESGibJXdEY38U43eINCcqz+
/qaT/CKaYpY5AuxKQXpjkQyAUiWkUSknQBar/GaWwsWAJ2hp+3zd0TQRx19zDF/M
pQYeP/sReuAt/wo3EHmXOahosg8muKwcesUxRNAzkzfGdpzdl/D7oJjwWXcJIBHA
PxltCD7MgQc17qJ60T+NbYmr2ux5qsiZQrmAeuUSbQsgtbrNaHz1U98MMLM5MtGY
hXnk2HoDlmE+XHXyyHN35LzgAWOyC8Xy2pMi+8oajaFKWX5CRQoC1cAvvIeh+lg/
9esA40+fsAwBFufs6O9TMfYHcr1QTozkEPCuHy0lrf/ZElvRFnRDi9vvTMOHerZE
Xx9ubt71sKBMJqM8pn9wFxYi8Br3rD3l9kMxNwO+ZBgFgVG62Yz0ixWjxFDFYsnm
yYJ/c03Jvn8acctX3DSpUKZNPd1ogyfaiDApDi1Mz+bZDUSBxgOamTb26HSInyeM
IwbY4PL8cmvPmkpOI4wIG8VrdrmgBQmxiGKOdNxNAOBp+t2/kuvOW8M80XPWLaG0
tHsOEXHVB7a7mSZOiUZfbtK0/QRYKdd2ShWlZ7NwguMAtTh386GFcyPPkKcJLHJD
ExtJjBNmdhTmq2mf4LVEYaxHXRHkYpb2luAtmCEDTP7qPzzYrukOmpJhkZkMBdQ3
erLJxISaP8+aVshtCDoKW9+8O35jW2Yh/rzVBoKIyo92S1zl+r8YmG22WgRyCAE6
naztAxy9W0dXPhVucchpIX42T0EPJ7M2JJIy85RXFivrQB0I5FoS5E4/IGXRdPNU
FM/uKnqwxULcJNR1tEhwLHSfMVDaq8gqgVfDZpKDW17VX2BpnJPNBRMogUHvi62A
1R7nRE55Eh6p8N+yCgzKBkdBt6WsFml+BHixDRbLhf92nrQYifTZQo8BvrnPDFqX
DYyDAQVikq5PqBEQVqfkLFffamtaPyuKtpQdUIWCJIHmtktfW09vtFMFK7n9XuHR
ZxSfPJlOvl1zUoB7GQoPdfV81999YtQ+IEeie4tlFaY135ayTJtmTwYXs4FjSLXU
O22xZ29IFrOthjZ+eTlDy+YuTeN4tjEnfLOGqbyIgyDEoAXrEiXnBMjCGakWhmIi
kJMsuFQf/y8WQd6IIVRZCoWe+ZhgnCCinLKl0101F5zgaI6xK+5U2vXnHToSm2R8
oM/g60+oeh8+TPPi2E7hAS/kQXhGwJLy2XieOdueV+xQcimcHeSvSGYvwtqe0P7B
+5bphD5lDSbDh6AR0XbEOxH5FDOP3JCPMahYjYuLZcFi7dvoLVleezMiDptrdRS2
XYVEQjMM65nilfDwLO2jtWGRxY0JI3+LIKzW+z+/x6T5GNXU4cRmWXPTdX8eiN0G
yw48JSqbmdwMWX2T/AbtkYSsoEx/hC4Cs0dnaVYPC7ia+CI9JDnr74ZdD61E0oK1
rxpG/E4eBH1+7Vhp3dedzWPEcNjJ+O9nuD3ZOKcyhtDtbzE827aT3Ql+Iyi6NyDI
DMx/xvXs+hy3qpx24+Jc2nX+CsZozzXVLIVJ95/9oVKGeuf4qE29GWuED8rGL8UW
EWROO7nEIyvnfOBaMNT9WaGDZhQLnrXQOLcOwmEQrDYitnPifnS5t8pVPBipJHMS
8NGu14rayi2Kzaboh/X+Twz+uppo4TUuSJy10mBC325UHNHxSiGRQpJdh3jpVFvv
C+q40q/S6KDWfQffGvSUIY/1+1FNMsRQSZna+ZqWwZKNZ4/veBXs3/VM91O2n7Yg
E4Jz5kfTUFFfYhBBGso/WF743zIbnT3Cd0IFpstnq2BB0Pr4us4BcVOaX/cE3RZu
ZvQPORlT2y8Ce3fwF5SVOy9hDiZEUlr/YFn4Nn/WpAsSRwHFl2My3OqqX1Sd3tIP
K9WMCU6z+waGYhHWMePGLb3uQq6/qvTN+461bBA1bxXgTjcFsTs7dnsLrC9EIJv+
q59STveJ/WEQJn65tYnXipgbQgH9GsznbVCXIxTImMPkZwYStAwwSn7Y6a4V7Hk5
S62BsCFhe+gBYNkWS0n7qbRQ8+Dpc+0VjS2JF1MwtWeWbwM/B5yxyIxJ1hN0Iuu4
LzzCrvUfa09bzlcRJtz0m2Vxzs1I25r5Fc+6pDeIL6fNeP56R3eCQ+7GnR13TWTA
VqU7MYUShkI0Ob85ZftcahJM+Oh0zLRYD0wi+TbVCIEIyY49X+DjyWa0wV9aBbNn
1Pzzw7xt2rmi4qJpG5cZtFzF0JfpmcgC5bG9YXKdV10IHZRWJRLfoUXks9nRPyQ0
wgT9cbBvPDC6kBWUhaIXae+snzO6CFlN+yMKptnl0indD8h8J1jvaKbPjO8ByL/5
nZgBDW7XemPR/1L46oD/9eDFkLG/3EKStvjyDQ2WEYL0gAIQhoS6PGngow+tjib9
cHhs9MWw7qKhLXXBMMHYpqCXAXXWR8mWyjHDo0FrhmPuphlO2WLN/0Jx4lpIBTAF
irbiDGlnluloi4THUXiDm2SRTM/t/bItXHOqWK7C8BgUsqQk0bQG1dOfhT+ULtks
RsDj+Fruucf+FaeVM2JEIB4xkcGh5RTcBHwgOp0W35TDeAuLLWpOooNXqPR0OwSi
2+cU43k5lhHrz4MCH4DhiChH5XV6wW4BFuSaMQ6yKz0kJxwv0ELsQkPSvmPIsaln
MtjI3lIbvlsfYkIvium+SZJkddW0dbgvOjqQ30SrDrtLlhIVdCnfLBp4H8im1zIk
s6UD+CQrvhWkF6unPHuIZkYh0Ggeb+nCDQFvehZ4L1GBHmX7su0Im+tid/dCmFX8
kwbyDdjWb5JpCRtiWLl3yIB+aJgz8UPftToz4DAZUVvMVYlXzOK4REYlJoa1fupf
4c5T9mRk7Lvbj7Def8Ri2UON0+CS6hKYbxy3lfL50Lc8N5GZLvwA9Vwag/6SBKrk
bog3gKieGaKeXgGVPzgYGWr8aWBG8z5paX+vfABXRzudMVQhYctxPLcyqiHuvd1l
lpwR0lIAaLVLOxZpizdvzWfpVyJCkQv7t8raniHQ5b4e6OGUF0EmAke5Sx/pxayy
JATxPd7o6t4s34hKC/eQB6Q2Id8HhRe9mxHQvLh+V+ymBVBVfL6NyS+G/nSueAr1
MRtNWdQgROVPXFtLtQVBIcsUzYGMDvtDWytclnpcJj+iP5XWQuT/fCQh98xrGZCK
FnD+JOPc/FDo4CgEUOqvIFlJ2s3KNj7C+zTUORWiRd5qgBpA2FL29oN1hcenAE03
75RSVvkxSum7od9AuxyuZ0pwNPBBREzznWXJuVWNPyrH8crvmhbbwylGSkkQnAE7
ro2473lZ01UXPEatvwECiy9LTJVdBSI3mrd584nRQUBQbFoj+HlLbA7pglV9i+UW
RViXz6OnpDqoYGscatqQ2XSQqop1YIL1x82wcGw7ViHCh1B9jHU6P2JF/HgiKzKL
rESZ2/1E5v6MJxPFaZnOdmFGrJCdNrb2raBohaF1NI5A0P+SmISFa306OIRzO4j8
2DuqOAOiYviNXEafpthUGJ5kypp8o4OGbVs8YQcuQJWjlj0Buv/b3VernkuHWPkq
JZfkmCDmJasPbygX6/20yMurG9HffOj1cWRW3xL5gstHN9+sFTsIJUT83wBxRbLn
SzKmJIhA407EScOxXFlbgk/LHqTpAC3KVAdkr4zpVa1o97gKt6yYst6HXQrgYq77
p2VopguCeo0qHJwBxc4J8n5z6FUJ1aml/Yn94Z5PtuVFm5Lez75J1K3YiianX27m
SCl7RKMzK47F9dkdTiId7sbk61M2SJT9k401CQ96eGu60UcN1YgnEwFm6sUfh3xF
2IrASf5oR1pgvuM+byTlm7o+bD4aznyJos+A/aaWGyM48c20VzYgTUKEbeT+Rp8t
0piUzDnKz6CopGR/VeAiVJs9Wo60pmdqdOuA4LD7sKFmgmiNnS+bV+DGcbNfCt1Q
QkoRS3UNgT5zhHSIA7SgiJkcQPMfmrHbiLEL9pSnfJ6WbVMgVuw9W4zAYcOFYYQP
qeXw8MhSSDMD9BPVwFWqtf1ZYA/bJi1vf/uHVi+cUTwhfAGKAKGOBqG0HtyJNvgN
r69pOLFZS8lnJR9kLZdIlfkZGj0P+hxjABMnSgUqCKZOHO4nRw5245g7h5deomXh
8my4vcAunild0OaseaXImPTN/yzCyg1IYo0Lxmq04gRq8QtqnAsTBm4VNAJ6qlkQ
IlWWfaPpEDTMrjrs4+7QTi+uyVTAOehmCKpWSzsro+WSg+svYTZD2YwKejWu1yR2
n+XUwBzfGGC17MvOGWWWraBtgMQdrxE8spQfsBwywPWEBomCmV1hhEdGFG0pGf5b
w2bzCgJi1hbwkLip7WcN6cIrsNA8PzHjTptqxWuTe+64HoUFFKLyKQTowAID0W/0
ijn1BKbVERgl3gMja2DOLR9Xb0XHmUa2GxkoCmcN3InMJ5W0I3e7Ry02aUVRcF27
vycOaS+Sm/3Rlk+X87qrsiZYm4thRGApOvLs1iiyCOK98bWkw/121yFYcIdEP3wN
p/ZX+67Li7++pKyqbRRHxafIRE0eat3zmbiwyYnS++n1j0gRcYe1Od1saQVxmq0E
FVMreehFHd6Ydh5FFxYadu3TjmdeTNcshu73/rFSu/1262wwhTOLJDoj+5f3oRUh
NSAkUAFmbSf4VsMaeZLDiwPKhG/R171Qkqp8VwrKXUk7s7Et8OskN3kKL6UrfnS9
ETag4IqpMMMdSWXrLjf1qH0ZslknBHDp7jfGOfYmoY9UjJ4VnrtOtZtB6T5FsT4u
5eyh6xOPl/mY/29PyNT5hyM4D667giOXrrjHha4Zot2ood0teJBqCOm8mLyC8eYa
opjyBW8A2gVx5eavAHiK1p33YjqafyMWDolGhfzlc2uwu1kc+kbkFN1HB+EUbKih
HqjG5Px3Hpls5LRy44fJqucHMnx0KfYWzgjH5q93tR8Z0K6X2+qo0Op2IrX1myUi
hUN6zbhWYekn43WlTwnWLaqSHFmVKwxNYZE44YbvGkyF5uoChaaJBIZiJMX3hNuu
qbHesh8GeZ57/gwhpANyRS+o6Af/NMDCTHHCZ1thPmaCfWr0tgLFzDUpmJzWFDFW
+fzckpp35WgZDUZOae0belXk0zh3b8W37N5cUkiyFqZblHVeX+eo9Up6//yDApjs
T66AcfkbjYrv3tJzKBaI4QcglzlqZ7tEGDKX94WfCoofS7Qjnvy6FmJEBrEiVPF0
em6KgCRBXblES864p5Ysuzg+uVT5kCIo+14Vfxa5YAhcC+cKf0joHyYLN6F0x7QK
2ETz/pk2xiRGShHVIjnCWTKSnld+zeADGHtCW1+uZe/xmzXH5Jd1mYiWm+idj/Yb
vvHZDB5hPGCoHRlwtsDkPL58hTz4jw/ewS7FWL9TpJJcJ4CuX1CTYXjOixSdyiOH
wtiFYuqWtlgiJAYYdz2H0jcM92H4grsB+zhUpfvi16o+gVFX1v1bGyBiIqMRFzaA
ZbpOipx4L9sBc4qtC9OMCtJxbdJQJeVWN/nfse+KdEjd/+pGUJ9yf5hk4jqLTxy4
nui57gnNyiutanAY3vh/ppXipJniHZibxNFVI+PNJaKkqq0Z+ddGtP3WvTnqI/uT
xe1KeDK6y9Dqg7HFtnC6UezbtQsrl+nn8yBPfx6YVGb/T6YIvRc5+obgBH8gpoma
0ahocOwpDFXWixVlxhq6GrABXWF6RiStrqfj4BRofNhPGVflSi5Hnvn9oDPWKplh
V/3LioJ6HFHHJJ0yDzAZNLfBLn70xE3h3hqEBj75EkG3DAvIvGcqNM743dEN0jzf
WCIUNVYWvPyt2fiDeDZfaL82sycKwoYMx9BVmZfM3GSPtWLdm0QvpWba/PfduWvt
v0lBSpYxrWEcsT9vdKbuknAdLRyYbl0/ubrIqzGxOCB5Z2I70DWZKRzs5lt3KLfk
XNJge9P3S4pBOF9s8lDQRVdPt5O+bJNs8UuEww7alNMKxveCBLJgMhRDUXdKsNYx
mKHlDjxvMcd0gvEFXKb6tmdgJyRSsOQLuSChtQCnjNj2DoBXJCSr3Pj8u3ZsJgv6
E29BVLds5keCw1Uxu2TJE5FRcekSv+YGuYALwJDmllywL0EzibTSXUqnndda5cKl
T1FQuo28I01K4gA+nhZRXXtrzjoN1F4CF/BVqXMe4ObfRK3dksdVGxVj9RBbAtJ9
Bcxz3GBW7eBWWfei8fIDg5YQ7Nd3cbpY3Ikty9lZVlMLuwF/E+qQ++T/7/YdVZIp
DJmV6bBlGmOKecjl2M0cIgZmBY0xCKl+IAI7IO1U1AKTQcD0szwIZKQ4ONX4E+UZ
alY7QOb3Rz7K0+GC7gfxp8GCjb64SuwJm3qC4XXuinrXFPRjMioWglTIKdYSdg6V
aq+C5jHc+tKshCXCbj4forA1BFLXzsQlH/eG0IagJvMLBFtsLmd5gwH/VF8wm2Nb
gOLVPh0SKzv802/WkqbjBr6U3fquJUoMy2yLa/O72/siTiwaDayYHQwv0uJeooDk
aap8+1jJrPyzzXxT28Yc+FNpmfmwcHoFiayNiw+eu0tsakWzacbhcFIfG/uV+/KF
z4Jx4muwscORLcgoimAe3EMx88qgbCQFq2g+5ls912MpjweMMgPe8Tr+t5xlN/9m
SAmMBi7qcddE+XmPbpKwvYdeaGcRct6cA7xPgrFLmoSnEUm/izuzUKS/apkdS8fl
jx9s7Misos0PQHwhqIy3XG6JjYriPWl8C3FwOrxBpNGfR/y5kbmoFjMMBz25zRg2
Tfuhs8PufqAOAnod3Kzhtazo38R5Z5jwTMk3Gh/I8Jy2JveYGOSUfWYXZrc0Opx9
q6PJbHDztPdVowhWXZ4fUeLfgFQfdPYgpO298MhmDEiagnFeylc+qd/WL6PHffft
x8HU28i7Asg9B7NMCPLC4249VaCT27zNd9UkA0PZUxjcvN5RQJjevyd7Cmz2yiGG
f+UHGWV08Bdppm3FLXeYuK9usdVQEFnKPjebcj8kiQdxjKXvLKFI0TO4jPTGFcwY
SoC7LFvWiWnuFamKm2t3kYVm+e/vkz8Ry1ynizxIO4jVncAVkLpOuQuhba2KAwUc
Cub+QIxm/Yvs14lvG9wMZbnojiM+/wqenoskwbkY+GQYqxCxxvFUmPth4pqThy31
om3CCuSZpgjXZnxrYWYbuCox4AfuMxidxkv/LA2b1O2G9Dra0ewaHYD1W6yuF1O6
9yWjbDmBruLqe8qc5s4fEMQkR27VVuHiYCFfuthnfZxQYeb0OVqDgmcL7wfDHeVU
zeYwNIH7ek/f343b81mjj8BTxirJUBvjYix75ntt77umieZvEie7sTwedRGOM1dF
A8qTI12hfX9O5UPWxqk7GAgNI2vPI6XPNnnDxILppL1s5Q/upF7NzXAwaxZ0Zf+1
+9JN5F2xDQDo5JeITJ16jyor/CEJfEWK8o6PmJllsbn0KOM5IBvHtRI8j2tBvoo9
15u4sxexUpQTHzPW02MXH1ySsFQsj5sO9y4cOAIJZCrWRUp2rzkhNfQrRqRYXMiF
V+SUtxXrPaU1fUSqSaLCwQ2rVYeept9Oaz/rU+HH/dCAeiNPffo+MpRFEma/Pjer
NYpAhYLxUFfXQMu+e2Hsrjbq7rtEtY9uo+8ZeE8TYknfW32kdBHAHZNJbvQc+iVI
VPRl1Zu2+qb21zFLUvw0gJChobhL1+19+Dra7wJFIjmfrrq62yvVisx0O6hHEJb7
cOPJHr5P9HSeRtqa7dcLeZW4Hs1KZM6AmcoS8pA8mA1++0u3pSiqDt7l6c6wWroB
HHBctihgh21IH5ZfsQNQP1JM7dK5fktJTUrem2vbGhZdcj1wwgnl6nb+jXKURHI5
PS0JW+Kx8Tjm76F5QHdMFNrhnVRjfDT8Bhgppi1Wcbnqs1A9jWBYW/MzaZjX4M+g
dKL12NUI0+I++HgKluZ6Oow6k79CqlLFanR2i8eFo5dR6/fnQV+fGaaLjaBGr8j5
wG3FAAAxsUJnP5Jw2atQ/wg3sGqWU+EiIXPDp3XdQnuPmxaz32+9kMsFbhxvvDcH
E5D6HEwnWBTvG2RJsYUiJd2WXmuUanSrifVx+tMOIbzRqOOoF/77hZJKsB/yJLj5
hs7LenB3kCSdLevuK2w4EWXX2tOewBDlquICvznosu9lpwrKyfF5mKxHjVEmYZvC
TxBdNddgXeEw24kHwFDBoJ0KO7UzMNDgMEHhagGYCkX07fUI3GPDZUeVv2BWD09o
qUA4L5IXg4MyNXR1h6ymAbmsqDBXP5ecKhqE7YJQpHGA+L6P2KYRyurdadSNYCbF
YGJ74ifQCSFpfdF96vGMl9aX2cBKfCEZdMtO0nsal04PA669NluyKyftghQksO/k
fjbI1NLf9EAJb+5uwigTLsp8xqDO0JNH4j/Qcimg1ZOUScpNPeQuf6xdpmMzhh6I
YizTGvRRQuHrckAjmEodyxpZgeIq1CzIifgILkLQXGY5LregKtL7r3hQNNE1XP1g
C0wGOR6d7qrGE86KIU7hkP9XYeMv63V1oIrFaEFPwZS6sS5vSZoiwc4cB0aqKDD2
PkizMOW+h6uXa+1b3/yU07CWf+YpjeLjEwXC29MvgfyUyXTzPVog02nfNM3sFdVQ
l1M/fk0k7L/YwfFTNRVzrqROOp40Tmaff2W9Q3yfdtSzTONRb7kwMT88wqgl0LHc
fbkEsl7CakvkH793eyFB7qqYPhimyYmOFLDeqFlfpIjH6uwgfa/wyZs9Zg2BQDkf
O7SHt+G9dFOhoDxixAjZZw1lOK33EesZzYDqj0zPH/211C+x0wCsFemg40OG2btR
HedbgJdYE3biuRvzZNpB0HDPoOsLNkJCd75pTNcj3q5S7RRznGUm/TwQjAei3CuG
tbsjYwq6lO80vAEwSsiyhU8jZsglDwHLYrtecjvQv3wWEtc2+056tDEiRfDOGXdk
VRmgV0Vn8fWwK70KcMKOjNJuGL+/2vJaECwNgpgf5hjLkTk/4+ygK2Retir9gGqK
rY5UiB563Sel2z4QhT3wb1FyZdo+f/dswB7TOhasZa/JtsTWdQHSYLTfnkAtLSFn
VD4r6EuF+1vPx8H7wCLCzxAt5Qdo4/FU6CvTLwzvMziRd39/C5CoDh+wN3dxWCoP
WknAH9ZEMkkbCDZcKmxpK8KqX++cALQHTWSFhVgFLJ9AIpWiIicDI6HYALaSpBp4
IBC9S1hr4J7WLwHIgmxdbhfeu+acfR7xxw1JXEALd5VjhVoBsXXM8U6tQVBN/7Ja
gG3ckltRyI7CJMb35eGqJa6dVorPBC0lz4ZE0VIKDVGrTR+klmaX2NrKtJ+DmsyA
2n44YC3hONn0wLVtZpE9nBw02s6dbK7cM6Dx06huj5Ba1uGH3migxHOqKCEwrZuE
Cm5kL+1oK78ntzU9vFKh9EkASlDYc3t4uU4RzVOgR+ONlUhkmXpR6kswlzG1rM/z
fT2elTgkSKJHSaZizHXpZbOb0OSoqHDRXi1xpRnAKzi4YgnKrcCyL9dB4y2ZGwCb
3mtBzuA2vPwFjOW9J2FrCU+mX485QvKatwIZJU1T3+dj+37HnFkWPgtVzoCOA7/+
/XTQGHQfO9ZMglygeRmjZ/XrSXYrRsIEHpFBOH/nmJjp24v6jsx1YE38sapN6j04
ccIvtO3f2WG2MUbQYAwKgekKts6u7r75ITgJXmvEZyW8F9L3zDJNGnYhDreR82oh
bG2WKhuoCFa0ZfFoIjV4/XV6Rey5UN0IqlvXUz78QUjb2DKvUh5Q9Mb2sk5uSN/e
sM6WaESwO9p9+fB5qeMOz26vZOmNJVvVGamUEWSEOWtvan4vzd8NEtmlHBiy8Spt
Pg+nVRgR1OJ8FDGiCleo1s37PrxKBf8L51aPA3XOoHLzuKkbi1DOiFIeR2k0H0ui
kV2VQdwTiR2KGGhgjvdxH/YhBK+UFLEedn/HQHhEJ1WGNpdSSC5+7TpwI1J+eKgo
tOXkLn7UEFon+mCxbnl6ZPPQZSictJQ6AooV0bbEVi6Vr/B/ki8e19A16tnPp1y+
PnJ5vhH7UM/UCLVRVOwklZID3/nzodDxbhm0dQj2xayzkS+i6bYofO7qqKFiNQGL
LcIDLcAZuP3GgUXS/7EsGZ8eeGo9TU8pXaI+txCditxB9qUGmfWu2WgXFCppWdQ8
0LKLeoK9I9cZfKk8MjXMYewN9/DxAl2Rus4aCrpPbz+wNqMqj/ESLmNzOXUOx4sp
1SvAKX2+eEAspLm9O/m18S6c11gX+rNWeSDOTeSO1cjYcaOM45GkhoJKwErmav2V
m6nz0cP0tO4RkGHxF5zfcvhountfhJ+xGQOXVTkXNcsbIQebd1sSlCY74b0X0Q8K
p001IKdhfjCGUcgfdDD7g5Z+AgvEKwVU3NPN7ltCkudcLThS6JxeMhNqFlsBrDjP
smROZQBQWMrtnplfKAMHdOe9tZ+Nr3uP4WyOC9bjlmmKnPi5DJQtznnpI2Gr2K3c
jDlMr4KyNtsAHmasBJItOfpsI2rixdd1RQJSs7Cfa5jmoBk0ZW/QS4NGzm2EKaE8
vvh0gLNw8fNjZH9rPFzmqpAxELvYnhTA4F+5Ozu1aT3IeOM8fvfzwakZM68RqtJn
S4G10fQvcVxpRjJHSikd/VUbZxQjE9Lqo7w2GbcXHyzzH1FIEOMpAhzzgbPd+52v
qlbqGy2rm6hPoLVr2f9XBxS27g4PNLyGallPmxHwR6FhBosIMzY59ATd2Igro1iE
fkiczNiL0ZAIO6lrAwUQsn4xhtUwrAAStLJ0J4jmVBtSRZ/NXeAYHZc7BAa+4PCk
3c3SmhSeUl7+khtfci+Jc+vzMHzejKuBQkkWqTeWvs8J6FjA0ruOw414zZ7ibkAB
/Cdf1ZZ2StDHY7aSAofVAa9yB/W3cBnYxigZoKnPLtF/LgicmGKtiyKN5+F2P0Hh
QxL5/xfxujzlQ1QZZlwg5lQ7sLxs0Qy980olCPpKJpBrQp+aXwlPPqbYhf7kKMvR
46aLpe3kNZFSko2xMYFWEfaj5uwFvY0hVE3xxj6AiEeVnJ2v4oZB+fzm8d0NhlEX
4BFSwDjrolepgM/Joo+/7It3rWf2M1WrDB2nPLSfWxCeOlyyM9pFtRoax3Ziqw7W
jReoIxuMse+hjSmft2tN/JrQIg9hBfxc4HAHFpv2nmRSLbp/jnQi0XgDy/zOyVUU
yl3l+QulmVWo2FeycKHPJ0hy5F8TjlDW70dckrbLFCsOJhAy8lfxhh7goY6cwCHu
0CHiJG/XWGuiJoL6cjrGuj7zdV+XJnY5i8N6kTZ7r6ndjEhiXjM+QW23XDLDrVCY
+P1Q2OFCX/p4i108rUGGHHaxBlpGRboIJ373WK5dXwbF4PfB2tfZgIvewhF0KsQv
r8yxZ+uoERQTkeH7Z8KvvchcFXgiXjTFy/Sy2TMrOe+y72DapievQ+95vegIXfe3
ZwD1vh0qSZM7bzBvtdoKHMoP6kBD2ZC9vaZAryC1GqdXzXTBmL1XUaXa8ivVj1iA
ys+AUyRYfGOpgww5Ypma5hY/h5UM35G8XCJhAvWDzRWzd84SfcDWnOUXBXDmCRwv
LPlTNmDrL1QkdDOD+OhB/0OGq6B/jcxNJgKmZbd+nxuwXfyXLkPHGEfWRy6eNnbn
Y5zX3JfeJrPiOd3RW8PJQ49CCiMn1Srs9Sm8jAdQpQReaFO7WFvwM0ZGrKEn/ifO
oBE0s49pN26pa9WV/IWHIYd93uzBa248MimUUr2HSaRPWOGX8Vhhe66yqMg12J6S
jdgKO/ryejqqSQeNU5TO/jorDsYJKgKC3psqq9leBrjNwJ0SDtQ/ts3x64YpIqg7
bfJcWi/Y39nyNCBwusaFsxCxgQRa+Y9L9PAymPmM3ItgxWPVwPzq813tpQkmzPKI
N5k4gtZNZcJZgYe8pbmj8ilaYQGlJ7cTJaqlN3QkRkGxQd9pILd4zWjYxG3X3Ul+
qdkaxi3Iy5yapeKxnblEW/d1Kj5OgeINtUevh9EsPh+flENfgbTa/5twYLYStxrf
bEs9lh/gN/8HHxrmbu6tBc3r34g8t3OfUDqbGzcW7xeyJ0/AmmC3qcNGlzM0Ya08
IN6k+w/HUcv0LpvvZPJNjBI9AdJMibdSw+2Q7dTHdQ0TAvKu4Lx/7HZHYkEJozGY
FV+ozBG0UWVtwBSby7lhU/9CRwdAtv1K0uck9HYB/S0LZaY3C1EEBrfj/MF06u5u
ZgdAZ1ahNTAot5/vPm9wYy8Py9dNN8nNGWzuFkL3t+AdBNgskN08Q1hccuIk/Fj+
5MYlG3JncQEs2lBvyrR3Pn1xB9vOy1Xlfhs9v2fS/9j2i/ulSNSgOKSE2wR1mH6g
Qrgzhm3GHo4jf8kpIRiE5+eHSZXCCMzevqkPFwsXzFT5K8WwNkJ3lrLp4Gyx5Nt+
YjaL1ks68N916dtPblweLml9Y3LtaZiX7Z6iCjWosmMUHy/qjKm8tsGPn0gcDI6O
XnJf8MzzaIEddNUJwBFLmtA9/vK8ce0BtZZ4IUVJ0+bNNHncyvp3mXpPtUG+SE1m
t3BS6jWjAdWgalPgpVRfROji9Y1+b6Sx0nOKBBlXdGyD47BgA55YA0Dnrg8AtuuH
JlFNVZptrpczCfR0UhDOGlyQ46uKTNo6E/+3EBUi/8jCk6SUH42vGBJxOcuRF9iJ
02F2KjAEYBuOvGUu7LiQGas+rEbotVJ4C9jV7IlG23ls+JWgx8bd2u3XEthEhdJo
RH0iLLm5pq9UqeluLAPJO8BcPpDttQbNLIzw+lpYEhKapvtHzPpFlRzyE9oBw4LW
+JxWwjSNYt6PqGdEqx2Ws1G+fMph/h5EZOMAQHSBpXTPEpIdtxvFTxq9Lx61zVke
FNK30D87cNhALMGymRMH4TkgGLYMszuBvVWm4abLuMi2HNyv+2g3cdgaIb1/qxxu
rAPq8uksrySBI66lKX+zTeo45aYrWL3u7A0UBk1sVpiGlZ22LhiCFp8SlwXC0xy9
WWxIrhpZ11V91WgaPnZLZFuMiX0DHcsKjHVPcSUjLg64ifnoRUDmFw1wPCeUKjrb
Ql/soC0i5Q4jMikMGcwsVmNfVkcvSAoqrlPfTH9UXJLSeoTSbpbF9qXQtwqdriGh
VHf2FgV10mriFMVUpDYvsCft5d5U7ECfb1POZVQ+quTnLSqRaPm9bFIw0Ckotm0n
3KYTxRD33wVCzBMweB63YCt9rzgZEn0uLwCLFJUwz7+2jJvyJSr0nht1Wpw1Tgf8
MUuGzzTVezAW45ngZtZBhoPq6apCnVdrb28xK7tvCGDPExinmo8v0uA2g74nhUbt
TzZlQUymtYGjK381iHpZq8a3gAXA9mZkc8O2XhENEGmXwX9f08R+DNVSEu+1pi2/
NOpcks3rWKafar3ykzdaa7u7DuctAnA2E7osm9xe1hS+AJs+m6uJf9zfi/WK+hUl
U3U+3C3CFSt4GP/VG2j/K47rekGE2aNEQ+Fo5DL1P5V4U3Re9Zmn0lRXW27yGw7E
PyUd3PjqoyJPDFTmPpLapQKG6ctr8NNEnjYdd91x+TNg5/a1v99t9F1volfLQBi1
h7uZC9u789MtfkxytKlUegoiAZKs5jEMfcXhzH5TCd7d/HxqLQ+AMKdjcZf41OiU
4W8zydUL1EAnFC+7wLxZAasZSKOvY4XuGZ9na7RUb09Q+rkjPxtToanD5Kh5msKW
NwEcMmSUGkvCTNb8iQNNI+GuG5hA9sVeTV2Uw2uEZS/q8IZLIweRz7ybiLMhkcMD
kQY8cNOsDuEN+/0c+vceAbXS9D1p6xneRJ/XPY6FCQadm/GvBNOtJV04z1WB/rOB
iywQbMnMXdA8WTzqYtBwmZi3kHJbamGLrol4DuEzAy3mDwsR3IKj218RvFCLWrMY
Mm87j2H4YmuDNbNLRw1pMw6cGbGBemRbhlTGQORWYASVEH/KMQyoP/2cEN3V7JP0
QEI3Sih2UPgGE2XOGU/DBeLMSAEiFer3lfnVF4/UzIFt99IwsBJu8bpeoXQyBe/O
tdG/fQzCl9XR0BpM3PBLIpj0F1rtVGQxwfJYQ4pA9H6tyF+n5aGR1DYFmVhI3J3z
0P2BG+WCcgCRegCQGsYQ5ldT0knJwO7Y+wJX5azSigxVQ1rfUoQZZZ+cabm2N3JS
STW6qV9M4aMTaWYfExSteOoonddPfq/0ij9m7qxji8uZ50Mku9SJwZZohBrLm14J
yVJAIruCe4oINAHmgsph9Lqdg1SjClPMhjGLSSU9xNKp5kPCC/MG8xf1xXJGo8Q2
sXzgAUuBALct347dHT4oTBFoPGtsQf5+3cwrzsCuO2f7NKRzR3nW1i4AIZ8z3cul
jYENpmu1ewLruwoPYw4pH/LnAq9aipjl+OkafKlyjm+FNpUP3UTc69uZWoj+CgyA
6Zm4T7ggnImukxieLxSBTRpWcw1sza3r3xpask10+Z/gsfYO2ck2L0T9iXoTHdDN
FR86HZa8UwstIzYujni7B07BrVW2vFDrVmtkUe/YXyCJBEnVPTQc8eZadcAYpxjV
zaRysCHEWgNVm2cyLfibGQleBs/fvV3fYvSTs7F7IfGwVVzH9XD8KpOj4mvzuVW/
efLtQTnvYQEzvW2esH08pXsRVae1FSkhDmDME2XqOJ+0LZLDXLUClgvBgKUkBaQP
pYa8myiqoGC/yc4ixiQJeBo3spTRbnziL0d2UBFpd6oJFWMVI/TnC4ZM4fvK3TKd
RGZC8yMJh4Cz0XyrupLKs1ZsuD83/vNZ41+6vkZpM3QawIMnNDJZ0V17LuYkJuer
78+B8QwYP6WgLQy5gldhr6bQyx9Egt3OAhJbiwRykQSr+cpLi52TIXfnKHYARvIN
JUlmtchT7OU0aaH4fBaVV2dtQQVRYA02SzNtXZWcwQ6khORiyMpx5LoGE1kpvZCw
ppiCwTLzvzJjRl4BzoBZYZL9tvSWr7WD7htvbAewfgIHLcZsrw/s95Ou0rPxKFGK
nnjBDciZuiqpEhqzGBrtj5m7cM5S9ALwl6p3CoU2lZMSOKv5Gqur0sBUU2D9/dUv
kb57X/Nj8rtyFNW9e5W0U5dOrMS4ibv8ql4izJA70WABLi3XAgjetn5NWrfzU1Vq
d7vodRvcy+WgpVJVTwH6nEH0hPDGMlNNnxNzFLLEJLrWcSgXFtcYhw/KudsICulA
vdKv9PN419IyytVKiEuxmi4haMteNRKOrS468YfVrKET8qzoh05v8zN7A18Xwi5T
RkTDxn52HbU5lnuUSib+2c3LN/sbyElf/O63ahBmMeaJqpwYxvSeMry18uZ9eqK4
XFnmZvzNSFFP9bVO84NL5VepjAtveBhwwUJegU/E15hd6YN3MY2eDgaQuDEwmXos
ySD9MepLREQpv073rmXdwwjXQD0F42VpLemo1vkaVRjjvGg/skgd9li6ov2Sc3dG
ZMbiFpZo1Zi2l631w/0I201WR/jgPVjiY5VZtOMJIHDsLJIhXV8WNsRBpR7FGbDi
cYarpP0OdR3rexhJbx7P9xI8JvqT8VY1eNI/4CpkbtTrgZF2YVRzCu1L2HzShgPz
ZoSycA2sYdeXCgcfI806JeONWlYaLYotySTZ/+d2j4/0of6HHxweJ9baOTIjrXBO
koHILAPbeLenyc/L7V9VgJEF4HF3/R60FyA5un6X1S8y3+m9oGBWxj5a5Do77IZT
ZuIPaju5rNYUWnrCI0bsctewEjy4BmKvo1KDmjVZl6hdQvi6YXe88dz28JQAcwi3
pMheanYIj+oTq9MVG2LeSOyOBgYAydijuqtw+b3Nkd+yGsZtBnrHM7EUdFPL81um
tcVn4KLtuqwoqBO3ccxz3CHFLARHJosYaNHptwZl7h447rQh6jnC79CJzuk2E3NP
RIm8J9A68xs5qcK2ns5KCdq+lb9Lg/BZuJ9yir8DaJoZHb9N8rGdg5DtB183+GUK
boBoeFKHsiz20THv4VLJVbt1ZQc4iyKhY5WEIGq9zhwe3DNwy3eRwWTz2kp0m0fz
qxRO4NIwlDoOD3yZ/amtmbeeG03+tf3wi4r+L7beCoD1OSZE27x88d5FwMNJE7SQ
ptj4cF0FWy0L5Dm4cc/c+kpml3KGgkQWiXTdvzmBoC92ToKQtfR8RXtpes/o9HG4
Hthv9qB/8ZST7I8S3/YZjtweEQcWhaLtHkJLZJBMkjLjtYtLUMohEstlssvMZJ58
AFBNFNcNJXF0V+NR/KGddTaNGKNmrMjn5BrfP/ZHiSfN/m5RNVglA0rQ9a8CJreW
bCPyfmdBFVGPzz7hvcZZRynxNj8IFr8cS3klxRgQO2UINzgBcqHrX7ScCgg7cCBh
QJ66ca/Yc2VinP+0o7hngf7Ah21FTKuy4u0aRyWjdF6Ck1Skyf83HB+ThdTDpA6C
tWtILcKDOF/b2aiCqkRye8etM+YNtu1FXfoIgwvTNya07OmO1QrYlcB/qUinShjF
PtioqKb1MhFslVbifmel9FRYC9uNOFo3gDm0HpTHO2RFiqt2nV9upBHDPz8bxpFi
d4IAoxz0lcw1bs6OQdOC4pR94togRC3Yy+LVYzASIWeI8bdDRjzwFLAWAYzJdYw/
D+B/17+Dd01napXjxjf1Ldv5IIMOOZM8umcHPimWm4JywQD4Tx9Y4VZ+HEw/SFaj
jqF4X9NXn3GeTEJg/d0pwqmTXxYoTXpIND6J4LHsXoe1sZd6NcY7aMd7vkSw3O8l
kD9bc+gamxAw2eV6oSZs5C1JgDU9TkPpZEm9gbqPqnaKR3NlvHwzFVd+ur+sC129
4aWOKTOAP5VHghENYvP5w9QIxfMOkvQxVF72Y2EQtQXlHLeFwRcY4l5yVPRWIp3/
oA6iFWkUenosngyk3myYSPNkf7m1x1lgLbdINDPKqfrjXLmIBWM1NNC5kxkLjthH
FhM62X1hMXrD9qxX/rNAhF6l2TRM8hA1j0GworT9id9ZKiPHkHHcQZZgaGa4VgqN
PfavcIRvoqSKszB9mHVSZ9wZCR6KnyGNNMUeUr+hpYILZlyKmY03iSma01LfRcmx
a/96V2DIsLlDCkliQ09vAhQbXFIRbWwn14B2WjHQBxxbmOauFGN5HaVRvSb15rz3
DomS4JtnNJim5fLs44KIHc45vgfWlyhQWCF8ZWquqXCsCcv06IwF2LFjG7SJxaZ4
zgVIxPfc977P36qFku1QTReD2bjpk/7Xi16WWB/FQS1DDogVGTAviqjvkC6aokRa
mA6d8CxJHCLalwNJ/twpb/BCF18DqTGkeaBDSJO5QJtZoWVzBZ8OlgKcGPXMAd6U
fxckqAh1VDrsQwDmRovrNHJ6uEiqr0A9zz133cG81uWNB9epA3fkKwnGWWwzYStZ
6nDbpFidUNo/+rFfh5vzEesyOEtkEfWB834pFB2rf00HGOy+J+IWXc8Sy7G3hKRQ
gddb4JOHwT5W62n0t+JWP2WaouOyyEv4ze+bhwxAJYRiTFxp0dHljvf44TdPQSJW
uKXftNALEsTLPD1dpcbdo1mqxZCUNwPyifkGXOPyNwzCez7Xbp7uzoCMXXRpsoRu
84u6wPJ+IVlxh/wRJP97R0NTg9MsMctPnrhQS2O92xGnvXUeOLF1Yr/BBsQBcLlt
Olkw3EHCzVcGbEN9LwlRPDHCenhSq2Qnid9kYDMXgaslf52KJ93LZ03PWzyZNKwp
HkPVAifFikO2duX/GW6+DlPIubNC+0Ng/KFtnmeX0hSdIkKps+cHlAb1bJJ/BSOS
REbdnxmihQkRmioh0+EKO2yNJPhNqkb3FrHutWbGgz3b6IgxJvXejrorx9ZKcYAa
XNlVNdogGMl0nHhYGbeP/7thQsLm6eHo5/zlATI/QEzQj8graB3AaJdM6UT5792A
m8aI6Jh0sHmuoP3O9Q/Az4DFzWYVMlS7Cyo9PaIP0Dlp2cfdG8PsFC1BUS4xYiZT
tpR0EiEIZbqPHhmaFuU78YnU6biLvraso3Gq63l+ukAe3JgLtpQ+xoul0wPitAdK
6dshP9/wOT/K11MF1Sb3d4tJiMkT5Ob7SB19unK4bHOL793LkAhoJwWFg5lFF0qg
IAbTJY49xiBDAUFawN6bm5w+nPXpgNy7S+6LsWMD0Lc2k+y1i0m6N8DFDLhwGIR2
LMhofCqLBwvDKOLnZpK7VjzKUJtdF1yX+hXBBTAnHDVTU2254v+RFSwelCFX77nc
jRdxib6imtDp0ZqZVwuhutfUSGhc0OaFvRjizz0yYEIyQQoJ24VLFrzVPrSMzj6h
n9kIrlYBfHnKoPMBSsvyPb40J64x5cTdcbziuzjSUb6ILF3QXV+hv3/W3yh+gC6D
wBRH389I5nQjwFvikkEXgS7g9XOpApj1KTsv8wdwOMGrpBtPG8PIDv1LnV++J6zk
y8pRweTd/5k+7XsxgFaBTCLpjcW1R6JKRBcbCHt8GSaUFOzMhOrdUyMnhSLRciwo
M8PUxkQVZZ38+hxVCzW8UxPM+N3mbXqGL986xIVsSsuta5rgh/BRebztoqYqHOyr
FFyQhiSTT0FSySYzbZ5wrQ2ZqKqBsOOjU8Wsg2TRwDGkeq440nbP2QsOG0Wya3/l
yI4Qq6s5BdXQLbt9K102NW+G0763tfprAImzN8ZsoiHulavbld3fLjAs3ILA6PBX
WDS3uFMXo7Jg/zFk/4IBOXhJLwG/gL51rMCpjqre2XkKyX3FdVnUTLjYNYIK834T
M5nxOkr2aMv5gTvCgNWe6+aXr/aRfTJ9HCsTvKyuNXSQjpfMKMa8fIV773qj7BxI
RPYyvnVwbJ2rJg81OeO+cnXRk+swhjxjZ2djvQBT+oQlJxaK51wonHIcRsiYbOd8
UREDkJwAwQGbriXgcqSTv6JuVOdE0D4RrOURhGnNp57ASZjp3llbXlSi5htcAL1n
gpcBGPO1G1Cxphmu1oDZiNDohD0Bijja0dtqJiWxXRyPWx51RbeqNYZxAwfCJs9g
MCUg54a2D9s3qidYygyStO53soOGU389+qZKXbKONGThNZQ/74kpnv+HCP8ON/ZQ
39KQjk8ZVnv98P7Dd3MNDO9sRdhowrksBqJ6eXSllq1VsjRdAdx2Z/MAbFLe2V1+
nfTaJTOA5fByAHawoDdBKlpJ+NUwnM9GxBDNKr+zNx3f61gK/SR5itHBjrv0uXTS
t4+h9l9+/2kbX2uKm8MFpbx8N0MHvToajoz0pIJVx5lK2EVr6CwktY81LbMW3WUj
KwGqKm6dwpwDHMYp4/MB4fOR+pCB5UaS9/Uavq1gxYBKgQj1WhNnB2iE6gIuLQrB
E8DXofK0L81UpXaN76uu/bKrEzwqTnO91ap00VrvwQlpZzfRNEb6WGKps4cRLqNr
UNVgMCz0vUPR1j7OCxJ1E2fuIYj0UUjr9sVa0fNgxR6smd6BiuoK3fExmWG0pBFa
21nqU2tbILmCadRx2MQE0H4aOqPIyQ+h82FVQKLWfgPpszyguVlw41moiXzodhW0
XdNq4BDxWuEEdojAeRMy/ly7wjT+3uo8H4GZlQAAmRmDYmZ5WqeHaTgNJtAg4doJ
QsF1Z8I/eZSnWQNTnGbSechcagdIFkMoi/lLQx7qQuUPsRI/zKGFshazpzZXSj6o
MFcqKYXsBnYn4hyK+DS1R968Lh6/z3RkVqpo1FxoyVVr91PQkXuZnq5mNZca1p5/
idXVEw/lMyJkoJmK8tZsFgHYBAsInrJ+R5m+0Zm0GjPkJob5VjU8lASMD49TS7Yf
6+Vi15TEyvu4uH1Fp3KCZ6onKusBwF5VKWjUbmJECjOJ937raHRjlKOp4BzHI53P
9g+Cqenlfw4iBUX8vdRx/v+JSTKVpIj4oqOCvjIojpr0QxUIB3PbOuKgp7vk/JN+
DobpCrZ9ePb1SS5nANkf8jtKeRGyuItu+bQDCqaX8B/N9KvNcnV0e3FTa6iDlI5t
FRyCGlPWsn4FT5j06TnXwOpD86rGQ9h68+SNJABSzOXha66Z28CoTK/B1nhM0Zzy
hwdIheLh6Mo55F6WOJKnJaOy+mQKLz4ZH1VKSs7pCE0W7yN/f2L9FNNf+VeAE9P3
smaHFELXuikeSGQ3AwtQQ6QR/caja0L881vAjRsDpAuD53I7a0t/PedhQTaEEoCV
TB+C3x797dCFfJhAnEzi+JoNbI7uGc1PQl+yLOHJbLZw1SQ7yr4EUvhKo4ouItDc
Jsv+YuWqvEcuDrisT0AXTx1fJXDZcj8JSJmywqNo3TKUioOSG794Dz8z5mCggrxB
lepdOsy8iZNzMnZ5aheqs9MDTLkwPqlRWWUzeh3wGy4Be+wwS036Kn9OEa7zZuOe
bxbTM+AZebMT1U2JWLKxA22Jwcs6b+p+AEShcDdbbeRZJQX+ojY7sOiFbCn/wzTX
IoY8gP/TcHvsOMB55jC9FLAMSTExzhDbF9YJ2XDVrg9k0BJKNB9hcaDr694lje/+
SYMD3rbpTX1k60pCahysZW/LKqPWwe8VnPiFi9q9O6OcZB3jzftgFJKT2GchKmaF
2pGLi4QdMKGuMWi75NevbGDesR0Qo8qO43TfkhXh4aqT0T1Ka8ilOKINyNQVZUGf
npNmTDKne+r42IpWGV2xqTxDJacS30X5sT/ewTqm/Poz5NIigRqV0Swb0R/9GErh
gnDcKTJSRl8VXIyQ8btZwf/v6Z9PkZN162Gwy0Yye7bmq13bcKcDwyPGgWo+iCJt
6LLKmYMVfFUc4YhuKtkCYk2scDoalrkdTjLN5Cu5HPoUdF9uOSseXhJoas5juWPf
AG6h9VhIGk8OQG9e/EdGCE2wWGSqi42ty4+sHkb3RkNHW7iWnKDpJzawqpqm1T89
1pNex6Uf0/v/tFcgt7EkRycqLB42psjfKeBTB1V99wKjySg2/rTbseicXX5HVD2q
CN8zY5z9mrqXCIxFCJZ8kFzPtB75skzNpG0j5AKowIPqmIKao9bucbAQ5ZetqlN7
c3G5EaMPTEN6g2DL8W9PTqDUmAWWbzpTv/1l5Nw5WrghFEKiEf2GhNbwaKoZ4zNh
m607G5F0PwdIxSCZEOGhxs8sNjWVZYpA0Cj7C7OiluwH2mUycrLMWjtNy3ScBzM6
EgLFXz1mkhzs4TzH8zVeuoJdP6DiIXhVpe05kbCBa1EoujKO/CapQPAZVqaijY5Y
AfPbYQYY+1+YJZb+irVxDnTHCQ4KV2EkM8wzECcO6qf8t5zbVdm6ULcAvNKq8ZrT
QYrZIXN3olA4PjOg8RdDtMMs0/15ivlU5GM2LAAxcGtih6oUHQIMQcH6yn2SjjzM
ExvlCAASvXGnsj6fDyTixokTKvK/aqtwEhWp14zmp3yEF8dAwao47/AODNs1mPPc
M8/lbMHhEm24ZJysOZAkOxhFYuWALWwoI5kOlarYHI5QWgbf7YazFCCRWndIsCa6
43p9eRfAdmk0f6by3+ukryiGOitvbW2st2L7undeZXpUlVub0Xb6f/91XX55E6yx
Nz3KFe7WsQhD1u9IXTGlgLGVT1mjoPGPSZByt2KxzU4w4aJBh2w9O8v9NRSbNmfY
kHnSH6M+H6jLwVU89hL8kl3ZLN2c/Z5VJmxDOuQNCDQ1/LSZ7vy2o79b5GvFor56
xBa6c0O3+8fuG9fRwMs+/wWIugoi+/buQhSIRBYjSvyPWSlsulK+WT5uzd7NCU3e
/sYdzdwc9yWM5DQ95c1689cXSSl7MWR4+yXHRviSMjc5vcHrZeVoJgHP9N2MG25u
rekxmx34ikMo5Iqc7niIxvxuIaAcM2hCqCmd97hbqm4Re5pc9wf0HM/zOZ92yGwg
v+awsPG8D9JrJOH59JW3Ok4fegEsQTo2/l15W9kK9tA5qRKaTPyJ+A9yRv4wCtP3
XiMqO7AgwyNtsrZ3ghcNz6JQqh4mYwoMBQvd2zGkjS/A0XZNOUhwAjQWhVV8Z5AL
GEAG0NNXXPiPH7uWBiVUuULQQWcaARRQqu8yOC7fj76utmQuRUuPMTq/Y0At77H4
5kUy2tGO3gR5/zgjs9tQvBAHdR2DY58gvRg8jCR0Kc0zcrnq3KFdDhomIjiWG/3E
5xTe8eMKzj6Tt+acBp+1cYzieVgmhc8N+MVaOoINeYzsJXPgpMCW9JgcBczUraEy
bxdcqvIUBlNrkR64iRHlyFHCUkNniEFXsrn69hcJjW51zEcSB9FgyfDZqR53QRLN
yodag5YeQG4+R8l1zgj0/0bGyH+CFo/PLaG4dAbrikV1Sjae2qZHCzwHmrFcaZeQ
XQazFy9eRAM2bQNMTcEWCnkVbadQLE2j5jLR5SVNJWT7DEgafM2YDWQwv+ic5Cwn
ljnplAxBs8PvWl0YSHZdkUdztN1J011pOszDapENEnsFZE+EJ0Oy24cauF8vXiNZ
+lyAT04XfVLcVq43RiqQR/nr8csHf2qIwAQSEUexHX6CN1DiHxYXj3bI4lKW/WwS
4KdCPH2VlCp1BidXgvRI8FcWalNSYa8jvHFRlmxSfeA3XDbeAvnvzDPkLDcGV5qo
oPdXdDDeq94YH5ygZxpKQ8c5G1lmJ5b8eXVRN68fxA+0mLGaXLqwtaKFD3avq80l
MQzLEskghDpNVP4agi8tfYLICr67SWckapZoFW5hJhfLQY/xJr6VivC9+e9+Pm6p
6HUdUm+o0+8+f3jxrXsS2iy2q4RpP56nOtSWzp2Pz71aB0RBbrpIdJkF6Z75/+Zs
UHxrEzRqERDndjDPpFNsTujzwwZtGBZPwCtxiNlnj7mCSqOiATMa6tIkhLbcK1XS
8u9FC+CQu3KVBZqGGwCsODMZ+doThElPvfxpQFc0F+ydYbkRLXpqBA8nI48QogpL
CXo4cKD4qbnZi5SsUJsMkaekAlHA5Ytqt1nFrQcdM97EiOVukzLDIA1efUy0ZLLu
odIKuUMii/gEi0gNi6y/1P2yHrbaeaEKKx+ZEoqkqj8ZDlS80GuCTNHcMDRXT64E
zACMxkVqCuUw6dOkT2EdXViwCfUfzY7e2b+OrvIJHx0cl89NaonhGaifFxTd+Si+
GMLaxWGbgXo0i2TEd7zXz3+LPxuq76yvFYz6k38TDxZaqpjfrgIg7XOosdwZxyiP
OtI3v1qEvdKoh+UbXYGT+39FWU/vlKO0ZyP2xNZ+q3FSGLOu69Mnvi8FLGGPdty/
+frieJnO0S6Z5zktAsnIZJ5l8K01gsqkg1KCjcHxlhJUJsLELxgCRhbeXQal0qcH
v5bOixYmvY78H6YYR6HF9U4B3ztsgqpIK/gcZs4wHTxqo88TCqXId49F+Ew1Gfmc
faekLyl9Bv9x7b+ywca1oTyuwOp6L5cCXV+OvUvqMEhlscLZX6lahZiykRhGZRl0
HbFaFMMd0ORw2nv/q3QKQUriX41r+d+yzzRl0l1MJ4el9U5dd1xvwdtgTPjOqXj9
/0lMXWb3S8vGw/deLOAJt+M4w7cjIXtfPvWHhYO3nqCIvxhOD3YeX9AoUGMUDJzm
9NMUigPOhH3L4wuimKHoML+aI+iK127Gh2jHhVyGKiNnHg8STHEEq86HGbkUSXol
/O4sILsg3Um3o756+ae2S1pWB+uoLZ5OMunC3GzFTcGjn0Zo0OgT7EOGywtjRxHq
NYkKj6K+fcMpr5Xn8GbAN+fzjmMSzMCwTlo0vj8EBFL/00QKBnag5yntdMsSU/vz
4dxQuj2NH7iJovowy7EJ8eEbc7Xiac1mO2+1XZwLTq913y+DdFkCgB263RAiIkmS
i+Xuc0Cau+PtTB1bbokve1E65fQjH3MYS/tmFUP53R2+sQAgZAOzsDZkXFXu9AJm
ino3Ra5Oc6l6z0jzIF92dLo+cmCq+gdAWthUJ4EHDxRM4Ezjemsa3149tIT0OaCx
XcWHB1pMhV4XQO+Z2fmamE8BwJrbZR3ruOZbhZCBln49EXe2xFe+pSYd6Ww15Rt6
mVMfht/2cwE1gEVCLCSXVon7X5jUG/I8ZmCkb/YhX95uDdL2IX6cWugvHleJ3e4m
V0yocceKHTV0RqdZcbcsUvl5BjdhLqbS6bBtj4s9V1Yps3pdD4WfnsshAwlfyx3c
WEvT+lyvfEPjUCE7/v7o30r6xq1MfG5y5cCnZ6JgAjp589Ia4QG46bbyBuqsu53k
ICXroXr1GUk//asWNw4qYh5dXD8aXmq51P1VIcMiHRxT/qjIReX5qb4IZTjqakn1
Mg+yrSqZ5FlGNnTWcOjtnsM+AP06ZkMm/0Z2rEpzkhe8lvJRZPLPOxACVhJEH3Iv
e1ZiJM4kwuc/wjbpOU5yQbV2obErB/j2YcdvdSbf9kYkceXiC4/UHH30vXM60Nq1
aZ/1DCaO7d2QsI+ZFd00ylDGfX6rJK+lLYTPblnJsvg/lcXbXkj9AUT1455I/Vh7
wY5x/AhqgNUU9/vueddX63sA0prsbjzZF6Yg5vWMNKJrYv2B2zGWxNCmCMWVhFcU
FuUn9w/CSY5RItIXHd7SQpjCq4KvqtMXExL4mKvNlrRnzjQ6iFPB235Zs96wgPAV
x3d59AoBPbDq0MtF6gDeeIEZjY6XUaHrbpicVklZlCCEb/+5RfrbAsu/drBz+g0v
0qpszY7UfZKsfvpFdtz6CGmhFo5I+FzyuzDV1spldLcNLitcBfTD6zpPTFmOwyOp
GU/OuXkk64l3sPggBeXxbLraMjxX1lD5+QyH8NYoha+wMhqNy7/SYTeXg1i5wnzj
WUA+YpfkW6Sw8IBxuHgkzNTct9oVoB6QvbzyfoIq1bY2qtOydGNSDjsS3R/0f2+W
gX8ytED6HbvtXqG9vC1MGbOxa5thMp8GIn9r0Ijehn4FDpVMiDuPt+zNKzifaWrQ
chaj2ZTpAB/GBmLialUT6PA1dPOiTh8jcmWi4k36HQH9uKiuvbgaulFe8QR984Tm
wYJvDjSRLIfIv9bgZ0pjXNLdleNXa5DCgylEsysdQbVTUGrQEhQBaXYgyYTpVvuC
TsuBl5oql65t5wEGkNGNzc91ZBFevM1hcaps8i9LRHZx5ZeH4jO4yWo9Uk5B3vvX
85VukRa7skewmcUlrXljn5fmM22HexDoFiaJSX08sI+HdBz490NmYh8oKgejdQeW
Qd/0XIxrRV7qqOrZnfkpFmuXOvvSEerjMMcxULqOdxKYzz1OtP4E/X2BCQVm10rL
nfD0rdHhm/3qLP1DYl+BzzKY0Fq78mWrvIjDKamWgIBKs4Jn1ES5yuu1KvVtUqA4
F8C7W5/Pr0mQoDO3/mdYMMow+X1RdlTXzPoNC7cbntKcH9aG3yUDAaqNNvzCdLM8
ed1n3ehkd6fF4/mtydm1D3EMc/vAMQaYtFs9KLWUEPdc0tSfiSrWyFXslNG0Fkzq
ehqJsZNMTV1TPxOgdidGXS7ad+Q36i27IShDVgBXLolUV4Kvt/OxcWIXP6H3WYsk
z0en+eNQtho0hUXdYu2wItxfzY1/2adkS8JiyH6TTSnzaCexB+PcZYYjH6ltwb0x
JefrZvvgbEby55AOkEX6oTX9keT930XgQ4y+llEl3oHfjusiR6Q6BE6QemJ+a0SX
+LFKkl0cnXvZPOPWNv2AJs7ByFuSy+rFbWewnRNqUgaipL2BzXMpmFCItgGLQGBu
3baJW+Y/m9M6vbp1gmjPxrVRI+3lQ0MAbqrNEeO5v8g1w2ASvhCt+v5q6nKjCeHF
dTLWb6qmUlAFexAglWj1UztnR0w95qDmnNYgC1yUgjMZphjWtOo9kh370VZ4GLRe
gFgIxfc5xs5NpW7Dv2HPp0QQvJwg/e2uNK5ZXTO74EU5tB/gRctOorg71CMApDIU
Ws3vPDBuAqI5OPpwDUsS0D7dh+7OShCJ9zBOsWX05bI6xk5kt08ceAE4nsoSRlIw
MEczp9zjzlNjxQZWt6oRGBCKH14tN3yKVf60agL/ADlwzmaKm9hZ8miLnFkC/SWc
03lrc6kYA6wx1r5EKihm9v4QGpFTvxVwgIu4Eqx9nRIUk0yRslD2rNr7NAqS+LyA
5Wyk6AX6ZH1+VDj8TKAKskjZrhDH4+Voojj4VzUZxtKIxTBYaYrMGzJ4M5HU/pUx
yilxNmhsZ7ZPxJDOGuIsuPcfFJlXFG7sIqLBJsi+JP+UdVwE7NC8Tz9ALNmsbRHt
3Z7dS4paVN8az46vxR7K4SrA0NT70oCNpy86nXyIjq7G6ebs1OQpCDQAiqNQWIGH
o7qm6XYtG3tYTVGlGqrAAR+82ZLsuaEZyu3/HSK3YHfIAo/FCvSL9emp6kLRcZCu
dPq/OoQJarbHS4JBk/0v1R/CwZwIvliOeyoBndDVNpUb/tL8zlzRbFmYmOOifFAL
ZKSsaJQOYzNlC3/aKNrptWRQCg5wXj00CvHsl7lZKxO6VhrcXCgMlY1uZFj2Oob+
5zZpD7U7vgokmx/OiBYTEDf78JzGqo82WdZRna+G0GKsvlfTCc+gSCmmxCO7GyzJ
1fc7SuXuukAHheMrntEEo5DgowRopRGIkvZREm1l+E7v1dyO+YGuwxDGL4PCuaIU
aAhTM+HRqeZs+tcAgxYdeh4jW23EXpZLxJgLaVk1qJjldpGMvLhohpox+cFSMy9w
4yppKCysJbFFDhpMlNWr7arS8hQlxFL0UqGsLfq44th4b0fa5GtQ1nAGXTVLuc4v
H4U6zX8SXETTSib2q1ynTdVHEiukinHgjU9246c7rbUSvZWG0qd6mzEmXbVP+fwp
bb05TBwKCIJ4lcOcnFvzDKf4FYZTZVImN8FeAYb+cPXmVBwcz91ehxTGtiCNuvvf
y221aHtgvUD016RLjD5QzTqLN3cC4Y1NOGsAuTHmCsJ9zIqCRqttnuj2L6j7XKqT
rJf6F0L8eCALhWTN+qiR5cSSvYd3UvYr7+MOmBWz4Y23unv4D+Tx3jHbI4Lg8ttt
g4D5cid5kJKE4Uf/1JydT+7+daKzy9ncOXjC9b33L/uHGDkM2EW/gFennsZUAuCu
VWZBqAdH5EPSoEK9dCXsac5YqiwqBCntsdGpfhmdze/G0Kyeo7ZDRRBKbZevrAT0
fODf6k2pLLwNX5yfFaLk+XvtMX+tkOs3QM1Fhp9nus/SvojY0AEVTV03KS9cFW1D
8P6t5yyg8MziYuns4ojilQXGNl20LMDwgxMaQDh+RVYTJ9do2kjehqre30FzK9Vf
TgQP6py2NMBu8Jxx9/OAEgqRcKPq7jdj2oFsyCcJrUmclt9fQnvcAhhWHeEbnjK+
eRaz4D6cpERhWRDYv/prXwXaYdKW2C4LzTP9wOEXn0pzJuO9bUaTKLWQmmuuTHnK
S/pFniK0/UpbtVPrac7HIKQHUxuLt7bL52UhSEuXYbqz1msl16PAA3GmvXFZCm8+
zCM8TV447NE0xdgV/SX744IDYLsDyljxBo0+u1oI/uhyVt3M+E3a4Tl8eHaPcNUH
x9lS1l+IfUkL2keXMd5Hh15hQrH97j44HS3mwN1PKTiVxHNcRDVDWV+uynRwC3n5
XTU9j3zNggllEQZl2FwzpaVNw2KMSUQINxBtvWwMH/EsaHtHGcQNn6JULhJ/z/wg
rlpwK3Gy4QE9SDpucuO4QDEV7QHZnp1oxrpEWlu6pMgFnjyY1jm9W2Lc71Ckr3aS
laFUbWB4ZQi0xSt2galqsnUk4zxdCgcI0cggYG1YqHX5JfIOX2tYErBUEhggmedI
fUfcfQXhuaAChcr0oJaoNk737yQLw82z89ZT2wQY1N6yt4mKWbY7n+wTekq8aQkU
Sr7UuWVmm+WRCphSyFCy+6wxy86DPC7IeXkC9twRyWhQw4RFeQdBb1bSblmmups9
8hCODNu8cdNGd49AAXZt7rFvsHL/wNEyY2oCAtkyhqxrPCyLO8YCScEE5UldX/BM
Ja1LM06YQNYsIzT8+TRBQbMCCpI5PFAFGcvqfqzMzoKF+sYH1f9iN8xK+539puSo
2uEEaiS8piVqwRmfoN5k2ZNb2WRMkHSTfg249q57EwChDjWcPKftqeMyhnGPocvo
jBwKdgMAkWRh0mVDM1/uKijHJi6JLoMTW4NRxoiPKqAGf7BIfjQyCYYFpBCB8vt8
BNt2DUVLDj9VjD9lgOEPOXEj2pen4OYmLyv1ZpXgf8jw4hZJk1xMwyWL+ZLnF7Zt
rH+xd0n+I21efrm+MJS87Tu1FNewFd9Lg5Ipoi+7HjwbSrqiUmMDHmd545T1Rw9M
utA1kJp0IBSdh3C+evePU1GbRWKT+UFjhw8gzXEtaU7Y9zLottEEx6mVaHp/3WkV
RGo8KkeTxzJcvO7kDG9x9mO3DS01uMzDiTCmTKhSscCp2wRLW6fyXbtjIx+6GPYR
GsGiatTdlL82BxjNeWrsmk8gWes5A4Ax5XyQt+FHeRQxI7P7I0iiFp6DR5UL4fcV
LgKY3Xk7bYpMmmUzxUulWPHSv9X6j7elAKLa23gO70z/Q9uqR3W/yatQnJrRQqae
f/W9qTOneFTJLhru98qaNJgxlpLQk9wJxctHThuFIA85W2NwMm4rQ+dExPwnUYfe
mSiQdgnOAecSB0TTfI/j1wAjBkd6fqOqqcbjXt2FOCsxgwOOC0fd5FtRJcuCMMbF
wb/bbZBNxngR2ud5xPkk0a9HJlu6KIL5iL8sckmsM95xxlakzUEUZGiHq5MQVs2i
G5rjCh4pUu11Onirn9hEasrG0U6EBpwrnxfK8ePHtvN5Y1u9F48cYe/XLTTWZcjF
/wzo/N4e4uxwtKvz86MoUS0qJ9/vVH5nKyLOAZS9l1KHqtzVMqnZRoOjkaEDCnrm
EQH3JhkWgdDagsY0juuTOAVN4l2TuKRSeM6LWGm3iTjfrZxWP5lZdPTXhRAmRnLb
nTslPbQHhzK6cfTs0SrPBTRooT24h5i3fgugRHKMGem7aMzsIR2AZEhs5yXmSVAM
9g5ezv4Vt8E2L/jKi0GZWYleK242gffkLQc8rZ3Cseja9TXRjp//dIciWYOvVnx0
76GgU0JCXChZIcGjZTOlmY4tGUyrowvFrQEcHAvR8rkSXnzKYkdDTpfNmXt5cx55
j/ntAa5TWGPuN1J4tjnhRfo2w+JAvi5Rxi2SmVNKR0MzdxD9CZR7GEMuW5wdyNHr
iXqVLS/LVdBbHFnOz7T/3agU2JLHtE+cj9fJaXDA8nqYFGtnQj6j/CiyWbW2l4dR
7hc5/0XZATQTX4R1upSwPYCDuyXzh+3A/q6I/8r3RV36iie5RRY4TXRP4N3ArlX+
83hmR4oh4KccxEGCoAm3uaZ0w4DFwXhxTpUcXzZc5Bc62POu6Tw39l0GhzNVZaP7
BIMcz++MDTQ3mYrPkmp/Op1uShlUxvZRzPBX+LKbUTERXH/PQiKWZCJ4wKPP/7YS
+cPJxNNWaD/F2VXEGrdqO6iffNrdDUkExg8llRVq1+q5yAKiKUBXKEn3N+KIyjsg
ebg7N/7vYyqEleXj8m2ez/5SbEIfqUClajuOXbcwPGmWjoIj9FRdBiNNf1Bsm1T5
hot0kcnzu5ULiyWHvA25KcdPQYMKLMVc4r9gCElY5/QMUVvZOSjH6SrvICQ//OxH
911fPICnfUVQwYdJljUS6awIVbz8bg9LXk7CM55KMMR65RKqWoOpI3zz9Q/veiHf
PMTj/rznH0I+ZRDXGtJdRGKfZ9vwYJyQLMQh2bMBk5AHsrrjHkkF0AZwe4RlIxun
KLnr0l/GgkLpLB3VjhwOZ9Z2iQ4hyUvhKrxkM8Nj7beRnFl1lqlBk0uJsY+G96cz
lfXLezXd5uHs8t6SyI/K0nOfqx93wfUz1Gwq/QOukH59TLyLsVSvbB3SDuFux2pc
DdLMNdhDma6PiLIFK68zqtr42bm+HM4rkyiz82uYq1PHoBpoS8iZ9a1D7K3u6r+F
Vm+BWWkmSOUmCnF1Vjbv///8gTKYZK/vCAs5bK58Etk4bkRUHYPhqYEHbAxx/obF
igpxUYs71D9wXP7JYKr6vgU96HhVTWzKFY25SrOX9QFGSmpqiOh06IdghXAbywG0
mR2hXRAe+XAY1xn862JpmsVdsH/paCgsC44rSn/nSYF3T0gKNZ9/p3iFJG4l1rld
SrsGJWMzILc9vvDEFQ6a6GFtkZrFyAgCGEvzpPvUeuPMsd1a0BJraVGyk4fjsYmc
SePT/Q4dnYzNLxkxw9u4a3D9hz5CzAQdVc/ofdvGjBavGNIIfuweMHMQXttr42mG
hrjkvpbS2Zd3VTygBN234l0BgHXAL7Bnb7DKmXTkZxSuwjUFI3F24fElcjM6mf5B
ogp0zRi4UsrVYH6mFaJ7rh1hvKB+rt4cCvhGUkxtpKN5GS/J5+cWq+k58GJqeAw5
lAT9GmPUIKMAaHUCXvp+kUHlvUUCBb58Mmn3iFuO59Z/oO5OrdOF9bwrmzHblwQK
83OufzkkRLKjIoV+InzGPOdIwrJku1W5w6ajheUxEiFmBjYNIHxblovmtVVy4oVS
cZ14cEsDQj+Xhmh10D6+Q09FJbcbV8jM+DGxiuGUS7/oLALJIj1dag9q7XoRiPj8
f1WsS+bMS9miCC8lf7K6WTo/dtdrqjFLr7IoCMNS7tQNLY09Anyf6JylOeSLcviL
7UyJOJskX1eRb/8RytUFUTH7+g5BPdpBsd+7y5pgxMPk4Q2gy2bz734KQM7kY3m9
RUTy63znlMXGy2CGafMq6KPahMbwtGPi7a5zWo6neG2tMR05qjGWLEXalPsQgJn2
adpN9vP3FrQ+hxj/k8VL4ZdVCX7MUapj+0oSNFB0Q/aNbI8KQz6095dFDExHtZTu
0GrOkiuoy5fBNm3zlNRJfqza2uymHV3Cmtg6KwZJj7A8EaJItNl4PeVZ+Z26E0IH
fokomNRnidXZUA1t/YK1jXVHmBrnjRpcrEvG9/SRn+orJ5rjIsjrr0S8KkwKqWPq
0OjVRU7qljmXBhPy8GBn0dYf3kijTTV02iUN+3x/ONWKO1y/bnm+fz9+FBd3VQpo
4Nf6F3vT1Wv3MLbaU7YhXRdmDmA0LkTeUGIkyHy6IBQW4zyqjnAF0zoWGTihr9QH
RkmPxz1REimf2B9ZcFMHnrM3ycLCD2vDYjWgf+kpKgQOcPBCjHxw0PXacq9Qy9Zh
LjGV++EfSHv5CCabEjCJ+gHpLtg38b3HEyVqEbqgjUBPDs8npLfFJ3m9wgJ8Ab0H
GYBChx/GvKdMoH/CbRbdNmK9jgRnRtI98M+But7FduRrPYJBHM/Q5baHjTD7CFDf
zoI9kumGDV7hIKNeHnuITAuNhWf7WSWHrOpZvToNLgknnmxbS4b30qwuWm9cdokf
/sAroPXtpwmxrDB7MLrbd7vo4yih6kru4iZP7A1V7zNbpdJbE9aB8MTKE/wj5MRT
twHHYOQjOfYtS57pF7NQgVd+HCJzcq6aEF9XXVI5xHFXGntiS2x4VB+r1f1VriUg
kkOOEomT5sX/Hz9rZG7NtydtzopDy1qw0aLbmNRW0X6eb15GmB6QwPI6wkiwUDR6
nJps9NSsLlYeFolcb6y0HERxlmR0SZsUH70z3FE1GyqGQ5CS/bb3BSTcGSMX5Gxf
WJqudWWmCjf+FYaVYLLMF8DFtH/MuFvUJuLUs78Hi/4ndtcPI852uo6LBXolYnA3
KDnUu3LukTdEKsIOwQzt1NBbsQCJ+rCyl/TT1SAvIXo1RviWl2HWZGDTVeBmXIay
F5AcpxDF36kOKgIGpdaSg6JUA3+ebiJluxSR2KNCFgAWHL0XbMBVYs4W792LLGcE
GShO6PnZrGNcElJohlGmEEH0D+nX2HIUz1MWT4lrR10AaS60aW0tJ2YL44kTMa4i
bJrjh4O7ufUzfNIVLw+dMW52i/NH1tgwmabnx4mBP8hW3taGBlCMApS3uUJpXPw/
gLD+oqSmzaq8q5VPVmgWF+cpOUdMI23Z4WualHv7Emk8Me/Nob/ieEwGvt+XkmB5
7NJ6SPi/5Q16/U4gnomIt8zNFbaQZFXENyVazZz2wkOLW8p9bw7y/FDARkOP1eE+
nGBaLuUrSvtZ9+QdCdXCF/a3dB2OcYPCFwF8AhBGSadjjXKRVMMuuiOQj0fD9HJU
iOZ9bVnbRsSfiK7soemJmgxIR83bd4MmtlLyPOVJ+iLmlrVilxxByqP+MohNdUam
QyzqpHowCyF0XFoWX4R/PWUVQkCKvbvvwgLtvzLHcrAj2W/YeMRf+S39tZ0ZB1VU
KN+40LlzhVJqJOltuf3Hq5ozgFX9nccp3jSp6yoWh7z78Totl6SAxKCBiH4ZQNZv
RXuCD6c+DqWE5lIwCChjJtdWcFMbdUYWnHdwjo9alprS7WP5XtsOjaHAAzeTpmKO
45Z5RhFiA2dRKLhaQXQbA0/U/mm5KWK0WsAVIfLzWlwaWoRB1QOfQKhdYoOolOod
bQGR3PQSU3NryCuKYE9pVqydljtHAOU9/KgSPfCpG6n9H3PCC71BZE3ifOC0W3o9
Hm4bxyxptaeLxRLRrw28mkQ4X/Toc2Dn8ufp7JaXx+4bezRoPawh8wEDL/w6j5Wc
PpyUSKuN06vztoyi4gnj5U3CqH0n2/NuERwAjd77ZJ9M1g68mWquE43G0A99Axse
xTXggv8T6QA6Ejh+0GAjMLaon7/epBcPwwYC/4n0f+L0S+a1UhAlqzGnA/BK+AkB
FLv4zGPSqfuNnNunGh/pN2gDcYAnOLMPV/WyuysEg8abnZLQVHPiie6IAOZOmdIG
fuun95hqA1FNNZuvg0STD2EQ3LXO5lQ6MxZJlyWhjl/9fiEQPYXd4PYo9oNKVkq5
52vE+YA+aasTzqgDzh9cR9MPgjV6h+0QWrpBxC/ZYSSC/n89SM6QFs9tS/LAsDiJ
wZHEKsNkpjUWDFeMyiauBkoSCuJaS2OY5PHnr2gDbpVGt0hrEET5qPJaD9wzJ0xg
5c3NyoewVcwFnGhq3X21ZGluWggjKTx2tmYtwxd1evAlHT0ZlR2qb/+VgeSGg4hs
SSlE4dkvuoEgWx5agmlzqr0CtCqvq1IPcq2cR9Ne+IhEKY3DgSBxPmYnVrPc6dU5
wnAYQam76PjLHXiB1bO48sHUUBVribND02SGJLhKXVTzaff/sVB0CKzUU1SOxJg+
LqoQiftLr082Lr52QlQnUC5pYkGL+CY4smnvx2RGzFCUz9IEI7Tg5pgOdtSy6R8n
dbNX0vCopzyp9mOFPqoR7Y3+5cO2FT6wOT4lyd1DR9GMKYIcim8Sb3Ptmlau1fa8
0fY/WvmqbxW8C8SG628SQnP1gndPoGCOI3IWIwVAF0jTMURjTzuygLjGJD4leyPI
Hd1Fn+W02tAUUma3G29NO6c8q7bB/ThdFxC/OxABujZ85GwaIqtDH/AX4zQ7uXJy
wKXhgcdqSWzJM2kh9hXZmHveGYf4iNjgUZavmRsuvTaWK8H4k3oHTW1QTgV/vjTL
Zw9xdomFqjry0+zE1y2kUuLAl/CzAJX7CJ+ra1P/iXI14EVvMAlgbIQyZS1MFOTh
LMgy/sZ7imJHSnuz4ZQT9XPTEa3gCcQJiNkgIYUeY5WIKX1YqQAdvUaJXvJmoO9I
Bv9OwdFPrm9qlrMTwnvk1o9QB3ThqSeuxtcICbX1k3PyjiBdjj7zfDxxljtC5vH+
7ad8aG7kJ+JBAHE1Eyg67pV8T64v9SpkOhO1q5/KY4CCtgRMjSPSeIahWj4fDi+z
DbIq96+l4GPUCdYIef/Sk3dQPRlLW6xh2XN6I26qmb0kifI0KMgVHRioVwGMQQpf
AaCwPPbU5hOebW83u5IQI6UEkQEBRsGARnkpCikTbIkYN2E8L0RNKOHA3i9sRjLU
IbOwkOGBIrr9fcQJiW6zaUn5FzObNrTcOXNEpRC3RPF3/986xbVDytkgjzAho6dB
H5BLjFm7vqPwQVgWe6VgvbCQvfjn3tdHK2kDjlXB5sURafxfVpytIkVsGs/yXsO7
AveMvifjp6pAB6R39cv3Lf93jBbrD5/ZnH4l8B55hjUhQQ+PbDXW+AHlo+uXj9Tg
l9yVb35hWN+obhQab/+W1mMMX/AKwUgY3/ljr8eX6GXdy6PzFpLhJ2dMzVyx8VpX
KMlkstUjxojC1rbA+c11Evj8KiPmCHVycDAqS6MXniWPtzgZbfA6Q3GjGyo4u9c1
N9Ec6n4nbi6kybjLr/E/u7nNZTzeAcDxV8Ix4R/sWjLA1/JvhJalQaQixYKxqTzx
6//K8b66i5PnjAUSZ0/o3xQYmFcwcckfRU8Ay+Gf3varCtCsW+mkHe83+DfjXU7T
H1Z1eheEKLRN1IYc1VLfA2XuUTFEtUFxOAnvLue2DdB8OR4K2zBJX/C6wgAjYPmW
4D0FHeVfJWfA3AeIX+kZj43abF5F6PGJY95Cn3KBa1LbXOyq1wPZ1HUdgECN69m7
9AIT6qm5WCOx+XNeTW1yxT6Shpgx+lpDvOg0en+5C3NUIe/PVNQ/A3GKczjWAxh7
dKuB6vlFSSfxEgbRS3nmZq2tEcAOniZZpU5YXL3huTSxkyULghj5HQAozmFQL+/B
9ed4mwQgWJSMKHZriOa8j4UngbTkd4fzP23mA+6TenZKDiRpBi+EisgOFx8hI7pQ
71tigfd+m4+hDjDbYGaDP3bRz0DOf7+7JZ/hh8nQe3AvIdQ0qkapgYDgR9+bmWMl
/UG2pTkcsSwOH+0cL1OPL7ak2SJwh1WJnlkeA8sUItpa0qEsuD161eUkxUCk8/hG
p/a2KUUbCJYFw0n1Yd9Kko2DDqRVWCQjtd1Yk/I5oGWTwsJoBr5Yv/Q3Z17H8K28
m3AgEbf8D5P/MDtCvcZLmo9yOQYR9qQUvl6eCxYuRGpmiG5pbRivUQc5A1ikRB+s
Zzr6L6FEA+5GjONg35NsAFvKdIco1QqPX1cmSdmM8E+HGd4CI5P2jTom+rhP42vT
yeufYjXE7RadTCPpu6sYmCZs93nhj3gtTCQg3phUzh4CfavRNpnJJk3b5fHZL4o/
QKijlAbfbL1vKEnidWFw/PHPWlBlsKjuRWPjfFvIa+zMNHq2W3jV6VNkdHgV/2+5
arFhtW+FlyY182xaST9ZYfl8G0/472A1y6SvpTuGucw3hB3fv1pYLSbtwiwVwQsZ
AHppAzQptFdJN3v578AG9OGV9cyNUn3n+XGGHeQ7J6eA3GHh8t880DPbxSGoCLt+
Ho0yZwtQNMx6mF5E9RyFrWMa1S4TrW39cFWGCyh4gKlNnWX76O8O/srMh73fMMLk
ToxSlho4aGgEjKpe4GC9WDjBv0LOdGT8Bcqpb9R7X/MsTX5wGmWMZ2DlCEKR0qEi
r5ptfphCjt/eiUBeI/r38GdGQbir80VpWLfLJYoc8Sxgh7pO3SstN0ZEMD85TvJf
+/r7FiZRMyMuSXRaEdzptGf8to2XRagY9B9UnDDUVuste7atDGSNg48g8j8HI+Xp
JS3xiWAbsdcTq/N9IBnrsfnGkxXBp8m3q4vD4B/6j9JmQnsT+wzeCg6fJJ4ctfr/
3SGDQSS7HhAMZ+/sE4zDp4oZ56UCW68b38p7EJuIBp7wagF+RlsRURNDyweuvqqW
ceMDPyhGeHdzNRS62iwujawVSiPmXPZeHYofwucPHWFdSG0wBfCE8oHT+RbUI3Lr
+mjTh+ciBWT2BozdcqBAVMfIcXr7/EMdj4DfjEorS77LIEz235Whs3qsCw01zLAY
K6bGcqcaIChpfCQdmQmBllBYCHuBL6UeXpMYzA5anSFh/RFDhLpctHLZuJJdjW0C
k0Lz9s1Y1RYPV06PBkyPxYEa/Mb1fK1ZCUB9gRi3GwfeFBynEYurIeBiqgA3K24r
MuY2IJPzcyRWc2iC8JXNY7GNvKcdtKIYSjF95WqeJJEdcSgUtEEi8gaZEXdWC/yY
wMI8431PTT+uQoDgs/1Bl2apd4OW0TVR7WLSOT/x8egrJ+BdPFBqYUGC9sgkYRpT
tlx0NM3jgJm5q+Hz2oOor6DNxUOycY6HEDv60KsihfaLI3hOXpiFEIXR2EsJ2VLB
Lv5pDzSV5EBXYi/Ubc5gtg9BeNkvytoUgQJp/n+Ie8DWmsG81ZLwqd3jj5Jd3EiU
d0pvS+izmaXkfGl59tJAAREws7rANKvroJYuAbrVNey+/Bxjyi2m+D1o/Auasbu4
B3kzkn6lfPFkCjyRMna8ZFpgXcNnmksEyXKRt7RTWVh1pmGZLkOjIPgYbvtrUhrM
1P9xndMEdchXPy7pkeaNxPkaM0zoQkSj3+3GRXWV9SI3pasTAJHLN5G10irxpPMI
g5MTdxWzYB5ZM6x9Lt0du7P018NsM8uTbzCVaQsNZZovjen/AzTz+78n0txO5Z1A
ogG3FbslWTTpKfBocwrd3loD5dIShZNcC0LMpqK5XmWpDYrh99YhGusp+WA+s0bD
7ff2t0btzThdEcAEx3aQdJ2jF6ky44vb0mWYfoaexjSzzrhPO6YEQyz2K2tWx7xX
TzBvqoflvNEMxBjx/1BieVnbAavYrnGWamCwatUQsuloaJQVblF3DxalgacdWny6
1mL8lTIA8jt6TqTJEl75Y7WTqwnh1P9hBrJJw0ExCBSyEELGH5x6g/q7CMHy5EvC
iFYuLXpgp/nzxI2Q6+vHNtRBuBoXiyD9eYKTP7H4DhYkKzDWnIJKTpfOJX06I8J7
qeOBdLIRFmQAg1YQLjMc6rQ9wauLLPHEoVR2RR5zXh8MIbZWfxQibWIIzrpSXouE
iHPpdGyOUtrPNv+91kOW6eSnjDCDGU7mWtVHNEvZYV6Fp9pYNzrC7qUyar100gOt
nKWD0IR42fGs6bsDNqVvWdWG2aC5BiavSUy605iDp1VyX1J8B4gOagYuiHoQt4pH
XzD8ppuBS5oonWF/ki8L8Xt8jGt9Yf0DCKTwleRm9kr/3c+ZLrl9dt4CgEh1f3Qx
yTDZx9kBD7xKjnGwW/u9ORpUyrVI8Y11yNtH4lIq3Vilj3hDRJRF1ADkeZDAk4rg
genZ/yDWBDVpic+y1lnSdN1ZL5m/OsDHeID0REOPv4gzAJOqKWkKwnbv+USCtboB
PNfKBG80/kHZWBWHzbn6pQPsEJ5x6NV+tNC3RL2k5yz8XdmwHkm7MlaCrNN6r1qA
LxjuchUD83cEHWnl++IufnmraNEHpnqp4+bk/UHEn8eAn+moRPNvIAGAmfzIt/f4
yPRHU7aAatOyIPEVJZOmL9eKdohsuedGHMf2+0FaHqArOEWghuENqsvTdjnH4ESR
V37cNVJv1AiVBYyZTbASQCRs9zU4W6l5Z1LpktjQzQioppjaEtvlQZs30fnEo3wK
iaC/fvvk0bfRetVgzYRuA/vNupgiDW21GXG2QPtAGbXeh3uKdgJ8BmJkAC5kKNce
posfGIz3SISE+uMNEaiWL28mXrtVU13PoRNqDyflELJOdxswUitKOHogPA1IbpFJ
Y9YPsI2rmcXA4avgbaQ2s+Ofb1au81RyUkbAY9hNmgejcT8S9fSEnyCa/OSCeMHY
gQpOHaDJRWDUFCIvR1tqpq6ikvkJoBn1SV9uX29E+pVwPbygIQ/791AizLO8LDlP
KieqqE2kGotADdsDASx3pFR4XEj6Tq2THyWT94fqqKcVpm2a2K/dl15qpMxEpy2m
IYjKdKN0Gd31AtTpXu94WPTbGPF+O1maGG7ACV5SZNpj7Q98vYNnBjZnVXdLbNzQ
eqvYBoYvbGmjqkdKsTvhk0nYWwvENin72eyNNaeW0sPuYbxDK6HcGkT/DXEaLsL2
NDTKfjWwsgTHarIbM3O1VPvPer7lPepy6IAb8dOf/KW+S5uKD3awe8TsRaDBevAO
DwQ1hiViITAhkkryPIgMCSdV3QKk3x/IVImdmPss+iLm1JKb2ylMYvKwUxCufrxp
G9SlXb9E07tHhT45btmWBG74NuGKmnRMMDBjsDDPz1p38goeJrOS5kzST0fax+o3
TQADdLxUrI4g6yTKlLuQ278wunG7GzHmc/3p7Enr+R2GBArM/78fRZ7hIu0EIw2q
KomgGS8mLq/hMfLn5sLS71UqTYuZ/1eZvrv9hgTbrdgB1CGXIwKB6dyscitVjm0i
d555DTdnNCKXfdJS+FWBaNa0omeMgORnSQNNG806W4OoqhciuxXuik1AVaB9d/eN
F9cnBuAySni+553js+Zqa8kHO5V40iOqaQ2L6epN+ibnYoMC5YFRYRVZbfvwjMHK
e6yumouwAPdwqHGAjrX9QEO8uh6rjHmRTdtnv7tB3nLV6DicOL/p+gDMx59BJpYR
7AsT8U/mjuQHXBCMl2fUcv8nYdyyZWuJ85Kh1wnz1eWYg5dxdZ495C/sgByafg6K
UXGuVTiAEPG/202mNjcD7XzjMi7JUUl0ZoVulHP2c/GyqyIyylPYiKpTp/M7bcEk
hNRawxkeqs5X2iweLuAPoFwKQ4U9ki5nK4fgGgoB+r0wyren0aoVBM6BJM1jiT26
wFiQivVQjLCKGlkbiQ4JQ8mSiYU7EXB2qJrDp/lVgs0YRhjYpDSX1HWclzFIs3wj
dhzNpNKtuUhWRIvfmEcnUg4pxAHi/tbIo6MEOURobucXVJU79FW9JyetYuo0b3oL
xkg5Yy+U731wKhfUZVsXgKIrLl0FWZWLctbTwdqDdjFSi2Cj20D/z4t1OKrRDzSz
6SKPN7doqWIRI/z0dS7OAlLExY+JWgA2n2Nqe4Hf2VP7QFobuXmE+VetoHl9Kw9y
aO4Tb5ZnM4TUghbfl2C+XAvrT5yM+NAGe6Nq/T+GGqFRU+Ir0LcO4PCQv0HMMi6L
LwYFUJQk9AlZhPDF1e2UmxdrUXp9D1mSKy+GNIop6PrEmTbkaAIQBeTHtv1vh85y
Y/MhA502ItQN6lDrnotB0t5usa/+NXMvkRg35pmTEocOIS1+oNmkSKxE6qOY6q08
Vn5VtE7CbVUMpqzps/2we08nTTwgcCWo5oJspB1yNuEmYSMr6bejxG0PvCity9j6
83IzMptaQZYQTJK5GHEMFJuslBh/UOAHAhQzcRz91WHv+tp6cLn40BoZseuB3ifa
BR8bWnIdUZHP3ZuGwPkCy70UDJWHVJjqOkE1colXh+1LYuYSH7ABjmeaL0MtG6d9
G7Zw99mop8gTAFt7t1sciqNJhZTWpLZnx0piXWWm3FFEbOEi3W7YFjDdfZPx7XjU
xmu9HBk47YwXY8rZo7i6ZjTVypeO1N5NmcTQ0MFmNw22lRobPxDTmdNlx4qqHZPI
bPUpv3jsKg3VknP9Yk/4vdmnprntEBDZGIvOcKMpVWacswdYK0wHdoTwjpAH/cvV
o3moZUHJqUbGZK6YAMDTJJsEqfiSVeSJ2DWIeEIbFX34lqbALOT6GOno6Z1fw4bb
mLMuD9zEpClQguzTIjmbEEXy9BHfguhhye30QDnUxMQ/dVSiVs+H43o7k9VyTgHX
sret4fNDK9b9if9t8UzJk7poYAevAT+/CM49Jj/vxI8eMOzY9VAItLVV9vNhLn9H
+l/hHbR2fbxx2p2bBf6A3iJTfN4thpyeMHOnwyGM5BnOGlTQi38q7x21WrQoYDPC
avtgD98YPfenoHXWOvg3ZZXLHSyG2C6G5CdTMndFYqJeh8ZUS5fVAm5OEklMTWlM
5oIip7h1rUx8Xy0UcbFG7SRi89Beeh+jKFxbuOl0L1tV6xMLpj7vErgBlN8fOi1O
WXQm38ENWOqiAgC1tqWKdYDqRhoSLAEdeMdzQ1D4EBerFyg7VPVzX3m/F9zuuD2b
I9tNu/teRos23h14wsgpZg008J0g1GFu91r3N3W+vwqLxTUkAx6mk+MWIzGhub88
R2lvCnkjAdXYfY3Z0d736CPdwsRVPBB4uADE5Zq8x/EE8LDMss0Yjukyc/5xco/5
Lt1JIMiegWIMe9JKjLLBIY+6SI5Swp++RzzrjGz4OA07rYIZB37UwHqhQuRKszAN
JdDWb/HF3Vfuv20FqpGSEobc4hVzN1lwz8Sp4hTFX1PCLHrVGOlmCVRyxHPjhdvy
IhuyiqNXtf9yQhrDa62LJWwMghvBi8co4VBnvAZloNQjvnCAvsB60DlHRTxjAn4D
lwjZGjp88IOVdaDiHtBl3XErkqD3dHd8IlFe98jIU+ZTfhMtdIB1RZl0tainFhth
KIKKxstiUY+OSo1ltLxhJLRetYObawg+f+48Ht2zKoX+22rSXl05Z8R9k4zvJ70O
SP1gSaucUzTXYYhdQ2dIA1+IwicdQiJk8UCXrMi7pnF1KBWAilyFAF33Bx6++P+k
V4rDg9F5M45cB31HZMBNR4uoxaRqN5vPhgTXwfChQdTIV7zkqp0HRqlKziEz9Px5
Yh7DpfYJETGvPx/2kl0l9VHWBgHhRWDd+L4USqXAml2kRVp5hy/bk/p8ZlHvGcGm
iNIvQYZaYKxYaiBogoeQnfZKVO1Q4FTiZDrKHiBJY3EE3t6E9uvA9FlkO+zEBIFO
0RJWY21h6PwA1LKiBmN8ob7ZiX773xhyW69YGZlPdHLseK8Df7U/vERj+RfPdXej
v8teVHWqCOUovyEqToymu0szFzaueF3vEbM54txhBaxRHS0NH3CQJ/TP5ZxkOu+B
OL3/sQ8jMe9YoecOlwReyc8q3+TOkx1N9EgS/ftc3Zd4yiIrNuB6zZa6TczR+NbZ
C44fVT6EwzpiSs3prxT8R+8gZyTgLPTp2YgOh8jCiLy6oI89XGS7L65IyXG+xEwr
YL7yQUUmyGwjKLTaceygVX76Xac1n8fJw2kcfvvZjn/+a821z0/tqSRAMVOpbSA0
qjvwJlB1w1JNLxhUYDVVJ5YkoZUQqP19XVSSvhkX6xIgJhxDFNGIlslwMwxweJvx
N2Kwo3DfVkS+9h5BJWiVfJZWlTmv5dG3dcUSDYMTS2UVFbWjLPtj+O2wGoGo7jhV
JCrsj6GaipAJUsPR5mQOBAfFhCVomNLCV9VxjW9OO13E9qrzIGBTliWEzTzDQVsC
hk07xdH5/2Vi5uoCcoN0zb8pzhZXm+YFrnNi9OB8p/arZS0XGii39MAuGEo/TI2w
fLQpZVSEYLDAmjTQMzRgmiHVy8RhEoM4wKVa0LGGLjjGBbsi/L51rShdTuDSg5St
04jAp0b4BQhDbq1A5OJJLLMVAK2aMZCTNAgg763TSRhHaAVn3sK6IRK/ZVXoFzkg
X/GBJnUy736kaxlHm/uClToxwQZyPyIIxDE+leqvCPOxyETleMedeyTrMtCpDT6E
NzwzKeeX2LjozWwCzrPnqj4kD/wU42+qtNw9dvl5K79c1SXH2vNGMua5zNUOkt+c
n5WZZxh+MhjYDO/p/QzDsbEVSqFnUzXZWjkk253RfRky2C9I7FxlEzGNDKxUaXOE
/Eh5KA9DGnJep7bFsvZEK1n/YuztEH4P0SksmMtbx464qfT1CWG91CGPmmy7BsCB
rOtuyj5qYz14icBb2YF/ut1rj2K+iRUbkKdUlRXW3CW1uT/NpKcNP3f3Irfua5p9
ihMEyYxdbCIMZfVuyH5eK3Z42e+6d2yD4gyaLTIAXXn9M5wdUzRkSCe3IoMKFOFt
oRjPqdbRRO1e1M7O00EPDCNnWJcxnLg5US7NHFeprwYWwZlyfDlDuJ4AbE3N+XWQ
0q/aXFBScE1GD8ALntw+HbQHYGcjFQbdPDfbR2gptPqdiyJuBPrl2rhSEqOK2Muh
wvd2sj6m7sQ/l+oKSYc9ybz9f2f3rIk5+wUq5w306AMMnBdPNliKaWFoOhO0Ohbs
61FUMo+qDV1F4H9A30auvG11hMDfQBzCh181ez6QnNd0ar+Ta11JZwM4tFOGpQMB
kOh0MBW5lHPTqbVrRaLFuuoQOXFbu1W0ZC8PQ6LgOkeHvI5MtYZpLErGj+37qzsY
e91j3OIrzz6doAOkX+r2Yakz9X4BfFGNn1QjpTDQeGjyBoCzwE2PqUF3xfbXqkGr
yAy7m0qQoZB8+6GtFLdiR8FFdpXjbzQPh+Bp1nuDtK0zi5Hql1f/PdWsmrrMUJs/
OQ+E6fIONVy7VYVoKew7Bfsd6NO1Zis+2Iga1NlkTg4EaEwNF2rmPIJK5aQC9e3+
aSABkpb5x/mCaOhtN4YMnfPblP0DazXSrj3o1bHGhiQFzjsQLesGK/TyVUKFOenZ
PsrCW36RyZUSP051ehhNIqQpDqOSbP0SNefmvwsN7kiX5t5O/z0QPNB/xE+50zNo
MNaFyQ0909IlJWxnwJc7gxUbgWVz2Qxm0R7WwfgOg2dtTSBoNkOy0oV6dFbX4Gjd
mNJtB2enM7YfocVLkv7uv/sa1fbTvlALD+21uftpLbwJgs/rK/1Y/4E1nNzV0mYr
XSdw8kBgAo2OQFsCbNcZou30tk0/bG/+i6oM3RrfXnPHHv/YafNNeCGBs++UgS6P
fZChU/XdLYoKP4ZJyUotDpoiQcxLWpKj2MhdZgEmzXfD5cA5jgXdOnlStfPU4QqD
ERvV/y8lpTXBS5WSac6GABwGZwBo1d7WjMdKagpSY9evaymjET9ZV2hxtjrPP84e
cabzdQEL1WWgsJHzJAPXodhoLKp5WAXxvIvItQOK/9qu/NyS1I6WsN1bhv7eHzAr
ZKa6WN8FkjaQBjf5SF+OqeSE978lrI6MlaLTB3tcCKgnRGEDA/gizCUGFzIheDmO
BFzKexf2dPaWh9TDnE+dzyDL/AFr+vvM5i+dC/lBinQ3/BIGm3Lk3VrIkeZPicKq
fHI3qeTXwlcfbYOdlE+zhiZRsTEUY9XpXT6/OSIdJMYzgWMVa0IR3pHBF8KuEF2p
GRxbNbBjHqecYtrciwhUNhVBQ3XsnGfmKNBOktqpn6RCtBj3wAnZULE4aJmgdOVF
mfwOOAyPFwMBxhqnjU0pAQlQh+QJ6wgmHq3Ynltg5QO9tLbG6Xsogk4f8MyxRu2y
o6h4IB6EO9WQ4BF2srVUHcog/RXQNdQ2fdBWrxU+zVu33iUXa5pXeA8JmdZfy+Yq
5qyhe1zTRG62zDqwPcDbkYCgIBpzX0UOcHG+2vUTUcl6MQYiQ6fVcj+V84D7a9R6
ffTbJ3ARki7JOlVGQsc+xM47zcGllrs+88uwvV4usFkw3t6BTGtYFPrWsGFSHvVe
uVLCyuH8Nut2iHUOdJdiEQZGMyT/myByP88+YMJOZiSnNVYO75BP4L0rCvGUbXLl
sVdQ3kvDCnQGLk2EdQOOGrEBWoVzH8t4CnIOG24N68RmofJPXgIfkeYDDrcuY3Z9
Ov6sF3fb35y1lDq0b1b9j7Cj9gQsujrR56aXuDNTzsST/Ee0OWPRnY5yDNQOwS4I
ul4l+akHqC796gY8xliCtxhPLPYLWWHv0+LLQA4LoDIbwBkrGbpQOp5qqwiA5WpJ
0pZcfOSoA8/4H/04b03N975GQ4+gVeSCSg2vE53zKvKUO0143aP+zKSWdO5wz1rw
6kMJtGuLiSM645jlTxMQaeSe72QVAs9nslK1F6F/2Qotjad77O18kqkGRN8mSPN6
+qVg1gA7/N0WDK1/4q3jtbTX+kIo6G4FTJlCjy0L85w7WcnBS1/FVsERlWpIyYYI
344YTO8UllBP4fRNfGbp7AZwetyh+G6qac4dciaDYqdEvpzhkaWDEqdPw0u5GNzN
D/yt3a7rYhgx7LSFkjZWdZl//kPRWYJfZkWIcGgwv9kWbDybCqm3T8hHOOQRTKNn
6g8zM8yP1px2IhZpxNYqzQxhXRqHeFA2lg8vbyW/XxUfCQwuVoTr56PFbZp1BDoF
0145uSnwa9e1LnqgHexxQFLjjMIeYk45eBuWg0c8gpE+uvyCo/8RYmnzWGOC47A/
v0LDw6jMSX+wp1o9d6RceOVVN1gspaFCiMRszJWTvtNxfOt/xNLQc8FaIXM4wr/5
Xyzlpq8lPvHylF7VLdKexV8r7UTx1Ppo5cUuvBAfUJ2GPEWJjFfoW88QICEkeH4X
xIyTu1FXDFL155Bb3y1g/OUHtQ7yt67037llmkGodTAS5Fo/mc/m/1N5ro67muIO
hWrZCDBKBCROWL3EYyFE1c7C5RoMnLAhdZUNLPnsE79gU4+UbjS8bck9XM6v8j9A
iEbOp6D8nOwcrF7JVhdWtI3Hzwz90a+FMj6MQV7U0KCdlPSMHsDwRaYKypDPd0Jz
Yd7Q7rDNwUbKGr/aCloxNFcfVMlu9xIdRpJ9SDpQqhhB8IDyqLEN5T5+2yWQO/st
tlwtiW2mpcVhT2kLPKNPl7Lc+tkyb5+QMgt+30QcgAKbXvdI27NSgCH0urYBiJ1m
2og/f67dIph9hc87YScyQjfq54FnVqjDxk/4fSNVs1zDtaiw4LfPk9czVduU0E/P
JW9Kgp65RNCfg2Cbh5Dn9tApEN40dchctUG3OyUihwpKw+mriUEzUHqng2/Pzn52
kTI/uPTJNT3t2+/iv/JWudSUkjyMJn13mNX4fzSsDjWhz5BWTlyBVnQELZljhDCV
njKT+eHnoiooEYbGSaoouzkFvfnRbSFgvmD2tTVGu8KYbZanFahf26z+mUZsaZ9c
WK0RB4iwiPCyGpg9sgp1mxTbhFXe01glNCOKDVy8y6IwUnEMaRTzKd3Q3Bs5eL+Z
+HVZaDj/FzA6be1UJcRx4o4N9M5+iH3qsgEwG2A2cgzWoDQoI4ngqRVGyXuQVvPi
6flFo+56Ssvln3zo4i8vZP9Kj/Srwh/Rckon4kgSWvAGwKAM65X377kh3N98/5Wv
QSCUkYy7ZetzRF2GwPcUpev7gUIZGQ6skWJhy5I7t9ENQrmN6sqqj8vg/rXcEvbQ
4tN4yG8yWXqH03mVhnO1lhl9r3y1vAKC/sm5S5ANyGRq+hsd+g/6qqZNUJtlx+Z0
06yOtgJngcobj1mb7/SQEEriIZMSQ6Rbhtm1vtEhZ0Ok/MwrR6YRGAalVPEdTZ4L
IQRUl6h5lzgX8cPL9kWxmHItZWKGh+RbFu5LnrEvoF1adeaH1VWtNUtnqNFoRcnK
p0I9ow9bqek7pIdoBpaYioyGAvM9CThZO+CrOdumlgdpTy8rMId6KC0sgFaG1ez+
gQzDBROLDgBcURsLIdy32Bvpc+Tm/KXEbCG9y/KtO9LmNsrprsY4S3hn3k/JOUOd
/vke6k13SIYdbs2ADNTcJRzh759UKdSBfWnZIa723qDMFHgrXOeGJsxFFSYO2AAY
cx9R+0pqgB7Xhc6rgNNvn5L9mQli2VJPsFPXWCvZLfzDUqxJGW0arRKxLTWo+49r
8U+wRmOcNjsyL5c3lwGS2X9JVtsDobHmfRoqzHL7cbZASPrkSdX8k5/CrVfb16T5
2Ft7Oopu5XuXta5kSD0/NKhgfceBDlwRaZ0YTdjhIFRHGMM9m9YBgwXRHCRgg5R1
q8vJYS+bWW3OuG+1IoF4u0JVj/HkAWs+wyiTY+wcXDcAwO2ZJaE3+gHcqvkp9xnK
iCmfHJRNcQns86whtO22pqeICAR7vtppLmUOL98IXWJno/6YTNEkru5x74T0Ng76
M00hTZIJxRNdVeObz9NdQyV87dKYIp1eEJBxECW7PjkhNi+/d28Ru1cfZJftC3OF
m5iA/qPpQJLOeoBFsRli0lV47OJZezYmp161ImKLZ3Ujhgq6ri1Z1YLbuIwWw1G4
KkOPJeyHQuIDnAQXFLAp5CTo0lUI4BVaFdCMyClllrC/Qdm3bxES+hBNrSukORzZ
FAzcSDa8jb5f8lgNozqGMeMSTqlkY2NJLV3SBFjVafxWWgttTeVwmlTo/K+5Qd6j
VorWsY3wATBPUy2wMXOHnTv6NrDzoOTCrp39QeQtC9Y/83Y3s9N9usz6hhc9NNto
Z8eDaP+QLUHXoWBaLNH9Vbd1LCXcgrVNxMkltajJOhTA3YvhiQZvmVmkYFx0QAF2
AE+dJ7puZM9ILTkt9iM9SlSEBfRh3Z80IB7p/Uo/Ut7NEMc6LL+cvQzx7/iYXHSZ
WSxd1Lfw4p/t/kdC1v2TMYjDxF7mbOaKQ+p5QLyEt6mDbMHGLdrab2N4QqbNYCNm
V+KBp82ErlVyMW3dan7CPzBa3t7eGfR+Ugg3lJjrcFirUCGUbodQmG+/kBaGiryF
fa64/bS2h8H6pn+tgV49F87FXjrVXNPOWJB5tuwofUga68YA85t3xO5y+W06yLlx
jxTcpwAkymL/4hpdVw11z7W71WuEk/pJV4miIOs8q/WMYAq7gaLAYAH2joY5fEgr
osMSDs5+/z15N9uBrjW2WLvMA/NWts0Pszn0Zz4TzI+Q2aMs7Uo/JmUawiDsJ6PB
1/6a9iPRYHYbZbAxvtVGTg5MpUirXOVeKnoPJZMOINGNiFS3d10Qx6EYKbWsg2SG
0ZB/E10KWHJ0Gf7/rIxzf25q25b9N9KmmOCeyOUvs9/AZ6vSO1IX0kWS7ssdDGYS
jEY56NYvGfdg8iD8Kdm98zlKH/6/u5teHVql69r7JkRBD/fQhMUUq+sts77XXU7+
CMdpefow5ax1ugZZd/nrwwS5mant/3RN55wS3RFPXNWVYVPV/zK5mdpMh5BKNkmJ
vRPv+l0dlJZaR6DzUwxkNBPyfDShkkRh6BkkLgqstomZDRDWmIEpdMZMboWtjyUb
jMosIMEH4iMyCrUQrR68+GY/nuraYl5gVAbVe/HTodnUrI9WCKiAZi9MaoilDhmd
0DSpCfLNGTK1SGJHWWiEtOKmkuNy0XFT1aLEIJf9tmN2cPvgq/I98vaVsP8TTdOp
E+MHKFxTnWRkyvYr9yi941uJaTmW+LnVTUxWJTeniV7mpiADrRt/z0BcvYhc+cwN
3MNfg7EO+PeI9mnUb7DchNMMFwxjlyx8VWFYn/Yy+GgBmy+IgPvLPxO3BdyDbPIo
aGf++qR+TViS6d2ifGxEe3AqYyU3cMFc6/QKgORb+Lsg5bwvztHu1HpaNTWJNo+5
pZkloFnpdUR337QdyRSHE4QgrnhsOzFYCHABIC3uqt9FZQFhW98/vkIfJ4X8lCEU
StM4sCkxypNcI3+qpfFZy45q4AS1MDw506duK17MibYMwDvTOLBKM1P1/iukmwRt
pLUXGWsQ6KmS45ZZqwgVrhG7rGkoBOUKumPjhvg/hG85CMORK4M6f0l7mqsJhHII
1MgbNaZ16f8bCqlNQmQSOx3m1OxCNkLz28nHQ3hgeFfcNmBKITyetlTxDd64Bisu
i+Z/3HB1uzo64iD7xrodkR2hnDkGsCEE8GWCVVKMSd0cGJ63O0uEvSxRHg11WRq2
7jaz68FbTkG+yu26e6FHsG+nYvPN6wCFRsD8oai3FSkuLhsC/qnyNYnoXUXB59c4
fcRL34SlyKe7tVOEfD3c/ajwVbXoF4t7VDhY9KWmDIRxpbzITb51IEUUUSdZNBIh
+Ea97VlCAjzSIjvKt9tLa45/Jcg+KJWImPEV+7P8XArzL/8ECkqBHiwcjFt/AQ+o
51KjGSeeA+dwJ/hEoc8TXsDLnghunsT13UoOgprhVolKRA+tlcqZ04TNKvHCnHIc
l1OVcmleTpkKBRQovGE1imbs/k3r/Zq3JlcbLzGIl91V2BUGIK43zHQHw5DIUoNF
fiNp/H+8YWHByUJeMbCz//AE3J86W2OsMtst1KS9vfYxKY/g5MWC1JQhkxBNmZmt
X2BY5nWDTYEETTEhY6QemJfR5bMNSTcSWF9uvKBbVVLQsCDCw0/4SX84QPapZGgv
31B0Z/XvLUdOsnKviUHPNOCx3yy8EyL/P4YP3dvsZz+rwuoh2oEaMVItFAcRiRgj
WrncsrVlkoVE8Lx2EW0kzZFJDLMp8w6n1y+UtN4nNJKqENn64A5W115RbVUY+YgE
HpB5M3L49eRQwed3el5cx0a656cUbp2Ky88tSqh5qc6ASVqEoy4bvqVgrl8JALMd
a20gUZ35dtaFaVb19kjTn+w7cgS8OtnyTYXYEez/nH6TbSonTVgMTJnWSdKAvur3
6Sjery66J0kl8c+rJkCUyMTDWZHXk0R0jL04r27atYNClTm8WOAviIA1pvY6lcvN
uqe80t0zuQQ1Vz2wFUPwJqEMHcvdrRnb2Q/gUWn14tats0k+5evEHYwSVkr0+0vk
lyrGYLtFovINgE9j/POSYSDTEceMcSbsb1NIQBJIOOukf2kKN5kM4oXnPgxtsqCG
N7AHKzZ6etxYc6UnDdCPwunNuxsbNmVUDP295AP89bawd3USPPBJtmpAlayN5F7E
SQvlah5dnYIZUZchcAOMh8RKNmn5LFgap/mR26BR722OsZZ0AlN/xY5oWDCS7xtF
zVp0ZKUXO/fD3RPYrbfDrjgoIJnTGW17qIfRj+lgQ0l0jfUWOCVgjjHicpB9v3+v
8AFSj/N7386niWr4MklW5gnp+t/7zDK6CftvucrhsIFUCo3ssNoscgjvxMNh4jax
wPFq/ALC3Q3da/vx2ofhXViD8CNKnuu4JOMwhWnmdKWktYkeAcujNO2vRkLWhKAP
0afC5DH85mzcuoENZS4rMOTsh9rO6cZlfliC4tU/G2e7onMfLQz7W2jQr3J4I9SE
/JKPZNdToHIJyTmj+nF8Xa2qXMoIoC8dUE0ojjSGTsTu4Nby9/1YrCGlmUuEI3Fy
ZQasj7Zjd3/Dt6UmjQ/Ec5GjYdTAPVzMaOfc+8veKDnyfoHKpmSE1sXlrC6VbvYk
rvvydqU6Q++AeEzZt+AYLAxlg74NM2ZTii6Z/HX+VyF9ApIxDP49I5M64rjlIY55
1dhyR9bm+h3hwCm1f0TqV5J87bVUH2iD0MCauplfhdipsqQM98UO7aVns1BmgjVr
nR7ns78lLzbC3R8LwxNLlccHfHnTAlGtUGmCiUHQ0lTzbmpMDBjWbBlNkW+mzbnB
JbtW6jpjhzewttVSSl/C8yK3nIesEGfjLeJuFCORpSJtVtk2drDbZUwPgr50Davx
pwAQ2DLGf8H+NpOtnGsZ6rqBEl0Yr+qilAc1XjHqW+3r5MRiU+B65K0TqTpiIzei
D94gwiJm3Jt1hFygC1+7o2jpz7210KF5YgfORkL81VP1KcOwae2kQBHU+rWJLEbH
5LToug4CWNuZSAGY4S+TCUS15N8kF8YquIbV0mb55n0p22rrbkN9nYVMIwv3ZcRy
IYYz8uOcHMqshZBLRj9q1Tp20OsAf7w6ompnYPs3mhmm8HFR1/QMnRihBYqmRklv
cd2F2USjwBLTluu1G3F+Ubb68guWNyv1naS5uaKORURYuyjwg0cT2Y/A0fesqjl4
do29M6c8n4O3gdy5D7iAmPq9SReB1QY4LwjIj1h0BCBesz86jda/yO/wvLEQxqE+
zDwDa5J0xLkQ1+abLqiWNp3h67SlnfppQ3BipXwm46GK0TA4kiJcyHaA0AcNRopB
bPgiGHzQIn/QybSoBkNJENHxdcEndvqvWZRU+s/G+0U4sY9BBzUyGzW52Hswghp8
ndp3u8KpVUPYkKTBU2iO9oAxW07gvLK2341TAPhFE10B/gzHAa2fXnEYVovzNPcm
PEkEVys4YxzCFxqe+lGW6xQjpII/GSfSxKP7gD3vMoq5ma6HlhpO/7RT/0YeGIVe
cJRuIEteBvFoKWaiz7uj6zeDNW1wGnFYoDJCwJXSjPdOOpZ5NqyMZaEJdzM8lPLX
orhZZ0oyswOob9hn12gXC7et/6OFcdcmDr9yarpT6TuVI5fN9CJd2rObMzy8lMfd
VyLhQ/XNt66PXnM3I+fSmGRyGIyOytOsS8WyN33mitTc5vsc5WMtqC3jo0rVCdvm
YqVl8BD2y3BJ++Rt01HglzDr/vIs18rN5Et7X0/bCCqcj/AxZQLUc4AbgCh5l4Dd
6PAuiBBQeKY7srAik7Q0crQ1QyfrNTCv9H40R5GAuCe8sDHiUZUnwSkwLYyKOYAq
sg+NO0yMbsXPCIbJN3oecjYEpbOK7b9P3/0KIuhosbsNgGzQE+lVJiWMNSiTAswk
KAaFCEW9PT5/ELp6Zs3PXG7syX0jHmrpSIfxVTKgwib1nj48FFf9uk03RqQWav81
e2VpS3opVSibeWn0AqM7TlIaj20f2IsVqNFiYLsyHbkjwbZE/CllHgdyNXXtyu4G
tWfXIt65vzYsjVFBiyv6FITdIkn+6pwlUNXTLfUSGL1Cy0MWd+H7PC1Eo3rZxLQB
Nm8u1/P9IPNSR2Z8Oz/oD0/3doae1TH4j2Km6qTbxVduTE93U4tcP7LlRekaxPyS
7T+s3enSerTi2NlEicDpvxtjBs3QmRQxrr1+UOmEA26cVJUWHDAulXkXGita8ubY
6HdSqetiOV6mET8ekVUUa10maYErP96WkQbeKq8J5xtNtC1rrIXm5CWGYQvcw8u0
jutd8i1l9A0eGxTMxRw+stXeTMchNkdcU5xifvfWVN+GY4/Pu5hEV7/ktBg4qp2A
R+EkD/KkV5gUmf1f6mj/ury44uJFcXTqm88he3dZng9HOK+lVY3ib9nfX/0ywnK/
Omt7XqN0euTpztRd8Mxph+SB1sW+h8ldRN8xDfxiNnQxdVmOb5jSmPsKnLzzOTvd
3zJPjYuO8gq2I7im5Wk7rkZhppF3n77n3Pv553BxvhCQPGVRvTWGFXly+CWHugQi
Jc3tIHyEpea5pIZPi4+vpyTXHrh310tOt0+VLjV3hJI7pe4xTLmvyBwjHNyFTDdQ
/xGun2Ywdh0Q2Mx8//RmmhLosTeX3cR2ZP7EsPNiVjRmZipcFuRp+GH+jTN1zm/R
tQ3CEaRq9mcf2Bf6lG7yv/QlgxxI5hHpM28u8+wP0HTfufzqqFWb+VPGeAX+QH+L
cCTdCGGaUkivs+8i1iTWaKvEAKrUGnOvQtJHcUCe5euTNZw4wcSSBicNjDBE3hGE
pdzhmL7M4W7RvpZMQKCB+xNa1O/nTLKE/AymLrgkeECkJS7HGYeKxfwLFxkA8nWL
LDWJbG6FlHIc5gX3j4pqc1M1IFEXNsjl+znH+JuXoUqqoxlo1vPg2Kl3NVXCP8GO
Gqz9NgT262k+l9ZBhFZbdkXwzIlN53QbFRQxb6pth6YxGYeTXl2HmlV79BXgMDXK
yuQ3bmBCG69eG3ihHYf3+DMlzmAgHpWy9nGQfLBlUmFnv2S8f6ElrDoa+kh4sFLl
hHSOPKWCjPzdsm6VwEqQom9wr8KOlPKIX5yrRbKLB1ihMo0zQPG/eibLY8yhorx7
7aWK9rFoLMX8fg00pZGhTSBgF2LLVdmEwzSEnT5PN/Y5bJtjcBGesibnpCBg7lhZ
WSDPHpgLW22tHOkeVpVbCCE6amA6erzLzUblY7Ir5NArWIJ7xenocsSb0M/qKQ+X
A1DHlkNmQYcHIdOGTI9EOMKrpQSlAhh2XTySrCQpnAK3yOGUZ7PFHaZILwzGzwKP
qFvgDweAFZQQ9UviiIMJrBvYY2M2GfI0Omf7oFC05rHm3LjNw+KFVDAq/Jr+VOYt
XuReK2LF0HC5GMWGfDNOBftmIqKnNB7KYcqUfIRm5wWhptOdeHkV7269XJYBhN7F
eyQYVEtmbk0vndntXaO7gZuhf8KFnYdQNvy5X6yHMgghnS/Wg0lLtPyhZO6opTMN
I85z+JG7dktAaLZ8oo7ahfjYKVoMHiaqb/x7ExiAPsZ/U3jnIqPkd+B445AafH46
NAPMbfapO/8bpBLyKOZp8u7cCVPdXGOlpaAEdRv18IufqddcY5pynwAnuWOjbaKN
D7q/nO74No+g1SAbBBnp3zC8b7Xn8oQ0jGPeHxvVCT7BD0ODj8jAnFsEJ+qkilzm
z2cX10iMcKcyYuQ3jJaFPl9XQlHIuMHKpRg7H+OpnRJrQe32rDr+GR0eS/cri5FX
dTj4h2wKG3ahpZazPPnnq8EzezsDvn65D+8HK4qm2HVxXXcvx392pIkdodW9bzve
qDIIgmlIwqkD4xQScPePJAC+eLSj5YZNnNaGhc4LAS3hr25G0jwcSdY09kgc3djF
fNJZyoNy6owhXK7bTm7CeSlhZxrha5IPifsqcFKt9YtfoethCBi1epntdWSGz94c
4qD8oIzwHmDMPP/on91t6HGkmO7PS041eSeYf3YUM+WJBDAMAghHjKu9XXhRFYtp
B3CcjwRDmfNo4ZZALS+ZFQ68ov2fI5I8DFrxQ+tyUaUjIe8IpqxmpkFBIFU1FwKA
dWP4mlaejyo/l6aMY3CLhB4KFpADxqAoiZlrIYWwQWeuAj94Q55h8eh0ZdBNQrpL
yQyYExIf5JZL/QpjBAin+UcC9IsHVY6CoUZa+AxNFUrrhYy14f4Slu88XjdK9eP2
lrbPt39xVSs9Z/ZbTHPTI8PMvz6PDcUjZ/ZrvW8F6QQCrfF4oMKWOPzJMh/1aZ2g
znOCB/Exe3XGYBrXx7mfLwdEEJiEUTaxj7+ZAYhtUM6CyUVylwBwhBBhhkwf0Q8C
H39FyBbfStat29y6mUBoIf9Z8mGEyYNCGS/TrqcW7fWh0QMLRTqKymX/5/I6rOre
Lazq1XPDPZ2R8l+d43uA9PF98mfOcliG2ZC//YCKTEpQJXW9pb+VnciufM8ULldk
NPj38uIKR7Jowa9bJ0GeguZxzh5gAGBAVLw2jGcKjoQuEVJ96lre/eAynMJlKFjT
5ZJH4H3QCAgteu6bbR0/eVI5Uq/2QRWfYkGVc8SSbJy3nznUbfyriQg4GCqj8E2W
7FOVI1DqXgtrkhf/gka8z6K/pl5TXujZp+mbrZC++wk2vbAlj7tBoKy+IOP4e9zJ
HZLgSaUG5i9wmITQ6RJG7dUnKoZ64duEt9xIA/j2w4RB5vKG9M4emSpul7e3xyKq
0wW9gISlHca+yb+wXTTt7dttYLH+H3puGHnLrr6GgOUFt8znBneUoRz4JLST1A6T
u0ds8kVrHkjPCemkMkxtMwbak9BrlhHAWOutPX+bmKr+8PG0zctuvyqO8+Parjre
FFNgRD5GkRlUKKrVQHEShL4lqydFrbgl+C7sFgZoKzUZMUzaSHEZVJGh9A8XvDh4
rzUDZJfPUmfbUYRgGs05OsL17SeSnKQLhZcfl2bVCzoMBdwz4Gim6SGWkkJFlEIu
de4Uk5o/3VyHXfD7VmRVHOBiY1P1wziWtd6L4cTDxV+a2YvbWXRZuqPK1HIGf1Sl
Hes/SU0H1dXanEmq+l2KEregSW/UT5NNFurXEbCpLepxuZbxTkN4Qjype6Fra25K
2R6a2+6XGYqCT4NL3DZyJ3w/Dhdp4jcgmZXv3dtMc9iU0S6RPoXCAZTK/6Ox5/w5
80eIJbA7Ec+lWjpVTnNzDfe68UfbW7XXBGi7qHlT1KgpSYecpTgsoKFH4IpfmBvR
TUuTNJZSvNkGFOovunelt35Ks5IRA/5A86AkmL0U0AF5MY7BFd0tz4FaHAS+LmpX
JQW7JJdKtjA7+atiAm2B6mOBnoCE7kC+10Lm4C+OSDI2pFwuhO1/g6iRIFj5cbWH
CLFJ4HumwxVninpsOCRUmkaYa7376pxr9CDAaARjQ2zkRnruCnEp7CgJHW1EtBrg
nzEh+KppAK2urrvP8TtnrytiOW8c/n7EDOGghrWCKS4=
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
F8+kSBpZN2vFIWU7E4EB3dneuxZN0Fvp1sylhbu0cSroO/Ln2U6YxUa4ngBDxJuM
VtTpQmu7oW0gFsdv8rN2GCjguOhYvvSVQ7J13oEsU2ClPQOHXgicVSh5TV/axd59
DbtuSvspxPqn0R4A/GSWDiPNrTce5Cj9J1blIQSzhwXjls2N6MWiZ+Gc3ISeiXOl
+1ZWqvOM+JRHbKgddcfrqbwCo2slXarN43nAhDQDIyZ9vUkM+EAWMwIi6E/anxki
VNp4OVdTXP17z7sSLBXzasOoh0h2O9CGCqTK8S6R7LhA8DEuSha15k4JH7IKkGSy
p3CwVSCFmdyc3VZxk4oSJQ==
//pragma protect end_key_block
//pragma protect digest_block
4UEcnSP24tDzxckxXYwuE2XWoCE=
//pragma protect end_digest_block
//pragma protect data_block
NY9SCTpboAVAuHhuX9ScH85IENmFkJoFfz9bo0Atf2KVHHbiYu9vy84tWjiKw8km
csbyx6yBj3av4GF6QxC+/qXn8au+GZg5RJS0RVCGHLT8bp8MYZtPpzFytmTndUPV
jHMuE/1XFmIePV1r1QDN4N482kC2lwULwKQbo6rX33hFuUcVJhdcQBn/xhscMN8B
+dW/682qK2fZDAsEJ5J1K8whqqbv72e1milrp4I50Mdz1KBVmlLBtvA0/4+vs1+k
q+xIeggZUTeLQDlY3fN66vxjm2vZmWiDWXr+e2QS5D1uke/RNxz3P4IZ0/Je0ThI
9V9nUbtleck01PxuTk9rDblWt1hnMpkpfeEm9UtEgUiUJ/bM3qTvH+mUUuxzC4Y1
+tgk/XcyVv+KpEwfbCsYO/B4BJV/YmEXxorcF8uxs4cmnAuj4krK4d580Buy24oL
ZQCaw3spsiDM+K8I2SDskdsBcR0Rv5M+ebJWNUivzc6MMdJgjB/H9eKZHnnAJ5En
khumWuAITa+lxtvZHzrMjZBA+kndpA93iVrSUgQMpSpHu33aipQXMQwQvtJ5OBi2
MPZZ9pNwcQfM0VLXEtW8TzQZSax540YsEOOnqk/o6rBb4MqD+zva+GoZlogDs/rn
NmV6vyAMpF38aI0d6Ry1Rf5Uy6zxHX5MTXlCDnFZFyY7DEk/urPlWl8bkzIZ7wvV
7Nb2MN9YmEzbppv0sxyFP6jCePSiYEIK3Y+JZJvvOv0p+H19MeTgEuYz/fv2n89P
EtZ2taINDvNwlcol4f9HRWAPtuN/E8hTwSzxrZh7qTdRTcFbcZwUC3M1MoQ5smC1
jbhQRXEDqDvHnUyOhawfkzuPNsX+Ou9fN1BGECFJhygmWKdKT7sBnbqPypw1MtJP
8xl5jTeQpPGylRax1ugsDwqBARFXfGdAm1SOENx6mqyGTcEFAmZV2X5+bH/JG86f
5rJicRlBHrZUHv5xcT/YbdngVONllBaC8mlLG9COmHdtp/hCNJSGsUNDtYl2xRmF
RR2nWLA4w5Kklpl949LdOFgC8AHSH2h3+bCgZVsyDN6YRr7NKvM0oJlWaNX4m2s9
m85FW/9E1aOzPPw6X5v3+esOGcZEE3EW5lvwXsNRySiqMfpHLnca606ykIwHw6W9
3wgsSOJxdYb6wI/vKlorpWLxNfCI0C8t8yCYWb2rtizdZ0BSTMwBba8dRXEPMDQy
Nd/nD6paByDErGKXH+Is9nqatIXsRvFeJz+HT1dwKAblRxHKiVebjLua/YIYfJYA
ODgOubAFMYOVYBbQW3fAyitJKZEh/wV6YeBXeoJ7hLozqS95yn9Lbl4RFrLPxF2G
5tRnL/PCrlE7MwoCF7vf0eBYvLYlwb/SOaGZDEXlGkFaiv6CHWAQzeCxFsRrKgnM
7QF5Ubmx9VztK1oLdPVnOTgz406Pg/x0b4mOYCQfFQ2aTl3Od77wwZI++GPiQ6Ez
jVWrJ1ryeWeFTZq9UCXzYUex2I+rWGaMes+V9jjj41dIUR/5ZDbDGc0i6azTWPf8
i6t1zriw+hqKHCKqm6E4EGuGcE+mKKAy/Z7RK147qZXwooLkNTRULX4K23GAVSx8
XuYNreCtvYDg/+aKBYwvmXqyjSkIo/FJo7LiSAD81NxYiz5bNOrnNumTyzZFcYGA
0HCnIRxuiWYa1KRDBkUQR4r9EZt8u3AxOD919sHhK09zwvpTDd3SgZ1F5dB+A4TJ
fkPSKWsGldkCY8/7+Hw/toqd/MnBfyO24EOzyNfQC1q+Jk9DUiWY/4nywRnJF+wa
e1uLQ2wOMd4v7copGSfsB1RwkUVwrYi7IzvJk7DC60DdUVc4hnIS6Tgba2HLx5RV
ceJpnyacY3YxW2MiWqolWkYwTQ5WJttWW+aELQmMEL48bbRPtK4tVBSz3kkTFiVJ
GGp5KLC387M1RiZ+hAWgmgGyGFVuSOH5inTZ3nBcB17PRVbevNu+AaVg2xJSMLQJ
GV6NfV1x1GBP2AfpXNRRFRl1k+BDxtYRyV6Q5nCF97zEmZcttiR9ByyAEjEZoM81
3ElwME1BPpimRm4trFhJpfwCtHp/R6HCAN1LtDT3TgWAyKLpCweCkroTc1s4suq8
y54etC3Q9X18b0b2Z/LdDQN3vhE+9AuRgfqQFrAzkwzRjQOZ+yznhav6v2OP2hd8
5lf9dWscw/W2nPC9HJUebhLB2LZJ38MzeNw4y/NiEGW/mZp8uNYf45O8EMb5qKJn
YGqNHwrNPBMbBS2vncfk5BcDdrVigmtNBBu0mbtVQdOJnxosFx4LXzHiE6VBOP5L
KZaOrc3BNx5tHR77qkf/CaSKRwh52nJi24oQwia+KaEh8PKYMLnwBxJxRnUBmpr5
dG34bbLSL7c5NKKozrJDvInmoiyVFYSI69VjRUBShnzynb3T++ZGNGqS3JFuxtoD
b3CrnuZE6R0h5CBfV7+NIo2ctjofzJBXjdBxJwbbEJenRn0pLRxZjorkjkATmjve
nMcz382ZVLZ+8PHUACqcWlnaQylsdQ5vZQrijDMIzW0hL2s8yKlszWqdz90rhI4j
sBJe103lsLG1I6Qs+uFPPPKTDOOsSN6yIekH1G27eo6aSKRc7J8SfDKLShlQgVE1
cwrlPA8HUivfxFEfGeNvDxxkDlMw+tUzJ8uvN//Kyf7WXt5u4jKlUM18OA2t9nav
hlK9DqqZSu9SU2tk/oUbXpi8pm7kZVHic0EwrxSYcUsXvaFO0IRVBbJYD8GOTmsD
BXqQFEAZxUI3ah1ffGZdn2xE6TzPOUD0tgbMd9amRyV1ETc0hLlCuqAdLTxPdCvR
5dJBcDd4FFY/n/Mpy4C9Lk4EGCLG4nsrxUVlQo8bPyUK2cH76qkmfMXCoVQ7bVJr
ENvHbYSFX3aGqHAxpL5cHTCzG6muPHymyfzzDLJF+oPhOUX4rQ0QuCiDvkW59hnd
7v15Sn9sUndb2WtyfsRcYX2vb97bSqZsj+FKAPlnkq4iU/EZ5PFWxHIS2JL7HEHe
v+eXv6iA8nhNg39111kjpcRNX/4adDmlBO7mYQ6r0xDp5WL5YYiMj0poLPY+ttUy
fmimBjAYWKxk8HUe4xAsnjV2uDw8ZwPwwAp94sGCL27M9tvKM0qiQ3JE9eNplReY
rLqYPmE5yP1k2bUluV+K4Atgsdeb9zEW7MhusbjR1bjaiuEEs8PgoTcXkzuHWojg
13rpmTOLhGrqvx8qDERoo4P5Z8mLn21lcs/zs54jI/tEiAKPemAv4WYXMFSTx2/n
C5ml1V6Q9nw7vRSkhYq/ok2DjZSCKOuLRbCK7I4MmSrjzpN9OWgtI8DLkUSggD93
AqPk0nRYo4F3DltSU4nta5SRSZlSQkduiPcjiJS9X73GKoLw8pSxJ8opINhieCZV
nTlIzU5o66dlBCHcSHRSnbSN5gSZrroSYiHVSiS9xcBWqtHsXHLRYnFTlR9xoAgx
X6MoOuYrWrZrSYuQVfF2pHeKGtSk3H2gNDAMVKdzZ6Kpa1lF4mTKeRFsRpRFO0FT
kU9zx4E8ZXSsFwRx0wYuKqKIwNxroKOosN+S4Ei2aVKWbKOz8xN7+Q8HLeTe1L1k
44D00b080KornqZJddp9Zq0gqTw97UV89iL6gQbRUk+KNqqQmvMAtjwO17zHsnc0
zIC7A8pf6eqHnfx9+q7uoCgI//ez6ETvB2vfZTAbENmm3W2CiWg9v3wD6Z59PBdo
GYUFGa3uEnQc7V6MEfCVjPxW4S0FRfyUUfSHCEvx4Ms0hMAU3wo03KFRTXtKvLQC
KyB1YjhLflhsestzl4V/HGHZ75kjnxvN15GqG4b1RjskTMb7aosaJTOyjCqfOf2h
GIbaHCGOVwtw/cyZdmfphxsHpuMMZ9Tl2v+mkWzLxIIoGQLCWrl4Xjs1h7exh5NU
PPO0TkIoVcrGlqVFMSwh965yQ9NP7SJEEQhRicaEfmZoGTjry+y9H8PyNZLMLmde
tbp860fS7ujZfVSf/jLRBb3IFoDcSQfCecburxX1xGcXH5OEVaJPfRpIx9X9Z7H1
aD31U0v4ulz5IGmCKCjrS5xM9YuBNkkqkUEFsrbw5Cglwi73auu3vuhJwFcFmDL9
ABgWPFVeEW0U4DJJlZi8FOrGyJoSDT5CJhA3ScsUwnXomzkIHLM+pDTwr79v3wlx
0SdJvXmMgn3xv0HdUMKD9Zzt93tnew61r8b1yWV3Z98+C/UFSJhw3jMlz+05OIL5
iFvsOb88wa0/TR0MU+kSh1V+uXbMdDrQxvjNx3NueenPKgRyS0aRT8QknpmED5t9
MowHUt4iQo7+rSvXW3Lt5a2C+DQw4oz08Wlfg6aOl4CGmpwMI15ZweTRNdFbKhQe
hs7wL8XhoMPb31zzdK4bCUBIUjCo3dYCgD1ayA+NFsK4pHoHcmoah6wa/7sWGP+j
BdCAJyzwXI7k9lPxFjIM1q1OQ7RCT++zRCG7wpWoOF7bfM9AnOz/7A66VEZ4fIZv
HQMDiUA+ojlp3AiUpFFRM7+eiF3Y5pW7s0f6cs+XwCz8NzAnWVbYRaEQkB3yLt7O
xTj8kGCpSskXWOcEeTnwU3NlNGO8y5pL+oHiTTYmZ9Ebari7fRBYLzN5vg6xVcG5
cKk3FzYIUpbVYYzHZPCrNgeAE8o0cha4vtYCP/vzfsfWntBsJbz2k+iOgLphjdKE
+q7xwSQsM2AAah+krMoEGNTHY4NcO76sU7PnmOio6Vz6j3H9U9Ba89W/8wFFs5AJ
VB3Ixxda5DZltpfXYgqQV1+bqu44T2DRw6IqB1KqB2Y5WskP6/+2RZukEunl2Nw0
Z7LLAwjtObgOy4UcEp/XI9YGBnasF/nzrRHcdC/qGvwVmGiWR/C3Ce4I1Zuk3vIa
rPSG2IMq3KdsznQ7JLgBrPY3oKHzlcGniyOEeAsZWs2gyZ6DT9AuTygghhIbqKfM
EMiwzD8MtUhiMkrJssTKq3leDmzk1IEf4N1aybe+uP7vUXe/TRjxPNSxIt/Bdkp+
cU9gJbX1mK33FEhsgEZYIUG6Dj25TrNUfaf7dhAbKoi0I9ysEaCji3Zq8Hm4SyN+
4wnt0usUpaxlNaVzqgeTt++9N59aa7XKvfYEoYwnYHPs0BeX1R6d3qUeyaoyPgBy
y06qzcLHi4b+Mr/ajMcM+u3bBXn3oMRBGzuUFSs33W/0LUsgHO3I7QbWgrjKKImB
U6TRyHGRun1PyKI0hFk/cwQ2Gg3ovfW0dccZupGy9oDHTQgtHzXsU3JBCiiESakH
vmWyvykpBBRWiLF5JbD9u+eqSw7xh4OqXK+h6yXgF8J7bap4YMEUupc2AY2olZ+W
SslENb5XHQB/LjrRFPGKh/23SLoqDDTBk51vexxtsLoD8RGlPaDrAgZPFi2MdQa9
tU4sTxdYwNoALORhq9MaB35nL4KGzqPFTMI7wkUEJl7w2vu09I+/Db0DPhlpjmYt
9YWePqZntXay9ItVfyX6TdfdmIRH4c2Hi+qaZ/j+j/LCTdBG/QYYTGT8YYNJ9FbG
rli51Zzt78B2MwCgrZXR70qfVVDh6RTWDtLhAjvktQhB1DIiGhj1N6DAVncJQhUC
sZ3NVDX6P/4ifeGEyaaFRJjsMVdDG1MkI3FBBaP6je7GV9M0+5UKGx5UwVuPax5h
0t3CwUmXUm+gf1bHQ2NRirt0/l0PMwXk4qvNXSdCOjTMScJuKicItFBJCPGBtuWD
auVwzLylVq/AymdquSJGnjirotxyqoHZzjfHCe+yw74wyAY/oaa35tZFOsbI4sCb
B3ia++sZJ7ZorDhHc3PqQF7eyt/IJXvxwoL/xbn9CGGi5PwEbtl1ba0BCTipwyRf
AZf6M/uVXn+lijBLSAWx30FthlxbBWLHaBPmXTEZJLGDc9oYkYRqkzFEOjYi0MGe
08NvSjb/V0pHG+cgk9PscYeqm462Oiu1dw5xSddVb+WS70cFIS0nhmR/hcYeUvrY
6L4AzxyUhLE3SNuE4qkUbC064U5V6LiPzjEvydL0F1yfFlJiWTn34eYTB9O0hvn5
Dxwz8+vjQreXQNZSglGM3o3c1EvqTLpLtk/I32LnuctPFGyLuw+eACSE0NM4CXfq
WMHv0zqwe2Bbpzmh64GvZQowGlP+WdTM56Xha3chMM99q3q2k14mdBBwxpVGXG7C
ghzG8hlhIF4P3wfiDcQGkYxgU/oheN2ZCyTWt/hasP5k9dUHseVOQz9BZa0gqMOD
TCUyaQXKRY1NWHaPh4dUf2U1bGOEsCCtYiEUd8aeyVf6H3KsMqf3Zet4nBbdpJ7Y
U4G0u5SzKc1OhuRHGNHCTYYQolU7By7p4eMljc/WbkYNu7kt+in2acgAfNrqLYm7
MUmTxvvjbVd5HqPJpIlyRWTDJXwzZlr8O+G+enHJRJiBGoZud2qYgX8a6QLG9dGX
PZgnjV73L7lo7wBpwM+vrNPjMBwPmEl16Ej8QmL4l8zIPPUl2vL4fgNdMm9of/Ia
QyJTLDN1AbQ07IjWcMcJPuA47dMLdCU25z8d816Om/Vh704/izCiiwzFrUT9RAww
cF6PO6jxaNsp70uxL4hr6coabyGOBhWnvmLuhiAusniYmSukJRam4gPv2va1Z8mF
ntx+ekt/umHZfHDz/YAiQ4u+SwUo2wDt8wPjXpkjWWUUbh8eVKP3jBoJ9Rl1ZSQ9
YwHs4F5+//ExbWx2OVNVdybUR+DrJBE9XKIel7TGxNjOGY6zRzY0dNmbsZ7qWhM2
O6UxHE+vyQIe79jDEpQMr3ZQn5L6P0roMaCR/FOrJ+SHcMihtgCrpPdzJikxeYT2
q4XWpUWmjBT4D/HQvmKRUfZrCDc/q0WEVFzCEUQ1TglkH4ck6JfNm9HF90HPYc3n
9NFhLy0GrZhHUYYVwqkik1ZefM71x/nd1jbW+zvgXK5bl6azFbnKe/mJwCrPQsWp
4FMLz6hnAqgTNelMBRpBTapSV4pm6l7QcgUEFWKRFkXDs+e4cTyvDYqvJv8eHVYg
hke6CtAVsv9nxK8W2xwfXsYsoSTNDWCcBVZkG4n70Ot/yS/jL/6bKIoasE4ScUSg
wQCXCNbp0HzQ0d2lVgdN3nmeNTsoinikXZAH0y9no4krMtzBUiKUT2C3uSqeULZF
iD68DTlXj40AQUGYWx4A/stRNahmwIf4/bVn2Sn19VRn5BF8NZ0+5aJ9KCW0Tpu2
w0Ik3NVtUWVl2RGTIlazgQPhezAYbojHqz/UwkOTaanPu4J6LrGwdndgsbU63t51
sML+aSJLf3/3K1YjjD5TZe8YTe0DIl8M97IAbTr4GH6Ps2LCmmhvdbSPZdCl8qLF
8dHcPji8tsq8sJ9wjpJEWu1wc8c7Ptn/vtcf0OC5OyecZgbwSI7t1WwGVlptsjLs
hgRuh1Y4vuAWTXIe9eGsg9cECUOTWGUUUrNl+tS/IDO2tyc0v65oSRpjHUtNaeAz
cuShnEX9eOWTDug0ODAChODApOUtyJgTwBY4H9Ufmbv4Jg4xdo7MAJcFdqFdtMU8
K4XfpJjyvaYlz0U5L9vcKChigZH8KCWo+fiObIPTONFZX9KpNuucCAPbd7JdN4Rk
Z9NjRvJ/cXYadm+OejbsYMRnubd/iUd1hQCkF3R2en9fRabQeveNVE3GsPejKw9o
WO4YICB4vAnJPEDuSxhHKtTK4Z4TlNY33UdLW7FURJWYBAk2BQQfWnpxrmEvh7Ii
AJkYgGiatapqjuRBsBf+k11iphkRlC8Wqhr5OPA7wURlGsp7PmrZIJcq/ejoYFlZ
XSFIFMwa3sNknWjvgL4MDBmi/3I24hdn6RAKtmbx75UoIrAakjrA5mCrGgJQGq76
pwfB7xCK58yjKtC6KiR4WHiQrnUhAdXxX0XJRi3qj7ulzhxxFIj0J6r7WmhStKH7
eLYbRygUCbJPzHrFOhkNj17RB3qclxByQf5ChlJAetpkcpHRTvs1yvaJw3bu5zC6
LHwsiN/zLBgVssK72eFX8ySDUsTWVbkISoPyO9m54oBIJcxN/BcnTuomuysKgYli
MiaXRhc9zTCxt6RQJIKe3sYegRq9P+iw/hwDUj1MQe0k6n/gITGxjuwUxHE1jn0+
txDItw3qYnn+qJT5+Go6HhjYaPPm4klIyqhmphzQN9nzPgzEpS4D6CeakkHRjhQ+
tnTBuSAsmM/+E7/yFUSOJ57izAfoK+EO5a7doSnA9lmjoH1UIUm+gW8k5g6JbUyb
KsX2s0K//6IUAtS6oIr8cnuHhRLS394f5IeNtvlGK8kaMlQLHk++84WD729NAx8P
WOFfNT5dQFj2HVEQU5P7LqA3TEhiKyFW+JaODIOetDCM584JCj966iuhIfIWLtNg
ulIfRBLxHZVWPgJUNh0XWh/jMOq8oVGnPgVngEtNcRp4NmMm5i7nEEaQ7a+bZuBE
zUH73jPerGm7AriYYN24nF8lXN0CwOtbQdGbTDXzi/eZWlhZTXLvaUsCXWTHPLgh
kemflrwz2DKiA8eyZ8KD7OLYBa6e/NnBy920aKrbyNaFTAKFfWjcAnxs1vk8pDfj
FS0dtjBNdQ2CLDzDs2/W5YJ/ngrKP0uDpalUPX8F2R1PwAodMpik5rJTzjDuRID9
GO6HpGrQQkxr98Xe9Qo3HDOz2ZLJqRe/AAzmaZe0xV/9UyTmwDEcreSPw1M5/RD+
RStcx9g/RS4ZZb//AcJAQ/gu9C2p5wthv91G+8fzcPat1Shzh1skZXWs6maeaAln
Ihr/mnHVeRRT/2TO5d2WI/DNHypsxe5XHJwVe2nre97tf2u51I3D/OchuBQjYk9k
9AYOsuntWecX1s8suJ7BJ/voRoxxCr3BZbzpcT+60Ct3h+zOd3WQreSKufooDwd/
/ay0g6fKX2plIk7h9KsLW2ImWf2CRJPfekycrC9bGr4EmdcVe8wQdBTs+hSWMLBD
WqWwUVGpDiwsk4Nksvgfu/MYrvCbn/DpB01Rk+koFwl3YvKvDiLx0Gah8WGKOptY
OMMGxv9UzC/KiA4y/rN8sgjgtI/FIh3NBnGGLSl9UwhJLydFOXbcfH2JyGbS4Fab
DVzCuoKn6hWdzENtuIrcEbjFSqOzKaysOwiSEmVk+CgrN50HfhmDXLEFnUN1/CMW
IuC8jnWro94wJ2GWrcxLe48fePwXf2AiI3qPDoo5hvD/oQnvq04ouDUehKPw0HzT
gYFdsRXQOHzONN5O0P2Jd7B0dcbiVw26gDgybA9okd2JbUG01ini9vD7pFcNh4mg
jEKmPJj+TM4Fep4RUee/s8MW9R1tIo0p0vIcQxwPFsYCbU3YEW96ExQZ/+Tk6xm/
YgxUYClJSaXa8jiyEJSGt2KKJpGKWF/nIWkttistcKph/p/E9xI5R8RPu5X8eudE
ksSBTIYdPUwkNnQaSBDnLDFKEjX9RKAmWW540sV6ZniKv/n2yfxkCDrz0izP1jqA
NZQhoK03lr1ZHlrBk1kKimc5Rjjmca8AjvAYGo5CCuaZ2yW0bFvWInYiPeoUXCV5
2M2bmf1EDJFVlr0QJHWaJmr3mPo2fKlvjj9co4rgo86EzbV191d/9lcX73aErIpx
GOGwjep+U4jdCWypfer7whiw9aoJ3c0/6XAidQTXZ5LfJUUtFE3L38EVUZO5LAFP
bDmQabgYHecsZYwL9mIZnb0lMLwg/BmiWhiK8qY42U+usp8j2srT7HRzjbQJ5Dgq
L+laVHqpjikRzt4+qzZxjX/coOB/u+BFaZJfktSsWLSZjygbH26Kwvp3Kq6q4uzH
VsiFO+RAG999tUlNvnqPJzW1+g1bO0MkHjfKAYPGqVmZp2s5BgdbN5/mftlOb54y
1wwECwMvXYzocJkOMDyc+0s3qK6iV15/AiqXlOCW5eHMSYO2xkXBORNcLLet35cw
Q1Nm7pQS4LwL4bhmJlyiGKJAe2VdXApoOHa8vbGnFAYf/MwEIeQVBi/71uDdn5l/
ZSRToAn6lWpxcHJdQ0Sq/LSEuSniRt4AAKU1wTIkCwExlx9a+MjYjkFRMiKEqyWA
nEak8hcHZMmg3RJGR6gKFNTAfae8QiJE4A5Nj2/1wZXB5YK1ZkQEE1xzBU1sphXG
LNLyF9sIu+tEMNY6nhIIPOZSrJxMSbuB8sdan9mWTg2hWHVRxgRyZgN7RtSNHGyZ
pYKbZt6is75oQCAc4NiAs79L7buE+egPqUGjVbpkfC4KyXPqOAd6KnC8eIW0denJ
2BKD/hh+VjxXsBKtJ3R5RQPDGnRAuVi1V+g7qEnd823pDtLTBE9qjpwWXszTt7b0
hjTVTxkwdNQ8S4t4IkRCjtStXP3SirMFhlfNNpH6j59Stfo6Fo82xm79xbSdIqpm
McF3PrFn1ssAuT9MIp8BsSe84+LpjqPp4JI1hhH2i23xCdLV8qI2mwp9DW98DPF2
J2eZp7t4iP/KDjdRxxRhB5hLBYkJ3/SYIuA1JgeHdS0P7cXUK/+npM52MTLke/+J
eSz91inO6wpj0U3838ha9BLeuhR4aHUp3S5T0+MG1IxtyM9aL4dPWZBskWZqPaSa
pMRLHIOix8bXJA82UtsZabiUBcKihfb4u65YNeFOfbXi4IafCulqStQK8BVEL9rD
SjLUHrV8MLKEbgNeid078gUjk59yfKnhJ6TM81Unjw5Y3REARbOZpwyh4y7Qem5Z
wFFuT0jtd8I/Rx3lRl0foDu4MUPrY8jgfQttEo5PLXRsn4JM2nuctSfhNVvDYCRb
JOvEtoXryQ3SeAiPRoV3MJ8JOZ9H7NRkU8JaIzWKTUkmRp205SDEHKm1FlHHRLaR
X0MpwC1ZG5kWpDZ97HvhPb7l0+xkjioEN+BLNJcWZU5RqHketqiIEAPnn/aWdBRm
ZSSm4RV4Ffh4TnZMgFMAVrPeZrfNjOmklq/YsY7KoC0cRY04Nfu/QjOoExUb3Hl0
IzoHG1mNbEiQOS6PmV5SRuYcbSGl34BmXYSnulRQMYcEAheWGfREjhz0tf96j2Ht
3Hr1n7OrXe64RRlIYs2ONd93USccZqmvIVFvMUWlvdUbSNgnTwUFDt8cxkc2cvjY
88bTm61WFnef2NmEDSgSjlkSrGlW3Qj84G3Jvsu7sH5GxpZViQQFAcuE4U31Gamw
ZhUi5x8QBdUI+qs9B7Bu+938+w2N+y3+cVM1eQPhOH2OR0ElbhnoQP21xtSnVN+m
It/x8Da/H2hH0aeyb4DMB9HnSruxiVpD11FDlILvGvU6NlPXM5ExhnWX8n2yhK3/
kjpD3iqv2qxWdq5cNBxodnyRCQhEjFp/QXu5GVp2SY8DX0JJEBDV7QY7fdDfIrHk
T5CaIQLY9yL5R6KVWqoscwvzuMvF/fEnKcTAI8v1ynByypOxEw1LULMDoQePOugM
cI/McqTFCS/q4xmSFdpyv9AiuM3h6kmtoB/Me/Rw/D5YhS8tnby7PNdY7Y2dPhgM
MHvhPJ9mTxkIjnPmQb/w8oGOsVH+TJfA4NKG/WZIxY55aE5Db1HRwiDZz7niwx3+
MheXsemCBTgTERYVEA805CLXpkrFMl8BFZBvw3GH7XGeEXvx5ULa4vyC3Ex+3w1J
2mSGEuSttImPbayXRJ/kl+K2/vkyvInMnud+w69r4Q56yhKexiU9beqxzo4qwf5V
SArdxzwkwDshNixYY1USEizEFYfmQvmtkg1/ct1ifO+AFyqyjEtloESc9dST0YuW
fGFNBh5qiIsFYEfKO4E5iIDjufpqq//ASiqDTGE38fcgZSo9Ye7r72aWTziDvY3J
hfoPZa15Uw+4gLIMKz3VB58I7/lccGy/eewE5xkxd+4keNwuv+kgutbdMbtXVrFg
dRL5e7IcYG4D3CEwPjtnRTq0U+giR3O9gs8gnG2XhNKCh758TbhbyR/2Am4ULeau
uDiE5l0AZSaaXKL6iQA1F40S0kwDwN3LdLHO3Ql6zhXkzjyldxnc6d+vyESFUa6B
hy5U05VefGAvMiv2sVav0Fwv51+fksEz0TlQynP53fvsLr6vjb1tWbR/45qYYtZH
RoPExSLP1nSi7LmHyXN1KtNmz1wzYzrOZ3rdnCE8a2ofrQVWCcM4HzwCtzbb/9yF
tt6AOQ2zPn8iNQ5CEYwMGgxRWMcfEZcj7vEHzeqfQA4mAHELNFJMuSKZ0P5vGycB
/VAvMn/PcU2Sq01qgMmZzZWcta/UIIGHsnxmgW8/4dOiNAb0WkNwHIEs3uwi/dkU
PCXVZ1zmfQ7b92NI+7m0TczJ2X2tw7AqrnvlefYSSLlIyzMW2NtUmA3VSjeqU/gX
CtrwLk2NOLor7Pgnel1AlrNwWbo2uDxAA51E1tTgSBYVvrWmSwMo6/vd/gNdr+aV
bJ91zSkgyBeNM8DN8bgZd+U4nMs97ldKjIhYIQOzxgbZYmO3ym39GZNxvkoSyHdo
sybNyRxl6qbMbHMimq9cCByyuzNnAcvQjwVbgLpxkW3ADKZwwCZ7SjNl9Qqc0Xf/
0cmIvKS6qlszMNcA3bbU6kgyinSZq9khunVSpjj92p0ak8foJbDJRaqGuZpWccuP
uhfZMau0Nc7z4SVaeAjZ0QTcWJIcOrW8SIoLGPw3I51FmDjxXaggI77B0k79LU0X
B0XI1f6Du+AI7bDULLOrqV9ih27fgkAP43tfboT9fkm+ZTNwzUUVDlDecj5H0XVz
MzcDVo/zExjIqkQBJ2X6MEzImo9r7jR0SDPG8A0oI9fk5rutCTIgsEM0QBTJC0nj
/qmaPp0riKqCmzOL3FWZ329uUvdysX+fF9uGBAMK/m4HhDKsuzWo9KRQ/u44IFV7
LSiXWVt/b/TMx5oTWnF7V4HG8wKGZqjszq3xkCvKjkYVh8Z+TsOtGYiG5aHFbYmc
6FB/4ertzq0oWz4cGj2pe42B6MXJod1b+2YvwFjqvkQ8c0Qp3lYpzLdb4mhO1Lq6
HtVLDX+Gi/2U4Dzs1GAGXOn8nIvTa9dquW0b9iianxSE/iZatnenJqZHMbbgIPky
ZI47G7uj7qhdwaeJWMvTso1UUhqZmgJfbV4aTVJGdwXRmjrwyoUMM6U6PZ4d2+Gq
tQkP/Dw0ZliDA10dBcFuiF5TNUjc+zvrIlWZeHg8iwwmOwxLCpq0IqKSnK5V5LVu
GDhvB1Bl7GhmcvEGct0po2oT4UJHdLier0K5rZOuh5nzI0rBYFwmERtmnr0mgAl1
2Pn+Pl+cSSXiMQGYIAfJMZ3Un32GWcZKUJPMolBPY+7OGC0YtW35bnawhfhhiJVW
l6fRZyXMjVp/Lm+I3BVdwpmgdEPvmtIFfs+RXIHnu5eR58+UhG9ENVdtw/tlp2C6
ZcMWEECWlNYOA+4kn9hgy9Foy3p5/CMW/p08fEwDMkJkHS3/imwhhFir17gI4AYH
14spP+h1HWoq+m+GRzXJOhFJe5vCKQPE0WQ4gOAjw196nS+yXryy/UJXczYqZ/1v
KL8Lw5KMISjbWgi41zGokndJ/aA09E6ZIbXmMxg54So0Fce4aKn/ujWe1gXlqOxo
h6/jKMZ3AtLDYeFpr/1iX1jh/OROt8BVTM27ibziFVY7wXQlSBocFhTtMPETYCrf
tuTvXiQMo1a9eTXJj4m5rfdwHNYkvwzmDTqTzkdyo0MmCJa2OMxlC9cS2WKImFfy
Ryj0a535Rf5jTAwooMhlzGUUMlcmllYKx9sxLT4HN3k+ScF+JqX5RgPXQX2O2XVh
tXZhi/jpthbQRtDPfi1/HZhsFgBwZGKspDqs8bgkf3Q3Xm/92PFZDMuELD6Hs9Fp
5eOe5B1y4zbk16gF1HEpJWBXDLit9Jkasg0VaQpD95SF9rjp5ACfGY3HF3y66iHR
HL+o4y9EKNJEkDbCNeareMmsV+SlevIzLy0QxwVZ8Mp2JSR6RsywCUfc+gsogUEe
6fhpjBSWLV2Vr57SbFuvakCAEtgfZH598N+hbvS1Bk7NQdifrwd7x99/mZ1Y7Yb1
C/W6VmRLbtfiE0eVTB/HiVOINBTHcxuB/137IuuBNq7K+zW2h5TQT2h0qg9nV3XH
AQYklDNw+NgJDBaQI1QClWOgeK9eOvw7VeoeGoHZquN/PjZatBlXUzdzKdQaSQmd
MugyT0s377+IYAow6flTrmPhG9s21boLkHao4ci+TM92MChikw3MrdIfw3lC5HBN
MaXYPXy+yhWDc8LaM0/ffPSk3THfTJZOK433zAvJLwH+yRDyWW/LSeIWmgr8Da2Z
JCurctsMYGp/tTbuBrhEmg0Z5J5A/yX9VnkiKgWn4OlpQTAGVRZdHZMZ8kEsjb93
TKNxggMd4Coar7K/9KpvS+c9DkMTsA4AcQeikwIRR9PqPsmKKkibfdmzXg//ODe6
Lv/Y1hH8wg3/YWT4icaFP6nmHVZQJfiO/hQDleKVqee5D1SRtjrmYdmqfv29XiYI
NjB2mWeyMjzJtfjlEWWcsH43qhga1R+eae39zGZdSfy4r+Z0/2J20FFjfiS6sVos
7RUmLvnFMqiUFzWZ7noOYDrJj1KB4g/JC6wNuoqYnMusx1U+JYlyHjWHlpcEXqjH
VCtGiUU+ZLCGdaiX4PERptVtxXlm18Oiq4DlCs1oR1cArboySOoRZVEzKSJnILOY
JvdSwZBy3GxDau5MjVX1g6ccq020RY9Gx5ARLhhUkpb5z4V0Mck7oJ1p01bpZbGz
XNjnqY3q2KoSMyl+eeHq25Fx9II7/v6oGJgKkz09OicCkfGHfy6j57ythMpbruuu
bzKQFCklFfS4fX/pgJvXKJSLKYjFfL6fUUwElQDluRjLIjKkiBmh7oNS3tipFgrc
OWhsvtroJyeZ/zZ8vpcnYwdwxfd7qSOXMIV/rLb48LJcW/Gji/z5S9Y1VvVYRvYF
jeiFjwAMyLjBmYN1e8WNwt6WWsjn1zfvPeiK68b56LzEWsGRVP1RRQmLdwYkuTQQ
yAPmquSMDaUyzParAktR9hbi5K9yp9m/w4shbidfvdWF/cISxCZ4Ye8JYkKa4Nlq
QtGWZ7bRtXtN0WYmZaCnI4YWyMH6fVrjoABVDO73Exz9VPqVlSSfVVTEV5SsqYyF
us4fu7IHzM6IWGcaQqRC6BllEECNqKEl+O8IB9avbfNd0pDP4B/lHTFLVjSSADyz
LcZTeoJDT84nuoaWF1DFaoi1pgFKqjLq5qiIBm8nDVx+x/8V/t39kjfsgkIWn9fm
idD0fpR5kJdoiKkvcODCDFVz7TtAT+ysRBPeUULdQQfsmQxKFJzy1j8ujfihKCA9
uR0MZJfc+0/8RFfJMC4NG7sxYRawPpJrLOOcRvWreKFKclsS65AunH/F465/7Ib/
vC2qJwEUtFmNjN70lwXAt3+wbI8giSaYAPzdHn30njimlCpF/yKW5pBQR83likWy
rD7hyIgmbklGAAI3P6nXn4TMEheDhP15ZyN8mnajlLS2TRN2/sDWwUvkLAJs8iIy
WDZUUcyi3nroCuljco3OgRDYTfHHnNu+E/oSduvcr/XysaYgvxTIuGgwhDVpmGFh
9mkkJ9m1lyvYStnHx/BJ2a0LAjTGMHxLep0jegUxC5waTFlaoMTruNAreGXyaIyR
Zf37JS+Z3XDKPBDSofiHRadmPht/KO99SAJ7Og9x+hNnovGApmgbck3ovbwRJg7w
V3kOvBlRmm1wSqt3VFN60imMUMhpL6OqniOtNnZQsNob2xBanoztVjuN1FW1FGwG
pra3IUxzyCFM5MHUSw8ATw7S/ay0ZG15ncU2PZVcKZNC8epdS3Um/+VPS/sO2Mue
ekIXyOCh2sBN8Xk9Es7OEiwppwt0/j+l6rjSAxlBrYJly7ep/XhuqYzoTmQNpddq
vban4dZL8VutGfu4xiZHh5cJgjuww86pIfvLtB1NlGLBvfjo6jVWsr91F5fcX7Hy
1mgGs3U4/Njmu+w0Ah7ph4bj7AwOtWMCAwkxxAKczAvjlNrkP8Vi/lh0pFi44iR3
VfjX9reUFN624JB9SSAE/VN55okhioZsGNh4HcDv2mJoHxBzW1byJBm7ajBda24K
fD8j1Hwf75IRBkpHtI8PbEvVaCtxPhLRTqdOqK3U4aCzMVOctcR9VwWRGM4bwrvJ
uHS+dNmXERtB+ltqAtph6oaRJZ4EWelftE8ZoprmBcYyRAhNuGgHk3GA4426MsBG
vsj9Lsa19fVKjGaTCBJzdNpc5dTk5/Pqy5j/3UAqznOCM3TueJTsCGVkHurkmFdY
/XUikt0266O58qxpo6aHFRs6kEya1YsIT65kdpNoTOUV5mTcAA0WXVJOk9bz2uqi
6QIOSaki6EBEzMAJq1Een+shlx+ZiYcnHriN00nORHUkobGxzuEEPknpOBRnjOmf
7uCob0GA1nAkgHzwkwU7hiltu4TAhK5MSCUr+hTYfh1ybPOU4MTp5MeEEwG9zHrx
UPIq7w6NjNyz2qGYGWo/kP/8u+LJ8X1p8FFpa4ZtgModQHvV4lEOeJMgn1qnbmkY
21lpwuyMsVPM/bKq/4hodQkev8ZFQUwHp5ISrhm8+YGIsvjwYX1P3FWpTnYwlvyr
eyRzLldt+rWIP50D4G+uhFFr0WRijdC3dQmpv09PxOH6yXLbFPiN4jjHuq1TSiUn
6Nx/LHl1x5yPwyYR60+JURTTMT0RuO+xsRLpqBcL2T1LnjKbCCUXik6ojPhqMBkX
ClfKFb2YDVfxgvju76jdBy3iasaouIzckw8Av1RdtDhg/k/SbySr1LZKdh2gVLB8
NcBclnBcsI628B7S+TRzo+LfLw/7B3G7qqjThN9XSQuFfGVd6uxSHvZqtQLYQ/2n
xRlIMvdfyGdGGhEqcsbOS9jrY9kxKbjdtcDl4wrNvonxIhbsatH8cxBfGNgXOV4+
dstcVXxTvC4X6HOFO9/UQ+dh2eVmXn6YE+/WNSLud7xm8cbGMk0S/SV8iB7VafFo
qb5zcB8jIWJqE8PN5RNgZELXdzVVHyP4FvzpdRygBKyhO5UsoXFIUYieU6LOI/+V
YDQsPNHuw63UI3thZuEDbdHv1UA7KDt6pKQK5eLamWPO6hTYdluD/R31wbRsFdvy
hnqCAdCjYs+d5cmkHPZK1l2eGMYiEHMSM2oyFx3pyvnn203U5AIswyV1pn0ngRIE
T/9zspAIggmDQSOpoUfbpeTpafEGh6RxAAPrr7cCqhprAFkTj3OEsRzzFlud3/J3
oJmXyREmWPNHo8RHELUYaKbqvJuxfg01BfgV8wy8tzxRzLeFxZt1kAdHRj9UvdKl
xHo7e8svLMa2StXElGvREZaezOQgeK1a0KpovNfk9aEVCNnU9Jhp5dKY/dM3Un0e
AYOgt/W+K6hehndepHMV4papRKnBhTUASFyjUM6GqsF6k0bT/f5sIATXBDpzo8tm
csz6MXi4XkEE3VUE8neiT5Lbke8lqwMUoAE/KgQQDcke+NO1LWGUaS8xYJj6+OS7
aaegFVpTVLdzOcH7T5RgJabp4Y6oUniCC6TkXW8iqV6wINdwDzjDZMUWBq7WwJnD
qannbi64I5e6/9giB3OjAcN+lMz0H1TLUZHSjgRWScFNogoGa3FrOjOegp76Ce9j
qgJ4BnF5ofmqWSrnkLY9XKmQUTYUAmCncKZClJ0bcSspjDCkjNqfarEYUxHEDuop
jvV9xvLCEbONJjDi8rhKcd2FiJchzlR4kBUuxZe3Kl7tFp8sq7UWXU0k3tG0Bsh3
38z1kONG3oyixjKIhYg4KWt1mlRNZvsXOHLfzFEcFQmqSO80a/my4oFtz5wpzKb+
aNqe2x8hn63eiOZYiUDdFVj1S+clnLeBdW8fw6XsVgHlgibRE/M2O+fDm4VLsH+h
zajLWIZFeTuaDf2Pl4yydxpgPUDAoyYTe7F6iNitUEBljhWUjvKlwUsaNDE4YGyr
72wgvQiTIm6Bd0EzptJtShfC9ymnO7G5D0f98+0FnHgJVyElfYgaABPDI4nrdlmi
jPMmOt/rGRORe0p0JCEfysn95LL2PFdp0ckLacn+8JF4EnPiibYtkLR7Lrzx8viH
6ZzordtejzdqeF2xFyhO1lkNLo2v8F0NgxRzoWmbFq9M/JsU9QYBttICoRF4IsUE
8A6sybE6nnbIMLnJzhptpiv34lyS+mPFMVL78X6L7d99cDVIwgNZy8fUvAEtCkVR
K5t4LK2VfBQtwTGJ6bfZFq2D7BFkIygDbISBHLft9A8/47yi7lxkPZ4PNY/puig3
00GCoodH0xqO9KMbueW0yGHMp3Rl9jUnUpCTq9FCF0jMpV7MqyiOzjS7X0gysuCw
kyhkhL5vnXH1vbZ/pEz8V8/C3ERuPCyvDQYxHOFuKQKEwfQPlZNgB4C5OzRXLd1J
Bf3i64YFA+qtZaV56uX4QIchMqLVaXndAXVj07vyGpW4FvLSBT7Kdz+m/ZA66egT
l0a1d3gBxti8yq0Q11LUORGyim4QEPcuxXNnKS1TUxCi+5xsGpLoGa3s2+kWnWlu
F11EkqfTrglw3P6rirGnT9bEHGQOFMX780Bddpoznoj0Daagkr7Vmy+XHbLuiErf
ib56dOEuwn9huY8Xy//mgtT8nLc33e1ObB0wqFOwIT4rJ3X1bu6BpjpoVoJEHl1j
oua6wBXRUvc5AYU6dICwMBmaD8bQ81ItayulPl5w2JsL5/9DG/Uc+3OUJ2CxqmDA
eqTrMx8QDbsw3ZlEfVAlK96gBOyo+RiNxvacgV5kAGzG/2DOSN4FkbM4OYZxDnN7
OHgInZDKVPWTJC7GOxOBqcg+GRxY2kGCfyLx3svJcuyjB1xSpEiCmFDu362p9K5F
LQBDwctlWeqSEeV7NgPWT3tmVhR8CwMtjnG3+rGY1aFA6/FpR7CRv6mH9z9oULKc
qpowFpc2O1St3x7JNUpbHjukObPOAmgXrVXt+fZzrPPdR4FCJcuBrPZKMBvw725n
IaBPz5mUA2kmR9tgnaHhwDDaIkXkN+KW6ULdPo7iTXujcnrgUxk9ZvGLtGAZSPGu
LSuTFfbxqNJTUrieKOzv7RsIXvdjxBdpyUW6MJzG5RAdZvOva7J7JU3ZGuLCo/7n
UoVDvvNWRaAnmEpRPBfMJbpeRBTJD+AFfkbcwhoybfUAjROwkbTHnR6UlP08zoor
oVR+ZleSCd20xeloBEv86s0FpER9hBov08jq59otcfGma9gSR1/jUWIqfnUP4lbv
Sx26HktqZHbICrLWbqq2ypnBn3AHrWJAvTNoF+weSg8wgMupScGXVjqNCb3Ozgr0
XoSWuq1cuvj3OTHgD1hiRpvbN/TtSDaQW92GEkfx2FWioDUPIEVCNQHPObr0KPCM
QjKM6vtMv5HJOloj9imTjTBDR1ng7maaivy3hBGk7bX2gxrjTBJbOyMOWW32jj8d
ylLNXLKIr2DSldSDRqoj6f1/vvc/dIYJZhelq5Jfgvam2UCCHT/QtwHX8WAljVQs
o5MJiLCJyskKoPXZYl8Oo+MTaoTuKUWgDRTpqUC1UmSlsfg4hM8p20SC4LBzx4Sz
KB7bEIRDw8dZeswILnJW4PcZYTmepL6dLp6k6Rw77MOaTG4JHk+96oxR1OC3U3ng
Vu9KEHp3mnHNMzAmVbTNl4ymNOZnbuCGXGRKna4cKDKgBhS2y9+4sWIwXlPzIs6w
G2PXxEXPXoWvctZPjdX5I/GzaHt7rkQurNxBWoqI/f1xcOTbjPhvCdsuZL1AezFR
bQdGpi44ejd1A4Ub2nDljywLfdza07QvzbzUvGyt8soOQ/VGcgPDYpdrr5POcXyq
2Q5aJZDuJkTIcqYU//6uXw/txuIntup7ZzYnqK9tC06F5/PBc/2+82FGg/fD80eL
yTrBuU6cokTTjawirWplzK3lNALGi0oJR6c45iL0IYlmQIaWM5aIG+fIQU6uUYnq
GJwHMGb7eohusdDuhPL9ERaIpw6t7S470lDieBXfmeLu/ac+bNB4ekJVtTm1bdfh
eOQt0BXfhgsl4fY/64s6BFazcXPf0jmK0ulgk2PrROMc4470fNdWYgq+3G+vJ7wP
Yekj6qkZn1BmzoLWi/l9sCJGGu4D6D4blbyqik51HIXbEyPQvYBRCuWOjVYYtMnj
Qs8Pr9ineV8mkvqmvThQeFAo5PdEjdqK9BJFYXBZJvmLw/JzDt2sydblb18f5dsp
dX7f+ZXD9YMt9aVYCRWoHAYNXlHUsx40LX2LxE97xh6D8LE4H5f+2x8T5LdWXuSd
8dqJZbN5ePPjBI2iDs8EbNNVWjObqz0xrEYRE0A7DrzFTY28TsUu0+9gNRC5rpck
0evolaaWdqRPTp+G6rx39FO1KhEupwtQxKgt1cJ5YcjS84Ys+7q/YZyW9mlubMZf
hSp96RYtbC5nluxlOZzK+Q5S6ca+57u0GyBfZjxHFIgE6TFL+SoZbC119y2Bptcs
Lu/ERfdX7EyFFr2/U8OQv3zf/MYfKOE22kEb2lcTvUpU+cA/vadtf5TsNk1wrN24
lqY2xjyIQMOwklAcNKQtu2eUo0uyR1vX/UBi7GcKrjEuA5bxoNg5aRDkl2EkXmIF
4gcFlUQJHOaNwal8NzKThhC38vljlQ5kGG+Zu2mwkT1ZKPNnI4SgvlSyNNK205Mh
EVkz3hWAwBCNGoIvipe/z3dr4mj+lzrSj9DXtq2Nu8cuJOd3hu9xYvN+TVZPxZTG
6fm8+FlZaxKJIEVjrnLrkynqRdV4BByC23Tg0N33/6Uj6Qj6iqV6tn8hKDK6PKf3
DbQpwToHm9Tx04lid4DiHIDYlGH4Lgj452iQ0SSOJNUCxHdmwoNyJUskCs+wNxQK
z3XpSLrmyKJUelQUJrBM9ufJx0TsDdLnS4HZfl/zG/mC4efkRRPo+/l7o8h+MXe1
EpL88NwqvLdOkqjRvDwsR+Sn7MWnGfN47qu+TawksWpdS+sPziPgjOgxjbvH679z
E0W3JOVWOMitQ0NHYE52MrXauHiPeLTPUjseWo+8QrnCbx2TtEToJUIMBepwkGxj
jVTnryT88YzbU/1m6Ja4h74y3/Mw7QOiD9ybYOHHofvKHRbxck8mcWhQUG0OFa1i
sx3GLLIutHOCceWqKf8cTz+G/aW4Y7XIZBNoQMju0dncAPvET4S1dp5fcXxHVbZs
Ik7YINwR9cGh0u+w0y8nhPx79R2Yc3XuNom19pFcb94w8sW7GgBBSz/Tr45+hy1w
S+TC2nhGY71l3YWmLJDD2VZ1geBG4Htr6p7MG7RBgeC2eSI6K/TG7ta2W2TE83/6
IcfSoBiIpTCsl2c6al45zNCrbsujo9HY5ehCyrKWIuhrnzqkWK1E6a8yh4xFsrjW
yrxjg14sIAi7zabPbHfLaqRkvRBMBpjsUo0VSJqQA+H9Jh0g1i+2v4wazoznzzDx
MCuUOfKhHBhKiTsz1kbaJtAO94oLlyixArHojGRy2eyFPkEsiXMcBXKuA9xzyoS5
Ko+cz3usxD+KHw1+0v2OTJkBZuorKpL/Xu0oJ8O9+okR2VULmq+SknKLgrg4SoFw
uiJBuBASVAVewEgcYwetN+bR1gboycRyrVnnDzFBIHFedY25ZsHFBdWwt3uawGd9
SRQjTOFwiNbbfI0no8S86SypXcriOVJ1EE9V5qr5mLoTjMIVbmFhN3TqdKNqR3Q0
UZjp+quRN++V+1t2ia0Dbp2igQdvszoiJWt1EiM3xct8Ut2yNxUAwJfxo3mLvuej
jfUqV3In6ESccY/m2f4Rr4Puqo7ruRqNKm3bus06uc5yFGguVdmdZpR1HxY8S+/s
QyAfywg+9Jtil3qvxEbNdPY+F4YsJNGjJJWcr92SQ9cAcVWBC7hpIENrtplauczE
BypL45hQq5L850CUciCJfXWbxnKaWrkAHE3zjqGEW/SYIvh2Zzj9ausEvg1UsAtv
cA4oZw6mRt2yh5PSHZyAizLKRy71BY3NS2G6QARKtpTJYchXiS0PFxGpr/iDnmW+
Yx0XkYi+SNCrCGt2v6EqfE+hKqiw3QtsrOwchlIHxrvGMxgPbHXiX0VVeYopxPof
uZdx4omPRYBSUFX3Fs27utmNPghGHMqoXFCgUu/FwlFMg3GooG2xUBNYKJWjp7N1
HuSrD3bnz46xuTWpBJgEyAo0JWRwQOw6fnYUrnSBhVruNAspL34Mh8R1p5d8a045
GiLj3wJxSWVHi0L9GipFRdnvycBLgKi0jEJAmeQM986AewKv11q0iAk/2l4St0l2
IYJtVwXtipa2zMIIp+K9boKkY1BOtIqmB66TmDhh+Afj2ELqs0TJY2wEkSV3aD2Q
y/FqykX2ZmTjUD/ICW3P73HGWkDub4mFNcvhsEKqCsZHkKQ1fX8MyTg7WO3PpOFo
q+wdie+sg2SfAp1jwLyB+VqCI2AKS/NOFbNcOJjtVXoKaD5zrdq9tMmEZrIYyZR8
bQpV7GTFnrb9Tsuuvg4fntuDkUf4n0bExqWDccFAg58F+hfTky44/4YCpmcdabLD
qZCojyC+dxNQNe0KUun8Ys3zlhd0T1mssEtP3dV6zQk+Ig3A2XrztuAMZL+8CPYO
b39SiohCNLOeghcYCC/yNOQo6QpFAtFojI+lcxnaa1km1ZzpwrhK9u8NIqO4zaKo
UomeUeVujfIT+0t9zZBfacVRRtZklfwEWjmi6yXrO7iBDXZT2D/W1pk5B1gUx273
nbLrFQs7GqwaCYfSn7sBCLhK9LB+FUl0B2lDcS4ULCkdMOukaEnqVymtyfgAawY/
hmTMgdEyPL1xNFmcGgmeojebnFKCDjMydeQiZ9kfXOgx074kS4Mbjx+rKOB5pzZT
VsH7aXrMo1GGQBTfatWkXkdu7tJykdmRAfz3/5/CeAYQD6D8q+btoXnTPinSKItn
rNoCp2Oq3WOkeEGHIJOepAdmB3Qk4JG36U050LormIUtgQo61GUI8gF7x1ry2kM7
OhbWAq0vtjzxcOe2qVxnDlgVPwmmwKWxDRXK/6zX22JAXlWRE1SAEj15oSkE/9hB
on+5ndbs77m0ORszOTSILMN9zK+wWcaZ1A9ctfQQvZpXJE4/HC92oHGadfRgR3Wd
xfBG9ZFCeBujNej0Ng4iwWaRWH3EriJOWQQHIAkOvPz9LEfeVBqqMAo7LxWfZibR
7x0WEsYJZHoqNpDuGKFFYiHrfEwn5mVfzJIJjW8DOgqAT70zcfOAhOAGY4E862VP
UqCMPrbQIwrO3RGEqreyg7zF/gTN13REKACqs+y/skj+BIZDYcDVsj20NuP1UXzW
nzLRd2MvgI7IOF9gmJ6RdE+jtJix8AsH9YW7tMFNBAB8sLeFZAyWDp8TW/0gI3DN
ogAKiBwXaGNKSDGQKau8SMz1Yg/2nfK9lzWNRz/F5uCHOa+9cRA2MDGzt9QMKpym
nyk9mtMzZupbYrctqMCXlXUb+NVSYeuqkgMG4/55UnCNZt2C7acJDWl4ZTrca/Hj
nCbsim8MWPgaTfiSWMGFsz0IBXliONer1jI6v3YqynIXdGY8yoCqiddw3zE9WKsW
O6LSIpgbMmjv551OWaBQSKuRny1B2XAnI/PLGDG4ohnuA/LkRBVVc2fvGmPrY6Xv
r4YaRP9Z7tTuXh6PN+1ytf0d2hdOD3+SnRS8ycdimcCkuRCYQOTvkoXUN8STCQyw
SfBNVbWviu8LV6qUxHq7bitpfcyV0Km8hca+7z+gnwJd6/Z4aDJdF1Ecsc4NqA5X
xQCD0NJijBkgoGF6X59X+FbWMLTwScC833iQpZBk/FcjyMEPboG92b8CtO5McPD1
UnortdgA975J/avwbHbUA+OGqj8+2uRJh8sSQtFVjZB8yaONCMOcYrNBjWHPIwo5
S8gOE2vt4k6t+mMflMm3M+4GvPrTbwW8oQyHF3fKmScyrue0J/8EHhjPrCrPZYfI
4Zlq4JSNZkSTirV1KDSP5CQjJrQ14YAR8nOTeBfzu9t7ofrCSbJzy9xS6IcKh8er
ubfp4dCwv++POn4k5Lk2B632l5I4iZh7xnLHXMN3pDLyp+LDOf35+RVgSw/mMkz/
XM/CsKd6/YQPaGxBDvI7wK8gePwpXm++6OdAlky5rilb+dO8/TVbdhI82S6Ol6KT
oIdM+EPk7kE4WcUclGoOrT5aodNXvHZBiziErU3rqYQymASaMKPqeahlfhvvNPQf
gYeYtbCZCgPbjWqFzTzU2wRtfdMcr9w4D1yAOl+aE+yti2XfTttF/DS4lhcd+Ayn
4vKxgwRDu//U+dtOST/5grVU7hWL+/PvBa/pb3cV/tdjK7ZW+dgxvjRcomL8REiq
Qu6AszOtOOpN7v6PBFJDnEWeNxCbMnaV8Gy0kEx58jj3c4kEynax2N6a7dRDyy/X
4B+B0vQSRM7O3UA45d2I+nYXC2yFELB6Y3b/DjZ9U3Y414ByUGT+W9UeQc4ZZOHl
S9wr0CbZzdivnoq1lIbuAtg0HFN6pqe72CW0hdYC0MOV7W4k0h2t7y7P50XUu416
E2GvmiFyItVAD12wwUzpd42rGv8tTZhza0BtQ4H1uQQSYOTXouAH/0rnf5hLpka0
DK6h9ZcjzcWdznJesWuoE5gY9XRI89Ew/tJYBH1+O0NGAbojYrX50psrO3lww+Qk
Z02xsYKNF+z4JionockZ0jfA/OxDJb8KqwOU2IuEg36g0/LbT+XCGwa7z2c6qM9J
UAzMB2AhAj8U75AAivvCu+RLVzakoI1wzk+BwlvL16pBXj8FK/2keBncL9kTlNG7
aeF9UMwUE3UQ4nO1VswBA8Faa1xOHD1uTVh4kIs9+yHRk7bPDO9HUmf+Z5EU7huK
tkeDhoeICKIrXJiQxxKkK8apFMnGM9stsWqmSRjm2cwquCazGMX82P1Oa1RUlRco
+tXifYl7tmPXP7J8MagvI6qC/ihHbgOQMTZtvTgH2qwIvymOLNU5wPsCFyrVQ025
QXIti9ou/QPpLwRkDJ1VQRdsG0R9ziwbtqHgpbZTC6waATxX4OBMbljlYS5Md3Yx
PCEZPlCJxSX0fa+A05byzIaNXXrp2d/kp0ej2pg+5PT5fk8ZNRtxAuyMncpa4TpM
6X551R9WUpK5DwTDLymJV10OEW6drVyc6/IxDLpy029pJ6XDImubnqZ9P3VuJxhU
bf49PZch39RfCeATjhr5ghwnkxgepUyn2u5rvDRXIA1/uUt86P+KjGfNPKaTnJrV
HNi1srY41zFqSUaZrdFiGVfEhESvQ6NTtSW0dFnWm1z/3Gjx3ak/XyEh2frt6TmM
hFLn/EGwr2JdawOcwc4edA3G6dTFqs/Jjdaa5n0QritpTFSBd30dUhPci6lyWz4E
nGva6EHKWfSq29TnRuCGGBl+msfiRyEjNCE4a1Fc0/5gVC31KcTJX7RLGnWu6tzf
CdJV/GEWC75MC5QtRR4B392RDXd+XfbjElvZXA4G821ntqrWFxdo/LQLc8WXKeLB
IBilYqySBm3tiJWwxKj8ZtNGP1GCpCOeyKZ0E9ragDRG9wTlbyDE/i19ocUYjjMW
V1CZGOArpWIZgUzlvD7KKo5SWRIsQtjOiSpV8E+1Ae5EE+a3qWm5NoeaC3FeaoCV
FNbizQrGZjz+hBs9l5VwEO3pujJOB0H5RSgUuDXn1T+PnyejISrmcjdx3gUw64Ss
EwtVhjFL8bmCkh48vI6Ei9nepJbycvMQ66Fp7hLALMc52sd24ks77+M0UJSDBHon
brFPND51f1tDfI7snvjoPEpNJ4x60LeEflJlz/qS03OyK5tVaSHFz9QcjUo0H4Kf
/FH7i6nh55uu582o2mebw27oRQG5o/QfncwBKRR5XvFeFwKs1odhLlc2TR1IZXPF
No16lP4pV1XJ81bG/Hfsu8SeDOfzSO3C1bKSrT3QHJkPLXlg3Wb2ignD3XAktXBQ
7qG3OGJN8Wa1FjyFooU3BAwyvtkwQOPt+dRPLS3Q11Odu+85rzE4FG6+5nBi5bp9
rjXyGWIWPwCRhb9ZrdZLF4bb3mLBqV1qCJxmvKMtE9QfEeFbCJ+Y2NX8a7BU40nH
6sLDEF7PZ63qtd63ghY1PTnLlFq/gWLcNsKPQ6fdj8NE+FOFyvz+bhxJjpWt19xY
8C1TuKmFACxwWzyhxXhkn3BAc1VDI8PuTBR4tzNPipRyLnpvXbXdHZKObgu5Dnwz
U/xSeBHB2XcSK1Q0IJJvfw8jOwS/qVXAXiKMTnaMto2PnSuu6pbNxaWZKt1aowxc
nAMK2uNVZTjPB9TfolgGZSNGJB8/phwKsAtHxcs1RF92yv0glYfxfndaKF8sPFep
zenmsKRzj7ffg3klRXI2xF9iYJD96OueQESsREkyY1XnJ4zOFc5ybhjxSHtq8JUj
urXOw9xET4iiVrWimsNiGx/hNADxRZlt+Y6S3hDkiYYY9zQkCaWHfW5APFo97qrF
HV/qVSkA6zPAdaOsTLHpFM9HXx/prla/I4+JrP1rz0T+Mk+PsMglAReae8Oiyv4D
wOGM9uIzVwDJC85tvd5wTt5ePIkA0U6qhnJmL1/el2kqQeKPJgCKoHW84BIk2xbD
ZViSKY+rVNk88xOLb6bwU14642/HZy7mIgGVtM/etXim/qyYylE9Thx///q/GbVx
zlCdBP6iEQPQBE/5S6nSjpf78EAXV/etnrjsQYX1ToYeTNaEDlXefrknH7VWW3i6
UMS0d3WSQ0jcqiSSBt414CCJ5b5J+xl+IZCTFugznFkTr9JDUBcM9TIQltkyXsC9
7MbBIPpxp8DBqjZem2vR53W1HhQZP1qhFSJVgzghtBjw275/F7vX9O9D9xIagEKk
0TGVDVS+T8eeh4bKFx4rAyCVE9joElkI8cJSXoLFu5ojU+hR7n8I4rx3H82h7NB0
NTuzR7rI1+mBLqicFFmZxgFtB35ua6+BWiC/C5hVcIGNn6JSnl6bGufir94miCO8
3nyoihnPTEidPdK5J0Hb7jrELdbMQmoP9FkpDint872KXOziClne7at4ORLASGMW
VqdTkNZvHRJBjhFbkAIX6LfyOULyJ1bQoV9wIiW474JtpBhI0Ro9ZPhiD0GQC9AL
LhrpS94WvdvaBShn7ZF5IPDey7RiynVG+AYV2q7sN8MrThJkZIsxFs84bU45/guf
cfv/NqfhKg3I17FPOCsZ5Uwbxsc8cCvD1i6cmxKU8jd75YWXvtcpy2Wuf1tuPYf7
T3qaHZO+MNAJFZSqkuO5HUX56EmhwWgltjzC/in2G5SjUDn+PP4ATCZ4mmdfnTDP
JZJr6zuviTQgdF8iETw7MyPzoxbN+1iAjKhSYtgs5V7HpmCH6OYf+KcoYal4VXFz
u4U2WuHzGPImc8KTrEztct31YjeBLEREXtEhtyrZggg5qtc5oqjjkMPJLWnx5X9O
/Qwho1Oh+QvS7m41fKnvNmtNojowAsMbiUkvkle3G08OsuQfz6MDZ8MOmhL13w4H
3jdy5bqYLTi6UNBhfkJ8cv8uggH6LS7ZkW1ZMA0S+lruXVs3fiK64gXy9VlKVyO0
TzVOe5XJvcfv0vYBfWAgiLTp2lRVvqj78V0wT6bzxTi2BK9b1bazNupyy0NnqR5h
iHqJtPIZeusAxQfsbo8lnviG7XWc85HbM2e82Lt/WXoF2ZRguCuTR1/gZETXfBo/
GEIoZQw57gvcFO71qZZTF99jXZJMvAVnzfO8AEW5uh8Eo87WtNzTXMEJhe5NgJNN
ovwdPAcwpCPmkxoGrT24ko1v1FwjAUhBsePTfPYUh8KpqDxf0IMsi/X1861OgsKo
CHsECu04YtXfLYLa8hZQvWteFNTf11bVwPkIsmZRjNM6aIimuH0c3SjOGInjs4Vt
pQiOqTrfnaRG42vjqUVu+w1A8SHEn8nyMHAHX4kQLLQDZysppe0nNQuYschXoa8m
6FAH2Pnz3vfbXczFkjEkNLsoOtNB0OCyrvoh9AqTQ4X3wQjg4WgwNR/jTWSbEtOA
7PoDO2WyDeeUHJW+npxGHNv5jZ/HVaU28BPYs7+t1y4s9uppc5vPiAwoiUt3uKK4
OhZuez4TNI1CTP/qmpM+HoiRRzd8ZMJDnuWe8JfY2fya5AVsbLCuX9ufDg/NAZcS
6niNoINafiAW/rZ1iBjmWPgpaitf7GGNo8EDJas7dnwJz3OXNur6f4Xybc3++Z8w
d6V9owrMmISqp4xVseCSLIG+F2Ec0s6rhptYCM8JD6oBCAtvikGx/PYpGoAvxV0e
zdJE6E5NdWz7Xa4wigXb92f8Od7XXooKSzi66CYy1GJUHTDDMcadcN0liyF61ie+
0x3WBy8pD7r8fj4IdVoOtIQ9HOWL5tLtSrXzDPGZf38kEtIz2yzgXFCaiFGvOLAj
DMWS5VZyBgyqqiWKqdQp6nmJ4j4UO4YrZ7afvh81pCqjTg3CTciml0Uhll0Lq9Zl
HV5Lz4Vf5/vIRIBTp4DbyYQYQRbnQuwM2C6lCBsSl32x/w/1sqlz+pA7i2DIoC5c
cA9Yryk4/7dkvhAum/MzdNfGUTyDIHEmd/iFntf/Qls6vMlz/st9FqolZgdrwXv4
imf+VaCGBYhEJb0G2ePRic/ZwuTDA9s/qYN6/DfQrJ5YC1g8aJELo6VTmI5ujI5v
TzsrD6yQvh7XogOZnpDMCcUmJSPv35qqQLpk1w3AWEs1K4rX2pWbtg9mirkK/fSr
XsNquzgwV23jYYC8IGHOOrVKRGt9eQJKKT9TFFJiyP9eXeWlYZkwhg0aS4GSsiTd
b0fg2VlTvQhXlAbQ0cDhtG/j6uEJkoIqS0QpUSyNTzOIS620p1LF5vOJev0vy93y
uBqIeDUKMxzEHXdlpcjLYEzaPgGsUIc9ZvTL68f+h2qyIStXLLN0WdIijd9YY+kV
bwOpkD657X749VxyBC2lXpRR68wp/J8UlOjpSPZxiWU3MRp+Gi76TT+xktqDd+gy
PLvJRvdLq1ijK3Tua8On5dL6HvGcUie/dczCbU06WHzQKiynX/1HLLMQ/LytqF9y
00ArtIDJdzA2LWQl4wEgZ+Ym+wKvp998j6FXrUBKuhkeTn23yxzTRL1SQQ81dTgP
VuDXxZCPhKBMG5wGhSbXe7RLXPXbXvGdzcNtOp9N6C2O7cZpnkVhBkko9fVKGpmr
zwwwJdAu2QV9BqzS9Bbb6rhY7s0ptd9PA/LzmhWoUEpByQ3AEQtwZ00ltmVNq7wc
aNmmQXtQj4SkXxICnq9Y6oNZlTpVoAyvIWKZG/fViAqqF4D7VRdAY4VHKsl4lFrA
gt/yMAQr8jEbXKZajLOw/+Z+nBcEkLY0vintfSG0JRyC4RgXZwqvyfQx+vhTCcvb
tE/YQbUJjh3BbDAi8z0eFUEQZ6V2jkFY6LM/LqOKfFIZj2O91TtURDSRxqha+8ji
dzDz3K7/QuqWg6jip/K3h4WvqyYG6WLbyF2EQi5U7tDy+mfee/cgSIl+UiFbfG+l
0IOzSDHqOSGR9qbPPRaFDgBYkYwbTVu2AGmXMM8GhOqKs+uTK/XV1EJQj7l/lGLJ
+bLKiMNfCYtThdCRs9xJihZGu288Yn+694+kfcwQeTtCxV3/aRtWFStO4RBq7Jrk
N5kBould+zUw9zO/pK7AoTCYKl4ZkaGdktDKvWX3roqnpEeiDUmXuQJE0K7Ozfu7
f0GzrdtRneyzZZ5AyC3xd5FbJCcO1e+CFhAlRzY5F5LS67ZhtS/9NfokaNXyZDWY
1oCPtYHcToVrtDwB98kwumcLQaHdxi7lj+lnZAQT2CCBwiH5+L6J7WpxhnTOqK9y
Fkc/88NY27PXka+5ShC9qsQlvxtR+B4ZQVC4P75Ztph8gqOin9nJnBjdWNOM51Dy
5PGi6KjrUInIBBHD5yDBG5de44c2sVMDYtegWW/kJZpa/k5T8PNgoY1UnDNfY8Nn
1VUI1bqfH4J8ameC/aUFoYps1Jaupq/uVorUr597FARDts6kw15BVnUpGj286D2k
EfXo6gXX9rzvPqlbLyXuuPp+Lyhl7ro2iK9GTSXpIVJv9NYacmcTI+po5e6NXc9h
xYMh3Dme58p4Y9KzzSSpdTqi7WE5edyLXTis/dB5O7thls1+Z+5gyuFMLXdxfV1T
fNuqEGhVaxKvljFuffLq5TE9UbO2CqtrwQv4vIa6aocUatomIBEwAlsD2mB+x9vq
12KVKlxuivCn60fgD6gQE+8zFZP0n3vqIkGLn/6kU2/8vD3m+iz3QCHEo9R/HMfi
mBB3ftwhLYZ23ieorjDQ/El1XAOnre05kezW33YC6w0sNgPBFyMBTRDFqWpocJXP
D17gNb19g/FFVJQKOJ6K0lCwSBYUrAAjfepzyjKXRqX3G47WgwzTD8InSnsqRemE
KGdjDsI+NOKhSGiCc80LIOBwetZXYIGJ0BnuOcNzXZvJ15+0v4XMknwex3lk1eIz
Xgbvp8CRyrLeJMCx9kekMB4KIm16fdh6TXqckK+zh1z3iQrCihymwsnn6hBahjsX
4kJ4erCfk3YX0o4FKHnUpA7gdCz1YJh61KCPtCDyr4wBMzL3PUW47qxjJpRYh4yu
pTq9mNVK8T078rFvnjuVQZtbI96uZrIBhSvGxnv9gDoiOxNmNYDKWz6mPGk4HGOm
WX/Oq3soSll9srL0gxkoBhEbWujPjtbvGGResUNOcZBX9atcvmFRnqZgcH+nygnn
j4LDKf5qHG2B+seq42LdgDjBi4YPwNgjz94rtmdtls6NgZGykJMCqwscdyuIi/kh
GC7iKM1Fj7O+4j+VskB8Ik5XUvluUz1skJONFBWi4WXGkz7Z3spabUOPvR3cXEWN
YjB/SE3sZb0aVuqwrTlF/meRl8eRpEWFftx0AF8AnRXWI+fziDh6FeJ4clzKZu2j
cXazYkY4qhrcos7i5iMAHsP17FtDnrrzHXto2rIeJ8lgRpMYzo5Y6XGJU655yw3D
EuxpKYP/VDGoOA16UJQT7aqijHwXyEtRBD/GG2RStDm20kTrMKma2B4SujMezSQ7
JFkAZue5303h3fUghXlWDFnpIjUyIvPRXC3NZ6/LOqD14u7SNrAlqiix9Oo5Von4
Y0sAR6ptVnKD9CSZD3TrvscfAwdCglB8BbyJH9OH3OJQDaV4MsqQkS3SmuxeNDBn
uPecX/xvINbr7VmrCbW19mGy6RjZMzfmWeBKkyunckfTiCtwqb7wcf5Rr6IgKmeI
6yl8xW+6Vlr5mzp04ObkitfvEGIpzeCY35XOg6QHboWIedxODU8W1vEZKOw2Vep6
FPPw9Zndp7/O17F1f/wSrNC+6ScLqUqhRKLTCnCfklS1XiTJDzVbAIfd3VoK1yPZ
GQRqS3gmir+w9ak6OK+JFBo1Kay8X6SmklxYdlcYgNaRGXhqJFKbJpMiCZZQi0CC
NTZRi2wVhU/rlY1CfSRVQVZxOpxieS9L0EvqNMFRTzwBhGzjxB0jxUBqudtCUsle
jCPke/bdfwwg5xJxl65vXWEHDl0XQB3IBA72oNjUsDe589gB8boR6Vi8LlDV55Wf
DEFly5Pr5RyIenaYAdRj1FLjMJ75cBFYR0m4rovvqLEnbAT4JT5bGbwFTX7QSWaw
sN+B94nVyNeyDQxAluESsoBmaC5akmcWv6sFE8zAIwTatWinY6+jPqx3W/ALGIo2
Ej9Kl7yiVfga2XojPEMjZIV1oqwHY54kjLAbUvQmZysOjXpJRpTEHPJUbGXhH+ty
Bs4yUioNP2hrnfdIaohAmFBiDj1+oAGNYa8eQrPAmB4ABTxxgxue75M9mVIwDnP2
YUUcEV9ZtFuKZ5+atTTtmXsJ/C8YxOV4wPCm7WEX4fvJPeP7aLiuvxNbvkcFUSY/
Q/grEwLI6YZOPYlS9nzbbP3wGfvmuQsyBn+adiAqh/MI7/O+qShvXRel2lbu46Tz
xvYlhoB1zvs082wiic2T/6YKlsxuykXjL4dq8dqEhOnS5GDbO/66CsCRliycqneK
+x+vwFCHDuz0OfYERC+bnGHlYsgju7cZKlQjFG5ayIMYQ0O1Mq6CqIQF9n79fd7T
Y0ROdQFxBIuwl8+WCgDH0Ua+A9tCJJ2xbYNc+dcKZLD2pdzscFMzirhtUspBkSiR
m4cR1c/PpvXC85iYmH7baUukPpn8eho3qdAXl2XdQQSWy3brLzG7c5bdPxxHZBcX
ParkoCfnwUVWhmbQS97Wh0ucCXncv0NG2IbxdlW0RQPj7Gw9pSA1kzfFGEO4Qr6M
zndt5asOfxMFkHTJS/ZM/TGkFg22E22z7MhT8ByubFM6oeZlZXdlM7oGgQNsqObO
DQyqm7m5wFyOWVQg4cK5pnkFlLZjiTn+vNBIvfNyHxyZCKzPEdUDLR3AXVSsypsI
Nh2bnU3GrZGK4b/UKruiwwoNVbrrQabHZtSs4jLlUZuwNab0v9kwja9c8UOD7xY6
RKJpPktuX7DRbXD0zPitRAr6lwrvYVquprZztgGObglNOiDHAVW7iFdvfMZ46Enb
oYaKIbjsCCgJ6wMu2+t7w6YLNd5FzWHWvj60ACeSkkM28pggUjwjQd+lSPrCRk8W
kIBkLppugQD8VBqOT1E0Ou1tHnjehm1E/RkTXSmemk+2uIU4ZNAeolAElV5abty2
DG5PdHJmFScC/1aIY+84YtFS4cOLBh9gZ/K+XzUXkkd5DTSgxkBxRrEJT+vZc7oo
FyfGIBcq3rXAuxJp76iavgzAFX8bAf3S2LDra3Wb3slpRGhvA7lsaMveZCXf69T7
MWv+d6fvE6uxt65w9nwgdYZHCjrVR6Po919p1TRqxrY5Q3P8mDx4tmy2jm6+St3C
P2CFaA90Vly0YGjr5I3xD7m1IVWY34F/v90EcCNsFRAJJ0b302wzBFAAy+JIgC/m
dXdPbGSbNW/9KHofpzFTS7j+Sdr/I33OLoZEHSTO3DtkNfyn9Jnz3wnMhLBLbJPJ
wmlNDsSJMtZM1zQM+RtDLk2WXxcRqut1S1Z681AaENWF1upiRgDLf+tOBBlEMJgd
zrSozq/YGas0TZ9Xrx32dYLJENaP9Z5kUAXvL+zA9QWhtEW4wdXAGNGxlAtjo6vg
dRKzOFlK4D8KNBDSaOGszWqMEn0BoFq1TvmzAJbc6r3luRKFsMC3/8KpS7jjP/Ry
GJxzgFXJWzRAjgWPMU/pVRxH7OMGEb4QcufRGgI/32hiX5+MGhBLGxyNBMFDtwox
a+BijZU174FiEdBMDmXPbx30YiPgLLFHcoXXLvwNTPvBzwcPoFr8i1ZlDdtuTo9l
Bt+UKlxxB0vyxwuQ4g85K/dt4tLR0/s32Uwa3/9Owy4UA6/uu5oByKDhNEubevC6
cmDPQ1h3E6I+mhH2pvOOnDOGptnPFtJcJTWVE2AQdENXCkVvTOMQVI9NujWWnkNC
vzLHFhSt6WtgvHNVr4VD0OMVQYDlOEC1SoyDlarBRfCMZGMCV3H+3zlwUZQ7kuwG
piiTafNwt174mI6HyGCNE0i2MRv7Bu/Ypwte3f2J/xSxytg/MzXSYhQJL/KnTsWI
f0oILiv0btwVPwsdypdK1VrvO+3iwEkodSF9U6m1lLqOHsNQdotCkAiNTTkYHbbl
CokCDtBRR/5StClNR/Jt+ksAcNOcB1AtRqWrEphGUH4KBzMjvG7bNOM0M2RouJvc
FTopQavIuC35CBJA27t2ot52opJu1Ui+d7aZcxWOlziAh+PzdmCAhG8qKPmyD8GN
5fYTC6rDemR6zX34OOF8RQqu+cN8OgX5S29zhUIKDjjlUb1CMvU+eDjHG5I8xZQV
BwgE773RX6TYO/bjaqRjExh0oDHkIvFq6KYAfEXHSvEd4D8+/GzkUPK7zhQmQLmm
vynFaorTYgVOmmSpf7phMqElrh66kIfiZzSjU45o41dHO/l+xJzmLvKgnL1butnn
uJbWw8kWeshVghMAMPYDXgDO2kFxQJ6cFfIHXiii2dCEiWwRW4CcbVVoZPdduaWM
7rspd2d/OKI9bMy8L9ROdzsrjtESJ7X7IPqAAMKWFBjTqLrd6ONhWTdD9hyQNoRL
Rm30sp56Ll5RsHD/YQQ9UX7ueL4Tv0dIBUn6DF4GePgcNtofh0KBHJAJP+WYJSKf
SClQxDx0Pf/bRnF5a3C4uLmKYvR8qFs8uEcuwSgL/jXd5MS2PrHHx9ZEfmbLSxQz
h7wW4zeFqO6CVdEMgqpyuu/8UURk1KgjKGlfhAmZkSrcjRXeSiRm8VhIIoEiYV4N
UaGBA/MgVmn7a17FWm34bxj9o/9eI9k4TZrzqd5SCMxsfpPvs07/ToSQt8fwIFYh
GUrNtHsWREbP1REThJn+encprremWllOcV5aWb6x5UZ4nN5m115eyGzkzLnnO1y8
WMxUoBHfus91qGZ96gcVCiH5rIDtl9TKte0IDUHa21xZfsjsfFb+qwZZ2JHLlkS1
NNl/zwpmdgh+9WYFc3Vkx6KIAQWayUvZWTDs+UW/+8zIGE1Ep2MFMI0IjTia8lqy
sWlECd9Mq12x6PE/1asY9DlfW8J/fIRWhXqFN6yYBdx95IivBttfEkH2KZR2Pmg1
GgpuK0EBmmJeWUSLDnT/MLGyM69FNqeCx16oO0wXbd/AerISDlipeFetw2ix3Kvl
lXY3gvRvK43rWVFilegIbYHIrxqznTvyvM8gRs1Odyme8FZaJ5nWGwJPrEE4iTrp
bdP/xx3ex4Mo5rsCwuKTzQJNpULoFJrWOeIJ1tdo+vdOYylBRY2ScjN503dWD4A5
NCMqdr8UD6YFZCJP9jPrktUDNt+rTJGyzdJAzJvykJGNgbAjMXsyT1ITKr3MurDh
9RO8ehWZxXxQk26B3PuQmc2v5umvSaC+rNch8j4A10IxvsQ1gdqd/Qv3DMbxVY3c
ksP+MMyU61CP43Qhh631xvpyEjH12Bg3JdUT6UTHBlTsbaURkbdrcflKsO70PZmf
+SZ87eKTylATd3OMAkU2gchxdoIVcp7Mkq05Qz7wwtQr3vIvraUvdijPhXkL57Ds
UxEg0OqaxzZZWZFPemDU+dV8XDZwx9CWq4K+apsBlk8mfzXyvcd9l9wZartEUug/
EYr3CiOhFhrg1SeNw8+rnvPfOrpjXrTEYZoqbRywGMWTMi2C8rat6LVu+uDTw6UN
cvhZCLjlJwM57WmSfDkl9PExNsFoufEx3lcvOR9mctyJ/PT0/aaacBkAbkZmqb5w
TBgegZWJE2hSaqYA6dWywA/ud3KWXiTCfrV8ijgwUQ5f8fCoXfh8/Z+xAFU1QfgE
Ycr7KCFSKwoMYlGcZ4bLuTdAKOanuQsjctidWWUxqOqHdJEQiBpDRHbDGAPlN3V8
RP07YYqJ5q06tAVb65PjRG6wlRY4p/fLpDkPdkiuEnfFjKg+YEihAjrA7wZRQ16u
w3KYZ667bXHdf6BH2HnZ+eQT19GUDIm5omnsToE4foFJ8he/cnCXuns9SyMF5j2k
kZj4nuloVa9MOrdWm+Uv6xC6WFGzBKVJ5lVMosJxKJTZlCcG/jv9m8pOOEj7uRxY
+32OXImDTocy2t70TI+/CxIfKjVrzgJNYg6G38sAQh0rDAQsBr+Qy+WOnqphDyyX
JWVve64GvoNDS657ZgKdPQv6c5r74PIC8N+XY0K9l1zZxL90EfyPiqgOtdOGYRHT
N7GGU73D3ygVDGRaiFbfnXkUgTrXlwWhdIAaIuuicqa56URpvryosa7iQPU3xkw6
VVthpOZ+uIZqtSiETWGhvfv0U/lec1A7WF846+G/YxCKijxlZ00xuQGpji27ik2Y
+iwsLzRGxBBHbXKlFcOMd/BPrma+cswbU3PO+MokJUMmrFLpz98IShNMYBVLC26s
z9Mi//LYmYh/dhrr7g1K3yxV+ATgMHWVhenRx6AYWr757sukxxx6/F0LgkKQemgX
wHFRaTzhJLJUr9ULgyTy45UlDtKBSDSDUPZbHqDWjhFv+uwGqyt3FmoZ9l3hpDRJ
DBL4lDsZIhgmdHmsuYyaKY7TBfs6XYdkkKTzIc6bwlASYud2ZPM2XziFNugXdKih
3BYRtwm0njSMq1UDBBaFb3/hBvu/uJChXRjh7cjuA0m3BrYaM8h6zZx8Lc4rYTFI
Kb9j9tl7CuHfOBSYcSmqjsvIZ7qTnw6WLzAJpULNfwrDE8F6ltMKKXBLMlRvyAu5
Bqo+dRGE8ZqOynuw8s0q5040RCusNKrLsHtq1iylQcp61eo1xgYeaIUsRORrYiKq
k0yGBUNygmGSKNoVTL45geDR5UYfvkDwwFQ/sLJeCUAGQa4Y/GJJ1hjug9+TZPWj
oicb3W4o6K3duK31aJ7TSX9HKtWVKO3TdSvCqZJCf8w3VaQcEXY48TzjEbpcEPK+
Er8On+d0hQvYzMi3XulHkzehciydFW0IlZJKJ90DJpvXGLfCT6Y/wEEbgpfaPi2Z
oOepSmNeE9m3hYOkcrZynWzBjw46KNYDPsTvbhflvMlrZoD6RKlk/yZmM5Q2bMxN
5lyZKxhnPNXv9Iy72u5vbq3wXHLHrLnq65vDZoxgI59cOqgASxXbgLLfcsbKaQMM
Wzhpas0jZ8KRh1VZGLGh//5uBCRvaPlzMbCpj43VrQkfX7/I2wYfrIumcUCX2EjS
+nUoTCm+gUnWL4bKa38AFMpHSwHZT9EptI7efwC5LGR4RG7Ijk4WiA5vkO12Yo+q
XydbAtarcbM3Tc/3t9Ue+R9b3MxfFY8NS6Qihn9mBx31jRweTh9KECnU8Axn01Hd
B97X0dkcffHc6oA3iTp9f2u16u+WCJWcR0K12U48mu3picMu74RHs4HQp/F4QRlg
8P82NYI+Yi8/TzdQRgUEVImVbo/6mHZq6Xad+sqgnIY2Q/lHjfSYWP0IzF70aIcU
zhMXPTF7f1//1hNBZqBFIybMdJGQt6rA0lMnu+TiioZVjzUKIPAGv7MEkP9Tbz2j
2t6qi3X1yoE9D54LFvP727Vufn3LnY/qVZpRNBQeyceTKndqj9Yz6GemxI5CLpw2
0rSf8ZnYLQt9yzDEpy/hZVIVTD7th1xgPn69h5+p+tOsWPXtfW+MVYW4XZt99a3N
d0FF3m6oLrgDBc83YoeocrCXzvrYln9zcnE74z3kjF08w3b1LjBdnFhntBN/vszB
z40abBLzJY9z5oVPaosyGEiTsIpXN/ljBrQT5got7GD10Na49Mn1o3dVspgjHlnD
vl74GFnBXxvqLgNzp4SaqIF/twciwgiiKcOuXBE0WVllm55Jj0h5stIP97sRKR6M
ZAxX/aSVJ+iGxYDV2Gt5tuURPwJHQe21j7wvzKe7Q0hJsp/YLP8pTBjMi4/9VLSB
I5N3YEH2gjIdJVD7zrplg6FqRpc9f7N2RvIWlu/DeQlyA6a6/yXmA4FRWbcE37G+
9wHlccEjdXpPKyxAQ0DHyqjEr9Jdda3YdvifXuH0dRqfg32fHzG1tCIeJzzBqD1E
7mKhbtZTiMYsY4IHf4AOJ4vxN+EvgHzJzHP+CJpvXkbSjo382/TsyC8v2R85BhU/
Qdd3VN28QEBe+/jYg8HowcnPXhMpEi98lnfYs4Dg8wwEf6jmvavmE6BKMcC6DQ5J
SMIfNDbiBGZ0k2Z/AsYxVC8BjLIYsRM+QeX/azwuX8p7hQfjgg8qDnPPYOtGC0Yv
xwyrkyS/2Iargq9w3o4aidMRvWKZNTOYWR1MxMQI3+InLcJrFjHr9HSVtgGKWBDY
auk+POIuT7+1LWbdpCAyD21S4cfkllLjFfeClX6G+r38v1UVm3cNgu7c26yncWei
UJOzDrOMXN7r/slkaKei5JBZMNBlsoJPGtFICUtOh9o9ITZvLMI1jmOG6Aan4knG
mYdQmsA9Fy4y5mD06C8tjZcbI2hBkxxzSs6KMIOrHVhN1mJb5gsSQVV+gpKHbMQ9
wH0zh2KJk/lnUQ/z0e/auaJrqQ57Y0pw/v3zrFDXM9oEAxvExyV24SnH4va84Fu/
I+9kolViAN6zWTPFbIKdbq3K5y4EjF20avIXzNCRnSafGEtiuMqdEYrRTUWRoDlt
gtFQ14Jv8/c9rVISsIoHUIoYA+wjC6yqJsS4BKOY+8qwQRY5/kTVzzGsIrTqeoDI
eQugpXvWn3oM52BW24V998Hy+q6vOfoe2bqvtsMebE7kdKZPC6FI7i16jA1SMAoz
9OvbaNXK1kotaPJcGFDofL8vCS8wiCdVNy3SCl04MyJuOakMMtOqBNFbeyIdAba4
ES2/a9f8IJnZJ8S57BUdf811wWZu6Z9LdedQxf3K0n9rAz9nHMem55VeH4N8CpTC
/NCHh82E/h27Mz7ep2xXyrURfg+QeRilSpAkGkTpMETlipOZX3PR46iMgGIAxWwY
uwiFlhcwfoMPymW1b2NYuroRTrAoeNXkWXCrmH65CBdPgpTrQDBXmDVLjNXo+aik
BNdqi716DRqd6B+0OHe/thd4aq+ph1CfJC03toc5uegwpO2RiIo8ekuRJTILBbpz
jqSap4cPt1svIl/BbBQ7ZfipoA/GNnsRSPuYIW8GoOx8mwR7rtYkScQERVeXKcEq
ssFUVU2D8Pw07oFSqAjHH7SEyYaHR/XrSgljYv/Puw0HJ/UEPFS/DIeetykKTgRh
JceccMRAcOz7h3Ve+Nzpcj8+jaJ6oUJBcpbvORIaVBeR1MLudkkZE81s/PEMb9pE
YODRNAe27cpNncAZdmfUtGs3hcORcS6AOL4OOjU84JF5KJH7lHixSn+/nXJbtoNJ
U0gxkkFOt5g9+7mzCw/PzH+pIiCLgZ8afWjutW1vMUqtOas3vDkH2VR9HNwM6gWv
2svJ5rbgDLrK52XI65kTl2d3G/BIsG73S+HGqlIK/PH4bREQ85PvDobjRqBjxCot
KveKlcHY0LPXY+Rqfo9cTU6fyWRVaMlBVtem6qaYdTnBwtKva63NsAdbQrYKVu7y
Pqw+VoY+8eWO15Bxumqg8h7sxUo+1ozKMuae4DCKM8Qj0hM4k+qG7R747itPSv3E
bjqVJj7XtZ95NlFtGoKpQ3kOOAdTEfGJIZldcw2GFZRaVpN1XSqa96rOt0SiXu6p
cywja1K1LeBZULEebHNZuT3jXnY2fHmCVKfv5FJro6xjxBCsHxHmh22jgPEsVny1
VBGbg6QofBfjOInqRx9ucDukUi0Wl0irgepoA2G/2w50WOPSReULBlKt6yGF0ft+
uqC07vKS0shPiq0Ql3WgmuvPFXY90UzTNdiywS7dZhMYiFdPB9a2AR14VtEPUuVm
KdczHVfo+QAHCzivZHiSrmgWO0gciegHP8VqE2UN+Qt/Rbsd0Po5K8AJNd9ZVC+7
gJSGQ1saIn3LKG803GcDcCu6E3iaPQLh79hrGoIBd2Je/amzAvPK3PR7En+0ofp9
TAbJGH2rAJnJuQwW3IySMaEzBy7uZ1t9BuQ7bpSEKFcH25cfZ+agAijXVpYuX9KD
LK3wkORIeIjWkk9GlSa0DRNrD4jvvmH995LbfMByRT0UZWoFN6/fFt4ENe5VA0sd
pJWURdfaehF7yexrCvBLSVHpJaYeLBtNiPxARopOvo+/yzh/ktitd7OHlGelFOH4
EiaN53OTEXvd8Q4J/QWDC9CvRaRy4hhPrDdlZUH77445YNppdDi95t4ocJFtjONi
PV5Y5iTA2Vu6EzwYAqJWJUtCCgwSEOHqaSqLLvp7WdkmixwqyralwzHgGZ/hlG80
+Lh1npfFPZOPHLXaPi4ZLyU9WmmD5WOsy4bVPJkJP/ArhNdDpdeqTsOqishJx0s8
Jp2LHhjaHXZL01DduewaJG6S8+JvI1WRmqGiCRh9GwbIMH0JCqUNYIyz5J2doSjD
VnNhgKE6uRMalELAvhiDADBdF3syVhaYn2RTndpzYmFpbPGMBq6sEk17vmj3BaGq
0vA7iYV3I807rrNz1DOz16Lf9H8Tjq1011BOKPR8g+R+0eJ+bJ1LyNBLiDu6v4Ob
nSRY/BsmMkRmLSeG46VYrKnCPwC6CwCujZW6nbA76GN+tX1bsfScCkp8OE1E8q1g
zfJQJSG6lwj0OSkdXGco5kxk74Zn3ehg8s6K01EHBefBdGmGU117d2f4d+IrtbYb
yCy4g6DRKU4yALYggqwFidBwqDgpnz/KxBtfF/vK5Phtt0FjiPxeO+AWZw505Jd8
NXcOAeWZ83RUXKsz6BO59cQyIE5cf8NKR/hNuX6oluNk4yALcB8wTORHhnitn+hB
jJthS9zoMMgODNTzCvrp7KiCjS6GLdCYHIoPHwQz/sX+M4hhR+4ft1rgtb33IpXI
q9lMJ575Gp9UuclXrpNS0GloHa0LXnf7BENDEdhnel9gr9lSiXZhif9kiAZkfmgb
L/hAnRIASM+qmPkUAt2mitGo6fbwfJDp+cdtic89A0Vo6N4TOQsot/g8rEmLIQcr
zaAZK7dsseDuFTdFDb6q5VyX8J8Yk7BDQlDfXIOlmVu7P0xF090toOOSJGiWR0AT
KdtHfPfD1srpYjoG6YGEDPVEUXgH4OaXWykXd2MPqCD9ThrNl6jR7udJTgkiFToK
i5FVXvD4u0o5uOLg+ujjgpEBI3bXi00rC6u3Vt2yCvbhhvWjgU47AKiryVwGBaZ/
+ITtzotyi/GMusIsWgD197BjbZn6GSx8ShDYZMe2YjnOw2WucqKNxC7wG+A5ALMS
/TY8EPwd54B79kOpQAsjg5XBFPkbbJbQJQhRRpqLdbpWJCwR9Cn57BGwbCUoTbg6
p0rK2KF73Jn5nFaOGwCwP2VJ0vcM1OFWExJNASeS88FC64K+m6xDhrWH8EQnuHya
WZQwuHeVpYRdmJI8uL4HChQ4CEsinMP9Qz/O/oPq+JIjNZ+DEUGC9LEVo0Aw0CGX
OPj+nU7/tNNCerYKZqzjpSVbwbPzDlbxDhMPdNqJm0ur5YlMeaAIve4RFINc06un
O+P2cBfmhPzDm9wrRHGVHrgZyBrMApTDGnF2LmVRaJPsiYI/7rVqkCoSAv4uXrpb
K5evnatkyQMJSF68c74oVKLoKtl/rpdLU25LNmfBunKXsCq5h0v4FWUzNkkfDQtv
RuPxDHprSuL9OQ88QLgfEp7/RFDMwztZV/IA6Vu3p6AoNgBzyUWRSETHKtP5FoRb
RpKvhX8IE1Iq9UZaIKUlNv3g/WfVZYGqsAAbAQ6dp/Eb/pTfmSRisb2lAQwaiJPc
r0oY0txhtkopAAhlA6QeKEtAaCwG3d8HZRb3xnHY4VoR6A1TjevNumddjotY7VsB
gwBfXg9LhNZmAnPwZ7E/32QO3OiiTiE25vcA8FwWYflsmthEZZiLvu3URIdgshig
00WElwH8Sm4I8Ug1N81gQ01By63YYsidQsM0RMtRZhpJxshn7UYQuUs+IJj1G5oJ
pprqia1g6w/x9NjZpleLM4y7yZFQVtn5QjM1heFXQqmC8aoT75D/t+ve18nXW+G4
0p6pEJoRQ4QcRnMI+XWmjSZW4ox+d925mlbgVUDmPEmD7ROCwfOatbN9496CS7ZG
aOAofJdU+iQZxrUiSO3ojmeZs3bX/km8eyPggImC9cxZ8it3MvA04PqKxP0qD+Mr
1Y/G695MgfmdUqZ3zfsjykflt8u8+RgcD6pcjVPXzJxkEhbk5atA2U17RoH3umxO
0k0FEIlrtSRfaCn6vE2n+3yCtNhC/I5EWOoDX7rDbA/26x43533eZXme/tLoTErQ
OKHcqhR9aboCKXTK9MKh1sLdJwmeDRYT77BgSpOWJkq4qBYkypIYucLOY0GrLcLt
cVV447JZDlFAeH8M+4i77uwy9OlbZDwiClzee4lBYO4J+U7tC2Ul9j0W3BDlneCQ
E45M9AiWoYUDExnLmBnMwDc/Z5cR2hwQPG3Jnf1TMMhso2qutZ8Zs6BGYYM1UIg8
S46oMAfWuWeXpZpY8BIq5GzX31PID0FOZHG3omiVBGf0Pv7Koi4IroGkfSSEtOW0
NetECQxd4XPKWd7JQvgvCTjvrf++v6wCiU00+PcCgZ010ifMdcleT4ny7NkLP23k
0JL48hCdpAElNyEpcmRpDzkp7PWXjNHY0VEfaibHQYj45/5tTgiyCjf59pIcstcX
E6Mu0PQLDLqiGQGYofkr6pGQlSZPMhClhTYlefS0SHQl3OJeNagZQLkLKnasIXbh
E3XZs/3qH1WI5b4ueR/uzwwPlR41DnK+LE5xTkj9v852goNImd4VuqbLSsKWCy7h
J//386+pe4z/9tmMU7HhXQydMk3OlYRyWQ5yLaMdJeSGFqnwTrmTxAplLzzf8z0w
I9tKWtzubQ3tFZzTo3z3Q0EESFbcGF7i5b3P13RU42I9z/+08KK/fdVtUe65IoG3
HSnWHzThF7MhrRlcR+lf4VxtiNfZOSCOvB0+9rd0JKSOjW0G36cvyO2Su2jnuZsM
7z++RGRXQxMAM0xUZ0uBUlJHurPKn6WBqaHcVUtNfyh1Cqzk1J7vhKIqbaBFYQ2d
iTy0Z8h/H3y90DyvuL2Nyolo1wRAs7VFwYFzP16u+oYw4Kja88+zqBrjXN2k0/T9
++8g4Gt93tRn91UM7oC2gtjfnAQjQL1hatRdILBC/jlfkqF3HUKLWKrWwFJcsLh8
maP+YX8uhENcwpK5tj94zQbA3bPfl7vCqOPTeSmOA1QtkTDB/89RcU3C4KuJkMOR
rc1xhvVirNbpV+A3MNXpqVmG04onCK75dWVOMZAjcKfSB1dXjpW8E1YLbwwyHTe8
7rKHGQfp1Uo3KheA6iFDxDrRqo9SrMP7VD+x4j3QeTxbvw4LlUmO0Z6NXXydLAep
dXFYIVbUod67+bTP4aZdBnPgphbjSydsdyajC278bxfIJKJFxf8AKezFE7VVCGNK
xNrM6ctYmCLgepgD22M26uvNL9Awm6q90W+gpxxHTtdmOPand+Bos0tG6xbgFECO
SJFGYEVSufSzkgiocHq/1YU9xBZysLPH4Xi1KheEIzKihkrFLIx0b39C5QW1xm6Z
t0rphBwT8qL3QcNB+i3im7tG55fdbLgUOjpyj7qs2Z7u5zJ/Wai9Q4VNOuQ6BcN/
WbiwOKpsxuaIjabos/YaG1D0F4feVikRbrkRPamb/XeBZkRV5p5Ua6etKjOrqwlz
I42kEbtK4n14ZAZmLQRjrWkdHW1G85nF7AnyDlekt7JONfTrSLF+mezjEWEsOmUa
qtoA5GWO1XY27JaiPsQXWzLh1F5xK3UcwlpFDOnkBl+RHKtSsxbDHkP/3nNjNdkA
qIjvwJ4fdpWLYKGZjSaPNgbJ3pS2fJ6Ec/ZFzh76RXcg9nlF9sU9hUOyeGhrQ23P
CZtc2ILYxwTAWKqFVcPpMbK6KLDvPBk3rXBJF5SbY6cSK4Q6kKzHcQRmoDZ/ToUs
UyIVdlYpw+NBQnz06nbiGVlxEJthpGWBfR076faJUpDZvxBfAUhD/29m6e8MbCti
IfAzCWF1vhhcZiG9+t8Rk0P0hTf5N/a7vmH70ergpvqiQD8pSTL4949wqU5cbbC/
1IJjsxDIc7HRfpTN8mZCc96IJWsmSL4GYg/VSdVKbRoa64vyj7wB5fL20qWxVXGl
vkVlrsqnjIQZCUY3MjJ/xmXXRBS+sFKBvJlCZD9JbbhzUH0MUjBGjV4tC7ToxDHO
Dh8p2Yi1EVJDQkqTq8OfX2npHdeLOudAoFe+GupHZ/kX/rmGeZhEr6mk1RHosev9
eCJXqr0/AGzhgROZD6M1Yv0/BvHhMEe5BHuxcGEOsJCfudFFFHeYmyYbeM0hkPJc
G7E8Hn0gPD11W7Aa/a5Ah3568WT9bn6CWUll6wIDG5V/RvPFfxDqr6FrooX+4l3z
up5+bGgimIe4JyAcRy9ppjmcpvBTtN6VPgd7HlDqY5vWTycQ3bb7NWCTeJKxcsdb
CqcBnWxDN1pzIgcb9D+SE/kiaJA4kdl912UWWieqZZIrFOtOaYaV6BZDj1nTgwGW
XOju1FxSz9vGQn6nirgSEQj8voNC4ufMTMpLuRVVVO2Y87tTuIPae3GyFuUjJSJF
sMkgsILCe4i93mIyVCToI90reiEoWuFg/LXxs7qHv0ARtrY3c0tGYP5UrIGAxQ7h
qIgbCYCMatOAM27E6t7IYdnYtWeK6Lwu7j8A44VMfE4FBRZq3JO69FsPrmg8gECQ
ljInp9YIS0YWmZa93xG61FG7WE5Cb5tWnQqUdH6ml4+DOKCK43HRs3hsLKeVRDRo
8dG34eTHlASPHnCg/EO0OIVis53+94JB+dFLfO3eoh/R2CvuGbO4JigirAs9AIw2
a0+SWYEJbxbZQeQYGVxZEckGzEAd/xaX1gmVIOSLntzb/zm3IBfHZgIUlMku/41w
yEBFbdtvd2DiGNZjIaecM490QKgSTcT1Gh6Hyq9QnXD74PW5PFpmbGuTggYIja75
uHFed1wSR+lqUmjrzw/9/pp2p6Uh32l983IdYD5DaVlhDdIgKC6zNRU/GugB5rRE
iryPXY3QFdcA5r5osu/lKt7TCxNwmuSp0ha5WkGc+kF8F5SfATvpt4s4lZsnYWzV
0Re6s0ASjg2fev8YlZ+93SGE0G0sba/xAATZyNM3PW7ZCEQtPzDbMBzuWniju0Kz
FypZEbYWYOD3gKEvrWewfU9gUJapTqE20RxNdoB3fs+7QA48qzq/FntcczPDYEmq
oRzMjp5Pu6V6NTEkQ028kgmhnOioPalC856cr6Ub9xjP23B28XpuWaWv44n0VI7+
Q6Ph/dRNQP+h5HpEUnj6G331WmwwNKqqUFF63DS646e6/zFrnG/chVEcRyGc82eX
QWjHNEl77nRcKfgD/CWLuq5WgtmuHDPcefOHFw/Pv7ZITGpVWzyqFCVHXIz5XYRQ
RvLCuu+skhax02zvtoFClpKYzRajlZzS6jfHORbi0iY44Ca7Rc6/3RmI8GrRTRFk
2Aiv55GhHFtkqrP0HaldfT+xsi28H9KHwk5Ic8zRKCSF7O92rjGkxH2E4TnDAvYL
MOHGIplOEa9XLeSDJP5ZqCJYAHcRIWwAkxwAHZCdvijJpYscRTBCNM02DeEwt4u3
zDDyT8GSsCONOQGL+n678zMxo9BiwkfV/XvXv9SlLjo+ve2M+Pzj9/UBRtDCRFzJ
pYwqFwiFQrra9k7CmtCWnIrwPP2t5qadVRIt+w1TTGnUsIDvDZM6O03n0nOzqeKk
YbJ8I+3C72qC6Wih5ZOe7XvOabdTZH2EhR2QvPExqvC40woocoYk9nFQg5P4jduM
/apEKOs8YXxta5Eb1DnNc7RTxA+ucp4Dm23Oui0Yzz6QZSBWXGuv5U/o4MJK8aN2
QXUXoDHVpaYuNgpysC1raqEfwQWcADuHWqQUXQSu5w/y1sYBiFa+JKvew6qYJ5op
JqpP1Js6Gs4ZNasdQWTigbyM9AymrtXkbigwM/vp7sChQed/M81BAkIHEbvB+Ev/
Y3eeqRIrs+Fxd1VuO4duGRV7nUg9ybXg57gC9QJ9jLkmayDRcR2J9bgWFSdp3Wfi
5gTWU41SkylPrOPQoinBYHU/Okd40hoWy3M44LmY6XjDBNvi2PcB8r/YbJJPnNpL
lLs66IhHlmlGxGkspzJnd1eYTKZHVo2XV9XOg3PRcUanri48k/PHmS4ogLZVHtPk
upEUJ3OldZOkE8PRVb1Wdn6ukU/SF0k//AmTLX3iB7GEHGj5C4sebeOWXqwrzVxb
Wp+Y7+cqYuJZay69Nz1hHpR09Uu5K1lbDBPjj5ziYZ1g04B7qT/DYDsHVfGVeS3y
tFOjuWuYMpbjGXpXUgB9K0xkOsPqWI9jZqf/XtK/4BRnr88XFiWw1VA2e8NfRDC7
CpipxytRzNdXZj5s5pjHw3rYEZzc9Fg8j3jKlBf6EZD2PlXmtIQlkQjXNXALqcyl
b1mC9nB3rnYoCfVZwdSfAmX7tp63AodoObszOwe5xueno81gcb4cxQj4uDiJo/q8
QDE0HUy8rONNwow/Cnq0+k1Q2C4Um1GnTO2inzT5rHWHoE1qt1kKiIpo9FKknxAu
CF1uLL9L+ImY4/36o52hg8P9OVDx06gLtrFHuijHBJxVlq3in8J6XGnqMrSZcJxZ
EgAk99UfQCOV9sVBKF9xpZRLxWkzWm1llUVyB2xFgqTLuC1fQck2BgXlFA1Iyv3/
JVveWfxjk3+7+Ee/JeYeAuI1g++iO9WqHKdxvScE/xrig+9Lg5NmsIXOq1XAEe0G
+jww7hm70GoWiCbINaEBIdT4CvhmyoSF0C78QoxA2iWgsT7jX2A0dx0MdEIQ3Wwp
6/mOqhcK6C3d6G4F2BHQqVAfvTVol4FhGrM+y+bIOFJuPiIh9dUzrWZSkVDOInmj
wGK9k4MqZSQ8dt/0vHtt+tgmcUth74BCiB1CVvVaA2xCAVStcVN8vVnUAjZY0oXV
zA+sZFktPk2CH34spr+taPRggbl855pGkCrgZ3halViLGzfW8xMwRXx7vHF10l/A
jd6nJ9cGFF3bGPYbkytGVDCrEtN0G16z77BWLG/eHuFPBLEDozE6Dyhlk6k9dqna
d0lbJ/JHXNOm00qLdMQQ/W11cMOhmWKk0EFm6sJKrK33MIIswoMsv7E82QIOMYW3
WkpvubZUqG3D2RHRNGaEn58ajthsCuj8/baBWwBVfKWeMmLeJ8vhTlJLer9pXeJo
2+fFCuOwOrQPBZ5JxZyYqAsjjgnyCOVwJTwV8KL9dJ/VXcK23abe5QS6r+h/q5Z+
AdrQN0GOKwPZqoN/RhYk13AFrux7JadnKvbmHa3bxqjcjbXnhw5nDzhCSzX33fKo
om1HKBIMODjQIY8UAM1UbCf3UW1fo7EPkEMZ6VOB9p2v/Hk8fryLJ5HM7fYV/r/5
YQ0L61ynb1TS8yW8GHd9G6+nT1GTP87BYTyo53028h/qlnl88pzW2M1FKchk4zQ+
B+JR+u6IAPmFWH51QVsOGO2HBdM7E5Ihm5AVxylkquCcWXpJNXOlBYbVDe5riGKX
0t6ZDPiVqD92clCPAUlPPkgedIcuse0DysMyZLtooCfRY9QqNxxMRTte267W8Vyg
Q/a1AdjHyAsHFlTmD7Ic1gWALQCsugxKII55SH5PQ+CEv/suiS0luR1fRXOsjl7o
CZNqGtmuQDyBpXHAiPMEGlOygqMsDLDez2YDrXVcsywLOWww+5IIoY/QWPvofeCA
8SwywGd4JlR7JluKS2aiZPu9B52PGXGYGtwz64ssKumgp8lVr4NQMnbGIzlKOgPI
P6BFwbc8aBp+abZQnjOuAz6CQFMIpHLfFjhofXWwHeEOsgxAg9JtmFKeUhDAGenG
ZFFS4oe/z3YU7dWtcwZkACnn5ITxDp5UI3keMYxTJs6fOd6DkQS8/LQj6ZebM6os
OQYLLzlCZa+3AVkWfB3G/WMmWk5KXKknky84UzhVHM1GYePHJRopJKwmAFE+5S+O
6kKpXWm9+dzFtKA6cUAsqYTRsZdmMkiVJlzSsYlfdwUtTJaGT4t3YtoUN/a+X/qk
k8rUrsXXcBHEowrP/gKKwIKhoHWVgagSEZnnRdsYaPA1jwS5PYIFPzPD3KgI4ZkB
yfWR5GL0bv6XtJuTb2MYDyw3OkletC/xsc2udiNd/gbz3DXZELr2H4x3RJZODy9/
spUG7wVyKI/HphFQMN03hkZJ2jJ82eh6QNopLyOZPOLwu9cyBB5K40cGGl27LDsN
+wtt7pmdNE7mrKDy+in8+ihbNor8QWuRSLGYhIhRf76gP0i8xj/M9lqEDBaXdgF1
LXZEnx0vRdMPnQ/JQPAyGTSf9vddntIOefUdALn/Pb0lMtpE6tMQMJFp2ecbDVA1
DmBfwmu9CtmtuhKsWtklu4Ct4QaoLyTv28lpUS7jSwT79y7wZvZIzYog9cyPl+Ac
QUN3GXFU1DIQMmpUaLDdLnKtgEGE6UXCX82mXGoQFsfI3CbCzusVOyaa/0bzs6YM
l6L9ZuQ+mheKT61XYJVtf3UMa04HQIIaZQ+7BQXhKlqBk/U8awVkFopAZon3zrwe
KY4gDML/WJxWqhzM1xQqiwbvHHjzwDcf9Qt/P3XMkiAniZw0gleoMHCESVVRWPP4
y2Mqz2/2BKPhJorf4QFYzxzk5WkuNoyEjalO9odwI8b9ttCeUghsUP4HliKkKDpw
1TEhpoKkVnFxXIsc6EsrzZHx7QvsQxnqwAB6+vedbknE545AnHcMUAmXCsDuG4Lp
joO1340jM9jOBJzDFTXm2TQIaWG2NnXiAw7z01+MEdt3jR+r2b+KHBv0zcaumXfQ
yHmNzaOEkVDx3eH9iPRZzJRuRHPfoEWWP3NgVy/u81LrtjlMkbq4AYfMUFr7+9zq
TNE98RtrPFuqh/2vwIXpAaB3YxTaiELgc9hmLP4i+H8lus2anlnWETtnC7BJz0cI
SyehnlQHkxMniWwwxlMye0cISJOaERAw3CKHTTp67mf1V8Z8bCNE/u3t4m0xVb/7
wOw8isblpT8kI9aWysOU8W2tIjRHPxq4If+Uoq5rUokH1SuLcyKdp6mGorve1Ikv
QmTzJNSl91q1pAynJwedMIaBtLPrdvPWozrulPRd3v4VRlXv3giKIeuXp/OFVInn
m9358mg76MVLR4HQZJSN9/0Iyo6swFmUbXymgQDyAykfl5MwVOw6AqAZxe7m4kCV
fekxzEuHMO62eB04l3kj6BYrvyeBDpEZfJh2Uelj68wjKhMlBDVuhVFX98QTXV5G
KAX66lVocLfYHND6JhUknLa1cYPuhSdF3bMNyCaowvZ+1/RbIMaVj6Wxf07CRECs
jKsV8sirKeacCIfFX+y+ZKxWcmrSaTCg55OVNaS6NPhp4LIDum9+Lj/2rJoSF6Gu
dky24Ijr6ZPSpT5WCx9akGLib1NStcyweyCCSNmVL9XYu60rJlRKfJ6wCeSORc0m
9LTrJFuoCiTsHaK4q045VtG8hdkgRRzTmK8/QhA4IuOVXVIMlZJAfKkZ/YEZjItG
tORduQ0ZfQgG6j+7dWFiD1VvfLq7AueCQWYAKjYNmpoIo5hQPtWZy8QPedWuXMqk
dvIjB3THW3yOpb4w8C9Uzv7b4rROm1ZOX0qAOEdwd0wPDeQe8YzXs2mp8jAkSZ8N
u1TqLiXUiS2k7PbkVKytGxq98+u5CyAY0v6x9l+mtO6KweuYzE4QU+Vpfk9SVMmD
cUS5sxXThTejOLtqP9mdzQvPUL9OLlOkjRWf0RJrui62IsZ9EhD8n0TyZn1wU/V6
mGJS03n8I5OwZMzmzibCC2DDwXQOxdtZFmeO6FY5wU5mf6Hs1z1bcxzwa2hJjhB4
8pReP7aXf8fWBgKt9v5sO/JzlTOIRJ3iB3B9Df+M/whglBNizDv+t6jChcFGqKCa
LTq/pMrY9rUCSHqrwr0LGWOceRVrmR5i4hde/2jsXrUA1HfEFPC9P7cRljE97NqP
acikibwU9NCwKaxpUUvV+xiWvGtnCh/MPTgxFvx0/rc5zH8iMBvZ61ab5sSssYHJ
AbEqGwoDeg781eFSjjeOHzTFfpcuuDzy2pGnal7+l3rHbJVmzT2jNmYutwJWk14X
0sfGMHzN1zNBOS3FkyH9Mr2WrJa/TUo2O/By34nVEUSj9Rh4xcKe2xJCkoxn9yA0
A1ofjq++h/FBKFDLuU10aYfgKda0yMyid+h5yjIdKtnhOg8anFK+vQ7JflMM04wP
m2KI1+cU8oO2jxovIp4YzsBdEZgGuLyw7sqPBdZFZQLATSEQAMwxJ4kOx90k2LQ/
ZXE0Nru21mZOBLeCRuXy5oXh5V1yCRnHRYrXFioz73JFAqOLWS9sHZeK5K4TaVa3
Cj7mN4fwU3G307zM4J8LXLl7n8QBTC33FoTjkOIhn16qphVhBh4uUhn65HOjprZI
xM6ExgO522pPIez6Nb+JzrVMbtToaT8WDWk4qNKDtKEOfz8ShyAUZ6Tn0DgzeXRm
2xQBAO7XBAzbtlRs/ZvlQt8/Lj79FtbYyGRZuakJtxOhYcR9SQ1JC/VtM9O97kcE
JWslO10y9dyqEJT5ydT1X+YBHvZH0I58quMBMrGGCHIPjM1r3K0Xj/mo3rLQA3TT
u0QNzNkHVD6St/OeznRX+694nYO/A9g9o99vohcTnyXEBOZjbH44TZ7CmfQXao6/
68e2WABeiVULKxxV4Gl6XGqc5GtOvenQhPvIGhn4QcvSmNPycWTp60F8fpoGUzFp
VDFt/K+6CsmulvvGMOwkSQwXCHDsR55nbNhrKx6mY9WOTnyHX+MxUeKZPjIvn1qm
q/gPz5Oe2cQmuAszhMg8AJ/TN1R+sQDwDsJ+VnWthl+E+xmHQjmiL1lUIC69Ksb1
uNCregzIL/JxO6BNnQV+M6v1RjmSBLKaDaJ/tWxpKE5zR2N+UmyKp3br5LD6uzUu
QjF2Gvko10pNKEfaInpAok4HIES4zgSTjjHartoI+crUgJ2ZY3K+LMclWakngG6E
wpo9AwquFw2RmwFO7oS0fGZBdAuV18iY0wMwdHOki2dfCCwalE14THYk2dyPkpSj
Pxmw8JsgOm1xj/fNocnHPtUUL2Ai/T3n9mDq3EPFiLvkT1EFLofGwl4I90nPSbjA
aj5RFXWx4vfoPfbQFsDPu4tR6vNnxBvFYAI4Hi5q/4A2JnNX1xq+zHpx5dewG6/L
4mDEIJG0UOVmduolyqNkoOhIouQnpWB1HXoaYdQvsXHq4HBAHcIsGzVQ5JyXD2PX
7nQE9GuQlN8KslC29+Dtd7i3aSh7q+/2N9k6CAKeUCbEvuIhemJtf4nEAmvR8BtC
VhWgvLxp0jg+LyIqau/uWhGlAslureRWQ2xgzISWdwX7c9C9kJfLSqVTcq4kbwcc
ci5JSxD4wUbwe/FsnIsfxcLwMrCR12VPwXwjn3sXnakUqqXZQ3lTGNWuge8MUMXH
4o0050K2tySkdIOzvatL+NeR9LOa33MuxrT5iSrx24Udr0fYldRJTfBWq6hHUkVB
pyP7s11NOJwizjX2IIoNDR0VVB7mjSJ70fKqkc3NChnrFvQvKld4S3ik/rKl/KLa
R1Ek0jxnBDXLcn5u/38nbbTkT2UG7+cabgFJyl6AaEpb3pnhKqfEfBN+5V4OBq7z
vgH2HdfdYjx9njvVPZUcmXgpNhyKQ4cWale5ARlQ3Ea39ygKZa++OLcM8UJ6GPNS
LVSpygtODo+4u/6U3a0KKjgtefSIqB38P09xrzYIbQkVs9TyBjUa8gWx2L0toUVb
FOGNyuET5ulh0iTAMu+f7KQlM/mfNP9a6o5LnLFQas+F27TYPXSD2aUR7Unimw8P
+DoDwEIa/173vtULRBzfeTvUnux00G1cEnBaLJX0ZA/2wAt/dya3YpY73X9Ei7+N
YvjZZtGrns1Ne9lLq1opQJgjPJfp71zwGUXb19pDmCLOr4AieXNxG9NGxWpKzFOy
cdGVz3RjqvbyYHAdWipIJpYprZ0MwoXCs+q7Slv+BVkQZwdpIYMgICP/b9yfPQUW
gFw+ENzpimBdomNw6Bl/1Mu+A4ts16+OD6T2TeeujeAWMlrKopnSdT6n7Y+y1JnC
UI79hsTJYNHE+WcwxaijC+bKMLVvjatLBaLw5HVr9+EslooBcUb8DSiIpyS37Fun
1BGklZNRN1ZNbCcHuULnUN3AgFEg3yAtV53is6j461HJRCdAuImlwk5zZhwBnWEs
rEgfEQdxs+LRyxWFQ9/8TLKj+cRLBCgp4n123iBakaoyWqmkmJGPeYGzHVlHyHvb
JUciVKcGcRqwSA5BAr+bUkmGdRZ0uyzg+XYjVi5M/fPsXFvUVV5IoFzElg+LwQON
3dRU97L+eP2sZtZH2A8u4FQNfNhYKLZRTQuJ40tvJN2+f16/3LMh2W64WasmbQ1v
5NZNs0vkfDfi7t8xKnfGwQ28pY1PKi2lpi1iGgDGUi19NatWoMRMv0ZW4HmRnf8x
yPRrBwDdqnTms5+dtau6kQY8tDkc1ixIKZvPJ4tIRvoSrtybDfDDVzU09EMW1efD
T6WiadMhc+GpQcywIV2sOdKrha9Ux0lOD5nkr5fQ2bVN5DYENjJol3mHkKmIF0wv
VGuT3HOYbwcOwW7nim5AwPM2/SMXJKmkK32EneQ7SFOqRd86vHS1tLZzr70lAhUT
8uIbXn8bIGEgVGLK0X0LG3ipKeQ1ihEsrb0b8N8nNH6WbnVVk9kJfep4/WJ81RMQ
ulqykLcWz/wYMl43JUnKDIAcsyvmRlIPzSJ3u069tP2HQkUc6M2NiKgwJhNxZpn4
fFC6z/5dGD8joMEJERVVWxslsaLMXex6TjjNnyKKb5odpgULL3f8SgCDPWmXpWLc
Z87pTUJ5lHh4kiSOm0Jj38QB4S4g2IEzUUYJaouhtFQ6qmAJVdC49yjSPE7wc9ob
Cb7inEGR/KyXf7ZVR8IQzsyJTvETI/sLwPlM5XcHbqhj0VfY4T68yurQv4dLuFXq
dnMWmvnBoYY/2oOEP25kORVCf3BHdf+WTMzgcAcDHGk3WPPUgoIe3j91F/w+vp6u
83nnFanFXQmbq/91vRmTHMhrxIjf/bFlkKyVjvPX5BRCY3nJtjz19gymipgie1nE
VJVoUL7jXBUbotIQRYKe/lA+L7B7uIfpcE1gLUCDz77DnqtYktXr2VO2JfKBLH1i
x8+TmMKSW/UEfpbcX7lGzinIK40655lJfH2QRHYlRUa3rjrUYWcoKTsEz+6ewbIv
HrAiihQ0NjKMuCuM1adhFD+TtqRAL9go94DkGH9t2ZYKXR4Py6y3TpzQwyRnPcrr
MOXbTuHPZGDIOLN+0bfs29nwVRQYJEsCD6B/FG5w6OZFRCd5YkNEr9jGCV7vLQnM
87VM5Y7DPzQhe+V4nUrEcbku5fvX3Gr9qIN2rESyP5YBjutHbzOVTWhIjCdI2JuB
2KkXnOUXfJQ369O+emvoRnqMYgWJGfSLyzNCmTzcv7kBUuBzxMT8M6McRTim71HA
ADGkqkBu2gU52M3k8Kzer7XM8EAZcCvo/YQ7jSoRjrCTPju4ArwZikbYmMrJEHcX
pg46rumeDxt95eGUJSCoHDOdibtgx+HSHdTErWdr8O406LX/gRISR8gXjQqTmOIH
qWun0Zr5hdEbsL3FHIBdOqn4rZk6xpUYe7SPLKqboD8JfsYgh9makUAnGhJ0cgN2
5n2FZ+LM/Uyn51ZpK+Exg5NHg1qRxRTlESMbCg/ZZAORmFOvA5W1Z06yGKw6oAqd
Sqbxf5+zEvmIu8gJ6zxhXv52Rdu8JFjKdDWGOREn5PzlAJMmpFDymafwBgO1DrZy
FHS6o1uFJGsnjB0t0mwxquAYU3Ywru1kk27NvczSctPTUtIEq0/DdDp3Br9XMK/o
yKUwPZJmdACvAeePoZWGa1gliHYqOWjgAGbYb2KJCgdKHxYRGhMFbtV8/sq2BgN6
6W/T2aA3vCxpIn9o2VOpcyfY3EhmY3DD0qgrKHHN0haRyyF3MUCg6bgLTszdrGtt
vhsta6R73VJGE2VrXwk4AVolYAqSZZrX0wEjfinE94RbC1uEkbmQBY2ZS7oSTv21
EblboVeQF3UYYwfUe/MbBP8QfD9frRM/o2uc5AwyYAm34kQD4K5GQ6InUW8P55Bp
6NshmtM4f7dOvqnZLWracGxhdr5hdCJhMmxlrAN1AlpswgRkhOUsQDdc/gqZr76m
QgAIVt3rtsgtAMU80w5UoTNKKdLGHb5shAnBLrRBUb93NJy6UcS4zwJ80ugJUW65
Kf/u21qmfT8+Jalr5HgRILMRBTzl2LxqUa1c4IVOdWvcqmZAZH7nrrhHc80M92sa
pHbnirQ91Wl9+vttnBlRh4cy32rhSYiUsNeItNTlX16iBZJbH8XVyrb6J02iFMUu
TME6rDe8H3ViGVUbj6BKegvVgYp82lXQqyXeiWNvlSDdbBbxn87fOlD4TP8+jvor
4vjvyZxrj5dEIO4qWVGm1JTbbAmwV8hHdC/q6Ki5Z37oY8M+VllZ0PWdnj6SpfVg
sjAKIMmiGQ5a+W4n7GYynSqXZ132mpKJEDIt8tfPRg18xg5gk0Sqzykk39JHSV89
Mw4xHxWBb6w8bomwa+6U/3DFCCxZQr/0lZXDlFPprx8zGYAjWUf3sC7xnZ2axW2y
O56rgxJZCoq7O5yQ8cIObyj8bpQH3ExQXG6IFJ4Dpk2gLaZnlh3amKIO6xYsjPEo
jAaJSoWwynaha9puta/VKp1aZYsRy+6Dx7nH0RvaV10SzShGqkp09U8qpYqyCIS4
voXicUF3pNwnXtJcGMiKMKRwqyi7qjz71Fe1ymm3P4KZylxjhmjTHm9QaLhLVxVZ
qaf2oRUG2MNsW8uvbDM9PAhUeXJqnHS/r3+4f+BlQfAw9RDjf26W+QoKYzlDsI1N
gQAImaQcoa+letJN7VECyS8hHpKHeqK6iJPh64XWGzgCotHvMevw+Cus7EMbvISH
h7V32sy4wgoi5P6aPJo0yhMvuZrYdhDM1w4QWnsDf6+wHImNzrchkQSyukW2bc6e
atWKPvV4KhaT2nR/SRcpw0ryr9u8S6CjCKSo4w1pZwJg7FVA4VARVEUYz+Bn+j7B
lVw6mMm2sCO9jXoTaEgrSWzPMXOYTsTiwsKljlN+maWeU+fTxAMIHaXho+QC38Sl
y9+0Y7+uK0sRp+K4fRgpRgkgYjnqsjHEUZtRwl+uqN0DbgoQJjyXp2XFGv1udfKY
Dup8l02/5P8Xh8oZNbLL4jOAkDvil3asFDl0qEvDKpdO364bqwyMf37OALxIAHmT
Z4Rwf1EB0wZFMZnyqW8/5UNqYHPk/KLFn40oTRsL3FgQszGnHK5ajOywBh3WXnHk
sOPP82Zl+UQMrfWwbPkFXQFAvv2zbIhdtCXnQRiRspkhGj8RRUV3Vtzc2VtRjiRV
Kuxt+n1d66bJXlJtNjqj3l3wP7nNsZuqcjXN1ZplSvIBGEeR6o4H/LatPDIHrYjX
Ivj01j9RyilzryAoHri+9vDy2zS7OYR65zIaZacxUEygk+0maxlnZLp+YDbfB6Nr
Z87kNip85zjDzD+nNdyccp62J9MNuiYi7Y8yFTPUdOIXoL6fMZzKqujTG1yT9JQS
vNCyFPL1a531iEKmWnDccQxQR0yuaQ+3Zk0SNdQMDKoTafhhMioOWrGpkTuH6UA2
+cTdtxvTxT+j3PM5Wt9HtYJJq9IgYTFKLcSxjW87x5c0pwBvEQBnViiM4e2DHX4g
uWulPfbRfOtCLmz21MAm095kayULMRdLuJS48IBEDpzE7IAh9Im6QzVVhy280JMZ
YsbwwSTCpmiE19Tz1HX7ICAaEw/jIOfHvhrk2AZwJKZo8XolBbbzFipfUS5ScveC
sFIMiyWG1j0ah9wLBxjv2P0a0JYmsXupMphcTqk5LCezfAvHUyhausPnBPGEj4KC
OD74QCtxqCWeaAHpxyNfepbfBTvjVgsySmCNh1iLJZC/NS78h4XSS8dqwO9eepq/
p7db2iKre0IsOHvP25hjib3d6tfmcsN0TxSYh+MEPEKkXd9AYNi4VPSVgAajH4ZB
NhrrPmWjoBxfM07Dy2Eevv+NZb9PY+uibCeHhYCWcZjDpK01duhI7lSpJoiE2C4f
hIiR6p3MVd6a7DruvBWOvVErddlg52jYXRjmuhErneXvIAZ5Hlq+qXduY0HsHnUw
u/cwk6xcBcBg2x6luNxNdPOpvflObFWyk/3LIIu0Dzy2lEl7P57HdI8XzkAmhnAy
JGleaTQrUM/ULnddS2Mg8xStNpFIHHXAVArOSy+0uGG9VlFUGtfOQDKuTt2+hhUH
6+sfnt0jXVJigNQDMZ8OpUMZcwnc5RniLCqgXPFumA3Cb5LY1WJVHWM3rRow9s6X
PQaTq+WHmpaNY+Y1+c9dS7y2iXZtS/DFVED2OFu4lERKoUen/7mGYp1DS7d6Wqeb
VyU4YY+IQNGgw4y6S5CY2wnCCzi8faF+OAljAc4otxTTLGjO9vZ6rTpH6vFPYqeJ
pdO6UjiFQrQyaBcaamEiNGkv8u+KdLDTke77mIStosHjjT1KjC+vF6KzNBoIugXN
9H8hROURwmes7pWtZVxB6MM0x8yB+tuaX7STIORKvsSJsF+kyL1NRJROKXm9jWV2
r8LojonZgVSuVMghefXSP6FUjruNLje27akO1qXAH2hbScf+08De+82zVpeHK+Qq
vfJjN42Qet5VQpNdnEjq8jJDc2A4boCaApLvevU73ZJaYkhyphcYcZCFigNchHHt
DfzvncaoimaGczojx4+Kwjf/HSbx63ESaRLBSvObrxDolht2HfqoxzdxWnlNoOdp
rl3DaH1qIM2oZN2R22jZcAglYjsI+mnptnZ9uUSegzJHLiZ7RbXgF+YgrB/yXcyW
uGsTC6eZcv2tfBvgnPSqrQQ26/+IwROi8XeIOvEo7U/xOJblqz5HNvWs33gLbd7q
Y9AOxREp98FuKEtTBi0lhRhkcQl+dCvqofhYbmKJbB7wnAFPKQ0Tj9YLxfqDNOL7
/Cn1iyVSPm8KpEKdfnMFKS3tUHgNVs+EoqZ0UUo/mKD1xYnn9gC3ojmzAkE/SLQy
WrNURoVibtZDgk4jFpx0io8nZ8fnutlV+16VGfrccG0rJOymMgF4CrsDtHmaZu/p
edGoXL/k35P0A82sVO6h3X6nce1FNh3BQ8eVY48iTtM8/Z8mx6W17u2f7kFxLQ75
NM5SkVBmG0eh9yOQY3df7zMus9huDUAeuH39qv9yneJLuIGIZOpg0Awl+EqsbSxZ
WQLKY0ufebDZU+FTo54uwsAo+eWR11OzYaQ4ZKzinw4Xb3urCCQxqDq46YE3qhIO
KUwGf3bSCllxVfO9d7kopAkn86dkhqwsMv9THE8oUVETYrOLvVdQ2/U0T+9ce9BG
lbctgP3SbiJ6Y2VcSUKqUSs0D4VP4/QNlTxOKVW58kRaGRDuJulK+Xi1/04faIC9
JnGwjr25rbnxZiPuIkg++9jtubQBd5QHWuZKvEToK1NIDKZHuvH83bSbwZ8tIXmQ
PpRutAMSfD/sukH/iKx9S8jgGHFyCSll74OCFbE7Dw82kSLX/3DlFSNv38riddym
81HoKFeGYVvatuM8gCN2iZnQ7iI1rZcQh5ospNQk33fERf4n5B5e5J0etwHhUQN6
/Nhhj8OpcMjJsH0i7NC56n+x5gyXl1IsuJ6WXsnaEZ1VSIpVYUsA+U+xXiA7JhKI
i8Ikwp7DDBP3z/41GtufWdmcIUJ4K7nqyX2LYrUXV7yETq/cQCuoKe6UGaCNXSW6
gGx3VwlmhIeEL6eiUkU0GmGVOSGCAUsPiba42p7bAOSP38PW8WYyrHu5aLTEKOjM
2OQN3XOv0xbtiy7Z45v5zQVf9CafaKcCDbdqHg8TTtT/PySiwbhPZc/o+ZZxJN01
BxOjJhPrT15av8A1z3l+jMpZYlnqGTtjfTsUUFGP2XMn/Frl4w9PeakitAp2T27P
GJEtrVvIHvbydxkGx4y2+YgaritVCt+PQwoT8PTzTPg5HH7Py/Q5csIHYUPVC129
vw4HbYzcZ2hjs6KxUOZAngj5culomoof+PRv857w5zSOFTQ8j0w4/8R1ecl+alms
M2jkvtmGeZc4HhqrZt5kp3OBCZWQbZNwVtmBslUBCmTOaJgIOhneFmhaotGP+xcy
+2+WfTko3EgGjYYUAH4zoleQSWmLrJlBxKiyFICwzaQnFZeJkJAS6M15ZYzBFf3s
RvAEBcpkMp5f2PnsiIqhlDV+SKj+JO+ccHT3EfQj8Wmf/iHt+UMXDPmsdkTTDcDx
uteo9SwRB1/DYhOEYphJPMKQz0agCGFozRRK04OHKePgLOp5MbUJcz9nal7jaJ2B
m3C3ZaGqcXRUmq0BUCfuBQQgRloZWxa6lr2wuDHBeAYTU5YfFZrcG8l+0YAsqbib
NTBJg0yIdnn/5/NCg+l6O1A4F8gq/p4kPMrGJofRc5NROFX2S3Rjpqi3xmk4zN4u
IlutpUMpWdLHCPGrR69rGmeBPLphNZK1ndvB2jg9Xt9G6udIF52hseDuZw4FEcOC
KidtBVgyUlX9MUoa+HQKrdMGw8a1Be75ZvKBtJLXwhUjH/Lq2p4EqDOxUmlwJ9Yx
MpjI33TxRRem5wNVuxv6jiZXUyHI85PIu0rZOnC/STGVHnDlONTZe/qwCPUdXo27
x1cVXeR00zhMrb4lRbP6hjzJNze3jf/g2R0j4iv3ZKX6bLxaTwIJx2uwy31yD40L
Ta4qDwFUQHuhicnCSdcRTZuwIPi64ZM6g/72fyUZ6lJ/8DrhW1+MmQ24oGWLMJ0h
aMVQRaExaLCUGzCQi9BP6sySd/hhTGLlRb2h2Zr58I6VHas19U6WP/ARTomE8xD7
ovkYxaiwS7nItpETGvu6DjIpNqv9Xl65ZYWYZlXAEC60Dw+k4leAFiCIqxjhkGzy
aQHucV1gSeZAuZtXTRSBgsbBg6TXYAogugB36wxIPonRGJ6X53EzNnymuWIJaK6g
W9t3ZaXUolnZfz/ZcAN9H3wYKEIxLNDUI7QIAb33jQgVquDkrSSGwzntYnLUNEfC
G5a/3i17o1juAIsMrbDs0E4skmwpbTWGAiKB18ybuZhBW6EQ1n47JW9ck8rzpMxX
xr5/3R9GUkj3VX4ZythCiwRb7NOP6MnEkOVrlTWLSNNAC47orAKdXqGY2RE4GDmD
lUnByyvSKGB1AY9SuOkNM8JhgZQybKhrJbG/eq8q811t3GIUVGvvIAdY6iJFxOnT
NI7wsGAqMETaNg4x5aOkfQ9TZUDOLKGyib3ODM+URZHQk5mrAF7JKAd+Uth3bVwa
JiZ6tsh3AtZHtD2KQfd0BbioTW6AXOhykUhjzKhszf0mlEw1SDkSLRmH3ZGV+mZh
z6Gj+GurdKsj0gO44cSCk5ZQiT+pvu8hnvQjeb2RYFaU+Ja6a1+dovvA8Zz6DPNT
oAHHEuRYr9zmrpaiFwsthKUuanoY/Dn/HozbJXiapupeQxVwOGiZn2Z6/JTgFdCO
WbxQiEhz/d3MB1cABJiNX/NcmpI/kQ3YBijS7u2Ob3f3ktQjePA9SduRuiRRNpuR
8cuOcTQjaVcqc/JkJC5Setw9l5qZPnmfJFVxECkgwlMLxix4jXdXD2zOxO0pVrlN
rU1BrQRLyTqaPbas7blnLVdTv+l83U1ePwMtQ+51csKUn5LgG9tT7MLdz7ol7aN2
AtJCHaiHiBF9QzlatqUemMvh5VwOmTlP1ApN7KimxhHYkhN57wG5843dtWenZPhH
/eS8lofRtfeB75qp5BZw0/NjobBfUPOxXCeRPfmFHYcnQwDt11xfOBa/6gDZozAo
x0VqPDGFclpsV3Y19f5QlNlMlixDrMxTN4vY8dX1FQ3hPJ02VwCUtKFgDdzNn41A
2CHUou/M8qwCZj5d3PNi9s+Lp3Vl07okzii/Awa+bF1wJAKX6tCyCriNRXIKhG0l
cU8IgeFRizGFXss66CZu7doB4yRNoGifJ/rEAlVcPCrUce/NI8ICb7sCazsiKUxS
mjIFLzxQJ4iNRTyBnMb/qMB+N7qiizlXs8RmoIT1gIPF35vxAkzsRmulKoyiBfBZ
eDz3/6jdd8GjcrlGUtN4t3Fod/r1uE5adNH+BfW+INGlR5XzrnkOVnJAz+K8fxlS
KQNgyeZWXE4d5+n8f63s8e3sQu9HDamJtEsECUh5B7J0XidRBam/7H50Xh2kox4f
tm0v6ksHFw60mC0uZ4qxiYRAPtcwS7rdEIiLUxNlL2VMNIGp2wD52Lb4jjeM9KH4
n3ielOs9Jop3d3YUzYGgiCUr1PTViEptAPnwavGNU5p6jL4H+cK0tHgTjuw3IPw5
gHNXL97KLNBxCwlbaHKTyYbYBMMIkHZt0mTwT8Vkotg1uaN0hM72mxIPBsXfh8v4
KCrXrRi4VgoznKujZHECgH3mI0p34pEEmP8XRnA/4HiL0enDVYnxcGtV4qO9yjYY
XIPR84k823Vacp9pfNcYdVC0xnLxhUTlmPEVKsnrYXPsIC00cFGliRDR5OTykRvX
8CQsxF0mzyQcCG0ylgQSrotdIznoxDzYUfmJIi9jIb1dIar/SjoT11jcCQO6kD4g
GnCDXfL5J0AH4z0W4iv1Dd3lz+dgWBykkkpyn3Ux1TrTjUKS1gdKoA6JAKGhfpRi
tzO2GAXXDxk13Ef/oohciiKOty6gj5viwMehkL8Fe85aibbLGkUm7yckxQnMXFOz
C0QZTL18gV2I2FQEeZ/nlqNvW/yfbzP2MhiSy80girRuVPI3QAgtKFs2b45EqoeY
eybZuSJYRRqcQ/4r4PPIebFHIL9uuryXbL8gM8nziJ8Vu5BC1F642lCvHyYShN5m
WUNQq4yNXvQ0FLh9EHj8+ecjl90ZyPZ4JWI1u/F2OrtShsFNYWtrTcBUu1SImiub
3XkIub2Zqv5vhev8j6i6dwRFFwtW5iu1uTb10inkkIxHl0+ALHIY8YG6KtL3foQ7
63ajcVGJQQUR63h9BakeA6mHWmnXwcux76367TodwdTy4xc2K4J8Y8YBiwpAFzyK
gBy7pldnThQjYETedJfOsuAR/tttvG6BQ4jYtgG4dRBVkROecXhmwi2t+zhE+0eS
WvKlTJIX+DmSCQpcIArmEDsDcOe7vTzarpwO2V2ZUDMCau7cOxwXcLdApG4/Xr5z
3dNno15R1ktP/+6X1CPc/srPiiqJfsqZYmUptntEJuYvyDWE3xMf45A0laz9sPWr
g8hdaqvdyVTkkeBCP+4VjkFj7pL2if7DQ6hkhESgG7yLnVdARkr+Rqa3Jt4Vpp7y
FsW74olJao9HFkDJLbk0YgACGBa4H25c3zK6A/pukJPGdUyJBl7kRw4wquxDkOUl
NBe52hATMfVdo3eD0m37KvqIJ03rtD92RCMsH+eurMW7l2doXSzncQ881KpGxMPl
oVpDN57UapPWHCfis5RKTBvebV1eEtftJhghOls1B7w8tzfqZS42LLVEOdq2+xeT
OEs/P8Nle6a4aRhVYQeag46hysof0cPrkN6DA7/OZUGL7fQXAZk1C8bvyg8CBEzA
x9UP1YEBDikt8r3Za1U4n51Fcv6TYZF1HjRHcJKY3MYWVbiSdcVj+Oz4RQ3WHflq
Zov1dm0lPWS6LUMVwPAIcysegzMfHrQuCtwxK2wUG4JiBT6NU+dBXeEJyRhWSunI
++l+hruzzyvbB6D8Xi70xAX5HPcQlA60VC4eJvgD+8yJ1dwy4jKo3gw6owlcLqw0
dQ0nY23FSd6/TZDsVGq7xgheAqbO2WE0qlnnwqQx6oCCYgkilYx0bB4yTa68ih9m
srMSZ3atxgYUICuPybv1ljC6XHx59VzTNFIxLqiM6S5ksMZGz4xpqWs4nwZzmRqv
5LGU1yqgOyZtRH/B+847IYZJuxSZtZDbSsiw/eG/Ty/8f5LwmKp4YdryhgafN647
uptH0tPhLSaRDDkRly4n/nP854PdTfpXfDSWGjaDedkrrJD/Z3dgDiqHK/KoYPXo
L+R0jyDMJRK+FhcpMg85eSILegMuG2tw/rvz7DhSadsJlWaz9TCswo01cLuuYziy
E/tgR+W+WZgNC6SZ/AbAw/f+eCyZxDqh1P61RWrYi/KkKe9UWCl5XirOZTOyPL9I
p+C2x8I5E94ERfOjv1PRO0t4GR0LSng0ojDBjz+I9ArCnorlyFto5fxnTw0kZn/D
mDpXS/f0kEuUehEQo/4Q6+kZ9mRiksgs0suNCoBwOfdrlB822JJs84sXT/ab9qJy
og+4LXe7w8rlp9MWLz0vHw8Vs0C+/GG99X4Xkw5oCEshSRGXK8+EIEIP73Ifxog/
KINPuJuhCU+pvkNMpRVD+YbUMeBmVhEjPkNCZ2GAa76qQrAfUcrFgASoG+9BXQzj
AibAcNpEVNKtZn8X4e/I8d4KLTxHf5b+Imjw3xUNhaXk2eTgF3H1EayuXs/Vt4t1
DQHe+kqKpOwm2JKHqmuq56swDwenKZlDqdIw3I8G6NiOMcDMmr4rguiK5UlxxIja
BEPEyNixxdg7HibE1TvbHWwvKMXKP6qLUiOgKqs9QF8/sl3PDWJ8bD41Rzx12eo1
6XjRPaHIoU1betX3cBdS1XH8Hw1sS/LzFTZCxpcCsCIt+FxfjL7RoJQVAlIr1bIk
VIPtjQOWMzbQ9lCYZmRToampI+Tbwz1Vx8rYI3NIgF08+cMVqL6wuqXUyhHSiDl2
ZWTifDc8s/Sd0d17tyKEkbnPktrQGMiboTS5VjcKsRyZr1laDJoFlX9OJNGisz62
lTedQCdBszi08PqB20/GAMrhHBvyUTtWIwFxh2JJcpg+1kZadFJVzBpCcELdMD6Y
iAbu3dI2NDdYJ3bUEiFTYiqtA1DpcdgkRrpjdqIocPTVacBCEywcGmSknl7fG8FU
gbrMRPPm37DBLJrTDsJE+qSlB5iDXhAI2n90mm9vgyROB9Ohw4KOo2YcJij6HLYU
vxRGAWxDUMGbcUZBg7HVH1nXjSy13ihoEfXP9n7576EsEWlWffiLI39mWKfYivC8
hk41Njm47Lfvw+Awcs5g/+an8OJ9XAmcnLKUFdkbPK/LRA+RnKmaI5ppl+KRvbhH
Y58jqEbr2D4TIjw9Q7VomGUu1/p4o5dkn9Rxw9wtUbi+0UpUP913D7uwq5Hbp6lU
b+yaFe26KfBmGn2CzH7GPSTb4BDWjz2vhIBSB4/CWKbg60yvtjT13OknGht10x0g
IKV63kFDCwraUl49tnIdqzjqHmStQhJJ0nZoIKN91IEKdvrJlAd4altPswG+p1oy
nGyQjFZRRa/xV+gnLVEBfPqP8RjeLEk4B5+9vpOxTJ6dZTICKvs4Zgi0dw/B/8OB
wgtk8pPW8EbxC/uPbZeqMrK9yFtStDW7tQLNbI4BpEom9pATdAxzW2r5bVUg9uUL
nEJV4bQW7lwW4cG/EtOQLM3tuAh06hn4IXVNsR/t982ZyXpNEPz6psW88WU7gqWY
1UXscWCIc3zoyIiwzzRG1XawUPKzS5Jh/5OFM88OKvRKPY906IeB87ZccOW45Pc2
n/Sv1n5DXfEqPAlsUuou2LVaUd7ARcBiMoCWs63FZobHdf7+rjmPrC0pquPNtLk0
jcDJQi80qP599Dhi0UpPDV0KAnkMUo8lU5lW96ug5o8uOCMc/8lGLF4nEVMWUHu2
AuJsWhFHAYrDY8Zp7P3aiD4CMz4hgbeWk+FosslURy/J9LrH4eZ9TGaH1JMJxVhG
WedxxsuM/oCN+R2ul7qn3Gba4vAWseQ5jv1JlSpqoiHd3SUGC826qUJluK3mlfrc
EWH97m5ruEPXx6FCm1Gn3oH1Skqk7JgzkgHSdo7hylYvr07xK0UUTknzNMZidtx7
k9EZGTmxGb8OC2CLANC+IeimTa9pIREmZpCiMbcv5CMfQYAWYdFsE6XM8UYpDKNm
GLNnAZMnjXZ8EeMMdVijJ2zTQcJSaUfXjU/T8EmsyiMSUqzM1fOOai8qEXc6j3MY
UNyLbQI3xiKQ22a2D36KfpjcJyaoPU5zj7ow9b1eojLbZvALyBSkgR35+WmIPtEh
fNKHuBQfAaoVAVhpOqvffzJU/Z8ejYqHIF4PPiwL7xD9v3clqOnyYQUe/0QXyruC
sMIa7Rv3X5am93a1MNIqVqiMaVIvOL5Bl8yes2JHUIU3UJAXwyJO9cwq81y7E4z8
PaEVrZZ7RI73S4LrJr0Ip9rXnW+Oo8fdoafAgPKX+NuTTyfstN6d949HpbOxwoh4
W+5k1j1kJaHpyeuNb5g04DjfdHak9ljjda5pa/GkJlSVc8NhGS76GxUHflsiJ1TT
9vqPItYK0tKzgB30Y57zXIik5/ZngXAWQtd7NHpMkpPTk7Np7xojNtA4+IO4PB39
NbRTbRYdPd66BZ7oe5DTHNJbY7GvRQ37JfYbKF6+7xv1VoaJYC5sPWCyy5TTmVBS
lOHO+ObF/z3KQsqI22vvTx/s4I17ubm1L0MrFKWitks6ZTYXA6dInyMY1Y/e0PhP
NMXuvhY3r+jh7GFyGqod2GI6Lpkt4AT3ZNkixjjEwmDYMZ4ujqA2GF4hFBFNIeBV
kVD+pcZmPbZBp/fEv8O818i8fWF/0hzfNnnm5/kwi8wVJ7XA/KvpH/c0eIaRjN/z
KUhvALiZLFQHE+7IUPWAmjkrQnUhQ0q8d40YtgbQyqdy18Y6crptAjnDDVgZKW6d
oeapU9Tzbp5AxhU9Va35cBJ2c0KeHOmjg0GyPAszpIedWAIsHDIVxrw0vVBjuTUr
u+vzCK4P6H3MF8y10IZv8W961b+Esf8J4mSW3OfTUN9TvyeTo/LC+NNEGoqbeMfN
krtViY+4Vm056K/kcnPSzqj1ls0CZuvnfCPxAQqBorzZkc74EZwJwhgkQGzfP/gi
k3y7GqhyxkETBauDnayqO2u87Vgu8Gsh1TM9jMJHyp0GX7AF0Bwr1vCm3aOh9Ya3
hc3z43v7G6PVvGxr3T9rCd92jumicTPMy3ZaQCm9vh/bRfMV56Hw8yPdpt9GazT+
xyV/HZfrz4gvdKF8BB2do+mY3r1qI+jemyWNIomqYYIiup7Bf/VKUx8tZf5NBwfX
U5kCrOMgNcZOv8vTCrpOVaRoJhpAIsle8xYbnAzMYKg+WSJTKkBy0KWfny0N2vut
84uqTIw6LCyxfKSGS7X162G84kjcBP0MinIS01EvSrR9JhJFQITRO+2NYkhsBSiL
Obkp957H8EXZFM280+BRHdkTNxnYocXcaj0qOQj9RcN9mySiIF/Lt4jwiVn5L4OA
DsKeok5a+mKjhNxclu71zHXLldNxz1ydyc5TpaHCjYTT+eXjfgO1Vjfxdt1XnQ2y
X40dIwySC7YEOP27HGveREocYGDUHwjHQNImPmsIqQA9JwsL4CUhxxefZ7HZe3Wf
E9WXhOn+XKVHpcuvB/esC9cgKkznJcdFSesp4y64H0ok/N93FPpjuTtj7oxhF/LX
Y83SnVzPNGfeMK9pqrtfPrrDV7O+hcV9wdwupFW7JFOQ0oUDl58KpmPrcXjJhVjq
l+Yeb+Z/S+4cRWvuVeFqQo/OUgCHSkfZBrgpbBqFDZ551BR83UFml2+yRtpTiifO
P3jrBm3JEdU0sjOR908Q+qSDZ4cCCGrmyeoBaQC0VV/NEOoaHnfFHGeWIO2JZp5e
j462i3zl5SDy+AVROT6r+PF2hOk6inxSz6wAbknqyIetaDmnILsDCu9obuk0VF3g
2cm3/a8G8JcZ3jTl1NwJ6ZOsoWgoBj5w5OMNHWTurcqcTTRlTNlxa8upHhD9tr45
OIDIsSLRiyyg6D8/A7/7Cpo8NyIWe8jRHYWuqHogXtLcXO8xidfbORXyUURZfbhd
ZjYi2RyPmEOMYRf484JDDK2F+94XE2IoQrA2tBYwfWqkvGZs0YZvPPkq/mwIvJdl
RmwQ17Aw4NMddpMa6qws2t0v6Hv2mPp5P7uHee/wSDTE9O2ahgFcRRitV0jJS+5B
y67T4dVllFQrSdj+7AfxvDD33jqWheJqLMfDMJEVQgtdSxCyW59nVjxFmXY4ATxC
//pragma protect end_data_block
//pragma protect digest_block
+z6gY0P09dT3l/Y+RcUc3X9dNwE=
//pragma protect end_digest_block
//pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
iNvUZPOVMd5Ch5fF3k/1zVqo3jvE/ewgZHia3SPVFL/B87/RvGu3+MePVF1wveu2
Iz4GW5podS9qFUqTKtmfs2Qxt8AC3OsUHpHXsFMUH/vg1dcq9dJbmix7824SQwmi
q1CnZ5F2ctamhtxMZxTyOS7EhH9imfuBcorCoZO+xp0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10944)
p9wZHuwMAz06dYmZ5rHwaSnM+HO3B8CJ6MNg55WZk+Nylz+fS3NSnRNEKsm/qXy4
5S9mIlXRMyZXkzIh1tdtb83zKV9ZjhNGlRT+XbWu03aKHWfXNliZRWp21z4Wle55
gEywd4gM5AM/isqTA+Ti75rsjpyLo327h7+fo/IhwKvw9pDzK6el/caLXv9opIlR
xLojQsowhuJfZgaqmKhmhxV6bQidLxH0OxGxovGougUvSA7KVD0ckxqQmtg5TAys
CBo7X2ZZYFxScgXPyfoAuGPyOEl8nWhiHjpLcT/QH67cFbSF7sT4nfMACMBFtAlc
hdjLTsCinqwMD5KaDsGL3gO4qoQ/wanAGcZL1//8TxTTvW8vhdInGbWWaR8u65IQ
B8DeFlk9NKJVN2PWJkpvz4O7xzTv/KnsObvyXa2BRbHKjJw25ZdV5cULRF8zQZ7i
aHG2QNIwnquBq6m1qHri9ShvG3SnaHkcl1O66yfltiJ4RhncbSArvos688xE/P9K
Vp3LC/owZWHgvry1omAZuV++HTk05buM0s4sthpITqfPWP4bFZWDOQsCKzzx+5qb
RyDo0OC9NpkUBSxHEMu1PSM8NdTknMg4Kcm8+2Vlyn4W6Wh/sVrrYRDTui4wIfox
jb2jNEOOG45XnvznZj/uVx0so2FI28lZW4x8k6FbFNyWYJSgUylwTn1jB31z6w4T
aam+h2TozDFJiDncCBzWBxjvf7bCVJ9NbY9ySe4Q4hLTEF3W+wY4nNB72jPP+e//
i5TRQAkiFWbLhko7oiFcOibtQSpbJRKBTrUmn4ymlEMlS93WFG4RCyD+bA0iTg6I
+KXcl5KO8Efgy5qmGdTpOX0JP/OxJ9G/UBJTTt9lj0Eaqg1iWAhdejGCGwTfnaSU
BsRw33cEJEZRk8bJzUqWI6zsvlXqSUWBmMMbW/Z1Km/ZzFiq4BQp/qRX1iWzqyTc
zpY5GY6OlbMdfVj+K4OakK3D97AeGDTlg9eiM49AASUdFgUQtklw2XgRcazwE3oF
bGQK1DNLSZdLETpfpgfhU01jn/cLqLIoM5/ri4HhFc1ta3ktOGRJbEDDZT8jmDCw
wOidx6CQlqB3KFr+KREnTP1MiSE0urjBnTXUTseXjyobAEut6K2TU0NWVbGb3r5u
o5NjBOXinNaWzaFh0gMZVWiqVE+7atfWQbmJpDg9MSTj1Xyyq4HZop9Vf4fTIECw
1c88p9hkyUEK+u/IoFnIEsoMf1w1kxDd++otxpf2RWSyCveS37q7bnz+28Pp/wlL
eJ85jxARgPAQ7GA0kdT9nbe9O6SxhG2Sy0Auso4UwfLNezA1W5vhHueAzvO5uJN/
W0aqpLl50UuUdyA+fCgcVcBiOaS5VncKjplBexd15b8BvcIRtErU9YkC8S/rQ5JV
2Ye7JzkBtrUgmPoKSLC/79fKtWNtCtJnGumwz1kcRu7D6HEIicdkZKIm/iAWDE6T
dNsoK+BKEeptGly4sVdo9GkUAivj2rlFwwADif/IWtKY/j2R3m/yhHfd0DMQ/QFO
8UpOWNXYoX53Q89tznJv5U4nJDt98YPKCdSmOTDNlzhRh35gbW+u60ulB7fxd/NR
JDmbxfz8EbSljPd36KB1jRvFFDs0GWZLj+JT9uZjcGdbGjeqDXZJFkzDSqXVTMzu
YLjvLiTKkbGwOF7KnWJ/g5gjs1cfvr4qdJO6Aec5mjiYGibE2fE8ejivPQ/x8ySW
ilOAk0hhoIfJzwq5dmqpLgUxlsKwlgtLTConjWSEmlJpEa8YyRAvF0oGNUCasQ1i
mEgRpIK1cRq9rCRfn966R4TS1tE8Ug11TrLQ4d338dHHXgfHQM+PnGqOcr9hsYG+
5HPJnogDhZaXspu8RtzQrpqbRlMKHU/amMx0oxdPFq57deR4FEArwQ5gLLNMxPoa
B++NqXuyfi9y/458SNWrcCjm12FcR2QGxL1lkvywbRzjJOmQHK9a1Ml+cCSOrgC6
fNGLHM1PoWiZQiJX5cBqC4QvP2u6q2kG5F2Dyp2NGQK702sEGi4jxK4d9n9kmJDw
OkYllESBJleZDI5WpdOnfVvdzvTMhyi/KZa3pESovBlZaQVmum4VPvsJLlK6RTw9
R6myGq3M5Jqx2fkj+AY/aW9PILvMJKULEyPxBowXLWlRKrKsWfhRP/L6mf3MYdYe
bMC1HqSV/BepI7j68n1OAAR09xYfpsvM40h8SM0EoJW5lZt13oHd3MuxVO/q5rNy
DDHE0alHqXU2H2dzXdRBtqqYLoE5mLKgcz8W/JWo8sFT8o6xyBkjXdrtYjQCvdb2
fpbx+nQFL+stpVwrLFx4KcmiZwzDIMCm2p0P2scv/eGlg2kBWFC6Wp1feoWkhf1y
wF4AU1qC+VICJDHOr6NG7lhBU+Z7QREgvDq6h4Mgykgs6YjvK86rgZ3cCt4W28fH
0Tkwb801hJr4l8DRUsmvdn8zWMWSla1RAzzz8UcTaSpYSj+oDZc4yO5+RkwE82yW
bPNbgOrLPPfK3N3wvFwD4+/krZhW/q8F5+z3MOC9hVfPcC2WiKvXMfAfcxSNAeKK
eqsZYFc+qA8hPeCvwGFVfksoofDxM/XQH3g8dp0o6XvfPXmgtfWumkh5mr3/mis2
udzrYeHbwjedXlUx2uSgnD7y7PHNEXtaXx38gxpBNo0VXcz8jSqEtFdm9jR6rnCr
4IwHr1oG3EMx18ogvyUCZGF22rOKQgxpaVSNUtK5HDC+bXFOpu2kYd9RMhPp9gIt
BxXkMqq80+XLusBDav8A0hRULgHmQgP1POHVnD9LJiYPm4Pol1tkNJpvSFx6Fz4a
HtSUL5EZXZ+/PT1MH91LkHwVyi123kLAxAOiWgiuOhrQGs0GMJ2fFViNH8krDvK2
Ki3XHRYmDNlnpwb9N5vEkNKA63ga0shKM6Tmw0Lfz/Lx8ofWwEd6kmrYVhMTNUNN
rvrvmSOpnSEf2YvioJz6WvlHa7NRRHuIldV5osZV62YFE0dniE+SX8JT7DQaXXik
y4zaIYCr2PqInN/KdQOaIQsXi/mfGtLxryeKd8sBDEqlGrWm3bqZ/dN00Z372hv3
icCeZow6eOKtgVPbB3NuUzzFsdf5iBrD4+MLdSAmc1SsgGWWuN8q1k3fvol4dUFg
lDhGlnOlqdAxzb+8ttPloVqsSJR5Z0yJwUWmUGhH/R+Mv+HJbWk51ELEEFPlBx+U
rwd+P/k7IpDvsh/iVL62Zex5W0S5ZH61/zqOEQncs58PrGYQr9pMz7ykkIZc9pzU
LeuuMCY6jBt7MKDORgphqsgjXU/Cv09RqIYYgvrzf7oI+B/iZmWZ439ruiDxumy/
t2Q4D9T2gUxgF501ohGUV6JihmmneCtP20CXk63MzMM5BdDiSC6khHvmlNbs5eSU
jxwIQ9/FjLhIHw8NcQpHzbkh+b2cYQ/4yG5BuyaqXmCLpZ1PY1lD2YWols4eTDXZ
ENOPibazN061QLfZLnjDXGoAtwBKaBPJ25qJtaENgxiL643FqNJ4uKFl8Of86+r2
7YUv2jqgDe1ozqJyPioX39wI7yILgoFYbrR+pJNMTunUeLqmelYuSmVaGSJx1D+l
GeYwByo9U3Y7qT2zWuBJ6WN379IlIbooAU84V2Vy5AFE241p+b0MTN1s+CU0aYkG
E6SKN6Z3Uc1M2MPMaKXpUHYp6cDTCLjyqIy7TrMHXFWkIM/1piTrHInVMRPIJfjY
mNm7u51KrvmKeFJgZgH51mRDUmuLHFH7y1NU8LKfgR/v73C8KT4T/+xkOsZhl4PN
ldbGruUFvdUEfqSeCHoJI5Ia6yqdjr/pZ/RwRxiObAvAylmk76weIaVyWB/z4qiI
gx+HQ3WGzj1Bs3cym/Poyje1+Q8b4JkLlGXbaQ/kMk0YuVCWhfPN5O95ZohJ0nOi
V8zb5n/jtBEZHCi7E77ZKZNrrXmodiQjoGvpQou2WiSDLrB1PIlbfww2qzMFRmUD
0M0SE8uD+UfaJjb8vd0Szk43L82N8mRCaY8Y2tTx1ISRfwSUaiGcnKToVZZIBfyv
4cBaVbrwl11i6jGhrW07uGqg/EG2OS1r4cLTlhKUwJaXMVoqFQdDSetNrM99J96E
E2cT5MLrUws5fAkS2k2qy2vUaYN6w2bW5fvGD4iuEd6jjZTkmPPej52HldcQx/RC
Nzo+iRK6r+NGPcYrX+skVdFde6f0OKpKPePBJOx1aizCKHSqlbCknOWLZoc3R53D
CcRMS3oQplKWKIoEIv3FCkZYmVqIPLYjTho1MoTiknWJFE7UsjHIzZaiL/B/bVlD
Jypb6iOlx3S5aCAtLdSfOT7SN+NN4Wiv9t6uSgL/Ij7ABydpDi2/STQdcRTmG8p2
eDfKOfP4hsOW6IaE/e48bJ6KpIUoPe2LnvpvA0uVQQIQINNOIAtYw+FZWa1jXQ90
KBE6N91tajFabhm+Gh9SLNPRmGqJu2tSVC7FkhIk0RowSR0GPVtuJNX4QkjVbPi1
eHIpyBvoz5u1uhPMM90OmJYT+gUSybRhODNOWmH106peQIoTwZ7+O1wF4DV1cRzq
r53QRUVyXFRF16+6UkDTd4RdaEDbcWVQBaQjMH9/Xruy00R2y/yimxPQhR+Fe0WO
gZkyFIDEOINvKmxdWAokwuXfdVTD2pcM0GmseUY0+90BhSC3+u89xVjrVSm9Dhlm
h0nwm1REnCNORWjRKpgDo54aStHfNDfSW4/J4jjpkw00VhyePTJBtg1vEhUji06s
ePdLvp1L3dmt/rMDyvf4c38xW+vkIG8CMx5QseNxZ+kI73dZr46y47zNgdGWUuE+
mqNxep4cLAD4f/BL8tpUoWOFpW0fs1FbPMMR67YWGK5KmkLqt3zifdbkVGInY047
NEShFoyWHOgFZcGzQssPj6r7cm3+1plVLAgHUgZM1oeMaKsbnXCjkV0Y6yXUvuo9
N/sXl3xlAHWckUEtkQ8SmFwjD99qJwWI1FILOF721A34ealrW4hTsoqe33Y0vCu9
3GMYYZRfm8/Av2QHsMJQ0RAcpTD3mfBxxzM7HqGdOObgO2KMbZtbBjPggBFA86QF
IiSg+Fwtx1S7ON6NqHohIXCKL/rv3QQsfpNUCMrbyjWUVJHZ2TZdVFbyMQ1s9foH
/lP9LPKOTJ2TON575NbG5zEOWXAZEbDrO4WgccjcefhYTTINNhQqbQgmTHXYAr/1
kQNeO21l7KUFV29dkE2IBl22D9gDJzQIArd9ajmzbLmOz6kKog+b4EpNugtHqybu
S9uQ026CQM4MQDfX1hLxEbpvCYmbyNzx2dlHbnbO24XNYXLDWpMoBljoknq3t2yY
hOY1H3jB7zQvQOTQZrj8k+Oo1qpGcQo5fHjaZsAqFlig9QyQysF79uNXk/1FylI1
7OaDOTplk0KYzs1IF0+RRvpjhABi2eILEoPcPQGKyc40PAIur6AeDNmGVtPPUTWx
EPraDfiuYyyseYpiwdoIY1z4JuE9AsIUYGY+FMGcAJGVCOIqZUkVTP3puC8PXXdd
X0fvPw494nWjO8tr/jqH9FGpOY6RQbR0TXTLGIzJb0GR3hK6SWwOZK/hIVAGVLO/
ky8QoukupwKyWV59OXG4Nbmwk5eef/P1f7pqNODQgqs7p2MbTKWmSSeQ9IMggniE
zqjLkxWwSkv6Ed0DZAWG8ymrdBtX5qsz3nenLvLxzc/3VvI2C2g9EPEykVLqzwZG
zM4icI5oGTCSDDBRwrR4lleYh/+MQ3UetzKMFeUb/cL87d4njyXHbygrGPIaBw0f
KAF+ojbkSxfIeMQA0Qxx6+8oycD3KJFK4/hz15vIYuKMyWnxNIuJfxp0FxdLrys9
b1w+BhSP5DukjrrsQSIfQw8Cjelpk0p1ndB7miyQUIK2WZZ/fTMIW1pqz62FMQGL
6445fNcngIJQMC+Qwg+Q2xs5IZ4lKX4lYLimVXEOVRW1vpP1gkzFAY3KVdPR/NMR
ZsXchDLj5+OU4MQ35MN/3A5wxEh6+eYBDZ1cK+yLiywn1tdfYf0UghN/3Ci3EqlB
eKgEEMU8ya5XYVgZd7JGBLX9yqWnfa/GU7cxxoFc1wQwczwjrpwc6WOY1jtwgkCH
bsvaUXJGsRQSB+5VMY5y7D/fngVXSWVXK42B2qUJB44ZK0p5C2zfpORYyvGAmCjw
uS/LW0aohjamYZj6Yzd5qqrWsBnyfXqfJlfwIJJhcVt9Ie9STmMuExbwNKr9crMC
V9O7H8TNxcd7Vz79JLX9Uic5rvtYfwFf57o9fTUrflc8Os+sk7qbp1MbgjonT1tT
Tx1tPugHx9l87B3vdnDv8SMKTJotXI/QTDqKtl31XlUJioS/4zBVWKP5SJwOwyJT
5qyygZRGkV/F5O2oVUQIeKrZu47rbQqiQz9Jn0nVMwb5dbYRzTv87PGw/8m/e0JE
p9j0r2l6KU0f3zjt/YUfwxySED5UrEUJNmWiI9NbM61HxYQ6IOatufLS/JzbwBva
f3lN6ANqlGm5N1gkRKM38juLMIYnXL6H0XLybkwN10WUiqbS7We8s/L3ippi1XW8
J58dHsxMFJiViTCcVblq81jEYPIU/ayLgkPArHKru7tYClaovI/x62KU8rTevB90
gqskY6QEh6B776/4qnE8bYhEHLCnPGJ7K5aF8Yb4U5OcBb1G+F3ucYmU/UAdgs/4
vIzAGqR1RSeVW7PcQJ08oyveMeiIiytGJZ+nI9QPPaAOapYB+YExmdtspmWu0CZ+
v0J8gZYG5yMY+THaxgcWOE6xZL2ArxsERubC6AlKXA1lBcnwXa6Y+oX8Nar4p6SC
NRhNvvcDY7/ak5isz30ctZdO3/CysTSrmTLcmRrILndM5g9tJLSJZqyBn0UiHRc2
0BVrZ3RZWGxc/GV9H9xuvglthvWJer1j68OU5vTMP3yLKazNr3TTmp5vLf0zp0LI
2c91Bk19RbVBj3cu9OP10elCTCrRxBJettYBHAM4ep57Ek++X7nCLkZNaJ773ZgL
9p8xaGVHF3T8bOuQds4KIRvDjse1MkTStmgd8QpfP8rrrni5AZZdn+98YN4hzbT0
LuqPmnnMAknpob0zG6ZtKh9X1QnZk/AO/F9XclVHTH5SXQEAZH7DBPfizadVqtkm
i3YxKFr8Do5FOQyIOE9y27CX+ZfjfxSBkXpMQndvCcHe2MftUn24Vh9RtmV0JvIK
RcWxIrAt4NZJFEmvcc/WInR9EZlrVYDtawb7a1GzhEcqFphGEEIP2eKWcen28cjb
D91+U4w7Mpr4ValbpShy0HOK8PU0cGmQe+dER8phC3gS6iNZjEoz+w2zEajt6F+f
tt7ZZ6D3sV9oygRdUwB5wk3DLi31kDXVCHqcFm3tiTpRHJLewrM5BC9oCZ5CRCCC
NmQc39h0bZc9Tyaw1yi3OQQ+qlu5LobALrxErLntnEkmjqyHCqMT+jgImqnFvZSV
xcfST4kNyM4f62VYa3E3JwvSM6bkGTN2UJgbnJAudZODXzCdJyFF8RMOEMZlvOyi
wssu5h5Wpa+4WBkWnfiuYK7xqUowI9ILiLqVWNWR9JOB3e5xEhkqW6MclcJCPWdf
5Kb3OIroW8Q2KRjtXs5DRFm/LL2+yNHdD00+2yNVp7Okf8XkdzwDdVgk/6e2aQnw
tfph6XzQ2UP06sNW8uFh4/olLk2FIbFfAzd+gpOwEVyTASXlnHFz6/ONS7WAx9IL
HgoUwQNRMG88gUppf5wAzMo7DvtuAjenTuvBgdtL012/8CfM2XxvFa/XPvK0RmKw
idFC/qUQTGJ+shH32BNLxUhUDzyhLPR4G591Wj0IK+56i9FZk5SA6PprYfUu4bMY
D7gUabifKQLckDQmYBjn7DljzbwNrO5L62uf+jgKhZyZ8E/hdileVgeY3t9gdbyt
3XUpQ2UWhirB3a5SeEw5+y7vDjMctIXaB++LKSu9f/cPCLiVVccMm4k5BLfRlEGn
eaG2Jh6xnQSJFqIwJ8+eNjPE4Qc7rKGf18sAQViesi9Z6OrWOqP3dvcsa2ohFKf2
PaXx6OZktFSyrDQLgkmJtQwo+2iDzSrU/ltsbHoEcF8/wsx0Fz07ktgGayKVbhxy
nyEsmLn/yAqYQv1+bRFXJNGvMYsErWOvyMTFKk5n2yU+jd1cEV+/k4rAm8qsDWBl
3d8aoSMT6SFB94eXR221Sc9BYUhxmO1Oqv8AEkxM0/0NmvUwSKQSzAv2f49mx4vy
X7k1zv42pmaR9MhGwot1dW9gB6hNxqwA8aPQ/5ZpsrDQ4fcUAATyjPiBjltrVe6Q
l68Qa/3V7VUzFGNaQ5YW+9ZDdtZsLXQqEq5V6IEHOTrjDyZsKYj7S1DJgG70lxu6
OEXErgE9CVFYr4GUjOrS43jG4UNfEyPSkR/GFBtjWM5O9vlRXRj3Xf4NRb0/9TiY
4eGHK2sFCDj0jm1OWmntO1RCiNlzBYu73TswRD407GlSDfZ1kkUQP7/V4RSQymLd
0GQnT5YwgM5gn4cAaiXOob6c0J3iP/a+z/DyVZ1CIMhqNYyAhNeOxpN6qYgRfwwp
FiU6jaPSPbQs/iC2Lys9ftEe3BsK9ZK03IZSJensBv4GjVNFBirH7ND64/Qto68d
UKBN0+pe/fWrP4kAVsj+xUB2aqybBQjHwOumK3uvTYEdqFWjBfLSe599sOw5DzP5
RUms87avu3k+bQhRUPaKGOj5uQMqfiEUmP8GsNDEOJrDibh08bS6zfg8nsquTik6
f4AOPC3NG7aX1vun0NdSDX6wRIfXVF9Ixcuxmy44xb1hqDCkjW0Zqtpe9kfZF6ki
GUVwlhi5Mncq4Uu1K9WK+yogvzaw6mi6bSMdc4233CIXy7FJW+2Oot4Y/4fSSXnB
qgR050eGXsrpSjS37xbzTPT2Y5KeoQgFi0OBBeQdKVcdRu3adnHm9I6BtQY8Lv9A
Z9e6Lpp/0VruW5BSlhjefySQHf/SPbuK1Tjr/YP67+3Wyome2ZKQBXIgs7il0xXJ
Ren548NWXO77iYYOxRQIyv572D/xYIJbEOLVMSnzHf1dAEPceQWvNqM9cmCQXkpU
6C0RTggWUSiBECDSNrSfWBtFRuFY7qV5136H2Eyg08WlB9o8a9wKcTuY8+HtfVD1
QlxEkoIlP7OaB/Ve9J/4KVgCbCO8fjnZ/zhImpAfc2l+lRDyB2TEwCmYSKRBBO8H
bHQS1ZszMSW9v7gjTISZHde+EFJr575Yl9Q3GtG9pP7Apd9Mx+7fYSkfpAcDBS4D
4dJgOtoWKPsYOiNmc5g4Bc+G0S1pJSig5W1XtOu03ywi54ZZMET8vxGOm2D0XnaK
CjA6G1jRVHj5PW9fb1zzRpL8M6Ug7U0z1fNOz+6Y9otUetbsvtYf3A2INjrhH1O+
OVbMlqN6cxreICWswQhkO7DWIyk26D18caGobpYtwQ+NgchUl7B3TO7hwb9yDDEg
lldVioklJhFa8ttx+UcD91ERlCsx17vGQXIhuyrZtjoq/xrhOOygAhHfyJSZ5mNO
rouHVz6vgzpyppqYVG1q2siDwmxh4p6/PbAw61SB1YH304dSXA483YRwF+Yfqhgv
6gQSxCUVxnXi0gXwyTJcZMlATc+C2ZO6qA6B+Ot9gdLFCBpEfUHpZ8N94IRd0757
adixB4HfXEB27rmHF6feC0R8q6mxdff+bChBrgejL7M/LaSL3pjLFNmxuOh9AvIJ
zCOtYQh41UCcCUnYM2q+vZYAzFvOTQFZhp35iyGhVbJichECLZPcH978u8ay+m9D
CBjoWJTdhwlxNI2X5PquCnR+2iNqTmO4+94RUtMKvrKzafA9cj1o+tz/9pIuuNiM
rxk77CHFTyMppObdpkLituh0ryRU++WWAybuJQ0LxOneMHIURd/pisax54jH5s/o
5edawuxa8TYDzwpbPRjE5dK6etm/59s+FbwGHNNDKy/TkWWE5y8xfmKan8jLQmpj
EStCdNv12Bqds5r0UboIveKQOFOCUMU3PkfReigHuv/kWAJy4SAvlEz6UQy/sQhf
k4BwxaNTFnAbNZUtcAfp/sLtbm4WZ4iVgvcq1nrLXxIchML1uhkiHa63L2KVvYPB
C8LP8AZwtuIckseaDGMIlue2rrFBh4UmqbnZGTmF1BGQky7M6Dyk/d16un3P96a5
BkNtp1lCaqDTGy1om4d2KpiWQxTrcn6RpALZDklldfZfvMgIZixolKEXZWKYegDV
U6LDhij30dXAu4zA+87/Vmb0pJOCot32ScySK2EC6GMBy89qkHxBwn1hzNTj9ciu
Z2gGQxACwP/d3KRegmJxpMG5FzvlpWyVJ1AjNd+Y5/zFgDcGj/JOVCAkb0tKvMvz
99STh/GbVS9JWY0xV2Q8w9HYqMo0C3PPr9NnW/zeWZXn+Hdq6z6kTABR0tumpj2D
QH1r5byrahEza7lQpRrQFagZBcNjY6mQAjdnNhL0Dy0doKk89JZy261QTx3gJgxH
GM26dbJd5c/m7/wLjNjs/uAeA/G6zpG37dnmrKE3DhyZyjQHusvv2IfqAKU5EK/x
roItRaWLyTBHaZ5XlDH6MMwfiv3bOel+FTzmXnLXF5g/conCZIs6koGHG6pye0lF
ruMZl1S1VqGhPbtzKzU5H46UDqSD0UX8b97QTuiGCvLQRlBgzZtiGxuTTmGhAwa5
zUYfNVKM8HJuIHjMOjybPIBZ+djj8nyK2iGoLzzWvyaPIM3DN1Uk2va/XbkFzgzU
IujjLYacgQhKbKbrltkZdC6Tc4UZYx+R6Z4UI3gvANp3efJ4licVWUokELy+udqF
QtiH9dlAoBmE6P+fspaT3vWH0d81T/s+yDON8mFXLZw665fY6OdCOsYV1S8mUWAh
dkVV/SoZxMUX0bKd67ITu4VaNi+QWo9idJzBcAQ4EK6XgPrDLlnTV5kschndgf4D
UE/om0ixJapBB9QmYTSttPizkuFFpctx2NC9Vd7GNrtXuq9ExzmByhnsSVBdHzbA
X/5wsN5M0PgawlhBJx63BF/7/EvrQlRK/64uGX7zQbyRzepJkudwKC9gHQ6eP4AZ
Kpvrt21abGBtOJoCOokogE5CJEB5b9Kh9+NEjN3OwW6CwBdxWbiU2DL6W88HXCS8
Bye9cZI0ORhX1OXQsTnXXID+1wQHTnuyoTdnXLMiIJo/BA0qic67jYWfU/6hSQHF
ziD5MQtar5PXGQpSXKcOuPDgzq3BXsSE48GWA2Lnxk+dGuydnbeN4HhJVMcp9Xhz
/kfTPsY57/UNFrchurOjlt7YUmDzddQ6rYDex0iZHIKAzKFicAeBNSqGZcKKznsw
jVmwWqaaf+ljX/lMA5ORuN5sJHHB9Jz6VL4bvdORx6ZgDLoONmPkBT/6bPPhCoNk
sN5KnrlYXq1eOdwioB4Tq8icXdC1FU2IJITuvmMjhXXDnkAKNkqDSWZ/d1zjQLDn
KFi7kBN7FqUOPLPsA+4iyKzUOyEOQrI6f06btM3WhcFOC1/WamVkjQxMrqShWHIY
qC7xmtq0ApMVJe4Z/gtABntAxpn8nyn3qhxjjHouxgml3iS+GyAAjHDw+VUcdq8S
K3WzLod04OmPJrMzZsGMcMtdpPo8iKTSRnMi7XC7nWLkCQgCxR9RHegsl0D4CuO1
xcYGlAzS8djUL+FNj0EgGqAoyfuULW9quSyCnIVveGhqOohhI9F0HPZoUuWqULck
ID/A5WQTaTwAVB70jXaDL9PnxCr9GNIja1Y+UvAomV3f/XOVheYfXe5D4Ad6JCb7
aSA7V2r1DOG4Tf1UHUGuWTwjybDvFI9ShszjwCPti4Z8wO/+H+eAJlPHurZcHJuf
GWWCS5riMYq2K7IPBRxZmOMY51AKLWv+EST8ltw1IX+5wln3+bNGOXCLnMJg+sMW
hEffyT/URMB87nTU+S/Jlqw+lfDyusGLPw2HlrrhFIsrAO99BdL3D2GnJeFhukbY
EDUOiUtIp78Qu5nTiq4RiYHZo4ijAKpbPnr7/A9kmMx+fogUuzokSnbE+/gADNcr
QNogXaB00twgjemTqRZo06OBP2zWIqyL3RR5Vnvfk73YYhVQe1Dg4gWbNLENRe8F
4Tv1Xvq6odhnUm4E1VOQeF2sMCi+26VnyCYpJIZlFxQY8rn1JCB0G83R0jhx0bKO
8rZNEI6fsWM15i9HhSNDdmFXnwd6XZeg1Ns8DTBox0e1kLhLmAIlFcGnwaASWNEO
aVJTfkssia583yomkTTM2rINlzWsyz//FbyZn9RwT4bfIAnyGWTVeaVhDUdPPOt+
zKNn8r0wqfhJF8y6t8ln3abrCRVHOj1/FawLxw+ADS1QGOxNIu+rXoLhay7Ho7eQ
vHH9p5XDOPLuDXQXY3f2sXLRqkPdWuvvmgFoM7LJwJtK/zN+IiOPEJgpgLFLZnrD
/wIkwrlNCtUtJfbUiwzk3KTPfaO7WvNsHCHPRzXlVCdtg6EQKxmMf2b4+R+6xdcH
UwAy1TUHNTe91AGVBnfn+33f0NA6HiD/6bOAJhXVJ4iSVBWuF2m0RVDn/JixhQlf
KQK3ZD0lAWj7yd9nGl0Yn1/hwxAPb6QSGFwo7pOOLI5oLgo9BnOH7LuuNdL8hwhV
kzkOP7rK1b6nwJ+KlOrNtdTlmMFlRbyxFhkPdudd14yYtXMGSc6H0iQqIrlIySOH
p0Sn+DSVhX3PwMiwywghi25n/fQkNxgYJa2DCUiZwvBwvQIkGW4wakaqHkRFmeHy
HWp3HCxyurjzjL5dgqVH9xIiHnTl5tupAHZBwcYi+MI+p2f+JIVYuCIHv7x5IHlR
C3k5cQkSj+IEKLCyze306SmFnZtwkwCKq5pQpIbRkC/2gT9pDcpdIsCI6f5x0gUr
kcOqvFieDB37p5Bu3ulRC/wxryyzEDIJ5m3cefAfbvJ6LzoYQ+K3ndTTIgcY2hit
CJt3coW2wGcynO16hf3R1gvh9gAj9bLY1QQHEUcBsDiGf+bmVCCC/XqxjUUBY+GJ
4ugo7dMpkOGxnf6udGnwU94Hd6Go6ztZAnU1DIVFg2TFAqBUrSaI4mWS9Z7MubWf
4ouXsHqXHipdaN08Qmzf6+/b+5VPnmv0wsQDbjadX0RtulcsyyIgrAacbalEoLFk
waOoeE48BOJ+NNNjIalq7+KiAqv3rBO2qgcAdPiHSqLvl/T8ov1TCqTIn6icg10g
9wtnWhxpAhDxgH19eNza1L9Lq/eEOPSVRQDEEEYsWH2HUu50NEfFYIMvlBBLktEt
2cSYwOl3yXSfA4z9Yp9WYfX5NwwR/k2CFpIZpxY/gxBeiQLu9ECoKYuYAT1eeoXZ
lqit7KNl33tyiBANPuxAdsj+WaaD8hw++VzG8mVnB1tGiJcCU9BzSTN3wImU4qdG
5eyxBgE5WWqRc5G+Z12Dd0t/OjgcfUn50pZZYF1JIPtXXmC6Dh59LHpviR6nqRmP
p5NSonWwpfwN7PDECTxwcwOx3yHomkeJu1Hk5ieVhqqmKSY23qXb38Yd91WfU9D7
9lKjLd8OW+7/lEgVY29Acg00WbneohpQX1WiHaJQMsAywqBTjPxTGIYuAX4MQ7St
GNkP/tr860BEPqPW0wl5L4kfHIiODBBSveTfuKUj5UqV4VvETTRFxYBAufwbvUUQ
1GijpGN/QO6RKBNDqCQhqljt3tBVeP6btNLKGaUOmnjZRRkrLi/UQK7wgE0yKE/X
T39XqFjQ59qIeCwXg1tDy2gItdlZwg/cXg7ZnvUclXJwkC7Tbqnf2kCVRqqApTtF
szZ63YkAJAHHQt1UgEXVXsSzlWd3tHYM70/n3SaZqnWEEFhFup2W0Faaob+LslQz
GfNAms8Z3i/0dUQRULcj+h2rAp2/mVjTy8+I+eLGXF+t4kBO1AwTGlzCrWlUKKAa
bb5eDK5wHyfhH4hkiYoBojPq76UKHJ3jXLKAYmEw50hqnTgMwjG2C6Vmew9lPjHw
vTroeGWwBGmYuoSRD6A+R/grvhlhxRjbbLZ41WoAXQnCRNKOL5Ed5jgAg2ePp3/N
v4zyxGSJET4fJOSDKyaJwOnnT08reGhLCVex4ClKdNomRVQk5oDtPa/o5yNFZIKC
tTWaMKeLtsa28k8uWQvm9JMhRjcQ64B0H+oqqM1USzOprLsKIPPCyY0pnKiek9Wf
YekEeHlOOeGy+KBTzgY7y3O7xv3xtPF0MGuNhZv1khjI+MSwhjN0k3w3wZhxnZt0
zmCCFoyN34TGz4ByexD2NhpnlO0WJ/R0cQOMTnvSqopEkVDucm6cZv1JkE0aZeN8
XZNbXMb4Tydn4A6YEuDY8XDJE8rflKHbx7c1TcBBWqUZMMo73FyUXhW78pQpzyej
8mSltc/jOZS1l/pJFwpEzvo66SyOSVYlZyOSuBm0GFxVd4/O7h97YGyfRKL1NmZZ
Pi+3MLHY3ibJT6FoTjDDnvkhbO+Ndikhn3sEO2QPB+OKLoLFAc5JY3GinL/3pF0C
NZ9+Lp5SuVn55xQ4UtC6Vq8PUlocR/cQPUY3Hd5ii08STJ0HTCMbP0x43ad7G5aQ
Ere1wa9TC6Ehx1Ux/pV6oAD014I9PjATJKHhjND7PRObM1ggQ5GMC+TaPtRfadAf
AYmt/KCfg0PheYtnf1w3iM1bcnG1gfCrsnMNN/Zojxbo+Wg4lMqRVKbofVfk1XCI
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
UDTLb/afCtDZ/Q9vf06UgwV+K4+p3sgRPZp4WdDVZGB2fMa6shpqC3cENkHo0tZ3bFgXLUliWq62
6OJwpkJykDZnYZjE/PPgo8c7lOxvtC0s4vAO1z0wGRrx3i4L+i3Hli0SVrssyDvKHvD7lHCm5sds
xSCwSrjo9jHofOo62TICqGt5qLiXBDhodOv94tET/+t0C+uOjjjGLo1d1nE9ax35boGlX6X282QH
j1yD+OL4oaIOBOPqoKm7CXKVRYyyy0ZQW7kWSgSxm3/kgXNKN7oXDxyC/Eas5Ey6gEVSwfKzB4OD
imm9TJNjKSHZ5ETtEwPcsxoVUUMsLCVXHiLm4g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8592)
sQKqjvq2rp42kutrChNXMBl2YxoFya/o6KrrPPQOt0ZiNip6QaFLTkHJTlGXnDUxFlRfJPG2oog5
p7vmbKxR1D1OVQUcUz72NHWBRs2n8sUbbOlEyjb7exZoM329vOW8tqxGO+N944fbHxWJZhgAYqKi
BjFBw+m7Op3/PHszAZPt+Jjf1YStO4/+aDs7GGXHeqk0s2QxM12NflxRsIHWnNdyu6QA6ZFmgCzG
F3D9ZtTYJ4JCs188z/jeECpyCJ1jTNMbMadJqyn0j6cOKtUlOFICtENTfmhS4jRo/VKsZzqz1n2S
Tdhk6rh9tKF6PQW8KBOPvQah9mklSd5QsGobRqX4V2VLZ4elbi4fIJdQIonCeO0l+aCF7ZhHhG/D
NPMGB190VmtD45m5Pb3n2hlxxatyx2AAwU/eoLhoGQeWCzAZMmSDMY9n5Ju7qTpqEffQkO3Pc6vp
Wo7PrpxYOAd65nqPP8ofYp+1qFWBsDprr2w5AK5WVBdUU11Dwh4xdjTJ8SKw86cZKOdwkIrEPqmT
fMKp9XAqGlJAl7zW6ieKzo84J8b04EcYzDMCUCs4xtH2g6NZGhcanYb1POUBu9J98KxGxqUkmX7O
Mz6+wYrhWDciXvhAkmb1Zm3pnEwhJRAtGrmTVxRH1mrFeeMssJ4FM5Px3UKKW62DapRIY97mllR1
k4gi05ufn2C0bvJukeULQGVSQUPSpSW91xvLLxJiMRkp0lQRRpB1jLMtN2W0Lup2q65aI/WTFlLQ
Sb6SC9gY0uay60zf/ntaPJSvI1+wExePqAzbd1ztcDRyNw37i0h8Cco8ubejh0sVVA5opuZVnUEU
VSwnem7cFSebB4QrFC1rJq2ixPuoNLCJhrHduGm5Cebbjd6BBFihruFMKmG1bzMzBSjpKM7DR48Q
xNL0ZX3m3B2gZjbRRJjcCdMs1O/kKvfWX8TLJFK29zGuvCdGsRFw5xZoT2suFHuao7/fQSzYBIyF
eyM5nQc5hlF8svf4UDyqEVnxs7Pl6GoKjRKeU8UAlaMOGVt4Z57xLMkOlCoihPTTxrWlfcVZFztf
qL6ARTNTRMQtY8GagCqFESaqQd8it0hnHPPZHXnFPHM8nNLqsDYrt0D/RTBM0R8cQ/5MbV/mUE0t
L24x9+vlFgkvmUZ8TNdWh++1gjdZbZq7VgeG7mAYuX6Gfx4eLOqa53hqX6vukEOoV8yZeI5sgLO5
MfEDYfWh2u9h6KIAdlokr4ocWWMsecrtP5nhvhX5NCrRlKb46R4dAJYQy10U/3JjpPu89lfeaX3G
hbUEDkkfik+ZSp2vntHGB3pq2wEWFO/6IGkGd8IOi0tN19klVLZyqoZdiWavcorfmFx5Csg5XU7r
34EEP4/RNYI6wSBkNtZkzDS7MXS7XBRFtXCHUdAddtMPBh8XOfCrSFYVfPD8ct4gQvkyhrYUAl6Z
yMjO4n0hqr5pO+6wqFzG5GnDyvveeCRXTSeulN2q+ENBr66bohL2R72qdlLf5GiA4JuYn+H4cFxg
cZDGNT+yI2QH7Txtzc+ztKt2F1z3ZcqcnNgjbl8XP1w3BeqqD3Mq3Ee+bobKJR8+TO2bj/1od2Ff
c/9ny+/DPw7eBx22PDwFr2ErvrJhIXFC11XMeIpfxI6UaZHEy4rt2Wr9zL3XC5TNDwyNnXS/bnQA
oB5GIRp7v8qyDm0ODdSyvyobla+HqD0smgu5N7IIxGte2yNPaTrn6iwZYq1FmYY/r2etukB9CAqC
mpIkKoSBaNf/3LBKnzs5kj/SaG9Kh3KGVgH1iRo79B74p/GacBzJs+H0uv2EoSGKSmIdVoy0FZIT
qJ5Z2TMYfSLqkJ1BGfayZJJiOeQiEzyy44Uiegtp8cNW5XXkdPQ+p1zyFXgsu9izS3WrgTEHT9b4
pgbCC42d5fjTIphU0buA5HznVpLT6yHoRKvM5J3EtqlHX2s6QtZTWiJ784drBufLgi/KbbUfhcmq
aRXQA8+WsBn15R0DlndW7XCvBhK1dH0SO+/8vDHA3xQHPeVzvOgUTY84U9pBNWH9xkwRoU1dgfX3
uDNmYWjwhrtJ+8fLaxNxB+3AIAVJWWcOpNCgCw3cknNK5/dNCE087BFZVdxCaObedpa2vIwSdL8i
YB09+kRcK+H6H/knlxYx6hTDf38IYG/U1Sf14GRz8DIJ3myVSb1gIiFjZvVaacUox1gY2n73QCBi
djPnTbFlUYWZo+STQp6WSFwnbEbfyu3Jimcao/Kqo+n4M75vKlA8WRKj4AkoXY6ojKQ2Oyy94/DX
I7O4JccjYsvB1/s2GVDkZGZfPrEwbuDmtZqhl22hKxYGd5oDtMYto5pBnqES8yNd9hh+SJjVUUSm
lMIIA7WNnvJ8Y2He7CrvjGQCjoJTyIGIh0ZwAAgsxPDjx7lDnf3JS3PzVFlU49noPy+ABVybynWS
A7wBpdJb4ngGdPF5xrp6i2ysJ9epVbeKbhm3WORFZ4lOE26kD0TaxV7XWs6FO6Ip5tTs9J0ORHcA
Nt3I7ANdnh5F/2WoUqHozccIvVsSnDCcXG6+0YTWIOPnMHFlyImiUVwwfRlpESAhTJh7guw8vgR0
T0dahtLaJaoYWfer5kQX4LjMxnayMNq5E44T29vAuqAPlgHryqi4wLq3OE3VKDnVt+VcXd/2sO4r
pd8B14E6OSOIaaltXnrku2VSnKp7kVzYG41HzN7KWut2HIddYNYAI2FEYqI2Os4cLFR+PWv/zxFn
3ZyerTYIIn8D5RGI56k9tSJNcO7pXPFlHNwwr87iJK6wCeiluesHOupdNdbUbaH8D4z95fvPSEQq
5tlD7RLnEwAsXIY3L9B0ECt185SyZfMUu+94XLAlRGuVINt4UT2QpdfQwtVgdeFwFjidzTgvhzyi
0tqlxD1mxXLluog4LYznqmddImsytorS1I5NxGaPrgxh2FVTwytGN2il7GY2BQPwZrCeo+J6mCuE
IoK6+ocnRiZ7BH5pfGRl3VLojeMa9AY6nVUml1omW2f0/NZlzW7RPiQPpdKTFuOvcjKmVVikEg4D
MIDPVraeNLvGjsMmm6+VnbocR8WLmqf7x3UhimxrmUf0/YEFJoNXMsjit7NGCKGj8T7EenT5amBj
5FlGn5jvq+kwN6SXgvMw8gqroDRFRFaUz6jtnh8oUI/MWqNTQ/nq/94Yszob97TZWf+cc1A63MUa
Y+ukZKrrD679LAIEP2WbcnD+hexXPlNQZxXrh5sycJgkhK3i6lR4onhfGvGMhDtAsO4iDhc1lCSr
/9zcIhpvwAJjXXQYnwG+iAs2EhbiGJ1ZkV1doHCCltg/0fBZbvqA1HhXBFH+b7drB2g/lhZg+dqO
GpAypop63b3oE8cngtNGvM05jfMg2Yai9rCFHPQh1XbPEe61yrGxuFA9CHPRiFUBlpO3JSmcqT35
NOql2zLgM0v8p4GLOM6CtHuvhRQgH7hb8dtMCLn3zGHCdE/x+kKBDkrlyOwRgXyo6UP4sX8/RulO
S2kdqzzmQvNZ2hQ1B8lUS5wK5347wzfEli1+d/Uos31qsGGNylOO3/xHLfWA6IC3EEYK671mRhjb
YYA0plsVa9MHLpybPMmw96TIy0zQkcsoUblwoRdJqBxeI1d8GKi2k0nB8k+5ovc11Mxo9+d8+zdF
twXZavz9SteA5+W6HDLMTmOGeY/I+WlEdTklzZzag1DjtfBLbXhXDfiZVrFbsKdaDchE+r7+xNyD
tKz8mIRcDWf4B0CUfYJSRb5drvhDa0OHoALLqpvQC9DUwA/HLLnuD4OHNO8e6i3IK3E5tXBHqjw/
SdLz/HFGUEZRpi+flyVs62V8V0Q1naBNtszEPYHrSWd9ptumAOi/379ZsHEVFR0rcaw1hlbER8kw
aknxR1So5lH8zGeq6HZ+IQacxiP5WwQ5QpuZ65kmB3YcevczB1jIQoGNPPgjlFq/yU34k2K2Yd7p
/f25+f6udHmtabZz19NaazUuidFKPOmxpw+eDs3Ub8EtctMZPhJEwFNRUzh4XASEj8VcEPn08SVn
9bVlfvg1tj1ZGW1ZP04KJcXQ0dRUapWHd2dGez9SywaasGYrPxNDqTZwArVLqcxCs7S14SPJQTiT
TrQ1UUBgzbiVoTI5ca2MBrzeZBwVXY+4NM38Kkruvq7ZJiJ4aDDhCeDCPcfOwdCa1o4VCMt5IOlW
xaSWxp+2OXOhffdr/uvRHFbJ7+E1vsYbHs7vIgDTUQm/bss0gXbA6CTlY7lrTnEdQ+dvymtryJRu
hf0w67AIzRw1B428UKUASVq7RIGSAS5P1vvPJzD0j+7M5JVF//I4LXiSbcypIpjb88JzuxeHDOiu
iLPPsUu63b5QxnwJG0PbR3gLrxPgdRjl5wzwDTJzn9BRHhSlsEA+CGOSVPCDpSA7GfJhP7YIG+Nh
EAvPnKZiHFj1rHp0Lt17VRFTNyyyb7cFjn2L2UoyIY2l2EyNNyYzBSyzzvqArIsw5831KQrZ4/tX
nYe2H5l/X65VPkD9VQNpVozcSs9Ml6I01V2z1NtH9wccbezCU0n44/50gTRtC4UJQaghnhBZn6ag
mr9AcGqg6yikomSd6QSE4oOqmtnDGATLjYikD4vPlaCRQmhfpDynlr4XVOfl+lnWPhrW7JlJU1Zo
5fDRn/mWDo7gCVCFR7eRPNiRL9rhD9cKrj1Xd0eE5qjZ2t7p+L4Rswffeb6Zf2kPoHrW/ImlBkuz
OgHOJfseG4nGP5QVRmV3mnFbGPade1MPpaf9IKA60kL//ojE2X+R4xvOr27YBaTe2l3T1LwKJFgO
dEo40NL2Rn6OfKNwtwHVZtpJb2PUbRqg67gj20qel9Hp9FXBTfFKfy2EGJIYrpm26pD9aNyCWI8P
PiVvJs/Pn0ZoGtsNYrMr9eUgaoghpZs0dEVRXs99H5bRa71PiGaPcgBp92YjK4VvryT414GZaeGk
Mth5rq8xsioCvigFa1hJyV7BQAYhhavZijX3RUz+GPVxUa/tP8r2En6tMEU7vqDL02rt1EZW4uKE
8Lgnap2N5UrWEiwUrStvFKkKrjYJG+cJLEIKBaxta6Vj6gD9AHerP1mG7957SqobsCMFrVcMNnG8
/A9Z7Ev3S64ZFOzV+DaYCCLnVx9/1GfhZBEkxpMZnAeoOwDNTKAHjTJt9+tBLsEKc6X/H7WL/goI
NhirHCP0VQ+OPgKjUr/eg6D9T4Ps0p7aMrjctWmBUmN7NfVJETloEhnfESJzfCsnR8fP5AR0i7Sf
AJfr7qqPKCS8WNWy4PA1cxamtZP3vUnF7JZWR7/pBzUAwoCRqL1pdjTWL+X7XgGANgS3ZjCV2MEt
E2abNzIt0d4CJ7EcgCGOKowv0LZMtZH/MbTaBs+pe9JExCTPPhrkGMUJzDNpwAOVVmpNV2D/gfP+
yX8kBMjCXmWprlHZaITf4b7OFp4oiEPqcAUxDiAB8QsnmeMfbHAdTTtQor1P1e7Bu6y2IfO0v2E5
4G7AfMjHwKbPDOupegvTNujlK08DA/1SUP2x24hqQkB2tZ6QeFRWeTIA+nPHBGCZAJ/ExjvQYO/E
/7MlQxwo6xieyI9v6ipmKSTc8oUhKvD/qHnDnaScePG82+np7l6ESmtITbyZUBFJYbb7nFYiTv8y
vIDnZb9pdyZWnGoOSACPAv70muUwBQs9NOl2jor0kNtOe56SwnJWKXGlzvOIblxOU/dx7B6drnz9
IiSVVlalsVG6kGt9sIegdNUxH+qWjeRUTXfI4hXOhBUBvWJqOHltaWBMb/PNF1ILCKJ61+fbCcfZ
zO1nyzgbqtcHrlsVgrQwHnxhs2mjZ1ZpXk4FAiJAmihZTyU++S5XAEix/UkjSfFjn8R2tG/dZaPr
IyXUc0JIOk0PnFAL66pmBbj2pCxsNwt8n3ZmSba7DjvRPyeTeOupCFiSCp22N7Km0+F7j06Rd2FZ
VOgGcCoGMjWJf7cdnGfR/cNOY1f2H1pcRv7Lp2txaqUQxy9ArDsOAqFzTFz6WfEmc8fxspwOLFUO
Z/FNOoD50Gc9dGpmk2a4Yf8da8iSEBC81YYqIX0O9CDoLQwDoD3uMGKMqm6NC5lT9logG33b5Tt5
p+PpnpyJ1IUcFwimpYtDxbZPxpM5fjNfAJ5XwJQC9UQNSDEIpFPtCqA1EDwmRTKnxPF8N6rPq8Li
ad/tnIusiZTiwf0vx7Xmmba8uETV4DCnRKClKHN6XMuuo4RLtfzYYl3ZQeXbGPgqYkVA+/LFVilL
zQW/++aWKJ3bEUWJ9sVzJoyJ77nDHyGU/wSIUGHnRkNGFlZ7yEehFcIvyzAF9Gv3ZnXv0ZqnpexA
61JXi3BJHtJgKWBLpMhiwqpx156YK3zzBrHhAjVE8DwUT8Ax2LgF89GKrwC5m1+6Z6NUKrMAN9YG
ZxymbiUfPUMa8DJ+43sshfVpAf8qePQHPVdWs0zNacl4Yxfowkwy7K2niWdZ2kqZtyxQfZJrdMi5
oRdwvkjWlRATMwi8Fyu+TUWMCbkdgQypHjYQIcIrD3LMd5XpthgcdNY/Cxa8azRgG3LQyRiKv2Rs
yPNg5J53bsTGT1S4TzA3F2yuTYxR+Q/NwRstMUNUXqsGAixJjuAFsnhaak53Nj090PdGDFEeJq0X
q3D7dODHq6pKld6owGiAgVpsnq+7ePBODHslHRF9ZszEu4RmlhEz+MC45i2klxo2P82KFY6wkJpx
I8de1FZHd39Z16XBPh/NpUWaAAso2pMh05pnD2yMQh36o/th1AeaE4MUMYyRFFpz7Q8ouzNE2J/x
IO59353pcqMm0dhHVSw/01nryCsr27vF1wjDxoKl2At1DvH4Eqld7+QPYc7W/mHr669JmC0PsBD3
fAQnyUk/aB+USgIc86ss9fUmLW+b2BuOJonsCJbMKgwlOKc/6R/oL8boM7/ZchbCAdfH/H1gitOS
LGtgNX/06Y9h9jMk3NYoRRxjRp2T6z5TwFY7tXq0XZ9pZvebZdip0mtE++5dSxprk2PVD0cFhgsG
xeJP6U9ITqY4Qn8DsDZcoDVSzk0gxTERgUB5557dpQt4UA5FxHMOZIiP1oB0K7MhFy5ymhhgZ9v3
XamPYXs98LnAn7CLpzktcFX2j9vX74H29CjEMH9pPzY7oLMcgc3RMPN+fu3NC7CFLZlWNrLmx7V2
iP5BNceG+QgbL/AeKCWaTFcba6vMprFpRJs4ubWexMLB1uboJ5N6EISDLxX0bIinbRqBy4R+6Jsz
usEDmxHGUup4iqzY2bsqBuAk+SYENmFhf9b7aFd1H51qwyWgC5juPJO4JFFaqiFTk5mQk6OBrliw
myiDwIJwHAsmDD3WpmOZam3gt1w6YPHVZ7mq3qckg22VXWyfdBCp+psh6ZWIW25NahoC1VBy7QaX
Hr3dYfEMJryYNK8LP1yD7aNMrqMYrR+pmfC0F/fsx7FVeSctpBuWjQFSp0Ml+NwjqyOiaRyO3h9i
VgRIChkQ8mtyObM9lcBc447OC5/0gka+riBucgxQY1VC1Q0qpjW3HwoUMRTUQUnKipJpqdvalGv4
Lehjk1BEF3Q9x0TjpBjkt4pp5HKc2HlYl6I0xOiAOY8h69A+ZlmfNlkatn+O3Gtdwh532gd7AoIz
Y0huS1jZIcUIL1QdUkqSs1ylxSHa9K32sXR9hHmJm6yL8RRoBqg3QhmLSlyiEJktiYCQ6fS2t3vm
N4YNyTyOdRVab5Nk8y9QkxmPWqhu2LW+dhEKdx90LASGgtuwfI6Cvr4xyChyMQrEdC3UdemxSUwy
4ziQucPid4TTY5LmfgOg2dz0zuo9qBKisCmyGRVp8/A/vZWAiz9AewpSgzSnJzRF5nfis7XxWaOR
cZnPJFyNmDRo/RG9U/WDqr8unfP3FD5QQstZ9H4WsPKwQxqV3L6ZGcIA2L5bBvLLpZ57a02lqpXO
G9nfHCddht7dB9goes+Dak9Vpt6xPl8+q/sXfjdhhDmTL9agVey3Ezr0y9PaeP9I1jYYyax+Grwf
KcwW8lu+cYCtxTknDrQfyACvavocAYYQGsw+rLWOCk1IQ7slthAS+7GDPie39aglEt5Fovva6sav
Xhk3GQU+8mHCzy+fC1wVxcIIK1SGXghONDnxfrVkhzhA9GP4kawGkHKJDNUX765/PClS6/t6DwV7
cdo8bETv4wvff9NC6e+dGNtVTj4kjE+5Zu2hQ8OUuF7yYQ3nfx0BaPKb8PvsT3VZmgzfY3hX74Hg
sDtTqSu14JRcqNXrB7l9P1m+VCkoU080OnQ+dwRHIYU9gSmnXhz15dE/vJ2KvFnbfyN8FMJ/fs43
ANEcGBJ9HxjISf7bdsfc2g0sSeJmFU+fUi5W6sOEz+MxN58O1IZfES+oVLez9aS6rrddCtefbzrl
hlIt4el9u4JOyGf3ND/b8tts00ZZvvSbgLMYOKDTGGB2qiJl3/AmgqXc/h88L3U3Z0FJ1sUhwsEw
3xZCDW9mIYffjSLgrmLrIkW65sO06vlehrF4b7DRhXp2+62X0XZfBjb+VsA8eS7qnREy05v6jqBi
KgQ4r4pbMGsgqkeFtMLKP8H8h1UREgaajFclVbvyzDbv0rV5hikni5biWPhRwMg2mjt+BOFOvtO0
MMuvV7gIpziyK3c3dR7TaVV/nafV9e/qKg9nvolcqeaG0rkaoWAldCL8VX540evGMxeiBYuMdCxs
s8wuLJmRPnm1XkZatxPyf0bpuOVGN7TSE/zf0wRhf4EUaYlqbtR79pI2Jo3grMiBvUxfJN/vDRPv
Xg2VPmlMHRmlqqzLVKEpeDs4OyNNrFaqquDxyqr0rpv0P8fmWVitRh7ZYUP0niLlRr2PZs0s2xqB
TJ2x9F/jDoqhTETtU2HHTamUpemNdJsbN6xYiwKyiF75hT5a6WefURJpBa5FJ332Xw4klI4YUgRe
BLAugD4haQjg5TeFz8EHVDZuXNxCu33EEprJEPKCu2/OSeSmWrA0YMwmQwk7SVHuuBVhYL+hLpKB
U4ob+v1CqmphYiqVVpaVU+Zq04XxNZ+1uG9l4UNwc7ZHElNng2If0a4cF7LBgRt8sV+BHGwu/KG3
y6T0ey3bUog6OaqcmHB9nogO7g0FwSQZ7JMMf4mXTxAfFmPjoedK4w/IQhi2+A13VOngbrpldpFa
VHZlWFEl/+7CXJ2NE5e/waomhanzwnDtEQT8mKvLy+J+OqXeCKaknzRgf16BhlAuyDmG9/reIvFl
cXP2Bw7I3um/eNNuHFOff+3Q/x4ofCkCGC/daqxCT1dnwa92ZHm7t6SYNEOoW8Ht/lRFCmquTfoI
Tbr2LSI7A9CNfhh3N8STOBF6OQVwuy1cAoFGJpY9XgfUo3Sc6P+xRq0OcUusbE1/+RC+jBcif5pQ
9ZWDUCxQODOHKfp808/sb8W96TNGYhLgdCc0ujviCV72n3Fis/MP0nbg7VhFQT7sFOj4n+/hAHYQ
53x9fyjMBWeQf4vcdz7BrESlbrN9cpsSJxv0xQjVLslRQR8yXWf5rYtusMwVORdY2Nzbl67u99qM
3keQAWq+L2H07iAEtaJgsAcwQ3yYC/Z8jYgUMtcNtEPQAapsVMp2Hsn32yguM76gU7YCKFqM2Rwz
+0zCup7ow25QMeK0yq6qE+ypJy/BksI8l+SAjb2e4tu4II6XYKbcRa2fIQrjPoCG9hUfSTia393+
7Ae/9lMpQa50Fo/XFjlbpY6UiSLSMX9DSSRUw/UTrYCw9SuL3RoJFOYFtNDkk2H1bzEwqAehTcpS
zJRuGlGd90moQXaMABBr7WuC931MLsYD8F6TvW7S0JWWgjhdz2A/pYXzAAqoLrMAqWrVuSuiJeiW
96aGSFkfyY1f62CTVVAA0hWYlf8RAkFF/0Bm10RQb/o3ucnmFRXZ87AcsQS2sTqHLXND1fgYvugq
HRGM2gC4vXCC2Vhxt2zEz7lM0STXZHiPsHIpCa3HkMBfAd6F/5TNYCgxHbm5c4Urr7ZSsQVuhbfW
27SqfY9W5dtlQIsAfPg7H3Zr1IVScpk4CeRjs1IdoNpEMZLNYh/38ONLSv0HsT/OC6zpGJPnkIRi
Y8d4cdqPBnSEEYRlVOVByl8CiqOAXGF1QtZZwM7Hk2bUch3NcsVAVWr6dg8XOHXrFsasz8ys8Mcy
30kVBR332IzYTRhCyNEjzW5rBz2nJ5wUdeUtQlRc9l4EazdlgA3SebKUj/QOOrF5tSCzK3uYE9Rl
poHQuht0lcnBCmmwuQ2jKk0q9Qh790RN3IFdNL86ozi8dmsfnUWYIR2Q561Vt/38jKurczNULZf3
Qh2zOvZ7nMTZAABFLH6OjFLqCdTWm3rNBEkTO6smd0en1ffpmx2qPeDnLSTIVrlB2E0ckwZmDB9W
IgDAQdyUaKzckHkMDDccapJjDzrtwFVtnAC0f2wtkY1Y42/fP2+OZDavgpR+85aboD8c/HCSJfcF
kt890vw2DrurmTR+jb7i1gx4LaGdgroHI7dlH5AxCMiW3Arv0hTFecs8jD3ZwrtklRM5ATtQC7l8
IAB54Of2OtINvkluPtJzJiaKRQjQ7uX388my0o6GigBB0CvzrC++UFRrjqNp2wa5VBZxtEb/Obo+
MyRdaWNgWMOc7bJXYhcxGUGdEBs78RsGe7sVfcJ1NueSHK+ly5DgFJkELRYp60JiaNIOBiVZKB5a
PKPShi6Xp3eQwRI+I3LUDCS9UaT2v2V4e+rmMN+GGNAeU+b/I3gDoQSJah4bdncsRvoB78jYOIH7
/R2p7gAFQqwQg61u44OihWLuO4vbbHA50MxfPOebiRk/caNaO+75zPLCSeWEs3yzgiaSvIAcLqc1
RUIofclEiHe81K+a4nIsghIsriQwiC13ZREwwXMPA44AHxNednxvr2WGvP8b0Lhew58jacJySN6O
LVRJ6NyjX+LtpW4B/nWYQPsR8lM90hEI9W5j9GdYjEbdHaNoNAYO7XOUVIKMb4OsxkS+Lw+jpGt4
cp7xXMeJQE+OD/iPLOPefdMPBjRi1sEHI/wXXg8o6eSa8Hi0++8Q6EZ/wTd2UUAhQHvs17eJdM+0
JJ1/64nj9ZucCIUU5JxWJXTGhcRCi1Gk33jbjSAAl77C+p6oPm5pKvz5r0pMwy1P+d3WklrfQdEm
DyPYoS5F7W3eXGifTlEpd6GTpYfLAn2oK1twhDlLrJhW8xDWu4uADKXNCLzo45Z4Y3oGvfrFfFjA
hFK4TbKkQhBWxUlB4rOKF8WnxS3L7Pr2zG8kNqo6MH7HthS7LR4Gf5XKdH3mqiYg3rBma7wONDaF
EQqxG9+ZKfa5WFSIR+WzEn4cGKWndQ30A8XFLj3naUUvgxvHmA+v09xJS84t54kOPTUnkB8gVEis
JDWprtQvu5sneVb5hrYW9U+SREZv08nrnz/Eb7BX3ONJTFtzoYim9QXF2uAPxF6Sg69dPsQQWPM6
u4heyRogmUzzsjIdN8YcUJIDt7p/9E57t5reMumHQ6HcbPEBUY6LZ15Q
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
haJyjSogfh2ZXExtG0c0d425MZA13zrmYRW62UoGKo2TuP460g+OpbaF7ZPol6iW
MwDEmdonOEf/g6FJcdO1ce0efXWjv4H/p5pL/wH3EV4kPwB2fwyJVru0CLJy8/TV
5K95Zjx5rLZcFuKXXMwiKqkwKOQKK7xkWCNVIxcNSOv0wT/sOSS3bQ7pHhYjFP7H
0gGeHxYFkMVRAHca9BkmpSbwtZujnlObKW9z8GeLCL04OIg463f8Qw8E+CBu+nxL
JzUygqXkeiFC715/oIIrEvfqbM19h6xsr9IThU1Y0lSna0m9FoceIKDoAhOI5sdb
/oP/HH7wkhBat2FFNAns7A==
//pragma protect end_key_block
//pragma protect digest_block
/VpXxf1kzveG5YEgA/4VqMOv2U8=
//pragma protect end_digest_block
//pragma protect data_block
0csh94YEsx73dDg3cvgiNmbn7sW2RgybvZudNVReu+DS4Wm13YXG8ds5BF1Ynoab
/jjA8/C8fwJv4m3BFUjoj51cyFXpwXqLiZOdRXqSi0o4/S4N5YH5e8f4c4qLbNU0
qS5dUHecTjLS8Kj0tK9q2bcz2c1GEUTCWkQRwux9WJkRuMn7R0zlaTYf3qrgaRV/
k7++zim3LCScP+JgeDYV2c2iH4IH0FyXkCP6kg3Ygy6Ero8SseK0Co1eKTDYjmRF
3z6+ZNssqG+JL95rA2F4DuhrMsmGi6XKZviHoCFA00DUcCLeFYIrChUwry0gFiYx
EicyxAzMe4o19bF8VRgIEttuvWzmGTosHCXBUujwK2/x4sc/H8ifhCtUZxruUhzR
l23UvmwP8C0gXq87ENkM5GEJiKJFv92ins3MJdF7CrtTC3Rz1eLgNe15oy9/pvVM
010rNJ3bbZ/Khuc0wPx/ZMKZAKV8sx9LSN63WXWVv8JlfPMyWFikb8c3aQDAnkMe
VNfia0ywjQexaQqiEwylHD0UeBacLQCtE3Q5wG9Y0Zfkk8Csiny5UJdf/VYeNImR
2ThHmjwn3qx8ElCycX95eVAg/WABt44iGMElBrNUVdMEl4AYkzA1DbR7gd4lKNtz
tplDROFATgaLxZhTB+c9nJhqi+t6UpOss34ygYJKCubNyhFIU6dI2L/1x4mBhVRM
mdu2LqRTiVZ6fR8Rw1Q87b3U4mGWWDbw4AbNQgHx1Z9de8gmaFdx3HQEdl23Dc9z
b9RyMyrx7zIh/4UfNZb2I0B/j4k2Jdv84SQZrbeuIw4mQRmNzasrY5KsoGRYW2Ih
iBhSh6Oew2j78wkdHfeK7InkxYtBqxSaRKFAmQXB4QKvZ/GqJ7//JS4K7t0a/CxT
pg6pPT83O7dXx0RIX5OYYZysLfDqt3cQHMDB5BMOOp0lulFO3W3Fm+8E4uI2TtYp
02lynl7mkDRbwvEFOmpLx0K0zJtHa+SR4PuC+ZwilOhob5mH8D1AA1Z89MrlXXPy
2Pdcq41vbHlRYunKRV9Y6RFsq5NH0L9jXujmKAy4nwLABhyi3uLpjFEhEPOGiKOa
cAhQZ2SlC2xZ1mEMqwhVNVTefPjGTj9Ste/gXgmXKix+sTs4rinUf+AWKFJLkAGb
GF3eJc4XZVHdDOrmNe1c5f4BXa20jbUyCltmFjg3SsGcqSspFk/UYGcnI4ZDloMM
RBbwJX53abG6C5BK71+qh1BkP/PMQ+aWh0L6xbjjJoP/QVq7675Q6eeEXRoIUNmG
x/D0WHfqfbFsdbF71p5cfPvdiPnwX9kVzuq3fQAfVMrRRG+qIbmOM1tvBiBRxjKM
n9s7Czdf75CvAYFEJnOlgOwfWc8PSQGiYF2xuxbnHcD5HXpqgJX4QOLBTtkvHvpU
aIVFezRHkr8qTkMZYcJAOD80vtRWFN7MSp3vs88Nrwk+ZHIRO3nLBua1l0KKvvlU
u93v4EBzlImmUHddLa7Aw/w+BmUIuVq7rihXH06T9p3dXvubScLspW0+Ype12QC6
DL85V0Urrl8hLwjndtitD5I38xBmBfGieRAaoJ18+fehpLybuMx3UVccgIqe1/La
88DR2JRVUUoLjCTqdPMG06/YPOQe4ARWvh93WPDrBE3Geno1XwqFeH1F3zU8xLUp
1PpnCPvpHMTm/aFdaPzyO0obyGmZE4vSxp7PZFIxmsxvNFoaomWqbifhm/3tojpL
zMPgb0PAnJrJ3wvcbCMwzZsOXjhD7d+DxOJs9A/yTF88Wb4A7GODz7HB/famqHiz
3WqmUg4vJTPxLlZj4XNG6nFrr1GToen/DcvSjs4CSMpEPd6j26PUHti3KvVhH+i1
kuQvDLawwHJVyZoF5BumjvlVXV5tCUeggxdb59wKTghC+4EZKcjo9awmJI1FO3Wt
ha20+jU6T1T/5BwWUPZVFAW06yLvDWW6AIX0WXSAm839ndZifdSNKGocELOj3asf
0TP1lrjZl5akp8MEEus8MF6ZpB2o4KCiG7VA9d5KYn/h5R8GiN+9T/m6YD/24TU2
0ZDDz4CucrhHWBzHTkZxmi6kwC5Vk39SYBJZgFo0N5L100qtW7hcIgGfIIh/tf0p
GntgnbUucP9u2HeaOW4+DtjyCVzF4wNYK9Y9HxupdxAxBhvbf1wqAb0Gr4hD6n23
F+UppDMia0uJ7WvU9Y05f3XECr7lNiF5XBpVgsblmL2KIwEsKnAkyKwuRYTcxgxo
MdjckAVIZfV9oljqBt5mS4wwtwgngDbkHnSm0GDpSuO5IymAN6SUJ4UjWJ8q9Smh
MGgUkgRU6F9uJ0tA1dbXHejU+F77Psd8Mm7y+WleqGGN9+eeK9P0GqY2OBxnGq0p
QXQduvysoXC0DIdT+577ddERmYtbXMqcxxKWZjU1FZ3ZpJ3vMGxfgnSNl/ryUNkR
cwA1uBeCBmpwbV7dfrJwtZ3kq4b0fKozXfC1Q4v5n4ZYfUiijjS6vgLGFZZ4Dc9K
/QH3Vc+BxCyKKRoeYwV4vqCqIbEdRXDrmFNgEYw9Z0fO8rrgD/IelmWICCG1X4mk
mUO5Wi873ahJBgcmeWbN4lF16jwRrYrQ5aU7VxEuxkX+hwXX1bWHEOGTa35Dd0kT
Yfm6fTcXw/ABc5ygsxHaD94h0kjl8yh6Qci6udi/xDwWINxc2KgbZdYWOe2/dPme
lTXHtPW+JAnCRVoG37RJnpAPYWYQ1Q/jA07zKVXPz5vIVJFKx/SAgv33IWXm5m0L
afxkrRTXbpsFuWW24NI2NApAvECqHhRaWj4OHZSRYW0OJUvk1Q0qxfihKUwmTouy
jdi2B5zl8S53X93M06glS7uy4sTD+nDrMEiBEq6YxZE03CcLWl2A7PMmr6whyd82
UomKW50UuIdx3H4glpxr1C0RxyS6weqh8p+d7QJ4olHCCUx8ZJMuvdxJMFPvP8Ht
T+8RG5lSTRm6fjb+CHVtDl8VVya6Yy3Ejm+ue+2bOI/cyrD4g76cAFoDmSmorJft
lhhk5xCLw+B21n0tFvkeaQbtgs4GYH/ChyqtX4LF3OGAECNF2St756gMr8OXY1n4
7Z+MI8yqBGGJG0Im0ooj6mZJE3ey68XXMduxiDyx7fjrsvFHpZvIYAZdAX3p3vne
bbDrfloOjMVOok9+XhtRlYSO1zKoRmxxyhfgOaGpLfF4T/4604ijWobxX6POrxBe
Yk5qRMA0IgAemRSojNz5hT+3BFCLqENphEnXrBkjOoBM5Kj+HAspGfqc7OIA8atG
WJX0bieU2T1h3qBMuDP2UuvRg9w888HezfaK2dN0qYNnYGsJHG2dF1QNdzhb77/c
CLpAXyJOzKiCv5+7+l7516uNKnCXxem0hTJOkrtlNVv6X1qelB1gJxyUJcVysxI2
l9z+hInhsWpbUlV5sFaRIo+ZQvY7zBBHIfL35WNpgmF+Km266pTdQHk+nItDH0Ta
QNOTVftyuZmeYUwsn67ST0VbOpnWEW+N4YLSE/x39kapSqbopIgcysbPaYI+URts
SEaApleguTjMq1frn+UCt7FY0k81hDv1x55ePhapFqIVjYpWlJHNH1/VnrC7V4uc
3HsUNVkQ73ewFrSi0UTZ7/sEEa7jyvN1vsb2iqetAzrg0wK6xWomf9rpqf7Gj5eX
ah6+ifgBzKWajAORwt+2wnwsiEwuQ9C9uhqzdG7rmU4VGbvAL78voWmywVvMDgNr
AshuXtDKdh6xVNngbtfVN+32zno4WAI3emHEMAp5qWbLF6vGbFlk0QNKE+ykyoD9
IYblCO93h/EHfPqqD9w4HIGMMdg62oxOwGK4cNviCmvRr+tklKqwgPAHV/Re6NaG
NaKMXtywJBCRVmmgoqgSDa98JAbfanMnNV5bm/P5mFj7e4+QsV1SoevaZ5ysId35
oxT8dEFaeFepQXuw1+1kU0GKKxQo2TMEZtW7rh4Zr8NGunxXEBzVr27DVcNAJjiq
sUTEtyjVZ10vRwiurSewd5aWjAb6ALZ3H/tzAW3yf428cohYoY8oehOhF9vhxdrs
GuDJ+z4kpWpANLwSxzat0r4r4W74uwBYOS92pp9ue4R24GmV5Ej9LcwFTh9mPnJS
5lOfuPKyJwc4bBF8OfzEyp6SoLa+i5A8aT5sDwRzeVrqsRom87qTNvfZRV5Io3Jl
XOnLQhcdyOf6vAwHYdfVv/cgd2NZGFfhWYEGgeJsp3CxJQOcL5XmB0yXJAt28xIi
GMuVYbYXVl08sGCoutBzmTzar+2lTreC1Iz6cW3PgFZ7lhEZzlKU10iK6FwDv0bd
J7KRlWifc6nRC9Xek5SZpiJTd1wmSmCCQHmBpPEL0boyQyYGx2cSzwmDd6hzE4dK
ow0DToZdXTpKqF1JczoHynZvIYjsq1CFpKNmmxMK+FSQAb5mMz/pFo+kW7Llyqgf
1WB0Vz4KWcBX3+6LnvfwfMEint4W6ReRpmrL76zGGAe4sNwNlbtI/G2SaBu3HUhw
OqMwGXi+iSzCU9yziWWrbX4DRzH5FpbuZwHCkAZTlhdJyMRqXu04ZQWIEIjLMiCN
U3DqDbxERO9/zp5qDbV+YVhuC1tyIRXzEX4Rqar7ra2PBJnPUsONmRCvyPMlM/8l
wbsUqWgQ5tHjjcTdJP/Hs698btdxTogZnOy2RqwgkKh20plc23dbeeDzjcNcEu4W
nCBJ5AeVpI7PpkECsoJAWG0mityT+0gGMBPxRP65PfVbZ+WQAOK2HMRNF95edUtN
RE0iTe5WO3W07ZqEly0h9Fid64ciZUpiy15YZvoLWRzCsUEXW5an73gQQ8An7kpn
49Ib59DFiJESYMLPDxcd/9fL06SD5EfmTXP3eJJshTtVtVDaAPdDl4PLpTAhOvXB
Irs8fE1c80oyYjaTDrkrpRwyHbdjuyqwWDMtP6XdQgicMLQeoGYxNio/Zjuiy5ey
WAmyjiV/GouDIgpkti1xanTswnL/MTcguJA5qeF1aPrnisV8eUb4yq3UPpaM71J4
azklFe9k/uU1SP4WcQREobZ55LT7/DqyBHv8YMCSDwaN3eUFDBtKmdwWA6KFAQVe
a4aQYDMvtVbW6ac9rBjSW+iDl1vmWvv96NiRRp+WixjEne/L753JEA7bdOEYPFou
6b47bEuNlF1C8/RvZDK8i3TzVWRnld/+8A++eU44/+NYMcXRqGIlWCfbDHTlMDA3
qDfLmL9sKftb0lHsVGedRCyI58tMsXqW3UQAcdMcJ/HNniCK2UHrujpny4ctrBfD
Xp7C8YHTUWmsSoR0ByHgSF7YX9mOkm2kFIaAgWfumh1JY+b7YMEl/tccPQBLU1bg
2T00Vb81WeE5I+vOCSvooVHXSWaEzd1OD6/v6Eqtbrllu0FOYipnDuBdCnP4qpkJ
//5qanusEvgS5f92j1U1GAnzqufGo2GHU6iWBS7t00AfxOlJ5GGDjpQECpuhyK8X
8oD30c1jQooBjGvxLJRl1xUIdwMA/5C5RP7Ta3jKfIzBCtoO6qQA+TPw8hsPAqM3
F2uzFR7HuAj+hOBI9xfjTCONKQunu8395uK5B4roedurMbX9PMzTgFk3vzhB+06w
da8yhkUY5yL8FnDNSMEQUBLy00A5fG4tQtdFbnj/SZIgenLK2R2XJRpCnB9KeGpZ
r44VhgpfL5pOEA9nT8jhK7W6tFCd+gQCsZaoDUdxvBWBDy32fIQ/1OnYzgdZOcZz
4e7r1vdbAvcYaMI8lVodtNQCN5BypUPH1wq5p7yWqAO2av0ip5M7evQAD2j0Gais
NOtwVYeNGvLTmom09y+b70kha1SPGQ71bGwPGmucVxFTw5YGd1xLGbviONjXnVR4
gpi1ZAYIrPquQCWTZh7RXgpYhKMNDw0Oz1CzhQx0JnXnCOr/qmhmEz+1tPLb9nVR
s863Z/sRbwtybyZCBqZL2oSPLHZmaig7QnP1hejvcmLvmZelakRP/NPgjstqxYve
BYj2AIUKTrr9UzgFkGRUXuZviYuBTx2X7IQGSxDY1KV6gSzSKJwOf2bt96uOrVuD
VtuKY5Z+KSOpPw07SEITr7d+CnDEkrfwjo0hM6t9xtgWJZr82EmMoDC66IN8qNI/
k6ZfbC+Hypv2da2muJW4yaPQ2gr76LYiMp3obHHpB4rcn+B+Z/UjcBhvJ0YKfMuD
sGe/dIfug6FiWTh7T0CDtPAC2I8Bao40/8Lw3x+CKwjhZj1FlVobuOx6kuelMUgH
nSm0+QlglDtDKPNeK/68dgu9RkV2hwPMgsLsMncVJOhzCH9wFRXq7Vtbfs2l3OCN
m+HrcGdOOaTosTlswl5Of6TnKXtJjOfmsVv6eyMsI1rEIptrVp7aQuEXBfv9D99V
7iVxzYHmcEa5DYZEEIlJUgY9DL16GyDMM1P8no7nucFWiHAda+YldwvxM6ldNkes
b7TBIzsbvVKi5SIRtS7r30X8O8tHkEzLVKZZHUX+gM9Yudm7aY1gJB1enV5VF+2C
0s4fLC3IrKvlfk4yLZro5ddVsf790lpmOo4HH0V1VeHJyaW4eoUpJCb17TPilG0R
4hPy/6kMqbNNhrMzKi/hbCWSSvDw429fZOSPiSzY+YPe6/nAwwdTe4yf2eiKQWDT
Kw8KTD385A16eEtWhoVNL0aY48MxQc4RirBoL7ghQPGzSOCelZAXyWFoO2CyFJKG
3YDBPnibwSjBEgVLFPhPwfPpPExAe66e2Ns/7/ntxGs/qF5Ig8SJCWbqELFqYplG
eoU1fx5icl9hd0LlyvrpRkqyH+4M/5vsAtO6x3F3vOQBtaFboF51h9jCEY+QOICE
x+X6iEluu4+U/b27Zk0B7fCiI4ctmk+iNZMADWYvDNlSZo4LrMGYztOENzuSsP1l
kCMKUg04O2DPoI5aabYWupNKDSumNKsFFx1D0CJ8UbEhFq1O1x3TLcY4jJFcaj4j
dXv01ChOnh7/RmNfS2NgyKatth+22ErbEMZMcPLGB6ZdchB/+Jtg0iOZdkKaZeuZ
om4BFViV7zrXlLhbQTEdn+Agc3MtJir8Xi+cTyoosL0OLvKrow0syEejuX7iCdww
Ro0Lz/CogqCy+Jqejqxx4sNU/Lng2Q1jw3ue2XClCKO7DQDDFxOnOPyk2lGnvBDH
+JeCWGSjt/SNz7LlKMETW8T6QwYq0WU0q6oujtBQ+bel4QhDQQDz28TDHiqUi2Bf
D9zEw9DYIGxFD0P3X6FeG8NgyOr8b1IwVgZBQyileO9KfhJ5dJ8k/rq34EebA4Ql
zn5FTd5q1tKm7hifNAXzN9fsTvu2eFqvDZOR6DmGL+akXfsgy3u0N5p2a9JMgHGT
0waH74ay2HH3UvT3EAIFPK/2HRtikr1VfLjUHABYYL2tGJ70YAdGGVRj0GlNQGsn
W2auBieg4sWkm8oAKBkUUaaPEnwIDxxfWjoZAnmxB1HzFkGsMfv1KyuXADzVbHpf
Z2ghHMha9QO19B2ICWn9jB6DMCulzmlcj4TQKq129hbOTy/pbSD8hytYkZ3ISMJS
EBjns2vjFifOYGkhgolQJ7fa6HkVThpK8DH5ke8AdSyZcTcU0WEZkYqlXanrxRK3
64o8/9TxFAyFn5LI7jGFVXu/f+tj6n29J8py6p9a6epF48XcOPWQ5MAlU6zkc1CS
+Mv+fq3AXa+WqjTIdLnuGX+WlJMkc/1F9v3wuWYjafSWbyLxt5LgtlvyvgHIaSM2
Ka9YdAMEm0hTmjmdsaDQRiyoRTB8moAiULyHObYomLr0BbG74IGFRSX4ZyQzIMA9
TKnvTJLEVH5X3AK/9MCRcX6hQOAL7zGqzvodyQebBKdT+Ih3Wweh8QrRe7wZiqdS
yHq5kXuW5whzfutIGNFN2D56ohlRzixo99/7HToS56CYRXuTe98RQ4W8mHaZGA33
yT36Ad1ZC1hCv0etMJEeEs1me1v6pbF1+BRR5g4tt3M5YlogDavJi8LC4eENM+D0
S7nbUKOb0Yb9+35VdEVloKXgHVSotcRSMYALVEO/tyPaIT7VGO9ncsWfnWy/feJQ
wKaQBRNeHXd8GftsZ436jSn4JpxgEue2hZwmyMLQRKhnaxpzrXTrB8sj0b97PJ/M
tr+ZcTvUfF1JknNubMl3O0sZeYMH6Qj2jezVr48ivv17LDh7EVDBjqi+qEhTIxPe
W+hNOPtGi3+ZGFk/DoOxVqdZEmqDhqiWShgcIsyIvrP/tdvbXRc3oE4MW1p6CDAU
akJUUSzE0R3Tt1orgzNNtw+fydKV4qqeweH5wBtjMtxhSdhojSMlYNcTsVgWa/bi
Nm1QGyssK0q4AhJQClnhbmmnKPEvo+eYsxogv8DoUvv/3ZGaNMmQi+9JAbRcBVdk
m5nKqVrApupQI4XFsjYxSQaLfibzcNULOVWTeklfrZkEzWT2CYnnlSv1lXn93mUZ
iMJx0OGF5Go8VeFNYxPGfrD+DDo+4H8wnzNkWZBwG+SsyMeDGF6H147hMRVeMlQn
IfcAyFybJvIpcL81l3nyYGhOmZGvvmWzlQ2vzHbO5CEu2Q1IBzaBLecsrQmN/Ic8
+B3ATXgPcfAH6QLSju7spG6o/yfeQSFtHcGGQuSaPOlyNdnA4tNvz4x3aJdxxlrL
qhY6xkXPQ4jZKR5I50a8H45UOabfr3b861dez/wX3/qaq+Yx8T/S9ln5HNJgH3PO
wZVjQKDO2Z/irha2xwIQ+cJOAf4a6a4at76fDGQGHK348hiD52M5dC0IdpD0ZmKn
+JXr1z0m0Di+J0dym1qpPVxmQczeBX9METL1PuUgE56nWcij71NQOiOaBBkX9YU6
uUFsA4/bazvhL9WGQtw378CyRdSgB24wCXtYk6cb+OBJurwVPE/1LxtrJXX9ibMp
ZQN7TPCDDaYfB7IuZbfJa+WZv5nuPehZMGWkxMa57vRh7Y4FrdoitEgYYG3d5raz
NJFV7y5Skvdys41nCpEiLdRvOjoQBLUEWJyRVytxCO7txHntbs97UsWPd9jG/K3B
SV0EE9htGDs7hewcBYXl9MpwCO8llNwYbJR/4QvyPX4Rd2cLAniLXQHGAyl/l+p6
1bhS8qczNUiwTvIjBo4e5zBb0QtiRTYYUdwKUeGww+fWlwb0IKC/JzISguDGZs7M
K7FxqN+TeSDPW5DimZ027SmOWaxJbm32hvfnoZVGC7uSgg9DxQK4vrq0mT13WCSK
m1pEM2d5yG1aEcdOzTOXG0IH4MoG0sHuQ3fbb6e6IHyCiemiOHruCsm5Uo+AM9nu
cCz0njJATAS7i7s1dliRDOrdp7zer2JeAHgKJACAKFdGfwwr8EJP72QT1D49mNyG
NaWqXFT3Rwz2lk9DKqE2saoBiOfmYmR6W3gXsyZX3GDeqOCHv2GHQl5ha2Ab0Y+C
QwfUb/5G+nDJM1N+8VijQhLzW5GTaB+0j3qr656WUIVvpHHXGhAfTGj45hYnA479
BoynNrb1fwKij3XSWfKfehDwBIkIZVnBHIq3ZJrOuAg7rrq3xR46Fxy6mtsj8d3j
gCknsMRXnZNivdIyYY/vVM4PjJ/Sgn+bbQR9qUA2KnbRqqKvLwAR8It6TrjTW1vJ
TcWTpIvM1pxsF1iduQDD4JoWmf6xinnLXG8jr0xzopE3nlKB27qiSHL9/G16YwIU
f3n85/5XPicAn7XnnNQQuhdJ71PbHiQU2Gz7++J5fyPOpIbX1wn8D+sefuQ6a5iR
o5tBN62XEF432BbL7XOikHShlHvJkoZs/cyX5tLPtscg1qm8VfCZiZZYFlLO/Gp7
BetvXJY9twk7ffKqpK1DVjcoYSjDQUMWKXxiR3W6YtXks03Ie63ijuQg4+o7y7tg
uIDZRxQtGHG0LedKAJYg/Bu6O0ufQepleJyDvxVGDJYv9GWXCVNpF1lEWft993m4
kiXHxOS4GFhlrf8uM7ACpWAZ5QCRgiPiZ9xvHC8nd46c5eH0b00c6kKQ4/ILzQOJ
ZN43J5WAnNGc2or0TA6BsnKZYmETIc7lpGBHY2Br8XBpUQKArSGCZ4TNKa8rmXzg
EDrFLnzjtb84pHF0j8sRn8imMRf4Qta1GGa3G+mULbsPxYua+zHd5m/5sMJHXAgA
1QOkxV2s5tHrgTDCpn488BxN8HED+TawRxLXwdbD7eBUNDxjVTTb0mzD10JDCDB9
fDFOb7zck3meVL5AMVB3bsdWS1G9MXtglUQSSV5o+VbX+HvQs5IAp62rg3qhXUnr
Xv+GILeNQCppYTDc1zpZbJB4RApYjJ39D9W9BP3TerGu2E5Pov7tdtXGwqfLgK72
nu52mQcheu7JSCfu7j1rzmef6ESLSS7uflB5meBgvPebQWr/VhGcnwUaOLxIMIl0
RwHefnm0gw+Je63E4/7KwP+fTgKsYH1YJrECVYCGdDeO2ym5XK1Meq/T0gIwMuKq
ezkszVeoz5NGo/1+T2qD1b3deta6MdVfjXsBUMZKg2H2zU/PjG+OwdzQfgDstvkl
RoA+vrtGN8ojufijouFw9LHshL5OPJ9jq6/G/yWdPfOT5KrGDIZ9/nrwvqiWhd8/
SXYIJ6nFynBswaADqwyiK0tqXHseAX8vS2YjttMIH/npbxyfzfbd1WfzesSpegCu
LRNsewwlgxDszBEivIVtRsA6gBzY4NMUwIuWWHEImnNJshk6iAE/8fAXhL44fxlE
OnXIKUVQpxyeQ64CtUIb4FcEwe8RiU2NC68/4Ygt1WslBNLBB11yQUG9KzKLHOpV
7GU1ZTbwERaXu0Ay9eklGYzuZIQyRe/rIBHzlqwo/dZLJtDtniDISE+uMrgfA+cL
nQVOc/aqdb1IPezx3eAiLOtYRytqVpiEOQmElLdqf7hfPKyK7xrlYkQajDaTwsG/
gtGTklkKO+ealupuhdePuGVEC/LgNx2WL7nZwgsMBjRt1S06Al6s4njYtCx0Hjqv
6GIekczIxL349zstFSNIep72R6kmGOvyFroSdMNcQEv69GgjRr8J5NO9ma0OTKE8
5isOlnANohKKpDHIZxxUUYdakJCZrT8mFF6lqyv3Z8mkKq5RvY31TbdjdsuYUGAH
dyU/fmTBiZdvCmXWLY7bqp+dg6ngHW8+9CyIImJFDhy8ASSBwncaJE4rN4IdIVdQ
vyKY4/BXVjGJBgy5j9dOhg9Fwpki2x5CXg6K1+M5ZPagFCS6areuh/AyC1tExZgz
9lXLVgfeTgxonsbZXnL/Zm7z+NgrLZCfMP/cWyxLiNFFlI4MVhNNAfYxuciqkw3O
3hlSgGWJU1ej4R6ocbTW8RuXCVRH45JNDhnHVtVG/17VLVuvatgeT7Qhv4IKTfwv
evlTWiWGCrDe0jw9LUU/ttNpBmXfZ/4uuu/UmXKLvzbjHBN10DcYl6mSpg0iso+H
T1AnM8yM4sqL0QYtaTH5DVHCIqonImvYaD191IyriovabQLiyBmMsRvSgRd67HtE
a1K5H083teUFyd3TTwGInNLuMw9mWFScpItMI4dH6wkarNLEGXn9Brdp5o68HlhB
4fUy7pSRLbWK9I47ptr3JhT4LUdLr0zGNVEQ2spOFxDPRinb2HC2gHSYSzEaQT43
1M/cKkh7hJxDgUgtkHqQ9Uw5640QvzMaJYspNZWfM4m0SRRnWjoynwH6QHP4H/AB
gw+O6BhMhSqmKOTSAKI5DhKEc2MVKgvYCSp+4TDPrxJjQqpNJ8mi3RhiEP3yqOxb
TT0S1hV0HHlVTfBv5JTOEdkqGGpYdiWuCb6GZlcQV9bRXgA6rz0WKuLG78NVR4mC
tJ8R2yQkCfuTiEf0kzlsBaA7EtomMJvaCsQsvFMn0xGNMamMqGtMG5B0AhYukj+V
oSq0ojLE7OjVoIDiJwjkCXVnOU4f+08HhwlPVnShPDRKAWbIGXWWgw5O2yPArYTE
B4bthE9uYKfVAlCtdeppmHnFbRcDiUAEHrRNeDh8JynsR+lTBZmndJVHlUFm9KvR
GkgP6nu0iCAdZdj3g+nahSReE3q24KgpCg92/MSEwPS5TtxcVGOUAsYxMucd7X7b
tm1X2GjNna+4fAhB0KcgqtAhKuQD9xmYQEwpe8CCNtcPr8o/bKrPGhbYMKFxK/FR
jQAn3imiDYwdnu/jRGRjq+2crXXW5M+qakTkfpVg6gfYmnfPonfNJV+x2UyMUC7v
74WlHYmC8pXyuz8SXaKzCn2bB2ZpgVH18pchluBe/tAUHVo6uBKRhTh5GqOYgZp7
LBTQ/RR2Cq6eiiflAicd9NSdqMns2j+QYQ3w1xaam9jBvBRkvJBJxiUReIxXAOPr
FvDN8gJV9VoYaAkTxee7osQyY1CbLZmxiir4NsxNYO8k+IJVs+YBvDFcp6SG5gXr
5x1Y8m4H8Wjw5Va7dpYUBlt/yFz8KCZudyqxqhsBZ3pxQTd1u8kFsc4mOTnni3Yu
EePZci8jsM/jhzzR5lzI0z8QDxifZGcN8pAsUVGh93zrUBsgZeXqJjrzfZ/hOPJf
qIxA+HvaYvUWXpc6rugDXBzP87377gyFwSYfl1aehJTb+iNKk9Ix8D3TkyctyEYZ
hPnODIe13JvDzQx+xhYaqOFnu8hU2/6pibclJpcrnDGaenmnLKCrjgOEMePHH2IO
315S+E6v3FMeVjCtx5m6wmZlBrZuJnK7+giccoLbvaI0ohFOmKR2AUL726Imi/8B
x4QIOWPMuupFrk+01IfQlII9u5v8no90aQw1D1JDVU5C+zaYx6XufoT8jkVm3nfz
mahp/j/ZFov/wYWdIM9rgmK8NvcZYU+56jFmBE3k3FU6BIzMx/GVWYXAV1bE77Aq
dmmhFYqsArcKejPo4GxgEHO2/b6BAph8pm1Gw3VyQS0dy4BnDCrtgRV0lEp4/4l6
Gp09P+fGoFvCYmpVy9/7KbdsvA8Ew5HDMndLDYB1ANH0Lf1ppSICqXrgTbrQvxUh
URSpWLQ2z5+Jdkn2Q2/WdQxNOYP3PWj1FIfME+eKZiX8Z22CI6EM/mDMr/g3/cNH
bCAg75yle6IHO7G+GSd7u6fprovyVf1xlmL+AzFZi1a9EikelMufD6y+eE6Jg8rb
U5REy8uhtYkdeIIoacODKtYw/nZZOr125U5wGSeeFZ0Ff+hXhTNOTHleIp92vPbH
agiwk1O6fBeYDk5bx8Z2ZAs+KmLe0N8ltYx5Sg+eEgAMO9ctyLDtKDxseyvTGyZM
4saseBIWXfenNs29Vyx9EEomgzPICpRto4tQrN6lvkYtg2zRWXkohOAtNQHfOBWn
WECL+jVPZrk7fzFsZkhGpOwZfaeEpgPt/KFoep4ivDOc5wGJOAge8YxzeSm5SbJF
HGmNdhFMD6EHezx4dA8GAbaXNt+d2MQbIa77VE8/nbozuFZmrdhF/nWv22MfJG1M
Pq4QUecDho38emhBHGt5BPhaLPkZ5c31JLLb3x2W0pH1wFIgWpDxJR8QcJcZEK0Q
2ETqk4QsyG1csh3v/w5MS25qP4ceK51wPIFJ2HT+/RoFZLBXf/TLVEgDizmJP1D3
+VuY0txJoVrtjmZ69pBVPBYDgCvWGNEEu0zdRfv1loKFgXbHqUhorOWlj2fgMmgq
lDZyf0Gm1hYW+TEo+qsC6qCbULru8kWVwz+lz9G9HynLZkxjmA9Kg5oPZeLsRSp4
tCoSM75GtPfs+Uf9yCgnP0FxttYYJ7kxPdlKhqAaKijC9FmPzpanhigB5lPgWmMp
26hT1w/iWSrCvHdj7/hCbVB65sgTJcKYkb2SciVeFhsGq1qnE4Xra1rke586Wn7Y
KFHE5fxkNWiWs3oKnOWO3XN/NnsMMW9bc8Jbxtm840ex0SEtY7PC8aLlO1/6xBQ+
BmNDoRVcaLMSP/17Tioar3WCptULWR+1ogu23FKnfKqKzfCiBwjQTFSOHZrqYey+
UEzgBl7iyAeFtGrc5PmBt9RMb1gXMIzCj7jqkRo7UIrndD0t4gRFuwwrIwVHPqEL
DEINYJR2ASDZ19VOPxDf36nBlTJwRyioG5jG4Rr/X9jSuaoKW1MYXSA7nBVgG8cS
gOYPoD15LnY/DVty/cHKMokZT2x5a455DMultvzHYbUiefE/KDMbvO7CxkHSdvSr
2Uzwi3CCsKDp5XQu9r762ooQgsPSrX62CpcTwlYn/CXsT/xA6MFWVFs+I/ttbN6+
6KYNrW5bDvcGBPgkWIEmOQ8VxcVbwksthAE6bN+eYIqGz0kQ4LvgdoPm6TICiOuK
LfaWmAd8TIoaBQrkphb0x5usfB1T8KoQPQTdyC2IjqZhc9t6iom5ZIU7miTd2cef
EJeEyjWfVqCxQdL4+CGUzJGSY6zfRL+n2roZivIvw9+utEdoI4veWr7+k1MXZhnk
u14wVFSb3EdGH9lgnsMpBBYFiQtMFQEXkp7CPrEUQDyIxeniVPzABQkuci10p038
P3TxEN2WoJ/RF3VF6BgMEIR9HWs7JwjpVu8WS4STYGJcpxyKMikzMvzkIl6cXy6y
qC10OgNxWeUCHF0vohhqCJQuGMPKSdFZ9KmRYPwPQ6Ng7ScCma7OANgtFxb/6m2/
VBxsR769FwvETggSjwaYL/R+fTehcr7aNpqXXyGIFKOA0zuyYpG7GTs9cmvBtMwt
1jZ0y37SSkWzKHUE3K88iMtl4C0vbdQRhyLUh1spBNxCqrNEKAyJwHEces61AX1D
qsbbWnrYZbpWhx60PtdtIqVIGlOyUJt5yqSfWKoylvOJaIAbCOiWqeZp9b9UczA7
qgCHwm0ChiS9Qy4MnGX27c4x1gNvUfHMzlVUBh4YFGVWVXNmS7+bPrRvwo2xnd7V
zVij+9/WXAl/U/UrvxiVkSU7ihsYXlAPKFBahjgQboSZFiDsYzwavtTgAPY0X2/i
1A4kUwtG7vHplFWHlmqMxOwhUsznh9h+zunaFtRXUrw0zfA6FdYs5h/Dy07qZQnB
vuiCu3RmegbNEmsvS5jEnMlO7csmSGMnKpZJs5Gq0bktI9njqWWUUrgP4sF3pIp2
XFpp2hRmhT+fD0LRiLfw+gdzlezL+8UIhRITtVLSXD7lNOgcjILpQgPCDQia8Tpq
yas6Kmf2ZEVjRC16jTJfBr3sB03Kqyzzmg2IGEsTdKsoRLnv2Y5pFWZQDUCod1Vp
T9wcOeZ52CHgZZBFKqsHwgwvnDNzpy4J3noNgsVfsVOBXxjh+x3UD8+cEZTSfFgM
HgcZEIaycXZBOUzH+X5MQyf0q42HQtPGIoLePlCfrGTlcHNmiTqd/2SaBFjGzq0s
0BJyKzrMrTNs5B9k+3vuD4l559zA8Qme2GNpvO17kp+EJwcnA9y/27f3F6l9vNRk
hb6A8u+d1ddlWgFwxdN10HB+GVrgJyU8yvnsvTW9Bs6WqESyiUfZlxe4a1UWPAlp
V7rSzYBM0uSLv673N7OVfOFopXWaOtM4nRUr3XjiF8r/JOSJUpFMOXMji/z0kY/s
nEtq7e1mQ8wom/wMy7ktJZYmTW+GPHIYGnox1ZHyIHoRRDvavQfcbAeFpPjsy5x3
iOFaiTF7/XCNe05M2B025wqlDhWKWEfB8fIp5cAhwjBd04s8PQwbrRvsgU4S4H6i
1E4mmd3ee0kolyE1rWiJa/BC6CPhcYJoYlGHPXxH5ArJ08T/7KCq8pv9OBNKtKK5
RO0JK81CtG1DDtmmv8DNt2OzbGfYnjXPVKJpMw8IhfR1hOq9zOJYPCXxmmV5GxGb
WxxAnrrFjX7bG/vdvMZNYIFmKkIs8jz2RMjlNhd/WQMb3bMi+7y8mXtHy1cGSjcM
FzNJVLInamgSRRaxFc/CY5UeUJsABJjwIcRg12FgpIWHNJeKfvklAD+9GxqM6gmu
KwztZGJzaJVCutYbBqlIRgfojcSOgGtwCqX+qkT9srN1nMJp5y2iuZH8JEtMGdFr
qiRWFz9DjtTWk7xraUyWzTqOo83J62ZbXikQ8ip9eXm9w8EPwM2dF90Drz8lAW0n
svsSBZ3IVDY9BjyuzjCaXU6uLqhpMUNxOIyG5DfWyfRdCjgiFik2PncZrPGCKNmo
JOIdVawsyk/nTkBZ21WcgzXTUeBrGeNDDp2VbUJjzyP8o/XO44uaXpII5oGv/TTs
KJEckiiWns+Va+H5mBDlBRiScUOjB+M7MD9AtQHgCu1giUybdSPoKja8cJn1iDVf
/aHMR/EWOiKlg7Mc3X+SEGADT0qndCo9aif8mEXGOG9P1yya7zEro9tUmRcn5qZK
l862ylGtnfgchnqo9yXSB63FZCXb2yb/RSwbPGattgZAa8U9M5oLXBvmb06eyG88
Se4g/kTUopDjmtHZGT/O2Joc3Prw3VJVvFtycvm42ibtf64LDdx8ttEQprnyMtjh
CPDFj4eYg/LUbaT0cWGOW1bwz2t6Ytzo3Kh7NO1by52hmTv0unBPRef4iI5X0TjE
ME8XA3Nos49f6o4XFQ+XMyVQtU3gJPbOlZK7+LNQPAshDkyWgsPRtwDQujHZtAqe
GVZb2vwLYXEfeT5urpW3tMsxaCGnDQwSVw4zy1sO73HRjfxTRY9bsTu0EH5K81gY
XRCytcmakiFh4cFXn0Ko1PduXCX9jeXnoucom2jgjNN1rsiBbkCjewkg6sgpD0Qc
F/te72yJGRbuVKwaahXtjAfZPSRgEfBW/iRu5AaQSfj+ywTd+GxWE4zzDiuNTr5S
Yfaz4Lsg8l4ZN2uATHttpe5euEkTQN1cfBVAjjHcKk7BNg8vqQ9pP4ZXtM3KGV3a
YebVav3kkO2oBksEBTn0Ou4FkzOX4kbKQjJKZogQHlrygCmIXCiMo1l+/5mnPqP+
TxL+lEfQzHdfVvK8TLUcTGPThF17EboSdBlySpn8kuc9nRrTt6AKNc8WtfajQXbo
s81T0iaBksuEc9UwDuy6xL4ZPL18EWIAcQP8jz4HIzNVJ4K/kMzuf3Ja3jM2f5OO
ewWSN8fDnI/xP8gSMHK15z/ruDKMg+IeovG53FqBwbVstMQRCjXQOvAkft+8J97R
QvyBBpzw8gAdC2vsTeNOSBOgmZpvxkKbG5vVxaHnfB0/vWuGGjJ+w5pyocL81LOk
/pos0w9KfI0w5PaEtf9LlPSA+NlvyzNf78fIEv9jrWaEKX3hlX/mr6nTP516q7+O
X/f1UkIMo3AS3a/ZQKeHwPXGiK2/Ff8WMjowOQhRVhVZs5VrDaFncVZ4ovza4lQl
CFk3zjz5RZPFKCUCcEyLbKz/E+HQZ+URCqdJZQ3ByfHG+JXKRzit16x2Jc7LIw+L
ELwbrjs4hQqG+AKMUJWJDxVl6ZBwK64TZcvY5/n/KN9FEv7J3CqPd8ydnOJDK9sW
+i7+f89LJwEsS9qCwUM3uQ1ICQY++phu3h0DNpI6JTc1aFFTHj6mXVAnI/fUYaCX
Go4D350KpWgiFz7CZRobEgTaBhcLHuERwk7kVDALuPVXFd6/aMr0dZBrA1mFVM3z
KDc/eKToQym3Cd3qctN3CVNOUJD3Nhf4W6A9ynBkhzWi+nBTl/cTJWS+CKzIXE2q
YmBK4Pfpzar9LBZYNo5xMpxOFgl3cZFyc/XaObLEPB3EAuFEp1Ju2OehtguN8Tgn
LCKFFY4W6EMqVNQTgt+ap1QSYjR2ZkES/T4KSVTqGLMfL/wi65lP957XToumrcwc
8F5d0U+v3HJCLdrf+PZL35cyCS/lPzfxQ2M5EhyXx18BrU+X7uUf1T2tyaMQAmOO
GfR29MBRoH/uPGm3Avq+cIvcwqzed1foIF1G3kTL48Thpgg+6xU52QHLuNQoCEp1
g6Vj5hcOGdOhVUC+gZBoTFClHbdzjLSCalGeyMUvPl4IyuZDoj0JGacoWm3VMH3T
UBUGNVMwPX1lPMalMyYjeNZy4QhgZpxA7WekRkQ+jFtr5rooXdpWmMCrGP1asZGb
dDftRwE4KlS3BvBGYD+rvoxXkdgg5GxwvVNIB9ck99HL3ZRdZ0e9KAZZR+ALrR4H
111vEVE1jIcFEm/ME4T1ZHOvtdujl6RvkDtHiKRBoEVgtN8sJuvqxLBxOGcCQPv4
P1YAem0tuVTWpfceQeu2A+embrF4Dm84Kw71UhyIf9m25iIlOoICGD7+ABnK61Ot
ERs/ZbshRQMuVR8H/ZZLryFSc7qUzhesL6mi0b1fyhsgk4fkH9BoNGpdS5I/zP9k
boq77b4zaCXob69a114qLply7V/4D+MJZN5b52YeyOMAORxnfkkpVzEDDSsabI3z
GW+QI8nkGo2CzkBaxIBkTppZIjXWcvh6GW1p+9EZzXY+TbL4oofXVKVEfQ1sagvv
mdZRiI8acbEbtzTsvER3QcikJHQ4+t2dIoNO4PKpKREFeXjmfy9uTTb1I9lKvLKL
0Lgu6MZZmnFDaoXIZ9Q0lNCGpi0tbB/Qt1G8AnPBx9UenqAvo12EWvhLoAKCGTgc
umBi75FtkI9pMBSz/HhwceoEu9vK3n4gQe2XiA/bUhe60E3wZnycq2NdgQHVZPfp
iyDt5+iGzdyXAgNJW8kgDgdvpxtmF1i1FYDvK42SOq3LW8SwN5VsUGkIjKB7fPv0
4D5GHfED+CVYKHyRTvq1J7ZjAHmHL5rcFWCEIu2BzgFGbJBxsA1DRtT6FXeNtI04
a/9AVcL5p0IIPnaQBWgYzmxAAHpaH36W9zPIB5aQG8IvLR72zpGTtkeI8eSqhHM8
cZMAvzPGCi5m7H21nxeCoBeeKmVEhiCVRgjIbk6vKpk29ZF+h1Aat5JIT5RBFxmE
0Pgj3c0JeM4y+pWLYjl8V371h3lUYoyTecRyy4NmuxlmOJN6cB55fIxPJFU2zAbT
mkElI5lXLgUgmkr9eJhWBAqlpEx5kMKTsKP6uBHeYIoATgysZKVUAtadgT/Eh1sG
gNcV1j3e+2GwA1nvNPxmMGU239XI1GquAjVyl7fgTilT2zwgOlgIu3+VnvyUsB0J
yi7A3PePrRS48b6ILb10ui3EaoV8MXSaWK6dQVYKQjKPl3e/1zLwhaMHa2Du3b2Q
EvUcqj7eHRJaTnOipbDGVHO4Tnps7+EDZRXJHabESHDZP3/wDhUUiacwsf5GXjHs
EmOjfJp3gmdhLs78S9jkIm8FhOfT0kS7qsvrR0XI+ynXWEymk7hZAvHEF2h8QIEv
ZjRcc658ot6ULQ0SSRYZ3m4m/f9j0XCsBjBA/jQoiVaNyA6oBt8A88OX7D1Anyql
vEvxhZPSuZWRLdbjgeBic2m3PDN0SHzUYQ2Q5IHmQ3FzWmR39z6WXTfXZA+EzGxL
E+t0o316XtA+VoyM+Mj20V+iPr6FXosaOlzuLG4eU9XIf7+PGGvLxmoxVNN7RrmJ
eH/KlKCdhzUEua8nqgmgamPN7F6EkOZkGnmehjbKlbqNDzrZTYOqDd3d8aFpPGVD
qnw8CscKgvWPnL2Z1XSeVk0NJcnRH+1afCw49WorZUwU5mVZE3yB2lCa+dv7WNRD
rmcgglOIJI6iWUPYKDPO1xvfpBmfN0SlzKp8j1MMJKxp3a4GipIwgZ3/0McaWS/4
lz7LZAlvUSJLjtBamSxr85KDZCMoUC3vY4G5mJbf41ewLYIdLXwnsbgVxkGu51qu
w3vEaPKl/j7rHYLVW+rADEBgSFjIsVXRTmG/zFFjOlAHMUaKQK6peIqyxgRfBPIm
6RQ+nA0KVvwp4C9LIpWwxZMCI8+DJUOm8oOdD5YzpcaNranSXsUQgwj/Mohfuyd8
n80yJ8+NTZkykEu5iKG86y7fDpVK5pU7Av0vJ53oK8j+bsGL5VoL2FTVcrrcVMX+
2PJyumHHdLaLimCjfBzBx2zIdTIINeQoGVj3hOF56ssflret35nkrP1S4wAyhYwz
A1DZcEMnrH64xdhPBcf3xj80FakM3nUzy89hTW8cD6M4iM3iAk7RWFffa2V+CLay
Py/JdD6wqV+TViRVxDlJwWIR2VDufurNo68dIloPcoPoIMPle1BBlEsJUV7pe4Xt
/fRE0piqBJKD0Crj9FISZC/CsTXMgI1qAByK8aH+KKnn7EQdMU0J+P6X0ufZyuW6
kuViUS+4g4JLLRAytc6nHa4w5aw0Ww6+aPwnVs33K0TJU/oifvENwP2KgXsoeh0/
f7pLSr+5vmDaOkp9B6i29f048F4ho3AIZ53fHXM8piXEE5FCIm8C4wJQZ0qP33eC
dJPNcUqpT+uweTXY9PrU7PcQQU8JUrkpIN6qOy7UVHC356Y2klv3WX0mercvzdHX
KOjiY5kdBOSHOYLrcHkGh3H03tnLbzfERl4r96rFbpyRk/IqZNQGm3pweIIIVKo3
L4DhyXKmZx3sMVoXMwyCJbiJjJIcjYbNznpagk2cj6F0zw1pUAKbj5RVsLYf4Z0F
6biFch+fHy04H26LXFVeN+KLOvLNb3dkefCZED/B0UYtcqC8U33htX37n2KfyYp/
LFqX0iROEQ/UgPQop2gaMMoEk5iKuq1SgLuYXtWlEcqiCiTGRl4XIM68ICdPofqT
VZikM8FujazKu0xAmffUPkvAYZFl0vHOF87pLCGZqZEkw6jgpCIDT9SSYbmcYvzw
iDLVJdg0uKkKVlnz0zSsJ62pFYGD+bBfI6GA+9jAEgItMHL4amozQdaHYrxB7Y9n
NCCEQibPvZLvyDJ2BVCaopOYg3hceCc1VGbE46ps1+MqPkT4GpFpDQ5kX7nM2D6/
o8mWuRLl6VcB+If3XSYFiOkgN5Rz2PeVKomvijK1kMtAMk9+E8IuSUfcXvL9gUZ7
qibl9W70rgjxyjpB9Zb/Pa0ZxaF/XrpGw9dEPBjjhv5jH9YPzea2wB7F+h9kvndR
Q/E4OuTftoKxrLeBhiIG0UHmSnUa7drtwQkIrRzmqQyqAYDBe8/occwcSNKQSvGf
4qgy/FI4KgT9sVqjyDS/FlozFuyoUVfO1C4RQuRsgvjm1Sc4Lfcbav71BXlc73gn
Gk2npUlQff0veqV2fX5EBdHnloICmyq9hClSqZsYrykCTasqBwZFfV4OLGXnFMpG
HSxf/vmWjHm6q+PFTeGTuN8IMPwfo2YwLONEsCNV08SXH9t9lCfxFUmf29eQAwwz
0Kvdpq3PgtepB83umds8xEpVDVrvPmwYUB6xKckoHgXN1NAXfe+uyjfCs/9FY8Cd
QRoM6x3GYTWnKLykRs7R7FZnFqd+1izG/SER31R4TjtTqNDRuHDdHDfv68eeyU4X
i19DbLbZnXRdzgr8YudcWtLreh8aQCHCZ+b4pvKK14oXZoXa7iuDeirK8NOjR5DL
61yCkd0nPqUE1i2Ug1BFxRMgnB6H77zlC38iO41rUnzZvKnuypv9mWMimA2T3JPg
aH1FCxCBP+4JUyak0fN1rsAiOy/yc95Uh/FPCbhARlA/evU0zy5MGn6049qAcALW
P0o00BLUWgvev/aDydmR+3Rwq6SeWFgCvI5IrgZ9dyTMeArLCo1oTLnKh8x8adVg
x+Z3duUb6ArBayuYfCyZLaQUCfxD7TD5s0tfzi88VIcPS5oT1sxsgjHjzOqFkOKY
xM6QBwiOdOR6PxD59teE98jxSvWMSR/G0pWP8HoMoTqzrSXibn5hKnuHJr01kAmV
Qve6aofxBkUuHtpfrg+hgOAp51ijK5OzKX/3I158ELbMpjd0UfqQKZFu0JwjKyD7
1GCLDa9O9BBwyLRKx5BXYug6R3wmJhHfIWwwSs4iIfwNC593z0fM7TIOWz8qRSWi
9VgncS1Xo+WE5ICEamu+4IZkm3yaVZECyhKNvhozhmHGkBix9/3MWGG8u4CjJq9M
nvd2kvFs7tjI1iw0iPC1Op5fA9qT4gSVMzvpSsGA0vuNmB25e3blzpHN2WuxmgNt
mJ+7YjnrNDc7x6b5q1czz4j0INNQ9hWGTARFS8LPSz3EDAREc4ZlG+tESk/vp0At
qo+I48IkvMMO0IaXVPj08ttmcc6lrlz/ezng0U1O3/0s5dvvzZhegflHzCKDJsny
STg1Z62i7EcAyr/MnGkcQLN7E52oFQ//rLAGOOZoqCDhcdDqrheBJ/29iMnogA8q
VxNTogWgRbataPBl1+uXtRZypcm1hI8lmgc7luAZga/zTtnRH6USrFd33Strp1TG
EYfymYfB2BFG95/fRDbuGFBN+mcLboTB1zjtX/yxhXVnVdtaYVO9C6BEG0Rdrgc/
vpsysWDJjfFjMKjdQd6J3edbfpQ3tA4PlcegPzt3KnySkWvkpGZrkSu6pfXhKjzt
hiYP9Bpxg8ifDnzCTRBbMCQDvIHhBMTKT6jBGnasvY3FruhDoZFqOZtorUw6BVFX
+7E+2sCz5xTtPVVyQzZ9P1vzo4SM/GOw+uIUUxIFZcjp+pbp5uSoAOL48lhX/Fc7
PaDfmdsRbSYLysMnU56+t60L/EBnjuhQsareg6XBE0HSwq8pVDK8HCjC9E2RdCvI
G3nAVBnw9fKfwlh4lzxhV11jym6OgsVDe4cyp9adtl3WqJB1JCxzF/A0DKdpNoiZ
LNXHBkMufOjhR2qnL6wwIZ6l6rJdcKbm5ZDo1deg7Cv5oEngqmBYX7poUfISh1XZ
fEznmh9239ZitluurGEwcMvLKOzafu3VFr/JVqcBc4bpDfI8WZZhzIrsUCt+wpj3
3EZFUWVKHlhfa39pKk0Mcpq6EaPjWt1qtyRcQ5dum1B7x16Dx8mASeX6OyYVM6jQ
d44X1Qg83MYvRSoEzlTQqlQdllL3EdgWahUD4dQfpbXO3KwBmg716pQpXsvmOun8
GeCj3CVRldh1yx9Ixv37c9DkHFJR7baF2kjpWtEeqcuRx0T8O65nxzh/PgsTHfa4
FtN9m4ZAqcnaSJ7K6wcDYRKGsODXMmnY+Nfpr0frNrKAlpnWNCU7hx/fFoUpHAeO
IuUdXc0+mdqIRC+mS6859CjdPII4xK55dHo0sDQyUQSqrWQRiqTTf+tKCBo1KEbn
e5A1ySN9S13IL/57JkjBY7pGMFxQFm16qxRxp7xXLiQOPIc0th9PApjpvbZtMass
BdSd2Kjq/+FC5Z72x6NwG/jw3r7IcJcAirQKDqf2l21W8tKhlwsJxAhC5A7ZHusB
EygeYo4u/5jyq6km2rRlfRgP61C4XruVz+V3uttqmQ9O0J8jj49pRf531H6S/Ef+
wUD4dIzv55AwH5KGP3Tg3qkA2Ug5xKmptWRLBLfDiRkBhOm7uueqaj5QY/AtV9hb
UHBaHo/1quja/sz8DU2XPW3reDymrjtaRs9gtVASFD0O7ttkIIW3N9EVL7zOSprL
rwCQcMsQ8XG5860GXCSsYQydc7rCCGrjiHpOueD83aEq8NZe52bAEiNfaH7+B1hN
Qa0jlPJU5+BKfeMU4fn8PL2cz11YL9t9jDRfD183fP0rM0fpK3RfuOO98+vqnHLk
4DJxYZaIU0bhpDxnsk5RTqcyMAjupyMcepDIKGKGpuLNo6tqMTrc0zEoKOHk/mNI
G/OPIuOL/ItpGtrIgssOkEFMSl2DckwjjdcqhIr+Jrn6SQKV6Vk50OFLn2VTXifN
kzemypRBUbUKMu/KPmRH8DRFPex2kgFlvmH/I55cxiQIo/lw2I03wIF7p/j6pmHG
2qWBRbYhLD/Fj1FrF5Sgel9DomdjtRsCV7zC2A7zG6ZxKZ/PfY73SOmnt28oCN41
fOohFEunWRQ++8/+XuisLOozwJDQHLo4w+G+wsAJrNiRXlOE3+r8qOy0IZeqvDqP
BkvRLTrZwoHHlWvNUC+JMrknHv17nbmmsQCV3WLDt/YsGbhoxNoUBaU1xDr/KQs3
HBeztqpCCEXSBKph4IXMcOHjIxtXsVlHBuh/Ikup28tTAwbZW4HT3baDmP2cGX3K
wD52BtR38md1TPoQNZL3mxQbkL8HQ3wH29HpSaRloe7ajjZipB3SQLY/1pCa1ZRj
Fp8nLBHPa85wLQK2XqOZRqQGKEKe+1w7QyUdt7rsJICoLBsREzY61Qa+WFjgJ5ec
0PB4f6GOEnIN9g9HJ0sBJHUlrGFddNme/0QLik1imBhx/24OwOrCIb6LiK8q6iLj
fE4Jq+CGaWmXeUuXNaipx1q+zfr01Zp9pkA9VUm3JtTPNqtX7R/K0Sk1F3H9Wldo
zdUANVQcnGiaAR12aW4OJ0XAbEljgs4fFe7FvCpYY3YKQ3Ls9EWe3KG+1Y03wZ3B
CFr8qz+aKyGj2Kk5+erfErDjve4FUh9tnQPXTIUt+3CqDchMoMnwYgOrcyeAG3YW
InlRrwSAQ5ET5N9Sy4wcmVCudz4d2ukQRdvdCJkIK1cyZeZPLahCfSzyfoTcEscb
AnjnAscf+8T1CD+Dxw2PfP1yO1DH/OQ+T4bLqZNAqltAcEk3lb7kw5V8x9hawxpR
L+GkuLHzhOSyhNlGJuAOhCAtatF4qP/KRAQf/LoekAXkE0Zz2Yo1Ki0+2WTowvcV
CcCSb6t+h9yLEw28a3CzDbPhCtIvhJR9a9hRn3eZrbSH/GQ5zzfs6Suhi/1oDgyW
7IuWLS5a9lGQ11i0NaUC0K7WJvm5VaraToWdpBEJZJfiAcZr/Q7NxxZbT+5CkCyX
FUeoXac5ixsQVaPzLEev84z09IT7AamqBGPHyBYgvwkgGReXxhdeuipt4GQHKMU5
XKUyIxIgM34C7thgRsE+nEk9WkPDZ7lJPw4sP0/q6d7w6JBU6xDmhOKBEVCPM6MQ
vcK40+kAat/L1SFsP2ZP2x27sGnU+CLQy9LYD/5S+oX5uDcqGtfNtt5h5T/HOn2x
h/ADoDBm2YfZDPkdKYw6z73aidlF/y4u7THEPEfV/hafgl8fs0M1XAq+BxcplK6T
qJmtYM0/k+jVPgO1h6saMp2p6fnARRameYtGo498Xh8ev0fhmIFgs2MqeFKAZBTF
CegpK7zvXKCadOA5dAifuEF8gkBx3hoBnh7ZwzsHKPZR8g60GJd4HRosCQDjeEKu
0aQV9xi3sRcSJMcatyetlQSCeMFARcVnMcgjQpQhmA0jEvpAbDEfxHzl8iKUDqAl
TNnkfY6zzH4Y2L+HEaCf8q5gfnPKspERdAJV+6CZa3jyhtyqgeJ8CP3UQrvlHhzx
Ti8Xypi98GYpv8amZdCXt8BWDaY8aLS/eF8CadmNp2HuhQEOEXLiH33hII/dy2V2
FKqT9yxU5Fz+IC2zB5WcS0O/CxRahR3/uEdoWP73b1iD4dDMCLBwe49+F90TAgHQ
X6dge1V46MQLL4gY7AJ+xMgLPQbmaVnzGkgJba8PfrRjLgPsNbB+D13IK0to+bVV
XW1W7g5DcUIKREOZm1WreKT1aGLjosozd+EPM+UFVfIHwC6ZOGgH47zDh6dda5Hx
Z397kn05mEAYoxl/JoXYY93UeAv/R+1/cUyqbD2hCjsLDKVvvrcQjJFeljHfAlxQ
5FeJBBRY0xHMOE7ksNhzZCM+YN6oSFhsCnXDiLWHOuS/ZrcOq6/aMJjVZhpCGRLM
aFAhPtTW9/1J48r8d3r+8k3OF9gOT9Ugq/wRxSphjhc7PYM1MGNH23N+WeWudIGI
/DFSGx9Q2kzTmZr8PNFyAjIfiVyQzQgt1wClJ/rSKibD0VdWwodXDW1ZwcCR4Ac8
tjeBDWECQSWgKIL1sB4s83/kkmmXSOnOqF2iJWvYF551kkqxs1RtLuzezV4UZzOV
Ld/1Xulrr/NL+wMxvpJ6MKRbfq8N5alIh6T0knoEtnf173mU19ldMAwU3UxwVH7E
IV825rpjRNU/Q/KEMWWOGUMWUYJu/3BR8gGpnqM8MvHKJoJjgcXsBpyWRTDkJORD
SqlbfKUHw6wegxFzFcCl/pefjRaefTteVc6SHTwXRsDoshIlUC05fwr4whXDlZSB
+AGa4jypvdMEGcT1fVfQS3DDE01huov4fciTMQwMEWguVogPYS8qHibwp6FC3DXh
/cYXZyiYgLUlrQ5XfrPREOhawTEw2vxxaDfnd706r/ZPjcxVxRPiHvJlMv4PAvep
uoIwMADtmFvDbMjXLYjrTRzbAbPacXIc8pR8GmCxRNC2RgXuP6S+kZ5TMYpU+V3d
+oiRn6hUQ1gwOdK96vSKLBw5ip6vUZH8qEcRw1RsT+k/ewIsChXt8P4OPMz+JrqC
PHjKSAjCy1bO5jGQaideXMVkUpFlESCQTKzOcCXreyC08FuOKV7TTQkKuZV0PHpb
NSpc18MSXT712V9qB5fBeuOTm8yPfh2sPdvIbwiK2uhLZ1VNr/epbTxclDvLz+zV
dPiepQqMaET2WId5YnI/DLyfl/BqrivpaFEPGDF6qM6Jpt9fnMqxrOvvefo49Cv1
jv6G6vkjYZ3PkjIS2FxAkL5XXkFpT/uGmQVMabMoI6ZvN3iiSB7XOVMy5OZ8H4Z9
gJVKUaqoDdDgDDl12Hr10/RzV8nB0Q4oV8vCvxJ9WEf/dbdbqRrZI+NuAINZnKcU
UsANA0rV6pHjxNdryRiLr6EhOVmfM2sWIdkByIR+eygh/a/jwRA4rVXgJ6l7C6Vg
zWv2AS/J4mUwWTuAEIMx6rpI+5GnQccF21uGBi4ST7VE31qeQNc1ihVcQuE2xrpz
HzMUEIbDZJmd02Nb5L/zu0VUkSsovRtiGMQwlb0THFsG0V4Hge3Cx3nnltsfDuo1
lEFxNXnyHxXAYWGFQyH5T5YbixpfZsyNl1gcMAarJpWphSxVaPH2T1vo6LPOuAfS
9LllSebzjAzEiyeTrqdH52GagZkLRe5BCEabQru8tECpr8TBA0/2Dng2HGEEr9wg
sRvgU9sHRX6+r5PcxJjNZuFNpiqyd6RV6OhgHo45rzGaFN9XPTAOAx9dxMFp1boz
feWbHzDZIyfHS9f+9UK3xc0HebK1X7oj5R/hT/Gll0JxMI0akCkX/9gqq+8wh/Lw
VIA36VfFcPkYZDv4egdwI36vkx7RO5jMN4btOz2zMEZFR5Oa1NQJpKWFhmDWPQ8K
GIzF1rhD+NvDPlQkX2oCWGZdobszjRr8XtMiJjOXudyMCzXAS6DBW/a1GMiq8RCr
X6ChFoFXSUaRoJ6r8EQ2FGLLPcuoWo6SiqgRxQXuGAVFf+f7dPKey2TzXi1LMQc+
PEvvt4Ge6UTFuh6b9UBpvsdogqTcUqkn2QTrw1Hfje8c/QJ8VokPqZMUaQ2fkBAA
JRqoXm7Jgdo979ACyMQkCZbv3/tBioyiGcLYexVy42G0w/lTngs10YVSCQs9E/zm
w+pc9PiqgdXasjtICG5wukCRYZyYUrT8Iq6FYang9DYwb+trXxVPNEPdMwWsetRW
Qa6iuZPrDTKaOPbcXirkJJyGlbRA7pmwvI3Brz9qjsD7BxLVWc4mhDcA1j0xmXaj
88dONE0wgbx+pPuX5XP/OaC57Rk8GfInbwWvVp9n9OpSJrQAxaR9ObTaDUUMN/qr
MyumIm5yJMt3F2+UlbaLTmEAi/3q3L2y7ouNLCNk/VibeJLPpPzNXQB695R+6136
FM5Y48FL/awixnzJ0Tx3E8RFxxP+BeABhGi5REz7DTspPwMNubeLsErSZMMMDb3C
fDjCoyec0k7i2gWJJL44av5sIrNKVPu3AT7oiKiab8KED2U6AAql9nUp6O0d1U4n
scTvP+7b1tN5RD0+knlEnnJcOqMP5Zn68Jw7BqcwhQq2PFaOksvXNmwATcgaYbvq
eB+sp41JAXJ20H3wj67aCMd/6xAuNPs8dNSDyLdTz97UO5rbwVpc6uNmnybb9MKM
XIE/sd/ZhJ8n5e6MkUxF+vvbVSVERZTecmmI/Jb2pEryjSdgWrfiA2aWKKNFvM+c
76FfTl2jMBWpNvnifsd+7Df7PZusEc9Bozb8ZvLWkRNqhhYSJcABDdy3l1+9md9x
ZUAbRZWH+vFO7X1j1HuXIBXh1GwVO+adLyunBtDt+wIiQzMwa0ekmykmLaT9zHMB
SnbSGVGNNJDVj4zSW9LlmaeFwDCZ+uJ3ZcOS2yf40E/+7LQirNIXBXnLdL2P5oYL
BRSsAoKUlgEp+ZgnaIsgCkCkcYnoyRkKbCAOu+EY5b/BRYo51WEyVrv3Epq8PUNI
UejqQBGsOAPhl9QZbFJB6Bk+nt5wQlvRPI4OJp9a5wMccaLfqhW5il1uy0M+f2Q8
+L44OEiWaK+Jit1yRt+rT+ADihtqhNJxpxMQWrzvHitoVFKfyT+Qi+nFHfFazyq7
6v1lHYglrXno8xGpvuoDLaR3L2aujm+MMxACNGbi+ggpGkhdqUG6a2/eFnbTf3N5
s9yELRgVaoV4paHopPv1Vwo0T8pAo3JovFI84OP8yAdZUWHiug8gd66NIfU0KdQR
AjssjB9HoJTTheiaiY7DfQ+YGqmIj8gzldBosHleI2Nv2y6NLYw63GUGMTVoQdwm
bnIotD8pWsUNdeddynpRXX8qpCyBDVTPLH7/+thCAZ3oOxuDD3mT/4L+OQt0+EMI
EdO4ux77SJCO4R2zd8WzqFbtwsUhFke4VpDb3lyFL4tFH9NLVxRlmqA3k/gOt0/Q
Rw2rNQ4MtDbZIm9j0gBAhTs+ygExJgse8I36kv8OECREDwadaUfsYCcqqTPlZ8UD
nmuNDJv9mhLpu5OQrWm0i91XP2xIxawObv3whrX3zcKiaJvORC3DWZnzuRlT9gg+
6FKAwOOYrl4BvEGE/SIDiZQAX6ck32J/F70IfOSNsMs0V4SA+ny9b96bwYP6qMf/
8FNfCElA6lUyoWefPSWpIFNxitS5GRvk+az4qZHvgdHG4G2YQ+odRy3SE0MCVTdE
GNvEl3mMxAJT8dlztgVNQI1S1j3MsdbPjuObAkSmonW9oEO1zl+HPRm8PV5NX2ZP
4XQp4qzu4Bpem+jxEYvtTdCxLJNvuA9WFa6vrmcQO/GU7tv5CLCitAMD88k84xUK
2xiuLoHmY5I4Oanb/0VGDF4La3XYmc31LQJ6C5pccsc3UErZiohzz7aw2QOprJgN
OrAOr9EAhM4CfCCIDJS6Um3aBXX4jxKXLyFOCQjEssEg6y/jOxk0K4RctLrpp5Ti
0Ur3WRGj2sF/+SK5JdbMDzIh2iiWp17dhDTnAlZhntOnGYdHGEWEETQvd7ecsNoi
HO1AZZyS+QhL0MdfDajs6vyKe5vL/KBuMWS3M9UTsnFtW+g8T0hhBazhBmqoITID
fKn5QuLyRSL1/s79l/GpL70mCnvYmMlpb8TYVv9fgUuyZUtMhF/UyPAp2hnqJB0e
dicvsZcfTvTV8uZndHAgCSiqn3Jy75esGW76mhhYGt1F0A4BnRTeQNM+/dNAp/gX
sYaOIYkxAuPtkv4CHNNIBuXR3vbzZwy/KHFYuHDAtZRnruP6b9pf7P5LWl+5J4h9
lyHvHCgCSX71YmC8jS2yMA1LRPdvwhwCzAR5/nARS0zTrfDERpbzlZMcszUSxQ5J
AJfCYEoc+2F/aqh/trG20zkFE+zsYRPc8tDQrQaKG+jzk2S1W4oIBelvzWBLHTu5
8yCjUCcyWhXw6cIhGm4wRviDD/9l3tuYT/gvNbq80UbRybG4yNGDnNfeEdrMikb0
8O3eoxOZCoKtL78hnNOucKfdyffs9h0X4EgFntST/GY6nzki4KYoGPr/nCjfL36h
uDlZV6ibKUJxmVeEwmw/VjB0fyQ7FcpDK/B9XrYKKN5F4TU04oOhvxa3/Xa9LBBm
ScLytei/LWIWbxLnCmf7WEYKHu1w1xh7S8XhvsSItVFRiKqPvnZ2JSGhePPR/xCU
M5vfo47CaJgLHzQSvzX+PgbPVWvoh2cMn0xLTGnsip5Paa7sh9WHaoyjKAHQvPg7
keRZ6mnIww8TiPjM0FTr1txtJX9ngRtqbEX4ZeeNHj5pWQB1d2F6fgUewL11nQ0V
J06n/EKq6Do7W71Li78rg2nsGH891zuLUcHoTt/cgv6EsUUcrRPgNPXUGXLYQNup
w3EfvQkzBym1hM2xxXrQ027Y8OGOuTwhVfw9nLPjcfQYXo3/G1sfptp/iu2CrAoX
FgDQ7iszZ7yRNiW5cuDIjl0k3mm5GmVO54LbwLzJlrW9rdJvbarDEiD88j5qsbfF
0cV91T4FMr+yll3GCSCStdoS9qk/IlN21rYS08D0KHJBpxRPUq0YiToY0n3ww7H0
F270iU/SHD7mglr7MOZ3Do8G73zTLTdGNJSqgVavUYiUQKpVL8uArVtk7bcpHVoL
kd0Bhi56gnHm7sehCuMOSl0fwd7VTUb/QMWvmqFH/2zztul/F+qoKzJ39rygllro
ryDd6L7tlSHjNv2AQAV72MO9cX01IjjByLQTcZffsqrVuT/IsA+A1zSg7DvlrvzI
NxPs5aet4WyZmrfK1st6pwIbgDa2/RMx8CMZvbXFHmhI5h4u67IIpIDJzvnsEeMZ
iJhuyfD+V52RyYLND6wUYEIYIcxJ6sSK+mlojKRVDOncd8jhSLqXRNeIYQCSM8hK
HKE80LJ8XuJ21PKEhYIoH60LqXXKcvW0V7GJBGJsVTZOakKT6E5f8UdWA228vB06
bn85isQSfMNLI4d4RcBLlZHw97j2WBZAV7Gp8OT4gVhVfxc6okq+YRK9OaP3ZFAh
7tRJua163z1qbGz8YQ0KoNQcWC3L+kRTKxEZj9bskPcZvJvxTesX87mUqV+JdxrP
houMkQMt5Ir57ejz57fcGaMFNCtvsc2Bq+oRKfTlVtSTXkBeuUMeHWAr1JBPtup3
VvBWRFkthDyce7Gfgol88yyHUNoOVJpD74yBYxld4/hjzbOZ6whwSqNMbg4do0IB
i5DB51HplNvpqSdqVfCysfE+fJ5x5f5QgIyVMZzJ2ex8KJpimLdSY6Ms0ezoSnq/
nv29hEKMATG4/94/wTJNo+HbgAttfLFKpTcSUQQp4zmkXzTW5GYF2whmDoEf5pgA
kwFL5fiJoIVPhYLpyqYiX7d0kLhr5ej3RAEzkfPvbITKe/BPeordmITrWngx+xEw
CdzZxXenuwzCM7BaHWLnO8LFq6ISqZr+6JP9D8fwhJN2LMjfeFjiA3y5hK4NGJuh
kuj71YCXd1LeTy0AFNxkUMPwmgShK1DIkYF8T7Gy5j7hgyFbRTvsPP2Q0aKcneWs
PMAbnrUalSPcacrAM0HtowMIGxWBzWZIPVG/K8sgopZrF8y5znUh8mJQxOug5OC8
YF97volJ4Uoaq/7xBsMZwLJIxW8WhAcH6Syuw51MDBTIeLUb2J3kDsz8JJPGEBtE
LBnEybLJLhdqeIgE8vLW03KBZUf+eJr+2Mn24P6K2M8Ft4kmKGaOInFVG7WrO7xi
+QcCnuGK61o2RUUzhhTB0d3AwqnN0Vd0IBIo0/tdW48WxiLwIo81yDLil3vqM8Uw
RS2g6fG4mAsZQWooSqex35qnOemW3qCpCsULQ+JA0l3SkDdG3vl7QPnIxAKqbZJG
llASHowC+Quy0oT8yS1RFQ9TcGuhLNuR/M3/lYd+gPisAh3OyCcVI7C912sj/DPz
UkR9kscxnjARvIRIGtdDCLeJ8KcpDxFUqrGjWEpMQH/lYV6k0Q1UQklsCI5vFK5k
O/dXL9aA/wGRNRQZeHamcAHNas9+CSrm1mHubJgPDTJ21TFvkQ7Y/HwJfXvpccs9
j/DRFuEr0G87aPr561oLXzrBnI7qrx3a4rEMg79R3GuJWf7ydbeeUJ9hAV+OeTH+
h8ip/I10wVPwLnL43wdOChoBMe9Y9BLGPy6UFsoiGooULxwE+v+KWmvZbECYg0le
bbjqSo6sVq/Dh9pbCw9PSlLK35frJrPJ73Na1S5pOBzEyEiFctk4jXfFnuis4w9F
0d6GcN2U7vPQMXtwPRhzkhBEl8jQX3S5e4IBv0lqqbTEHlOSkQOHb+z+d8lmrUpp
xFvrq+uYzybkGJJx3cEUxuIu7WnNSV0/cyRGTkoQrogItIrVfDmoK9Pgfvc9OhDE
CtURq72w3pqIKdkOxigg0g5NEEV+jKB53x0hmD7x+/kDO8DDBEAoG1QZJd7G8KTn
p9QZw3S6DkrxWxvUh4rolUQmdV6F7Z6o5rTD66EMkmNv7iK5f0rgeWGnOHnzsB11
3HWq+rh6T5qoT0iaKaSZyflNY6ICODGjBOej5dr4icBEHLTC79Nh0vQSq6BURkXE
EabPohmp1i2/n9DZ8zTDNtqpZkMKN4chppeagCV52Jnd961JEmJ4TmhoW5dAQW+P
TmQjRyuGsG2dB/SlNVBFAWFEcZNcTZacf0g4ldXmDNPfXHabuiA75p06+L6/Cnqe
DyGeZqlJ+ZVQlqJqfSQVYLdb6KVvWf9BAkM4IAT6bOiXMU5V1sAth1tph36hEIIP
jrxLHXET2/8UmQjoX6e5W5ExAMZQreE1Dzk8r5wrO921EKUna84oi6/P5yMuL2AB
KWCpBb1ut0FbBIWK1/poBXAvxCxCQcjj9iYlWdAN0ymADide8ttkGjWmBfOZRiI8
4XHnRyqEW+K3sE1KhaOwomzt1WA344W44u9adlg7LygqSOCISWzhT6eAF6ivH8hZ
2vH5krGIAW7hbrkv+MIgJ3Ia2XagdMOGStcyTdRG40O7K3HbY3W8SU0Kj+95ITP8
d8+Fq7IysfGHu8ne9gmUnOavjR8PDnt1eyXZImYse4yTKmAiVYkLG0wvO+ewyDV3
8Nj96lrIaipN5PV1mMTKCSuwkv5WDnFFRUxWncUYq3j2zXFve7+H2Tb/SWur625H
pcKugAVnC92mJV8X1e+ZEg/I8rMl9c2LwPZDU96sKNxkXzx9qpKHT7dINaGT8nZ5
lhytF9dtcyMuszV/FjQEOJvB9f5vq123714pGsz2eF8XpxJzv7VqAT/DT3HXuYNn
bSF0VTXm++kxjYgs6th62HsBBE2OXvqMznyCAUEl7p9keif1BaRGQnj2oym0XwUI
T/Z70Dw4p45E6wc1XEqqAhP0nYu0J9HXPsRh1qE94Wvz7iVoJ3ujnTp5tI99CGTI
eO0HtUoMYiF3DZdvzVIWbqtONt5XYEhqfuVlxJ4YOjAUcJbB1tSAef39tndt8wXF
eVeJUoiWq9958uuYLV8EUwwItOl+RyzfptjAqbC80VIuyTbAjtEeHZuDialBgB1+
3GRUMNZ0P4m+Hway8C9HCX3nYpqbvLj38x+3VojO2HdTjpOabDqjaB4BrYL1aukb
Up4XajJ/GZOpv7uXSHCvv9IS5nu/3i8IfKwnT+vUhVP0VVYtgQb9Mf6rF9W7TI0L
GqH2wvRSBN7t6l3ErgBYcwy5RbNQ8fRxw+FDBmmaTOctTni4VgE3mQBQLdaxoXOG
XlrICfUZpcmubMnUPPkEdVkPjpHB0hcqBSleOKG4qkT1HRbBVaI0iceIgd6K2ZSU
fO5fV/n3MwFp7q5A1LkrUuGWTHPuD88M+fxqGkXFggDBo/KvVHGBwDgIDRXdhA3K
KFxdY3PWDPx3cLFq7D6CBealZ9Ubde3hPctT80eGsy0ps9u9ZzSc3HDw9kToxTeP
gh7LqnCgr2mpI7d/nSWR/SgQSBPyAs8OD/oPZrzvGJwuEOvi/wdGoPKKaGATJg6t
JwK2OAI/18mnOk3q/AhFQ8SUlpLRNqeCFsb0kJ+l4vmWOZhxWSUuEO1/otgpot8A
eqArpY0qwNEupS5jYL5RWLs1FDD+18Yaf/OMsBAHEfeHh1TwqJDCSyg57H3w9QdQ
HNnsmcemuyxBsU89a2jHu6h8zit66Gs1l83AL98GTXWNrrF6TA+J5O9aTarABs/I
LNVg7aTG4Qds31Bx4BoQ1Uc3jjk+oQiyu2ti43gQenA7s2iDN3oWPLbhgklUk3QV
XTh6UkLpKFQDZufgZqjVXjV7lqPtUpqeoih1+h75YNGUnEyMtECdOy8UlUhlyqUc
2Cda0Isr89w1xfBle2WKWi1CyOFc6TImX8y13YTKxi7zo4YdX8bH2pOVDobfVLPy
/LGpFEZQVcLbY26h3/ZDYG7C5c/ypVr3TFgUyxWmaaae1M4hZdog/sdoIFVLVUxG
nh/+VlaffVGVZ/bgSMAwWnGUHPxbkhlyjVdcG7MJOgOOJV83QU4moQQc2LgU2EQo
jGdNIy8e9mxyHBqQLDXmv+9xJgNPY/UtuNg6PnyKDgYvpWNIQqy2X4XnOfb+4jmW
mU3Alq4+imXD2pqbKwbIxE8H7PMCDE62OqLfWpUfR2HVzn5hPb/YuYSDNwGV5kVJ
/pxATYplxETthnOBl3tv7DotGRilrhRjRxCyWnG9SHoEOgS8l9izwC/x0N2CHqaB
AUsNod/UrO5zY1C2Vr+UidgDZ1hfyU+T1kuCiBAmqlcM1H+qLRW5lO+2ti+9cU3+
v+GxthTd4ZC2sbqZ/qDJZ19yO+nu6cLxJPFcTcqQptzSfQs4uUCZTUfup9ETGLFX
QdFaLPTId+X00qrIVeGkN3dCBkhtZY34yyiEU94zDALVjtP9tDuqoIUvdFNwYhY1
GVS4ZSVT4hNLqV2jZbLbsgwPNU3OPSyU9AZisMDfQzezVEYieceT7n4OKsFge2mP
AUw2mM0xSjXQSaC8eMJcEvoTSuP8wdz080uy3PvuSXk4SJeYjUXM+K2PZ+S395GN
aGeIuj3TgrpXiKBVbCNsb2FqLoNmIWq3qPFmLsY9GDwg+BoKI4kHv3i6wwRxOqgX
xSU/Vb4yaOvsy0/qQ78fSUcSLzGbfBdst/LYGlKPsvrBWz1n4cXmjxecy7l2YohL
4HplgSw9XthJgz6tzrHV8pAxmxokzH+oXldLrBCtbh9wvAzSwg5bSndfs9ctIkIL
CxsQib7v0fAuTZpqMGQttoH2aYRwmGjtOpj0NMokEPe5gim4CVqGOLqgZOo1HIIA
MBmgP33+krPNmQpuKJlpad83APJ6I+utekucEigDjfqXKPFC5W8c2WqukJR+S5Ch
nbAkV8uMNpl9mKPIuL9xTaqs459NT+RziOcIa/OWqnfWF+2qo/2nVTRwoSutSKLV
qUqwSDiC3UAJmZVAWlbTSbgis/qXBjcy+D4ujyzC0q1BmZ0ceDpBGZJlDMhzNZb2
3G6S2nC38CJR4ynRF/kIe2cumFG8njxiNO5T5Es4p/33fVIgjevy7vzD85fQH1W3
cFknrAqUzGrAWZUkfCRX+VVaHS/mtFBCOSONNl4igTRXGkdLNA3DMqq8Y09zCQQW
6Fh3g6vly9LjnwYKmXsQGGq8CdQpE2QeOIYlapLS2/AVoxXkoZeSrlS0bVPQiKTO
74gmRm5S7OqAxfMf8laN9sEeWiaKLdp6J34t+TfUEm502S5eoixzZl5cFFbt5oSf
ZaWOup31Q7PJ9E/4WQWp0Gy4fl33K2GO91H9Qp5gL/dJgRf037SaVrnbckFSVLOR
wFRUssHspmPnlm8+EmJa4DwgUPKkUbnhrHOfwftKp6ZfR9AkXUmnOHABPskPSJqc
2Hua26PMRjvce0fR+flpq+ztRd1JWqShQ2/zdxXX+AW/NHog9Ndm4JcEt6rM+Lwr
AkKUQlAXb6m1cRspTHFNNJCZiMI1fKsaLjC5iMLYgdgUZw6jlFrZqPBaXojsr7sp
1HeJXuzvUgddIudVHNzsL/wf6jRE3RKLVOwQudV5aYSlPdxGpAHcUOStbtcR0Ba9
/z2rd7WxcA1kw+z7OVsJvb8/DEdkEWc1v+pdhtw93RqfgEX+NqqoCS4wP4vbvz9o
vpok1e/lBXbky9eH1JwObGq4LpB9KDdKRx2Aav5q4lu6DU+Jf69pL6oLaAViwDNP
lf6nuF5+Hmp/rxEcHT6Iq3Qjh2ERCaZM3eZ9BEkYbGiAyKd8CNIPw3InHQKbyI6g
4awgvEOQMPfwId2cGtAPspvqTHJOAM255WRnFq3EVsScoxt1LhwVC/qsjSZuStNr
dqUf89Y0fXS5V2UDR5nBWl/ARHN/0/r8mgoOSuDrHipOd/kaO3H6pAjok2jiNfzv
eHiEvaefR2Gx9lj0QAiRBQVcYgDkJe6bV1VncOv6kELSiOh4ovl9nKo+YrFybtAD
AbEBaerylGwgxA933CbYyu9M0YrtaJjb4kvRCrn9Ys3V+RC3TApmMrR5omqcFmB4
onY/u61U++GcqZVJyCeGO8yEOx6b6FZOzkWXlWL+DRFKXwdPp1iRXMkxCW8S54sG
ahMxJNDOVibSewGzcBu8yxV7Uj9SQJ0pYl75OOqHUc4PPz0awL+2BM7jgfzFlfuG
L+6KwEG0KWvWNLeKg/alFb0AhDiQsTO5VSSYfvfHWalohQAEtFHxF23OZf2Z84Sq
nC+cA4lQixT+K6+jUzB/LSp0zkvOxe+j0IeZNYP1BBCRJOI/CguO+1CCP+gcpPW4
nRY5z54SreGJ3XqEbd1NO7ch2m0ta2cFWT/OU8T/Jv5nSr2BQ1x3KKOqq8wzQRDm
O7wjcNDstJe+4yjwetaGyJOq22OnfxzQ8KTjGomJsuPGw0KnzD+8cCkQz06E4F9n
f+y8LNSppHdYt8kU2GM0RJWDJzRlxKcgYAO8DXEf5jM3FRTp06iCrg/5X81rFTrw
xn68zg13VANBzoXYxTWS+91oM4+LmmK3l/rFZzI0XAIjpNru14KJAVbzD6hBVgfC
twn1iA25lwKKzNSKuoiuOhXNl0mxWnEzJW5i4emor98mttG1XmGZrjhWWO5kNQmC
MjerI/zt+uQ4f3wf7Jzy1AVuXDSVpktvuoz46tKZe62S6bTgm7JshGSuU//ezCsp
InPWWQdGlTVMmTD45yeK69S5qLX5eUwPYc2XNx/IZHQM30dRxwPG0wi/8hUWexJ/
V0V8F6y0XzAiEL3+/xfk6mmwFMosI+Gs7wajmtjuvf5r64N0nb3VndprDMdZdGZb
or9CR+mkKD2tjgZUtEETOUcHExymHljAnf2EH09JlFD9fiBPSnB3VxmdI1KXAwEI
nvzPPI6H3HAUIv/T3aRyFK7tgoJHx6b16ElJC0ihu21yT6xay2T25I6QNIP2hfQ1
+GIGwKqVeW//3jGXgAoDqkZJq+0KouAsXb5OLXts7CAXY3ClYsrTp6nMdbF/+uEa
OzzRQsQA70wRpThG4JOuJM3CQjLSpgZR1z0rvbNGPMWNOED0GM5mVvIEv4A0WyRj
RUC+HD/XO+hNCywo4nA8puH842cWOWTbBeVXsfu2R/3kc+RCk2iwPJZWn3f3YcL7
wNkhbTqYrYctRA2rSmHMtLQ/LScSsYOo0nEMfu0bwaCnVp7MG8S9JwPp8p+r38K5
VUeSV0sh3Vh1HKyqdi8hlChaiddwk6gSSgAdTIWmAl2CLpfuqfrnn22E/EI7+pK3
f7rjCNtjT8ixgGOGuxSqg2jx+rqQkbhzeZyADvAxHIqwzbeabDQ4pHEYkUswgXOm
kPkL701h2gKKxCJMhaXIdhZy5pFd3sGAKtKx7di6IypYrxlgB/VD8VHli6ZFcMk7
SNFbUouHfTJbb/gMEMdQfJGSRm1rfQ/t3XCL2jgNfHNpb+L/FwY5MdUwXvAbC8QQ
f4OeZAKEs7JYEqqFUYEvSUHnmS2EKWWXmZEyeU31hn8iZrpmbzuvbd5XkyB6I471
+NXFwDbvfarIlVVAwLSrMRE4d3UhAvIZyLMJ7NW4TXfjkH1tZ0XkeiWtFe7a1SKZ
We7Eciw7+SXP9geHQ7pAkoe5R2LWpk0w4pPSnkEs1YOBZuXVNkKpm+Ks17eAOQl7
pCRykpYqh2U5XPWfai0kRn9qcK4lVzqmFjx/65DxV5hTaukMyqlm/IPvTwT0z27U
eGyY9Rw3uamjuGKqsAIgdmmMxOsyvTrRcEl03RkteybqG9JEkr0X6wdbYtGDHSxh
W/h9Ib2JbWaenVXAXY+kvxgpKYm2X5ePyVZptqgOechTRLf+PJ70jmDmFrBxM8AC
XVWkbQa+QeOfMrs3pJ/4Z/197gJun/HIbDeJyi7Z+SRDezGT4GfOEiwuOZvoi5Ln
mYYRxZtSOYBNnu3RlMC3HDsbkHTGrKDeS7bbcJIoT22vkZ/serSpVH6xEReR+J+k
CGqJWrhviaLEdLe4z2lrbL6zUNGPxqKP69pVXC+y50K/JpBy90Lflx7t0ehqb358
98JuCYhL21s3jZM+azWEob2YrLGklFGyijtwfY5bSyu47cHb1R4yg83a4Q+AePZK
Q6Qds/UGXQJOyBZtsUgIj5sYhxLAB5uqY1C0Jdk6oJXhixRVnqUIJ/71HYc6AScR
UH+DSc/xKAigtogxh9zY1poAk+8GfEJXfP4cNdnm6d3QXZM7NzNIzPxTRdOUVa+B
TVoWQmP+McZ1fZ1Z2bDFk2yMdq1jE1dRSWdsicYbzinAODksF+VtPQO/sBuTYGQh
AANydV9bwJfAWJhJd0erLEmrEyaLpbeZAqPAU8lzs4i9AbbKVtpsmV/IEBZAusxV
gcMSLe+UtjIIxXjbOBTV+oDTLCC0eRCw0yu1cwrJC4VypicKqAsTZrpbwIqm8iXX
/3TgpZSnVfdKRNbbDE/jVYQqqvoeOY+NSu3ZmxMME8nVWDg7Be5dH10nqKuI97Fg
NYR09uBwEyTVkdQtrj2KAIi7RQmaM00oMtZ7PvKBjmxot/cvfUDVeQ4hyBrFoDd1
IAHHsFA42smlXiw84+hp6gW0HUExt8LWlLMFSftXNhBIiM2bNQo+oV89HGNWW8wE
6qE2ykeMqejCVFPUDNOBEzMe93GuCrAL2ZYXBcGtsrH5VQJzM+C+WPadvzJpncjC
KDV3++OsHTdds6NbwMhnbazF9foC1TW6dxVKy5udRbZefCxz7VnSl19Dg3p1omrH
9zUGZQYelgBFvRpTBcedNRTxCTG2FOVBdt+Afkw9ruZie71zmolOM8D0H95ypoOu
oKMGEv+BsldTLLjsJuUs9wUUiaEP18iMvm2PKcyJLxZ0V9SdLL75Xb/NmqF6PwlP
MT0dGH/NReti2/MjJ09HnClmDs5fwMU/cA9qTmgCVlaSUIzahvaA8UQgNcJCiBlK
BHwhSIZ+SedyOu3psqGuuzFDlq6H7eUx6Pak6TdNRsqsMjPVi+OQhYhxg+KNg08i
jduyKmmWR+OybhvtFEfXi9ydsNkMS1PmGQX7PhB4ZS6rY6dD+nwt9fTzLjkkKm2b
KcpkU+P9b5Cgy20DM0Z2vBpw/M0dWy4xlwsohaACU2MCYd7X8enNEcnXgpM4QTuc
Kc7UcWGEx//YJ7ncbPJFOUuy1M25DXciAgxRdfYchuQv1e6R+DNRAuvUTswGJqLz
4CO4kHXLRvCqUqKlMcRS8vb2P/b/gJxanMvvqEYWPSj16ycLZ1fs017bXjnwWw39
bGIGQUyZqxOAqgFhQdfGj3Fwc0l+iY8SaGpKDS9/ohyCE5KY8dzrc4Lj7vo5X0Ub
3pRFpP3hZZyU5JgRvG2YkNSz7BXfEZhNyOrfseFh9R/xXsRaxWXRR8zdmBWF6UBh
IPP23GsEPbT6nglhhlDpkJNLo8lQPQr9A4z6ueudZaabNf5wQrapIIYKMtCI/0Zs
ySX3zxFX4OZgZIdZSiC6ElTNFPVy6KW0O3zJadSQhcGt8w17sV6sz8XvA76oTgsL
5hS0h3C2lBx9FZH773jpVe9PWj0NjUxgDsZq+wtCO3mK24br//3UneSpWyxJYpyi
QzwhuoRa+81TXMYD4vYqj76g0hy4PNl/rTQOgLR5NVXEhW7j/jB6aGSOdVxG0X5y
OHAXCeLg5sqQo+Cip/EXkkSPdlYiShVvoYx6qasp7LUWSfd4VdCIP351Hw2V02Lk
GC7xgZX/wqvBVejGLxdzoQep1UA3zyXutgpvHM5rgvYGrQ9JY8E/tPIv0LCoHuhD
lZTFJGz3sELO6H8JHh+HYya1zG+RHURGvPBIPBrL/ixD+lHVUeevF+ZfeJqMY+Hf
SKyZ9MfZJjYk8kTm8tGv+Ua74pcy7UrKkhRE3orYf2Gm5NQ8HZhghtoiehhdYAdT
2Qreu1AwD6VHGTKloef70b/lGazjZqrnAYWFPgxGcfnEq3Go3LYKU2qDb7P3xFsu
DvtNm6ApMzlcXXVZFw0p4q2qU8w5juojxqiwwySdyP3bdpX3PyJZNLVe2NWVOlSO
gSwCHjyVElX2mEfHdp0Vcphl4Sp7B5TTg3latjnNZ9AbcITRcEf6D0TwIiM8v9xK
AWqZp+8bT9MBBeeDPIais1or6E8O4kTq1YT4qsP5T94Y+2ZhHbXPGn2Bp7/4jVFg
q7qMtFsRtjrkurZ8qZ4LuqmFRERn78nQXmYq9sHbXv+tRuZTKQcEYFbQf/JufLDW
PN0AD8corWj3Iqt0xmxIfkfqCNNzK6rmCtS2nLYdcJOucCzDOj6bdwM831HuMgpp
I22D8WxNL9Fwm9S5/0otHUiVPSgyXCkjwsBoqxj+ix2i/WiBin3nUnT3x944pp6H
/SDBim3b6mze4oK08rYAcSxQGxU4IYhXYO4qzh82DYL7gKd9UV4L1SY3P7XK8N/T
t2nD8+EI+6h7aRUB6hwh2JH9sWfQiUljDPT4+CsZMF8S8tpb6FvjKfrFM6v+izo7
GUwr3k+/ekLqkJ03SuJWer2whEwM40CoqjHKLWIBt+5Xu6w8nbCG7avCHzBPdDHL
A/yDsMR+nmPnzNPYF998R/V7vBsgv+IKhuuUN9bbi2Frl5DD+/uERm6o6P9uSr3O
ICR0jECpDsZwFNPdNIYzvAHIUt59UVqkpSwiDBM+nUipRR4oCRxMOdqL7d8zg5vA
WmoRfCFc9u3gtSEPSn0rsk6CPxX6+WXCx0IlcBoXaIqBjoA/D6Tbu3Fb3iSV6DxI
PbTzB6lkVNTXzrp7CaCvXsrdLT5hjF7ebW1ebtcOzg3GoxUxcQgQT3CSjZef2CkJ
QkUfqy3Zc67YlaFYiBvzQ0qSJPnGVpvU6Kr2hc1DlUXXO2jzLg2evo1NDjOdocWE
z0BDoqQ7ydET/gTqDwUZQh7gHzIUrRaLIVczBV/G4++spCK4OTpy/IwV9wLW4FAr
HJwI9whLN+ogdFoKpjQtmAl9Dz/O2cwGR7b8aydHE+C7WVToEilyKaRGDlqUPejX
HGO4nrw008XwDiCSZDeRiISmoQzSi2ju4U2DlqqCkUMJeySo/8x29brTpK0m9JR9
FSHJQL7lMApfJ3W8VTCW8llgqjEt7Twulah71CsZpBKy5nmRa8OLL7Og+CJXP6Xm
w9yvVfTWC8+o117Mtcr7iudS9ibfYE1ZqWgCUZfJqSX308KHiFAnT/h7rWXhu6Lp
E8yd22M2IQ1yRWOI66ahNcewQXdktFlPkvE0LleoSvzbTwYP0lsvqRh/20EFZd9i
K4d2cuVjiut+TW/Ow0R+Jg6tli3FREOupUJvzKtNq93zSN6RaZTKV+gtuQ7HIMpI
zsG9aKyCLuEGtlIda2JYAhRJWXrSr2D7QLrrbFcDlnMnzgoI5xAlM8DvuQ4hk7bH
wonms566FGa+MkeemRYQZP7twlxnN8U0I77RD6uwpKEtqqmYSuZ7rloOl4f5BDLA
grj6uK9PnkniShxUMwg6Vi5OzIv0wcNI3090OrHXj6rhQAjF/z1BlKUT/XKfghg3
vNsvDhG3TsQAGEsa6dXDeqqGiq/V20yoVWBJx8mNnMdbULBiH/hJkFWOPRVQgYnn
b3pljvDXDH5XQw2vSpK9IiRjlTaQt75EXLww5vVrsX57NRZArkxSXqvcRXcKitMw
eLacZgmdPj8Yup1t+qNAA7mI3MMM7aa2BML/Hz8QGHoxCw5GB7xT7UOcs+Nevlb4
r4uDlb1fYbNjXWiygl4hD/rAzFAbG5M2EZg9qdaibIhN8+DP9sJ9Z51rAJFDwh8K
nJrq9coDRf3lVNmC8Hy562OzK5qx9fP1nqRJuDQiDLszKGE0I9JbMydBaaGXjGyo
FyV7K3dSkHZMv3yzRS3FNUwrXMIqk4sOsU5poTFHZZW3LinWQx1qdnnyBu52F8/l
tASEJSL0Wawx3GjUPXqBhuCp2ko4doRpKRZp+uP5iAoHSjn1i/DpJ5Srvzfj129D
ViAhbHbpNLbEByi3jqTzMGSmNJ8amhwfZJ5ARuKhkCp/m4LwdkL761GB9ftJShQN
KbJVYMcryMw4DDo1lTuBBPw9yyS+KtFYA8tpAqCVGHCN9RCSzTDxN6oVyfenv7Se
pkcrXAJ3H1mKGb123leM0Gr1NrXT+bXX24FqeaSeOSN1l3BjiuldzSQiBr0O1m4n
ZJ6sRIO1qxh9a3imh43J+B+Fq8BoqfAEEUQ/u4Y9lQP51iIS8hi+m2FjNTcE75ac
M81HmfVTD+ZIgQBnCtsAHyYc+6gr+ejudZmucJGvrTynibq9ffjnfQeDpSB1t86O
uBmVjg96oHvSOUg2kaAId3dokOfYodicF72w+QOe3x6GpBFfUNx1OcfRKvZopBAH
NHJoAz3rmwXEsq1ex75bwQyn49UBvjGwBraUiGYJ/KsvTlnr/FeSe+p+BbIONYKm
Usn+H8PNhoyKCfmY6/0cvic9tUoL3an11jUUor85gWlUefYzLPv85UYNr8xthB98
eTs60bjQj73BCKtNNI63awjSyZjIWuurAKJRCdWrxUUIi79z8FedQ2glx/EegQj3
1XGSIQgWGS0qxun4E54klxJhsdOTiHYphgxhOsOGA3E7mTIB3VgLRLFyERvpiNaM
KW80n3mBH/V8VBOVs+WrCMkWvg9BODMEYQ+nvw7dcSYNlRdkoYJhx3lnnSM0tq/q
D4Lr7tEKio7cm2jljBxnjwxlQ8ef4b8OChkPvYSgOpoi93HIi7VjLJlDAa/HlKnD
/syuGQd79ycU/sN0kQsJ+t75r0a1olSaQA++8r1f+4ov4zKAzrqjXqxZmVfO3w9G
84K2bhDxSCJpmtbYo3aL/bDcC1JaAH3topRHMQAMAPadYeTrlOGNoWLVN5ximeIt
BlL4nGbYzJBz2F6ZBiutN9pVRf4X1+en2Lvll0pMsXCkbUiRyCm47HWFdwxSek4v
xp8IMxP9XnvFTiyeW1hGdazh6ht/IUVXU1Ma3SofzJuDWh2p2wMlcbtIES0raFaI
U6lH1On/umblBtcKy7TpRL4jsbxctG8qNSlp28ttvhxOPIqt/oyymI7pZ4uuihBh
+WG19aUn6NfX1rvSsdrCUBigkpZOsNc08BsV+D1R5MQ9EMjRzuU45OFwGrXF0UR+
doszSxmy9ONDNTOG9FBXHO5KSS+feDUkry8ATSL654DLSG0gmeFFVcv+oE/1+hu7
FIZO/+UhKtH1u3NL/dbiie2A/NBCjmBo5nFann72FndnuaosWHYyB/5wN+6jPH8V
EbRcvWd96R5497WxQzENzo09r5Cv/sFBbWz8L76ySnYEGh/6aczMMsfd2c/geK7Z
ggI2KaVD373LwsxD1FNZY7UgLpiq/O1l7sr6rrYkgq9m2+cuOymRaS1EZrn0TVXJ
25OAxZ20/RBtFC8nb4hEcQNt1MrvUXTwI2nbMV2UqPHfRjG9gGCZdXMXuU550moK
0Me2UyigBvq2FqV/SLioQsG+7f0xU9HkijZX4bk4Sq4VsJ0enz9UTSB4OVRKQDct
DVflCac9xveiaQv2EkqIenuXXGg9wsad37Y6iooX+Q8z/hmFJ34nnyTKoLTim2Ze
4egZ9twkXwmTDAU1HxBuMRgRMtFLPdeDBaKYCZ9112I8EA/xvvQlfKhtHeHvFf0I
hrKwuSnmE0zOT8tszAlfB5LlRYIzgk31CMY+3pGmIOEDaIMYE4pU2v3Q6kel/f89
hPXOQ2TFHmiB4IhicZGadRcPOApybr41iVsVtuaH3srQaBny34GqXQ2n2VZgePmq
bR/skLqfQMDr9eDkXo3cbaxR4fWvdZXn/ASfnfwshSFtyRz+g1/uPsB6TEro7Yqx
hEw9KhiZ7RDA8JZ8R2tGMz0ZlXoSEdoy69s0OIgaD03M2TX94Zus+2pliKVz0slR
vd1SDFDkwefsfQWvvY9QyfqQ413HlsBq1vT1XS3oMMNdLZgkvAxQ/ZL+4aWaIJUK
XA3YqD0NUe/k/FrSgHqqI63mkqVXOgfCUcolPCDO7OEK/4b1bFHfjxH6yIYRZUWW
OMR8Oms0WPqmDD7Ep1Om4OUrbFrCyW+ylfBWK+fvpAFVnP8O0Zi2cKP2JYKU38oX
KY7jKbgaoeCB2WR4ajY0S3t6fWESL0iM6+lA0RLGp9GH4G5zGKiRD1rsJB4wbIE6
YitcXVDIQK7UI81sgvsynpRBhUuTvn8SCWuN1Sg2bFOYTAWx9ISfkYV3zUkvlINd
R6lDzZVklC+6jAyNIjwsbLjnicgFuQ37j/fZUmLNXv3ArgKe8P75fcpYfesffMNF
n2jTSC09CytM0k9OhXaKTM5EQ7bXxsvfzumVNA6dKPf4ocqOHUXMxsCXMsC+Sc6w
mRyNyC7GNu1K649BKOWA+LePL8+TVq5mjdE6RLFCFa9YLRVT4CLEz8m7z161s4DM
5xXXuOaiy12NDSEqiyCf3CDuYgbQtuUPcdf5iowIvV9cs+oCboQCKmNwW9gu9XI3
CQmX56ia40yJm9PzF0MwhLAZqBy42bBOqJZJr7F9KQFxFtuPoFgMhWR97CmACz1L
0eHCQKYp05/1031x4lsFFRtiQa9rSux7sm92zJryxzUik7WnMJv6HtemNVuQZuBA
qfG3fIcZDy95ooWwAsGeGGI2F8u0i6YQ4RU3BpeRUKi6OgZWkKd+s0d62am3dghI
8XIeFJfY/L7B7vfjopGnWvyKaojLpC8zzUF+94cjKzFV2714wrN39WS0a0x+48b2
YOF9B0nfexzWjwT2PBYwGXzALBJYD9Ty32iUptsQWXFXXxu/AaaUiM50sanK1VMZ
yTietpZoAuXQrkBEXa91bFWVk4dh9NMUABcNaW3LIElqMVpc0UtN8AvxOhuwTGUN
Vo0pSg81gfjYva2F+LASWSIeJKUY9VoKOC9srQX1GqsQ6P3dZnzC8IMJr6DR7BFA
e2USDLxuSYe6BpPct+gKAaONFn6Nk/SH/gGiV1vfdnD56oZfB3RWxBZDLqPS+LGW
d9qHgdev+rOW484b3ObdY4QHRAJ77cxjHF0jbk/vX9iMKV9kojTbqZsgH5Rvzwm7
1Zbz3Kk0jOVo8ErO+uVr/zgtlxTLWuDGl4bEWdQTYdVfbrSfPw4o0VDePVYGqiET
L+6flVmTQtdRKACYgNmj0lZkBc9UJSoHHuCda18x75Tkt/Pxx+zZXu+XyihevMJA
i2lPKBPKgu4rlF6B9GhRzDXx2vlE6yzi650JqyS+k1OuPeSOWlLeHFYqEqlp5479
E5MarDdj+w2tHg67rWRatiZXPfybdKE149ajhaQ05XVtJK90JMBz6xVEYjvAruk1
HWTt4O/O4fkVIRovGOfW/NR03woTsvDnRmVtwrokl8mYxQiVhXqwsxvFjsUhHM34
v81cWGD4JuIqtkmXZWVn2j5OhwnMdVRj1pSWEnzwwd8SSh/FJ5606j2SJNdZRDDj
2al5hC2hYQiVHvGOtwfLijcnfJ0OLZ2QFWX1Ipyv3quXHkPK/vSj2BWXjthD4fXC
BgUqPhs5+oF1J26OocgF7h3J063ZsW5Acf84upM0IOHfTCcnfedHQ/rHIzX/Xl07
4QP2EbkIzfbhJWfcVjdAte0D93x9cA7w86Q2qZ1OQpim2OP04/YsGfkKP5aKNlEZ
h/S+xPd7fAnZkTiKIaEYuEeGHttYEi8MDqD9/jhZJVbe3QIc4RwOHafojRQQoe50
y1Nz2GSOf6IixV4oO/nHaFOkgjpT1b+Whmc/wH1EknZHOJlSpqp1Oc6FSoG9PWlW
fbQa+9AKvPOhtjlnC8qlO20MxydeHtibHmnalo5HCnhcovivjfrnMjPnJ4N8zwrz
efbruSQJQeBnKP4rNwqeqZBOkikufPzmgYZPapCSG89d67ygAG/CJVOpwZf3lItv
FyvOd+1jZqVg0yetLcZwkWM2QzCE9TryF1Xd/VOL4/fCtThjeXV3hqef+AC/qkmw
0LmXUqYhgoaEjBX9j+zFqojZsnDJDgpSpwGA00/SlHLXcyRInsW8EYXcXtM1xA/G
wHEX/p+z2h0L507z49HqqS1eQ2qeZV+qiJ7Zfmyy5AalHJOyqdcHnKb1YRrYAJkX
hMFf1zxFrd/9cyIcX07D8qpVB9VyINBMxo3zfMDEZwDirI4/hR7qIe8YoaLTQkhZ
uZQqKaQL5XNdygHxABHZ7KPRyre1XWr8PUHooXYCbaF9ALo4i/nKd+mHCzILl+Es
LL0N1XLNqSktPOQRQ5AZL/4GpaJ6iWH7pR/NhUWBcBztZug0AJI7rJAB1UIAcdGY
UZPQfXITqU0nkMkJhKnEJCMOjveL0LSgvvt706fWalNiQ2EuNTHvL/G/hPn/ieuC
1nhEAv8OfKeTiEne4jwciXGaY1z3uAVwxkbNzTWAjQQt/KlKp/TgMdcNn/asWPky
M3RFQidLp6NcvZxyliyg5Pr9K/KGWs0Tnlbvac8TDfDZydHJPPJL6iMwHBi8TUaw
1F2wLmITtJILKEjXbw3xyPRDYr0HnUmpS3ReHwwPM3fbCRDeW4tuD2sRXWXo4GOt
vw3S/JTapcKowlWXqKYifAYKxZiQZ0VUDSJzo0Rqk5ZWyXf5HF9UO6VIfkOz2A7+
k4oWRLHTHrfi1WLw/sVAgY2LX8vOU+2efSNkEgbZD0MOMis/4fWFXION7U78qwDX
6F9EESmAdbQcKrStQGcGfEjtvGMkR2LShzAZRqjjW+egrlhCP1Zek1uUuPmOH+9o
Xjdqx7FbX1pb157GxcRMo1MAdYwEkU2CnTpKhBpoJNrPjzYrhccohjlFJfPQmSbN
S1AFL1cQkf1oiI+bV1iZQ6PjmyfqTQJqd7qNUz+swaTBP5HsCVXxQyRLu3bBwX2N
RqniJb8w/nhkoM00Bu6zF+QgbXrDeWR7gLeACLiIy7DOSds60ZZsedL9PTeY8Mce
luzOhzBqvGvBkqxEKs1PEWZFAwmtAaOpMprZAt9bjSITBWiTOYP1vxKzsKBqkJd9
MisBZhwA4UbMGfrdNn0o70MkftYtijxZTqjx3FCOJ0nQWQzqIj38UOeiJh5ttxYn
qs2sanrRJlqgarUsucZmBirLLuIzlwIFZIXkjNmvtMEbt9utWgi9+NYD8wCnd3is
IgR/zcMqcEuB1/W417pemppvZG+ziIFDt5MEqI1A5dnLZcZ8dSRoPS/PxQGv7t4Y
0hApm5+NjoKcVFsyrrGiA9Bi08odsogsHXHCcHTHgTmi4SDy+5RpXVWqSiaUQ++C
CKNm5OQJLAGce9hpVT1tPQUclUzQlLI6jTQHKRCSu4OkwiCYWV2qY0bKLaZB6ZO0
Wg3D0CFGJj6AvW+P0LtSyj7cmQmbeq1Gyyd/DsDb1D8AZuBbKzn56yFfo9RMOEkq
I1KDSyOwFIQcakHfX+4mZWtfSEvFruVfArqmFs+eWRuTrVFcnIdPStvC+617JDAq
EKlLfJ5XSkfYOkKmcanmlm8hU9BTTPevLglJnbm89oUMVapiE4jqxvP11kvVdZym
S+lM2XbEw8QgxCkHOHw1w1GT6gcJRY1GQngEEwv2ZhRVoTtemhSTZ4FR1SkkVM+Q
7ROIQryj4CftgFUpwkh7NsBr44HwuOi5VzAmNPnyNcbR5m0n9a+RmSubYyyPRN6R
o49ctAYQ0Uutsz5P46ZSoDtvdd3lOqowWQg7usDda0fWyH9036hqFTR/D9lwG84M
+UqrR4wDuo8Iy2SWzGb9LNKzNFwZYAlSo1Df5RSrmJMvKndWqnk2VOtC108DRtAl
JdjUbh5Pe5aC/E9mnQeZKk1v7fkGVx0n9SyeliH9EOuVhSAmCAJ33OTSnY+RBgN5
PJOxo7EsBnrmEBJc/J2/tVcNSDyPPLzf128TqE8BLwu7BULwr0wkP8NM3sooSqa6
mNYxQhrMPPOUGeYHdgigagO4+hNwIRlJ1EsMWhKHKRa76L1eUPHA83TiUgQ+J7mD
BmIeQ4QzM7xVNwAcc2XGkP9XzRcyR/fH+rrfGuQEN1ruQm4pKgfJaHUAPN+TFHN0
vZXnpOIngeNb1E5CpaBeF4hNDayFt0uDPFVpDq+PaMZM6afnb3oazzeiWsDCWn42
z5VnIGPCSFtTMktdM5UFCNEMKBaduxGJKToZZmukjLVrNyIBvheVrPNLqV8uxDVB
gWo+TadGc6l9sKYy9p+c6HqrVN+F0SZYrMF12wkOLkAqXgkkdKaC3kywHJqyfCHv
U5gmdyIqD6m5pZchkLZ7r1S7pkwMNvnmi9CXtwkzVic8qg8AgIXmr5UOG56CK6mA
eOr8hqBD7rNhdRcZJViSHKmQqLT65avOFKsIDbM9C3BoWuDBNhNwApIPNrHj/ppc
sYliBYydFGxoq69oyk24/V/NPtYbX4ddwUsDEU5VexLnyRLYHAp97H44JzIPG1Qc
+aZiyAOA3EHIsbArEDn7Ri933dJKFdbJc34LzkSHNQcT0L5GNF2eeBaJMxxhiwh8
jouYaa4tx7KeUUNJcKQCED0uqeBYwa9yKcQHX32XG6kO7lKCWw5Fn7KEJpQEZcl7
U4wQ10sL2tkJESZ9ENJGoUK5DDQ7jCfoW4It2A+dO4nrlorqArQ3jbC2dtT3QrZH
yaFgGRkLgjLqRTidDph0AmXsSZYT3vJ2U3JilMiq4Dy3zbQs8dRBNJubAwhcrIv2
XrBKKsd++U0OnjcR2GvXH4UKZoubk2L65cIHs810CLY0fO5km7HxIVKGK163v83I
ChIAiA//eg/FcQSQx81a4h7FgVAhrAHeze3d3bqot4Otwl5aS8op3uSKdJff+Gbm
53hJ5+rMRUvU8bTHS9xDlBAgZW4+zyszPbCDuWtpDFIDlZb+7Ki/OiROjChKo0Z6
BdoaA9uBrLx/yAD/s1+GEkhykutLQKL5cLsWDOL596s0CS6DvSKK+BsTuqO2VtrV
c7ppYec4hPu0OoGKG8UKykweDYhDPhSWIriZPZkb2vHcQyF1mErXr6PReifMBKmn
dLqeLnn8+gqrr8suzuP0Wavg9WsSyEukG48y/JbUZ9gLtLwjhCw88oD5kYeUOZj9
Qvhn+5Cg8I1lNqYw2+DkAsXejw78NdYNUT4Y0TI2yniXiekD+//FJBP2R0TXbtiH
IGfP+3W71gzm8OX1HWtGnZpbhLZdZhwsLlmDv/nPtPxr/QTi5LEapJ9Jdqu7ABX1
mX7fapvURd/IA5L78XfijJbqksAnmQ8PdDmIf6RTCNKMPpNA2e2+ZREmOfgaWhZN
EES2DB53bKJB77YKNPLx1FrOMKCzzDcln4WG+TENNllHhRSsfoZW7zDu3F4mD7uJ
IzVhw68c8NdsaifgYI3C/kwiYRKKyWMhhojLCrmJJ8R4rSCynayfeS/lk+VUKWLC
uXWnDMyQ0EZNHwp1pLDx63sgDBN9rcYvTRtF/SazKDkSjA7pgjEkNXRJaC68ReLP
xzsGzorlIHjTnEGWVtlBhpp3BTrYKOlBwbIY02Jw2tG+mhWgTIQNUvzyr9fQI8/r
MmU+G+9I5Lil5Pdhzxun39taN0RcqzXEJyxgmV1Ds0ruBbKfsHBOA5xl41mZmJAZ
ei/gqJAIEzTRKdweJFeVc82zBqIb6pb7YAXb9fYV5zZncMWjiI3Ertc+Yd697zNS
//pragma protect end_data_block
//pragma protect digest_block
vQSI3srmZi0X3gimfNyE03VjpQ8=
//pragma protect end_digest_block
//pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
nb9oG+BunXzpeKicQsYHftL8OuxGQfgiflwWsF+bkKcDI88UrCM/NDi8o2br0f8b
UhzY3crm73KFScViZyHwuG4PuHlHldT0w9Db6IjgECfM9SI4bR57GXEKNVLYbxa2
XwvDVWDvamiueDFGJGopY0ScLM9cjvobzLAtzglFyca9V114qHYJXvPTWSmF62DM
KbcON5CWxB8XnIsj2xemQ8Bg7EeCZKJCxYmuxjxKm21HZtjTnF16jFypNQeGZktN
PkpC9ZUHIGf6RZbefAFOKwuEQfyykuZVeZHVMCEjRNPim0otxBC/OVShiz5PBbWt
NDVFMddmKfZ6LbIysUgvrg==
//pragma protect end_key_block
//pragma protect digest_block
cT4XO1DEQp/R3n0e6x47n415eJc=
//pragma protect end_digest_block
//pragma protect data_block
OlthMht+0tleXlnA3cvYTMZbWiY/d4ckHyHWSjuIEZgY1XP7JV+cf3AjGqQv04ms
Eawtn3wSEMpgRxJJHyJzS2kp2e/Nv5xUWMN9UsqV3EIsVfl9u85ZVAsMCCSEkEoj
5dRU5/4Aaq+CE6Eoj/OKCRgkJH3RW1Zmp0TZjjo3KUql7H6sn6sGE10QLAoaoW+e
EEBU1J9joAT12b+xVjWgdYN/z2iqyqLJl+Q3fTMVGMDLb6ViNFrgjK9CEJ/tFSDb
rpo3V6ZVOisfZV/P1XUe5IKO/GzVbdaoWSaot2O9wI+LUqk9DTfFpQbh1cB66wbH
9emqh7XVtk3wv2R6Ac5lA5WpoFfbSYDjDa+XLkkM1rer0/vV0Qg1c4eKSsUOX7BF
Q3fkBAMadhHPCFmVBqstoZqKwbwevuJrF+JZBrhYPyTJW32+pb6jga9zDJNmLLbQ
LqujWsKt1Ksam9QRgKLG8ChC/6CIxzi8dUdljEs049Rsfx+NRZXY9Rh9pSYbeoow
e6bI7X//awqZPRklbm2TJbL6CmSjxaRE6GLlThgUYHo1YCKCj35K8ztZCMaWdaON
TyRYOJPeVFzdOmOuaPvx+MoKE6PwZ5nxRfWZnoIZXgUUeuC1p6QRw3ddlFxp62qe
kecsVziFJGJIxkLXAY0rO0M+FlN9wrXXdYhnCS/hceptAfRBzQZuLhAPwBPElGJO
EApIQlyAJxSsGJJw3TLoEwwdLZll4P75xXnW0w17j3jJJz8ryNpxRMehAIFjHHWw
EyO0OTtsCJe4lkTHVJtbiBRNP+xjHRxf/VLmGJvHh6c7Xea+rLuCfWaKoNmJiqhw
/JEjQ9U4nj/3yKLG5h8Fj+L2dE52n41R8V9J7hb7cgjvy5P0NpijnZXqv3EKzrAb
Zr1kB1N+4kRLy4eqfEdoOJA5PzMj4iAZrXxsYjknJ4b/yGCXdCjdQYT+GckMuUWB
KLKD/eENu5EmupDHgBistl7XMkNzfmAZq47Yq0kY628HsX76RnR3z1hbb517y7X0
ao5GrnF6yNebAfjkNyeLsRs2C3GX4qEC/6qfIy9QM4gmBLxSJFsABZ4w7CtcSzBI
XlWA815atVLAFkpuOhB97Fl+NyLajkLJafNmCR1VzpSTjCmFPjGv4ZmMvXFAaeAn
e1cx09hBAB3GTGuJua6DdzWAyNTPN29pVo3Ht8lapZN1vr3eWD6iTSfW2JkgMDP5
VGC6MZSsBz7iWq1JsmePEKsmpzO6ZUdqNTngl0ydY40bOJANeoWC0pnqhD3gFCAa
jxIpUoSHMHUbUVzm352z1+N4Yc8bHpXwHZ+w8wwsnktlC6wmo0X5NTmz4RfX0EYh
19EPVOCEb6UFKZIvpEs2BS4MUBtqWWHHt+n53efOU14KiXLnozpFJd/Np/lIQsyP
JukwyATe6tXcPOdd3J4rEVUpGYDkOlYW+KxOWJk4WUHN84voYrD420iMkYpiKaHS
K3RlaPYVylmelJMvdoY4VR6C0jXcGak3t3ySUW19yw1qGDzxLLEyfDIeCvg1Yt37
AJfMeRrRSYQCZCjnXJPbFNXArfJ4e4holRDtrcZoRD/rqMKbl865gxIr7tbTZQfM
n6e9sFJDNpx9dHMV6ZNhLsKRoJVhjg93E771c52ji+JgVvCya/wBXwBHzMswmsMZ
NTI/IcOG/E/mvWGG9mdlgWsYFTvZasw50mjSefgROk3yiJqlhS2/mu5mFpVNWAfq
ijYMmyPLrduxg68vYfVmhVM7xmIClyUIFkir2mEY8VfnuiR0RF9DXzpdymfqtAbR
H45cCeqx25ZT7qcuHzsnYry1Bf8B2Kzf6DJgNzJlJ8QnMxvABFYqW/k7r+P52yI2
pWlLdgScrkk+Na13j57ZOJaCnakIOsxOhOtZPmW7118V++2QD33Ei7N6AkB5t1aD
Ouuj/s38w9xiPaSOjbmoswzJ6gUTwQlnDhm+VtBr7e6WWFe7E0umaaxxUAS8u1lt
H6aTrr99wBBhRt4S24TKOXXkfVfzub/8z8iCoKMglhh/EeVHsEmCqCJ7+WShtPZg
ezTGXARPX0YM28XXUpONaoB+yquGA+/TWqnbs67G0p9VgnY7WbUCrk/fbJ/pWmAq
zD88ZZJQvM/PrlQYQRbC7TAjPgWufESVKtRdvPnmnQfnXIA1pyXaxz2QdO2iHO6z
JEYm8nydBT07GqzBbpwyH7MinF6NSu7DBjlCVG+AB+R4F4/EZ2OaYzPP/4JbLqqk
AjUSQJYhs/KpGiDKxew/yiMEPw5vUAy1mJfD3UseyvxzwPwn56WCNVKLsQaN8neS
ZnPEPa3ScqWpoo+HdTdsS1o4qEWynprmV1Qd3H1Lx3lOu0pfE7RBKvAUXe0AZwJF
WK5FUNGygJl/Vnfy2m4detfKoxSBhRCxRKK64WVo2am4AGEPiwmQJh8YHG16p4es
N9C8B5Bev3U1kyBcPKAAcJwytyIR0Riqz/0SY7hroxrAPU5GCxfMP+VPmvnvZbqA
eR+jbWxZ91wqHBCslp28pmFkLFRSzN7MneLgDnmtz92/AwN470xCh9hvn/L+Tu5F
pZyR/CiqBIQfdMJqcXnQ1KCbGCMOpHVXwoBz5oJGjPmW3SKHJJweAmFeZdi6fanD
3F5+aJUi8yf7cjac/D9CIUNEtFcPqGWgZ4c2wbO6O1tKa5aQ0ODdovkhryc8EXAg
oGDJIpeGFPd8T9fRvC6FHOf3PvVr2Z42hPNpgnXzEYLIVAS7SXZ5k9WJgUWocJUV
z/UJbA5Hm+2i1b1LrmUCpN5hUNoYutwm0BUt/MOd9VpOt8wNlwlzVYmd01l1cP/C
Z4Bs2HzhymwONYyY13nagamKOfE65xFrNQV4YapGJ7vqDYnrASdhbT0OHULOGxWx
tZLDyel18EUPPgU9Yl9WFV0e0zSRg6DiGpL0QqUzB7tp1n/CZBFsBnE7xMEuWOwM
b8nUuxfYfM17eUy5pmyJWhzN9Dk0pztRnlK67Hue+3qlIoyEWrZnE4z2uR4DL8V2
F1QOfVrU5xulYspU90M0Ny1t/+iN8jHb34Sxy4Hk+nPDuahf+AVm/212O1kOZvHj
Ew8loRyNBPXYHIkT/ZL6hPEbCUqj8DimYIBSsj0tIvhVGvsBR9FTxWYIci32eslO
9smNkhiY8GZQ5XzyFLCrJu9sd+/aShmzT74qdukATPV0whm8fgRpTx74djFNRus7
/M7uw9jVa0WA8eXmFdzW/idZ0mGT6rrNGJ0fXfG7dLc7SjO8+F62kEnN5CoXzLYv
b93ON4/Ks3wy0cHctkJcbM1nZETbXOgTdNF+C0xrPlGRHnOt8wH5W8cEdNYAirzx
XvXO/dPkGI0sxFT4ugzTBECltQDmGZHqQO1eIleJqMtZr2OzwEFHLbN0Mlr8877t
zbXZbdOCQuALN93LhnqCHPLc4trhUP/WPftH3HBw7BqyGaEk03lX6XSYOL/YyH/B
mhi4hkVNqXeXMuiW9dilEt7EVgKwDcdZlSVPu8pKZOAXRh7zcNjJy1BcpQJxhSv8
ty0S05a3CwFPAkHotAsjAjlBdgpqO60b7EvYzL2dsRWOGOXbgvdZFn59wO5M1fvn
W+JFSiuab1t97HJlDO+u2z/G9xHBiDR42tHVDQIIZwJMnLCtr58nk5JNbBd3yqri
b9zEJQJ5gN3kSzMIpFwjl92XSZOjYMSuJN2L+2ikrRX66bE6yOrY7iLdKsA+PO95
hGhiVyf9d7CPmokZ5CT/jzMef7mQBlkKQp1GYaAh7BHHIudCoqDFoHCRjaVEPRw3
dpWdOcqIzyeOoclcLLg0nZ4CdMyEwXI0y2RRO9LSm4qRxyf3Kh4A1qUkYo8K5veg
3t8aAh45aE2auVfg5Z237bUzS9nVd2KJTobHGzMdnWdeasHhPqD96bureFlnX4pV
YvpQT3xiBjN9yznhybftBVbwm0KQuYb6ZwNSHHUusDk05qZQ2A7XntDWutG7Dohx
fjvRl4TWxwgKZLCyjotHpJQalSDFFgYG3fX+qP72nl+nWstyIZ7H4xyTfoxfvfpt
3pA4XYSjmqjv7c1lP5BLEcyffpKGf6pOHfhzjjp9JTfY1Oh1A8eXgh2F+p0yqEdH
HGm1OyfWwMyADT8AbzpIidYI4ZELkHZ9bYqPnmVq91uVPg7AvB81sd2fUBS07CoJ
u2ziPMFP1rKMuuG6RacJpkZRF1Lf0hmGq0DmmwNChouaLLmMiegVQyYCB+xXNPrE
EJ8UivCs37vbg6gmQTM1U19JM3AY0cFgs5lY9lY/XqKHLQdHxzr1m4QxCRp9I+di
eaW6NKQJ/r8DrXGif9VYmJwv0arlfnqMMx8oBN59ucIZGGTBceWSZZ0uoaYTTUw1
3hYZIjo1k2EivCglBiPeCfaL+rbLIotFfdqJI9ffzP7nihPH1ZCe0vkRUjm/MzY+
t08yo0wRAJlodEOeWea18l+P07lW5yQE/cdYLl9WGSQL4AG+xX2tVnNxI9vvgqlU
E3koLybCIylijLnnqR9L42/3bU9gzFyRjKoM4Vwmk1demgfkG4NtreZWPvywPm2y
0C0R7dZAsrqXnrOeYGkJLvt9H4OuPZ1Y3wlVLZtOZhl5yc4fFw3J7XEeOZF5ViOM
FaW+/xnM8ZKlhSsriie7BMtl4rEFqEjht7tcL7iywcZgubAATUH/y5I3bALA4Z0C
A9pnAGFqDMFSVQzObKJLDVgsrPQxl/TqDDhKVkk7z5MUODZoWyCr02avg/c33ea3
bdHk49Xwx/bsMw0NdqckW/WuUPeEu19i5OantdsxNLj1PRSdIuXzJMovJU4H61JL
t2nEp5z9ejbDwcV8mhziw2tx27R1+qFBIfWMxIbWOvt4RtHyHmjky1FVRi//9mOu
KX5DhWDNg6GVBF2MoRAJgCR6X20d+irvlSIyP9V/Ju17iPdi3bSCr3gDfuCd9sKP
1TMx8imCztSdm2GX0/sXC94GgrjI2d4+LLwXcbaQP3/as7pCAZKO36AlPKRC8k2G
8DhEHv9zi/XKS9jf/b6l8FP5w5zm5yuWUd1qRsH1/jqxoEB8a9V2mlJLdSNWqD1W
t0e4usZOSQ2jrhaEORVtn9Ymu//2oR/u+vuEJ5pMrMck7ef0pgvidjBlePPehIea
91eI5XyuLroFFQUANyHnZs8mz25SGgkMUWI1ENVAKpnqH6U49MXS2MrK1SlnOV/+
hXsGAZBhYNnhz248NdaMDw40kaT0pUccuTYN24SiWONBPTXKzLfWm/dWmUoBVPIw
ynkhe6sz7oVdqYePedlj/gzG4SXIbEAL3NNGWlUyJL5WWgsGfhzVI2JxSGDhR1TO
+woh4JojCoj7OBM79AKXkq7e4bE0n09qmkBJG+HAZMhNjul6rcP8V1ihU3UhB53q
6T+0f0kSJOa0egj1vqSDwE+MQByUDoF4EmiIWcekiZg7r8/fr3HIipjLzR6muf4b
PfadhoSwGNORyUT3neZnXCZ9eU03T9zB6ETSldYjm2s0W1s79QOgmvOYhxyk51q0
Rng0xRal+0A7SG6F16iv5TaHkiNPKyiGTwBq6FSPKWSwNB9C4xEwKcDywWO6dymi
DySNpBE6S8omEfaWP5eThxVGf6LDoXnUcUDDH1fXkfd9FiPkyQyRQOWHE5rlYI8x
m1WbJaTJLxBflWj4wV6U1jvzcs+FGY7LoODcUEJXKkNj2NCOG/1Yv544JD6YecMh
OTGD8/i+Tp5NMpcN3H23jyQqoctdUSSrzPbIhj4HQOpPawKGiXWsOTdc8oci6tRJ
OzC2KMZ33H70DmPFMiXMVZr8mK3dKH9BomreV28UDTz87416ELRt0ITJIJLjkc5d
eOr/8panuSLsSrWa3TyUQ9jaiFUwzblsw13iaPtCTKpmKu2QgjpaAM5yoadiOoFN
H+ORDVCrIT+uC/b6pYWX5CcxYYuTjTGjLVcy8TrEykpYHS69V5YAq8dzp38oPOSN
ck9OvN56hdt3NXiQqTAnoEuu4XsfF1LHWOvCmeLIm7YpXNmB4Wx0WetOGuA+o2/x
Lxo+8lV5fsaXYPZXY+4sC8IS7LCfEcWiJQ6ZaQbXW0rRCb1iavuYkzjmckFIRWFL
bCN3r+yzdeOgaS/GHqIc+BlhCrMCYIAHEhTZn9AdKHXDSDTmu+GcbLRFQK/4ejcn
tQFAcx2TZoj2ABxUIyFAtQrJQBw945e+iMpMewxqUa/Vzrxb4hFlfew2JMq6BCMx
LHB/tidiabeg4I2XBknoOStrsUPkjQpH6FY50WWRxuGP5+3V7MjK3egcLwJu36Ex
DruVwN69pRRf937LjTc1fxLfpacrzULY3PewADuzRzv6ekurT3a8jLrlmwLl/Ph3
xhp7o5w/nawNNffyjiaTpaKseXHviB9f1+sRyKw7m1VORlW3yPjzzrcwbKXfcNTP
qJwLFKkNTdPSzCZHdFBbB5LwyAB7AOdiQCWYt015/PMnwet6Q+52IxCjJc/uCh30
3xgB4EXb/mVty07oTH05EwK2D9F0+OCQvskyu2vHLkvNZr4NNusIXjJfkxhftqFi
qtKD5B0arDLq1OduHUvyImGsVOxK10v7d1oeeUnap3+THvRW+96W0FE84xqEBFJk
Kxq/Y1/3SFJHqxgLS7Kn3CD5TDGx9zgI8wjT7TUCDq6QST4lFzaxibkb4M/GLy28
QpAGQAqO9kqx+U86/nUaLTt8ISQwIkQQjAYSnugQ+SUh8r5d7COyZeUAbSYp9pLN
0/tX96pia80pv9v+OHS6df9KnEyM+ldzUOMLuB7jBmEVVPU3mTNwjOy8QfAXGS2L
fA7w/oV2nWCQK7b1/WyCKQOhmlUrnnTU+hEm3dtuBynXoYljEBvTLG1ajBR58No0
4rGhjICaVmUBlHDRYXxr2eOPuVg2/q3myQ7OKD9LHxCLFWsOCBbNM8FNbFbsIf71
ScmHZ0cwRfCPb2CNiRl60Oq+Z6jgNrhAA2xgDq7mkhWPz7D0aeg9mSZmTIfuslse
NTReWqVE+fpwl5MZOX2RNJzIvqM0uNDkyoWE5VgRHAHJdcdCvNzVEmYx2kPCCyke
XF5Bc7UX190puh/bHrvQC9fTi6tYWT48enxUjLsCXUumarzC7lxDK0N7fOsgt6Jm
46Wh8nU5eKf/AWmjAJucvy6eus2XP91SxBwCKC3eRl+kb+fuHDpNpdgVmpOcUmjN
5GNDSaJtJ3n040BpxTBt3h7ZFxbxuXwBS318QYYMxlgKxmLWthkvfKkOolXPMZBp
AZLC0+7/hioGBk/mkTHe7SA61upEC/pmoTsjU/l2RFTsnNyti0os6pKysg7rcQ5M
3+8R/SdzzgIA1clqxgsInJV5cSVvOkadONAycklHrTO6mWmOaIAxytceSLzr9vmc
AZqPkmPR/JZDsVtoxW4cbz4AjwgxmfUAsVrr5kGH5eMovDNfaK00Pam++PgYpxtM
R5zkxryXnFYzaNyu0VaQQ0Uqu6GxMB6e8u+3vOT95gCvoXQAiVMpnFB/4EV6jcJq
QMeyHrHffRPJbYp1mayge7PHFHfUBbd0j+kOaHDLSmzJBo5MFCKiWyBfNaul3T7r
YzwS78dxlPiOWSZSHwe3FqC84GfFBLbqh4oHwbKVhnozut7IgsWxo+Z7cryVyxDq
9UASYZjlIS1yI4O0ZANusZ7DHlbq/4SliEEecyrZBIbI56lKipeKIZRsaURVajgR
3toAbRf9Kp3QOgQMfbH1Hq1S0itHZ6bdOfSxqA0Ta1rJqVMlNA3DOkzj6HbSkg4T
8Tf/szb48I7/cPj96Aa5CcuEDQEyTnF8r5esw/84Austu/cfUhnbKPlxdFmDaVq2
oNrUKGfpWLdMfBoTbsvdZ3OVLoD5VAulxPA2/Tx7d1O3vpIDVIcl4GpoEeyzMaJj
NB5OPFS/oSYXpBqYSL8VKDeynPI4RfepSdI+0KjBK7Lzeof7ZLv5VP9/vJkVAfp6
Kxwx8MJcxgvvJuMlNL3SobRk1l9s+Yu5e/gkKIUGBo3f9q0HjdehuCSTAxOBJhvA
Vy0z4v68GURlGwewk13DfkhbPuwiolwBKBne7gkuezRQacfPDEDaJmeKGEiQH1/6
n4vqGjIVp0lBVg2lWdg/mON8mGrQnuoOGDI0PqRo2TBiXcBAoi4u8dsb4F6b0qiS
ckt4MSBCJkM4fpLGqkHxLyTwQPdMzW6nhuXtI8yWJvTawthAWGaJ3l3AULHWAnHQ
b9livczwNgCA+Q3mhRN4qk6FIJdWzq9/QXQN8kpzezNWOApDFVwZ2Y/dikCy7vZw
3cqJTpdbAju0JFCTQFTvz6jksXV6CuFGaOjqzcNxmHBMzv2O48i45L0T659UpMI4
74MR6IWq9EC06+35raP6+LxWsZM//nWV5B68BftTPDgA+ubuJiUnnOjcLuj3t4Ll
gApqusx4RaCBGLUEfi1eo4CnOkIVWljqznbqa7zXlnGvZmMXahNoJ+jUHh/X396e
sb2QM/5cF5Zs6014Zk9GZfryUIBm59Uoo6Oj+avC3g+p1EsiWDqkSgn/34ZfUIdJ
ORH0HUDjWprrpeooNvyTzb7jWv9gCI8SKXZpMe4XCoxvoMG/XNaVWyiUHZoDf0y5
YRM4A9Rj7ql5fQRC9+C0DNA8pm/8g6sphI5JfhWCfxEbusfV4e6kpBu86gZCBzuh
EcDjZqDIHA0c3RjJ/ExWVovsBbcZBABXWZwMoeZXAfIsFaZRjTqVeDhi6sZfxXJR
bG/ZpXidOKLE7gpgfWetzoffLIpBwbPuhPW4ovM77xHodvtZm3o41ObpNEWdpQXF
9l51WZTNMEie4bpYduhbl0ydVq0AlQLr+XIt7+Nj8Rluu5NX5R3j2spYxSB/B+WX
J0D3gCVPaPQ0s0Xna9pJOlB11b+9TMlJ3Nvpf3wii9pJqcsLUeJepICqDrsyNvFr
vybnfz6Mzu9pTaOvx22x5ICSr5uVFFD35Sw/1RQQGZN7EsBXXUSaGH68IS2qh12O
Sdq+giOCz4Ywd9BMKVJKGh7BYL3iTVYZya6Y8+x5XerkuwbHzwCt2sYxnP9OOsrY
8T4vhmPcyCjnj9ZmTmXyscKW+G0qlgVVMSI4WPI0+VSmjheBrLAsmsFh7H0LSupj
mLRq809m/78AAbjf/7En5toMw/QhQJaAi5n42PaS7C134c7mWschowgpM74y5EI+
wtExO9EKSD0WxyWVb4WlEwYbYN5YPQc08T7RIYbBXldh3iCQIK/uGzxEchUbDog4
rrnECyaN0Qb8vAoGWG/tUMRtQhIO32YAKuPeE/d8Phlah2wMJ0xfiwiG9jBnLMgk
Cq0J35vxd9jvGyIAk53gsRIx/tM4WsGgQ7ILAG8gaQRdD8J7ZC8imKIGb8+lUJ5k
plJQADrS6Q+JP4Idzle78gvNAS0Y0U3xuuERnJoQyIjw6iFJPsM2jPjpSBSYeS44
AsrtutU72DLbvOtHk+9hYi2X/0Pb6qOH4mjm47iugzGCmwKHntMxAPFksWtCTIHU
IFjFf5oKnYAil6IuDvWRPMpQ/iMYjIRyFHgALbSISJ8KEF1Hn+f9BtGC1XwzigIC
UMFqiXOx/fACgv71vBPk25zkBaKf6ztkpS4SmEd/29yvZrstd4iq9LGsadI+WVqP
surqm0+8UjyJ6gLWALG7I6O7Iid9uvVb5dlAQmY59SBVCxW2bh9toDH2Uyk22nI4
ZhZLcnbrTlP1DsuYwbLogS308TFFgBzy2ZQ/swFW5XNgnR80ChEWmQBp9FBU1Hxf
O8gtsMasWrbZnQEL9Ap+Q+vYhXQ159jo68UQbouUTyGhQvhFGWN9Yyg3qzYgRnrU
aBDg47cqgcB9KPak6IlPxQ9NytU+nrCxgs9rNm7OQpyvmnJ8mmmGMSkgmavZorOz
QV4tcGOGYLZmqDDvQOpFl4pbz7oqqMPUDa80FG6xFAuzlid1eMVHgSh2BHCAnum3
i2C5+Y/uoGcuEfOQq5BoVHUGD1BcEffhu2/N8y+HRxMmE+qaBOYToAr/JG6b9uYC
IQw0XsKUyrOftD3C61EFn26CsASxCnt3yddj9z3SVSl9XDqii8mmXqlWHmGNd4Xd
O/J9iyGwgn0P+1FQ7qp+Kn1Gtuvjwb2ZzfUl+KjxpU/hrtNq1/DTGJmcah3/g4ig
gE0zAEepUg2g5nudBTvQXXuJXtUV7k5qe8YCZl9Op6l9tr1khhCkUbLq6koHRBKU
B0DPJkm4d7D3HItrNvKUwnC6oNAgr9gzmigLdhUNbVukr28NP5BDhnNrlvwWLuhR
Kbeh7oEGIbTmcsSa0pmOuYZ24VF50SodyxE8WJxi2n6fJpMHSXkn2hGrn6P90O/J
xMg6p3EIRosoBftLeLuCGItUoDldqBUSHIT2DF8mh5cxLQ/CATuzEEKDdaTuZOIQ
TrSF3ssaYEipueJ0f8VZ3d7rM693P0WR5csJxJFoQGZUGKaISpayWWzbt4/FSITb
wTA0PCns+gVS9OvxSnqGYU6bkD9LSWeh0cDsrGF+aaM1TnfTxvD/6H5ohU7eQRuT
0fajohdd8PKzqdV4g/AOG0lH4uPHym+Rp45nGrxP1p3hou15XFxFfKaNZ8OXdr7K
r7HF5V2n3dOGuORmKVw5Gsqk41/3y0C6G54SIQqZxFy7WcFoqPoNyRsdcSR4CQ+O
teQvgxn8vxM5afMmjWpCjSzLszuJvHA1HrgqWPmLWU38VyaqdiCe70wFIZIxNfrO
7fO/6px7d7JQTi/vC0n2JOxbdKV1FkKFr0kqaQ4PicpuMqBZk9wcLkSeDh8NHT/d
WOSgUt9GuwsS/JDBwo5PoxPvNnnTuIhgtIhXhJCBtz/frP3wAVxb0ET9mH/SCY1P
fqs69mRw64ssplNfIyNUsRMx3JLSnzJxL4usgfYIYzoX9B44eLZciOg23V3J0FCG
7Nd8jFGAGT4iW0yTscVCatGLqpbz4PNSs6FRQZgZZbBj9cirCPkQJubmQM0MgKb0
30NgE1lo1ts1tmqbJ4uhTf8SBZBh3dDmrxjVuJQsM3poZSoMjNF205v712VsRrqr
kS+Qxa/wc0ABdhE04Usc6CkJqoJjlgq0jojLntdkohhH5iwWJjKiBOcY6tSWEmb6
qABibdkXEx5NxGMkFMenEMUQl9xCsd7mO+6UO45X/qhMgHAvyKaDeLpzBBtwAX7X
Tq3WofC6H8ZNMeQSlCuS3rndOmyukDOCzmHpe/kHtQZ64FLrcu5nx+66KuINPMZP
jewPNsAC52Js3/8ymDVpp1p4b3HS61hFlxNDqD9thC9WNGfw1Rlrd8iCoA6FY+hT
w2UTtHN0LjM1nsPli495FsgroV9ukb0GoI4ZM4CMGdYVIP8YVf65nEaKb8ngle0f
xO+awLxoMBFoL7hZ0afekAcNsehStZZuRTWUi6sJBbKh/mj5TDgfgPsed1MXXlT0
3cgsxi6TyXXtweG7lxiPuZ6KAvzpWQ+mqKMV7hLf9ZZYKac5fbPMwXt3WavQdFk5
/fUFdFezU61UxwT1X9cBZqAoKhqKcQ6J+I025OkIHjf0Q3Xp2l98Xc9YR1VdiBuE
D/loptyLBFqzBB+kqe5cxnH4gecgQkn4xVCKkqHTdm7wMrRSZ8NZGrfQidrgjayJ
xhY/hI86DC9epWvbBTuqCLAtYg71jnb14Bq8xEpqTA4NwvsrJPV7NWdT7BxI8bvB
tjdvgIJ9lR+h0XKbCmLRAq/+2TsagOVKj9Ap+KBeRnzF/elR5ctgzw7ACpf+1jPS
qCvMYS3n9QSYQs5yMJtHVOupe3GlrvBvTTpFrJ0TONoqwzXmrN9j3MMkll40U+w/
buCcZbWccmYEubU+/xsa2/s1BQGH2o2+7yz6lnAN576fZ04G8n8YG8tZbVQn5E5E
1MC1TKZPT0zgXnjtQiiRMWrmyZffD5eGfR04goF09cXhDBiuTX95q+lM3LI5pjNZ
DD43TPl/dIM9Tpcmh32qtQYA6eYVfidaRdVCphD396TT/5HBHzbVX0vqFrAZ33sb
5fEasP1NH1H6UrK/3aI+W7wy2DlF7yTgQrIwz+MEZkJ/1Pj/xtNyrfOFUF0DbsDI
QL1ibrzh7P6gHUGNKBrJ29F2C+qTaG9umTtpmiWUNN4lrHiJ+zyP0dWah2WyD+sz
krHg+/NYF9YkRMz8zxx8FUP3sji3Zf2FVBK1b3kftFun3cZWztOC3JxrdrjSUdrW
sKr4+gL+NQyfawXxWXMxOQg+ih8gTwgZF1DF6H+CmhBK09xZOrN8E0M4lpujXahQ
O6E3+2S+dXPLV3dJ+HoKJURhr5RMBhpn4bJNEaxzXff1/6j+fnz3LiNmn+bs6bVw
wqezw9lC4nXV+uuQ/mLxkEMboArolEgvTZfjQPnVrvaarxrigb5zWq0mxm82psc9
+aQBeN3v/HnLBgWV+c+NFuC4v8tZLSD3NRXWDP09WPpStpuBV2Uso7vQfbnCgHSo
NGcf4HUTSHXzcjjlBdczsKuEkTNYGGHb/1t+q+0sYhm8u3x9kOSm7vXEiQXCvUJD
S7aPfqjZA1gszY6j8gDEPkr3sAphvSNlTPYFhTxFCG8FtFUshqds6DY+L7En1Wh+
AFuFhyK2YEiUPDSo+pqF+xhFyR6WUtHi2YPmJC4JhBoQ753TSGRLggL5gs6yl3uE
gU+vkhxgNByWOcgvtWyfnWws7GUgmQRuE9TiuuNceJP8CiwpkcSYGzZw2g8RkpNP
OQVskRz3ERHlatf1ekaqjAq/1AYiZbYXvZtquPpWMPi9rAidz8n0w2AHAAe53TcP
L+29OsISIfmqG/kqYqT8VYnBj2SvjCd7RgWgWGqB0UinJgCZFliNebSheDlZn7ag
e1Xzd508kGl9ENW9whoLqw0HZVQWrJEGDOxrusNnOywKMebMhPAEIp87GCCwQOSf
0cKz4P3p+fb0Jx2TCSnI4G1EHXiSG6ZMjfJEgfyxhUuyBcA1jYwBgyHz+/UyTqpv
Xw8T61DtVpfiOXstda5WfJQ01L5Nac0IzLP+8ydDPxtR9z88S0zNMBtoBp0BW9Y0
BjbrwGS59Wntkbra8WlIy8Ul91BddPSIAhP0OopppmFYHx/Wvu/0HQh0CBDsYDVf
IroKkqfIWvvpYTe9ERqahGm/DEXv4lHnqxb57XDi+OvemVUX5xb13iDqQb9SkWEe
YUgz8DqS2qxDRBZU1PFf4h6ihGkVMxzFjK2SoHb6oz9Ft5ijw6SnAp6MAS2QKX02
plMO1DJUGGEt8cGLvQvq0rbgRhc8sg7oP3eOIHa8zVtaMQQY/ijqfCQQ6uLoU4Z1
c0KdUX4ho7a2mMH4mq44OOH57wvZt7zJAIo1tAklPwfiqwl+pWTUNyGnhEs9jrJ+
yOp8h/i3LCSQ/Fey+S1oW9mRK4Hazmv5juijZn2f+LVKj8kxg5piB3bjn43YRDsy
33EZr9RokdNUDTGtE8vQOTs+OlRKjgtgrNgzQAAoWDag8ey+Wkws0Xm09m0MEQV8
5Iy8J2tviBGZ0lY5XKDLO8zmRG4+h+3KPdCXEwskAAst1+Ql2676OBjiJx3L26ib
sK/O6zRWWItI0mGbdmWK+lOvub53kXsiHc8vP7BYhq741am8dKs7wsRQt9jgtuuT
aAvWwUV3C3v0iKmFlXsNtOUgB+bqs3qJLeuZ4Y+x3zBNJrVmlDZqhXfq1R9UifKs
p+IRBgi0jz7LhMIpI3/EAs4KscsRJYoQ09tRuoG4ODLajU/88YzG6dmlXnnm9k6M
GgSZ2MfPor3K5DvN1RadVEknj7iW4pfZn19Xlq1xMul8c9jGUODxcoSeT/X+oqdg
6dMD7L9l6vSlmWj85T1c6+GFN9Qx5uSn0cOQSNGXrzVmMSFiJe+HHFpUwPiTij82
NuuV74YhTiDZG//eqUKcpzkDoie07+qBknK9AAEkEoG3c+GR6hil6oXPtuCRClcK
Ho3G5So/tJABkbGwq5c2TVxMDHWaxBtZ0IjwHy1o5Qm5l2gjaOvKuAY81lLsSEf0
Fsm1FORAvhmbBnUL46IVJcJQ9te1XvlBhe/N+iIvZqPbDb+8t5BomHoLkEymoXYv
n6nQFqQiXPtkTxttzXtkNWWIH8+y5euOcA4Z3NJ1KIBEzmff7XjwhzFrhuQT1bSC
mR2axOwiR8eAVdja6q6yzB//Vs2qPHKPAfsBUe3uZz+TM30Guh67F+Em9N0gj2Ao
rC/pUgcdDeeJe5zhRIm1kTzowcglaSLVcE1XybA/qkh5NFLbgAt2hJiPvtts9hLi
/+d9xnBEI8eD606EseXjWyTFqq98YPv3lUmRjndjLqEp5baWvar6BKjeeztT8UB5
sH5YH9rdXX2RyxsdmxDde6jJZ16mfsh/vno9KKOU0sEuJE12orRGz4amBS2Uhbg9
fWN/JGTVJHzTh4s7QG6PDVypmvYEBlT7yyoZTVtBI9bo32kwSSMhVHxyBLFlI7pd
Jh8BVZDD5KpPYd4ApAgvlk13v3E8VvV6ZGr7i/LsNIKqhomGdaMCdDMPSk58djRu
h6RF6X8IkIZYk8RCEEvmK22I5DzUJYccJYhk7sQWBfd/IW0Whorv6/ZIKSujdvL2
RlMxAe4pJH4j/TW2/62V2xzqv/iuYP52C47iGbiDsgeUjEfBS6YBGqLAJS0FyXRn
iw8HCmP14DbnB2gTgLdaZPR21OTDumGfajAHECTnAbwv5vFbTYQfOTiZCHvgZnSR
tkUcFsWniUQyUcODIuu3vRTbqoAmQS81kJvCDHgWDZ9agVJBssS3aK33asnxJZmB
mFulRulZ/xa8LmqV2FmCEge0aKAirBFs+9T+Uq1FdwdpOCReTYneh24XJMQAanpd
m49Ri+Ps12VrRJefzlGQKZAxYDBytv+jBg16OrRYu59Vf2oamuaeFroJkNx4gzYP
jN+JT899nlwqp/Ss6q0qaVA3a4eep1s+Y7K6nGHdexu4TaKZHyVjkGyz1OV4i51J
K/Pn3GJ3UmT42snlwwNlGgRx2ib4NHV232sIPk7zdJEFmy5vlPmywcU8dXO7r7CD
cjwcdH5DD47Ro3wcVIxX1n2b+JQmIKpMhwXizcbRfk6Y7lnwQJF8m/sX3E/pUYXq
vPzPQal0SYW2herfZVdL3rVjGKsWT7LbzySEle0pmlRRdxvIeF+kYrxmOn/hwCF4
T3CIBp+7QxT0MT1Fx+xSpAszSVSA/GWoejqUczUrbWdU1cR6FRZz6gmCxETKu+uW
vDEPoHoGHZj/EW/LurgcdOJ26BRTGHWUU1TuMHbHr4bZNieH1CDJPOJOyDukbeXU
oKoQW4dIB4dzPFRTVLUhHY9fmpMya034jcT2srpC3pgpw9I+jFFq7opXgCDBRAlY
GV2GEStFGbm/rFa96J5iDP77AAeFpUssV0/i1lKs1iYzg7aU6m4JgtMSeAQyXZ6R
130dnQ0FT++7eC2PLnzA1Cm4PYBjcyXOxf1Mp1y6PRGOAJwBQjwzpcvq3i/y+FuM
SS1xsqi1GkRbdvOWAJfuJzBXhIv6cUFAJZ1L0PsOHZHyjxwB+1MWFKVffuWZcKgL
hyH3dsh1flUgARkko0KZ0HZ7KvnbZV3LDGTLESY8Uy3yC3uMajxnOvdyRwe59FXd
WtxPzRzojtaMkoXLOWI3KXvsDAx2wNXlpnXDsejRZ53FTwei/Q5rxughHu2Dwa2A
ssBNdW77OOOjzInHuAHPXWIHwljJCfPbzZTqMg+koPt51jbXAQJWEfd/c2ootbxF
YKA7oXMa0vP5QooJiGkuQJ+gv3uoGXc2osxyPgveBfkgMMPrghMcD7jtOWX6I2Ys
MHPFFHPrQLi9Dp17f6d0/yDxtslwqBb6Jaa/eSjN49pUwRg6FHRPYNFEMZJJ7Pnz
HnwyUPT4bVkig5//T3rIkv2b0L83RYkyLsinNJXB5cpMkkZVe43W2iEBkiC84+ur
pWdNgfag93juMG1AUEDm4vj5tQbmezFnsPx1WdoSTFrHUjb6AL1Dh5BxnsTQGx9S
vWnQIuUJfK4bLWsFFBlTZUNfS8hB5MjU7iwRMgGH+NazL+dLjCa1ffZO5N6MFgHi
cNDz/vNdf012cBhCPXFubsPo3ZaFaimWQsVg3ZxXgi+HP+MrCPIrwGSSWpCXIlJL
FY1GDgju7hrVrd6+pmks1CNxfNFFJVn28mKhG0tWJYPZgfdoVSZ1ocAm/RLhVPx3
jta6ADB2xUSVgV5qZUtHAUsRCVC2UM4bM0QDBHx9w0JYEKw42DsFVpxTbbZyr9yH
B6CXiZt3gE2PePYPT+jrtFzIjf5n4fjRIbmAT0Al5tHQ+/b8kDsfdDpaYNDF/fym
S2IpJC9DZJQDQlxiN9zd2+ym/icSwQgd9EkhDTIjgIMRaHKccgccpl2tJWT+mZRA
ATOuWiAny2OW96Ta4/4+wICBqjiwW4U/yCROcuC63JQGLb3OE5QN074Hxfj+r6wf
F/sj+FoKvDNtFIVn/332DZlPAODkPUDv9CaqpHMrO56ZlJyRESd0d/HerjiT9KBP
PWunpVnKCPsrr5+id1HCYbf+NIcmptNssCZcR5CALooIw8U9wzyS3EJbx7x30rIX
aG/uSVXeXlhP8usCQVOmi9he0KrOKxwIp2CfLZx12FLkAloYbLoi27mLdEgflTr0
d3drA8IbxZEOumL7dW5/r0aBVt3Z4rtv/YxHDxAXPXxHVJnlqZNYswx5ML28IZTJ
oBzByUJAmaHB7oS/duaRsXbJIewO2NijYZ4hq/n16dKpQuQFYrRCSebNpkzXWhpl
gtQ35eRy1IAqwhaGa3DFRSBAb1VFj1aQQp/sQL7qayDXW2YtqAPr3SWQ38C1bOD/
lWjRPNGA+VOgN1s+hYi8F8JBa2dH2qEglYaPvVdO1cDlpGUhAGwcgndhMy6FWUsX
XIKJ506bBv9Mj7f5e1cDB5LXewruh2OwpBryoUPGakIPcFCWi/y/5CoqNsxNT7/s
Wg/UG61ESGRY8inDHUP0WGNXyH6zaxtqFW4h/ChEQjyodZlyt76QA/6nhbF3kj6q
ldOm3VKTEoxxnNCYpNYlGSYj2jBaN0R8AvP/wxNOSbPlaoiJ0O2f5CMYrH2At7JC
8lDj//fwirjS/DLQNo/+n/TbpMxwSVFs5+sCRy+YIkfY29GM2igdJV+oG+hNEfkL
yV8VPVyPu8SLX5C9YftmqlkG2nTPzL5+btulge8VxHLnuLlPMPm1LT4/BPLZIlWf
zkqm8tyIDdCBS8e5NU2ltQNTJ9RGeEhL/Njyt6CDBt+nwcdI3pR7Du27dEOn1nI3
maZHW1IAdAkj7sweOVCnvXOBqZXsnc8EfIxn2QzifiATsI9dOyV+UZ8nwseUdpNd
lSwmQLbJIz4j4OtGmjwPKy6JgiBLLtXZS9SKE/XjDaQpwmvsobqkKNq2YwnEaSwS
Uf9T+hcaxhU0d6QRz+QccMLuZotwZOEAsig2FTUvsH04auXGySxGUa6Ybs1AW58g
dbm8gNyObr8txBEKvJV7d4qoiqmHP7ou9nmGkYTCvuDGkNWbA1pc6fZWGD3hH1pq
uz/oRGRIc/iLhWAILlPvE0sUdFzEbVXGleoPaEyZcqm6XhzlfVIfmiz7jcxiv4T/
FfuwtwDm+Ck9nwm3HlUenRLAwZ6NStF4HENwHX/CWQhuGYh+h3arW9a/HWgytLMl
FY8hRzlhQemqMBTwDXkrDMRMKAZO79yeib/OW84M/WTGhw+gIxQwjbP9kg6ru5+1
IIcgUDTHTJInHhWTP3nEV7b1jEx3bekRf760vvj6L1TQEQ7bQP/mxMeHHvKxDLlm
8yVTRfnDoeHIkyrDR75H3C5KgSYHXYFAB+86Bhqq8u0FpqMQEeOTE7/oMFe+1l09
03slfHZigb/YmOrUGQMh031buaCRqNvUqKOnySEUDbh0grb7Xw7+LQMLb+3dMDK5
9aSmqpYlRqlhyaBWxI8NxhBNnREtA53ku9Cgmfb1M3lmASaVl2J0n8nvVRYR7XQH
MS3jN3LzUdSczMyvyPa2WGpye6D+dQmya3SrZAso9z9pDdHDBfqURKkAOPTHu7tq
C8HcuusQECW2fkUQvqmcMI5GHUlDzEDoCYEHWa1dFoiqnsapVvln0pkvV2fDGBct
AJi0msAwrZjZdxbE+tRraTfngbKQn0szF/lrOwAbAO6klEUeUNAU7/PyaE9CtpRu
HyQZAvYjH8F0GEBsdSmEqgNF58jxormo1Mj2IPvT56fDmEM4MVzKwmr3JyqsFQzB
0wKp739rW9zb/FAb0Gsfl3UAYQRKqpN8C+UMp5S0Eo/GCp5Z8obzLcdR4zUa5Djg
WZ+4yGa2EyWqFK1wQDWqyYSuXIkSN3s0O+ca7qI6TpxjERRoO6AE+QNEq+9L8q7r
HFtZKw60ay46spdtAtZ2WAkbdzXvEtlk35F42IdkhO/gYrraxKqaMbiaUUgw9sG4
ncHUKFMzAh6/yLfnPh7lZAe9T+mZhBLFChQun0DXIVFGD/p+5HlJqmbIS8DHG0Rc
7gADCLebh1uHOpFPp9s7MTHqGBPLH5RIiFxFvuFJXln5pU8Rg8CxDnJ+Js9nlIju
HILJF5ZxrKxVGCEmw66HRUqG3cU3Thonu0DfpKvXbLEO4rdSTJU702LqwmNf/76e
/Tq5KkDx4NHIys75cx1qeOj4Z3vSfO5N5/LwqUWrHrYXD8hu7A5g337Kqvzn7EWx
fh1gcYRmSjlYQAUegYjh3ltu6yBLV0rbd87noMNoPY6HHUVZALqhMn3c7MRgWkrc
Gb2ZygKq+PxKqOmbmCBnYbnHz5U7OzzctHm6PKg/Y0LbTkvHzhz4cB//tsz9wn/E
jwZVu9r97y5ublV3Qy5oRQq8gvYOU6W5ByFgA+szNguSb44bwOr6GMgaFlFosaq1
dZo4Gd+9J3W2Il7KJnq6wTIQp5TF+bR00Z82QolTfHH59zWjDQO7jj+Kmwgmg5h2
qp9gystUv/ovVSf99h3XzAVWUtEQIvFaK5z9MQzy2f6QCD6i1uIXzjt6Xi26ZP42
yihUHnvQHl5h868lc/wZMaba/w9LrpREVpLJ7tf+NtCimR3nbGeaOQB8w22jCs3c
FZsaq+sBmFe7Tb5uZAD1loePABe6m7XB4LiNV99qDo5dPPXq/qRNZqaI+4IUAw3V
FND+tSZWqmsK1SQgMqiN5XtBkfnTemUwm/ZzmUZUq9gOA/ZdZtiLUwsPQaImjWY4
wkApuJO/QIpAa83Hnd8UVc5O2ZulpICpDRmve6J2k8jK9rGKtEFiv2RDRl165JN8
9a5GN8ZWkKx4DsWKsGJzaoOnWn7YUbSxOv05CDcV6vqoFP8lmDRyCBHyNPdmlrVC
IUZjgYxiCiVK5yAhDZ8Vocld/nY2vAMK1Td8rxYo91Khib87yCRJV72NPQV1nwTT
836XDsR5AxjhR/hJA8L8g0pVwdgyUfHGlHVxdCqBBDOwLDitfEahAFRExGqUU6Xr
qq86qKJDwuoeYwwZMxzG0n6nRiYBQt8Z+JpWH1h0iD2j0bUGM/A5T3B5I6ykuZIU
D8fRZpGOjVPSRWuSRiKWkpQKDaIQDFII0WSuTokzo5jCrhuAc32roAKvDfFXIPM6
wCC6o4qhLf5TIjWN8+L4zeprmFaLbtnuHAlNGAErYtQNnQwPf2rEwydAI8UHtK6D
BY5+S3QFU6P4vg8rIsVv+AeIfA0peYB/lvcsFNJo6J5d3sThyHLLWHJPQAKqXFkq
ZPzP8dztTpGMi3/ktr+8zuPr22Rf7IBltgjdYGM/e4RLiAelkrxh9v3JCZ9vqumH
ISi6yAPUwqPEc7fxUoROA/PnVFZyCft01Z1Cfx2//DHgK0V6qZSKqUBeW21TLaRw
QK4UHZdEzvkYan9Zg1PcokxBgvzfXbNCJlRzH7gIkGYNPfGHEnP7lT7aQEnS4+vv
IKJ+HEkBSLMFtOi7SEhiPyjP2d6DQBnv/jOIdGfFhWHWBejXfx+9MPH4dH8uVGhG
OLiyndW8ygUCoKC3YPyr3udiXBUcT+4zaWWcje0sXQUytEuvAlCk+QdTfEbkcobu
zprUfVCXbXSC27AnnaT/2i7IpZUmxQEovZO9JgBRkwJgW7tJOpJVfj1n14sdMGcr
GVvdbVdY+6Xt4gspnQjUqFbEl+AoKRk3pLno4JEmULskDMz9eSn5g5NJwfYgc5GA
c0Iafrya76JN+uZVK4ZZrL0MUsRoe8zEcNRFdKsZAzR3vUxdGLoAmZkxFeN95WMz
n7ZX3ZMMWeLQsyuom7/+NOksvMg1SGrtsiYf3Vgo8jTjTJobzWO1qHkRaPgJxi+h
I6LhZREGQyVlHP/kfhLtlEwn96JNe3yZRogvVXyzUCtT8PcIQInLCe6iAAmJ76oM
kBfPCmseedpjzF49H1yafH/hvbECYOQ3K+EvUUm3dO0Av30n292YEBJur1HGyMVK
87mT2Lju1j3PxTmxxd9b9xYo/wtqbKxk8FC6s3SvPTbp97/Oiji6LW2mi/1F7taS
6Is03D336F0djSGRg51Dh0RAybtDKoK3Nwk/rEVdtcGB6jqXGxQt+czd2MkQhHzp
iMXq7E1AnNIoJVEcuq+SUZ1vgMJh4hXHQVli73MQCSAbd4DrKOb4tZDh0p5xTrfv
Jjki/X8zw432PprDQWZXqdkWpF1FmdicbgCWeKoZHSsUUyIAXQy8OhIAMIndfnYc
IWP7acWd+6wRNbMjdi/RcFvM23Z5foPmjcxlCqdvRg7EWN3ubfm9oO6roLuyXdLS
cKRemRT93WwSsVHVCezL/wTE6HV0FS7Q1lzlEA8koOCcOZoGTlqqNeqxj359AFW6
4axAgRvFxHLUiEABQlL0xhED1Jf1rWTW5pEnh1blMFtxmB/fpH4p3+BMfQH+3Fri
rtnVXTIG9D3I4nezivmYH7gLp4oWjoYK9dusd1TT20LrL8VEVJHHV+NLaRVab+Ha
LCtHYUYaGHczH68jZup6q8itklr/yFO+gwajIV3T7hi0aAWPDjlBx9miB16jO9bF
/cXsX1XHqv4TrOouCIYuSRMsbAkwdYIqsfe013h+YlAFNlW+kJaOiypqKTMr3mZ6
gibJuu1XIXrBATYhqeH+cNfwBtGA7+N6jJ8AY9gQYw9SBuWDw9jhLSb0h0wJjz5l
lFmS84rOc/oFQqrvpGNdvDbBUWZYi0Zk+uihP9mMeZdoo44xlwDSnlTqySjtPgEV
UYUtOZn2+/eXtTNIxtJ21ZQ2jjjjxG2iFPmiTIYdOUJZByLs2kJY/BB1z6UwM+Qj
equco5JAcOQNPFgYR64kT60l1HQkMC6U92g88wSR0MgLqkMNXIf7WsXswXJNeHUX
DlVnzuY3zYB8wn70Y2i8/rKxzPrx5UDDKX3ukt4VgZN3JL8XZqi+5TgodYMM0oPj
Y+HBACj2bleU+X0OW9VsFzCr2Nbb7d8bWeAgDpua1kTY5isYEGyubN3h45FOElFu
QZCvNKPzQb2uO4p/z87OXQSfq+7I7u440cye4Jn/5CQM22v4vMzq1HYKrOT4I1gq
YnoiWayIpkaV5728NnDpkVU6VWBN/PUO93qmMvdBmzKKwSt79c52f8Q50vZxJgfq
voNBw76X/Ke6DrT/a1tl0KbADxjXmRmXo/sNNFoaz9Y7YtBVmiAjlfIpCsWkbhC1
Ca7LeDF87e/fWfmV5te+N7la6pKXuFCzS1dsLIL/nCaCliq3nytHEIN3TAL0Wylf
+TXaIvxpHFXG3kChGdsu2FDz1LnWVH9FeoJt5veQJMUKkIdOk4pVIpmTkqldyRvQ
pSIXIZZMdKLUDQ6cBpdgcTouBI2KGGyQP0d6767nP01sERMnOAi7rNaAyQ48JkRo
zdEbM0my9KezE+A1xoz8LMKCq70G5PrXUggETPtRe/C2oVynhjuZLJjlos4v6s0T
ZG+KtDxC2hdhdnisJ4g70YqvNHkWXTeAt44mkr+I7uCG3lyGL8GrEe+HImmROn/S
2oaEQeKQ/q90aeo1iPU4wgUwx/MQprPXe5a5VAp5QYlHyR7SBOq/Ml9J4TUvjrh6
vzpwzP+UKeRovM4yfLPCaRBq9TBqvo3Uj1LmxEFyWhw0D6fpWBccCS8ReRY1Gxjr
wHURiHSS+HDMeCc/Ztk810MBi184T4ZhPlS4sfX5/OR8+COTtNXG5Undps5DZZ2M
KQn/Ix2O0E3KWwjdTlfjf4HD+UnRaEkmE3dh88kIs034sfdUNgjD+I1NrgdjSoX5
epMvGk9tNTURUhWwE3tsVuOCXoj2WrosKq74qU+2JUXzDAfwYXkS9buWnktjeZuh
VuBTvCfFE7uvnCaZMaarebCe3EM07FQrp4xyepCOZVcTJKRA88pnX+gn5BLAPYHm
2yjUY6icWcxrThi8INR3Me8G+rfTRv95CtR9H4ef8Em5csYPTUiwCSVFGHjgFOKB
nk0zxH32aFW3CH2wowmjLNF0RDAMOKQPELyYs6pqRSBnBIcBYWRYGF2FYfIXidPR
6MPv9xmy+qJW+P5E2DRhGuc/xkZGkWraFmFkdVz/NxtguX1zi7i6cWUnJFCj4+Xi
TyJxSv+tRUCXqNr2QUW48qYS82rNWAqGeCL4womqyfg/x0t5+oETSWloWeE6Dq8D
KwxUe/9Moh5n4rWDLE3wmtTl0nJnhuBbKXKBtba+vnXa/sAiCp8f0/pxf06mCKmK
LtODe/fya7eBwt/tlNxzTRW+FXnCAWC6Lle4mm9sQu7OhJzCS20prd5nw58nfhXb
cogoeEXSzUd0QvZOb/Gf7wZY5aQ5StUA8NrnFeFAtEI3msJszV3/EBHMzxkqBzS2
bS91Q5on5NwFVC0I1AGJgV8opC3krD3BMQSw6WdIhbBLubomOxzFs3FmFAJcfe+C
zp7j5sONRBehOATTNeNwgiHHsAuwl9vsPk1ZTeQpXJrItZ4FJ2ifPlALQoLmMAF3
acWXgveCx7CTa6N04YSxtMLiptcdpO7KBURhhtSD7iqZADCVZ0qOcv6HcimNeXl3
UiBvSyKFS5Tjk8iVNZpeUWbLvlIkCE4XSPmuCQTZNnMV4+mFWjY83GPCnB3oaqau
U+BCBNyojwynyXfxSnGrW18nD3U/+Wd7iIy8CQCp7ZPZl5O7R41oVFeEIRcz6Ma/
Jkrp7JcIHhlFFjD4qI2uqcKoqWl5zvJfqyaMXZ3YqOZ+KfvkrWq+2CAzHD0gqX/j
53b2aLD/p1YFy/wG87XpTKL4n7sl6pmhbQFzkD6mPq03slOMhX8SmykpFjugW02V
94FRoht6gqzliPXURINL9EDc7/P04to7E9kHNBo6mgeGZid3ffMQCgZMGjqLtYJW
dOTaPtvtcZmrDSvh7GUO6AOZiglGr3O9JVPpbxRw2D3owqN97HlavOH0ldMGsTQZ
F77V/cLaH938OUVy0pfQLTxClt9/HzmUPg4ujhGXAaEx1YWvytaXsZD1JUc2kDqd
j7Rxb1bM5c4JT29TYt91KXgfSn8wW5HdNcN0IdFh3Y5QUeZ4Z5Umphq8VJxLAImI
MGFKhwlHsq9dNo/RWSIC0TOx2y8/K80mJZNY7eRsk+YOec0rsJU+vXSwlhr4IIq7
jJUy5n423VGSYSdi2V4x8yAqXOOGal8Pog2SgkFo/9gtMu/9Nkmp9L4LPYtjcece
XDWorif+NKNRHWNdsiYUh2XdM2QQq3qGRJ1TDgovPd+9K9cNpRqNU01UuTFcQyaE
h73T6w+0CCwiI7Qi7Kl9EK8CaCXLyS1dR7oVhSpVBMsT1LCdWWg5uIPTi7hYmXxH
BVmdo0UfV6VOlshRPVBsn15YSzptJ7jM7/g4TdaLCL1KcI8xQrSqRjC9JX0Thg33
X1Pry+axXksM4fbvLuATaVPhQtL7h7wYKXJqffv+MTahuGJIv1HNXhjvjCeplAC2
BVka3CD3EsomSU7gZpZdBD5bJ9GEd6rcuYf/3hI8QVUg4g8+yfNU/xdTGCq41NVs
zlnM2TYxlmve+b8UV0kGC9iwRZWGuLCj5StGUTSPOuneQrrVuP0HEqOXJeTXGzk4
wFPxfK3nUgfq4cMMrosS42vQTGtVuXmPT1NzXQQkY+ys9F+4SC+/E/K4sU/1lHs1
Fi51S0xb6eAq2CKy/7LpC0wlA5cWfyhzKGpMgDbJMtSuDRpreyRqKurX/Nsx9H45
4ZGS9ERlv2ykl01AzvFO9qOCGQKt+noXrBDl+Cj+wTnFCY6L5hskRI+t83jq19vs
KCWJBLweyCI2EfjJi7ZicuH5fmsECQ9njjkNs5tR/f/UA11IlZd+BCEdrZevciIR
ql5Wqzgb8zu1yukyG8Kj19orU20klJDLzzrwo89qKrYiiGH3fS5rohrL7wr4drNY
PKosjxUIAJ8RJvniSTy7tWSsFh3t16X1rUu8+K/pxZiCOXtiLs/mev/X+hoTTbFg
/nIJHniCKGTCAQk92i16WFoGf/qgLRybEePotIlaDh9SmIBCBtqi6no4XHTkD3cg
nXhKACBNn1X57RU7k9wmqCksUoE0XRF7TLBkSY3zkWPC5R32Tr2+VDLMi7tG0A9Z
ng91zN+cFvly26gtghf20VWB1ufLpSEDmaek5+x1FEaMTOKKbc0B09K21skWi4L2
0WjuCuMjYD1Io5GcxfTGewoKPv9LABe9hTfeQhzaa8pK0WZpO5Od0zhkED7RFHau
e/x6N9jwh7lADLEIlNUa4u7kfPXf4doSekmELgsd48rTV+H54zvGRmYxf9hl+eNy
l6rYf9YrfQqnOu0THz9XUbYvjfUkn3W2vxOH7ToJEESbnd9bryxiMI3C4ennPISq
Jy0+5dgf85ergYXXnDjQ9+fR7KyAE9QMcbyhWldjsJR7SHL8oZzxMiIZS8AN2M/b
TYZeMZWt45DdPWF2OKIQFEfzbLCGdLn6qpv5b2l7WLawA+zzgwFmCA3EgoQoCQF3
n3gppAqGg1BkayjFd7YFXMegBDWIX7+JS/Hiqns5tA+nk5BiGSSmziBJL0zXBGXQ
1nve6oDZjFN1EcV5OmjtntIUdLfHswbWuzRJOZPNmcDVj4oCfkwk3tRmlpaqmiK7
ybsO2/LLyfeM36UvsqJnLdyYnYJH7bxjkZdVZR3/HzLEdJYnIKptZF70E4IWMco0
fZPmqqSYdRllOsxU2kexb0SfyuiN1VHmVYU7N4OFp66oHgegDRr8vEAou8S6ITwB
hnQu4ADJ7JxyE2p6w1JAbOlw1uBudxNEy+P2TNjo6RDEvMS0LYDDwoWkpy+DBhKf
mH4HNptkjBb/J09uTVh13kUP0Km1T9AjbnDxzv9sKm0OatnyEnoZXAnc+3ClF3pp
wo/kwgSSbEsI1OyElw5vaZjsJxoNsDesPQWS7GbEQEs+kITi9Sd1jHzDrLF1syY/
yfYPItss/9j9P2SA3eeJ3X7pZKPgZGIJY7ClrumxpDjeChbWKDpFctGj8COuHk3u
OJYtbdke7oe00UCgqSF5YFjyZDh8ImpYDY6Y7JzlwUZDr33abL6kgQs2T/CHLiyP
FCXzotEvJkhJ7wqolu/xvc7khSVEElvO0VazPwdp6Q8cdYtDkANDLiGbeRjMhItU
fdwXf15EiiDQ9MyVpWD/+3mMd4bQnD9IzXn49Oykg2zcRNEJQdc4IOqXefw7yMVM
56dKBBuMzLtgxOpNXIHJV8B4nntxgkN+pHi5ZPojtL6nU2u9wr/3qT4/6z8X71s0
ghvmjlvUe0Zijb5C0KnGEC54SYzXJBJ2wwNoiOM9H3Zt7cq4keSAvu8huZcq9fAY
tjSVOhRmJ2+vmfhkYqhZ5DYb/pWF05+THo4uc9l3/zUbl/1sQamrTr84PTxfC1Fv
7Fl2ATtNEp7XKPRe95zF+3MLRIZcFttkjOQaCAfdO7IRlYvv7wquHbDYHD8QGGEX
thfna2itOxHqMkVhr1gRTuigMvqlu/njNoWbjfdMW+2ccTSYEq4gbEriccwC/omT
wH+tBr76QqgkndZyPOL4OEXebnrLGftYstKx4FOkM7c7ANyvbP0mDxOgD+gSpHwL
E0R1G5m9IBIP1Z3YL+CP9nin8T/8LPYxs+11lEhlqRPhHnN1FwdTNswUa+4T+o7x
mFJ03T3W9rblgkfG7mIJfhaarj4yBXSAaJFkWxtXbhvISTj5kQOMHRcxJG9yUVc/
1/7IpzQWnIqPbdH/qouOnEwGpH+3M7jp7JqtCge9SuOAbdMzHbeycRMRnBPkfvZm
wbt3rMewk6Dor5vlIQuf2S3JewJve0Kf3OL4W0tnONqrDmRiHI8gZruK1bG33STy
HCB3p7KPP5oZrD46F4J90ZMbLad3kQVSZ09ykyOahR8Rzp61Nk4ALINvKhpzoj0D
i5e9HcNaT0BBk5xUV5AUW9z1G1W2puvhVuFRZ9slPlIKFeSYOPvRNCyNOHsGf7bF
KHMBuEPbKA0Sq+HwiKIJm/ISW69R2MQXpoiRKyACSPlf2CVbxpkCP8tBgLHYz++m
TQFWZooIK5pXLNWKOMjbIvAFK/urgkPkZRg1cuxlZFllndoMams4mqvbv+tQuTJp
/JHr0GBstEgwoJkwuwYqDIW0TyIQm6oeSwEHuxg9mLDOMeW+WZrEWJiMehZIoOYY
MSJwT8OeCbxe74Wvy6G3aVOeZx13+qxQZWgU0e8uNIMvz+e9FszG4JCzyYA4TqZJ
RGzeRVK4XlMghj33ptfCS19aOF26nduGgjahg16ZqUM9/52S19XdSuNrvcMuPp/Y
GhSrMkLcSWPr9Uer2R0JUF2LtW7zH0eX1dPoU+/QR1FGFW5fmGV9NotnoqmThpyY
Df21UHDiTm8NvMIRWQwNxrPDNRQrQRHfmns970CCrDzLHEfp95LASALHZBAgAgbq
vWMDm5a1Bdj1jaGVPHf5+aplZMcFHC3ESHgXZEmZ30Nmf6XH58lOczuslrlCwLyQ
HotTTkqUoqR9MxYvI3lQxI591YtukB4/3Pr3aPopfUb6PPVzoKNL6cKuhUC0y4bo
SRJSG1XHDHMIRwptDMUAffPgO75AEZDZOGFBGwoYLuFMU5jRBT9col3m2u2+h5d2
uWABOuKwdoIUTy1BkaotxUbhThNLSKwSEJMCdppbQk2TxSeM5u4iPglebNMAtq7y
JjoewHDWvvkoZMmND13w07NsuP7P/sKRsJcqGX44P4enGFOkBhSMK/lHRUqT3UF/
AVWJnpqpEwgaiZUOiG14wjkcqxL7psLB75W33PrWrmWjD8OzJV6y8Os3g5Qa1AGu
AOnNkT5D8cxRh+SI90RCBESFVJV2fg1X4p5/x1HDuPf7EpvXsQxGX7VV/YIUiyO0
OdSDdy6wLMM3XVsbcyxkztFaShPdcqsu98Sv0b3tLO8gHKT8P9r1jnEeFxRItUxj
yhdDnOd5Sa4ygh9IAHGyuh3Ek1FbEVzOEz+9n3OATGLl7lpAgSc6rsG2BGiGRp+f
kUJi1o9pT449UHl/KNE8bLYvAwxKFC6ZyEiGvbDrrB4Am3PQrhRJcOoLUu+dgetJ
XjjVYVYDbMunDzA/VopTAsjLscU5+llksqeI8Y3hzZRgR2ETiBQ6cyN/TBHFRLfT
UPl9JZ+IPhJ5Loh+aZx3fFLu67glEblLsgQAW3MtKicewLTKXKwK3LrMQTXPjdWh
H8HxnCD98t6mofBzKBJS6ByBO5PW9DdFs05kwMq8r7pABRoMpWA9ozHv0vFxwULk
WHOQaRGPQFRiXqd5qppDCBz7BDBkUOAToX09Jh0PHSbwlIk8cSH/dzGyGjk5nbwN
aUSSs3O6yaHsIplKxkpqMGasyGldqpHlK0xFWUjYkW0TxmxYEjWckqnIg5acWajR
hd8TaRTUbCsbMc/tuHOSGxANwuIHasEVMp+XDeFooW6fbr8ezLgbYgyLPlgIv37s
pCK1S0yEEfngDkTyjr9hISeByngHQh81eb7JcRHe4sktt7R+RyXz6DNJU9SlP5FI
kzX+ZAVyLdoNpSOTsb6QWmuio5FU1ir3c/9PEyEwirVvmNs0V2IxfB12JFLQZY3l
geJvQQuKra9E7rcd73y+rUlO+tu+ojRWKl7ooolObpL7e5FjCL/tpoHHWZHmGTD4
MtOfxuXdvtuS6jcgiOmruvCxi+qX0K27m1shItgbUF/2H59sB3c9xOXpm4m/J2Nk
HxP3F69BMJJ5G6FbyI5pCggc6d5mi+E+nJ8rnZlkpBMFyecjV63kMzI+A7EqXrWD
jbZAAdIEtE+4Kmq6hLhiYiwnnwfgoFIJQ6TSq8vg4dA7o9BNaId9An7ODfsuEEIL
ae8ipTQ99Na9sR8h7sDuEjgvp+RTQ+Prs3uEbmIx4N8oxNuMLiOKFeafgDtI5ipV
g3Ew875YTp39hIORe++D/vbZ8fVDkcm2Vr05ZucqcxQDtwqMwOPTh81O9YfImhh7
SMkVimcryTNV2qatKZcihuQodWRAF0g9d0I4c24fV+47iIBVqX0kO4EADsneO+Ik
5fHmfw1a6yE163SHAjxZW8P7NE0KS6oiKFdstG0OzQTaoDgs7yqpMU32WYHvcrOq
Nu4PpRvYiiFRhRRpEL57Bb4AnfqZlJB4Gppx4mfKXBl168N8cB5EE2fFu1vl1Q0H
Du6RfUG6kkVSsJJRraj4hEGkiBKSsJ1iac95IhWU6YpERSuqCaV78rzVeIqVdzHf
sNZeRKhV9JVxPP79A4kVx8794+oFz6fh+6/uC9S6IWi9DWlpz78bMznNxcDZMD9/
dGvbrNyilfa4tw1eTr2MvRabIP/4iUL7ZnZ2yKgjpkMHBOiLBlR5+KLueCoaYC5J
bpRqzz1ZeqPVkU3lsTC/N7tYYuea5lpnXphZsJsVHQ3QAJpLSWgHyf6C8B71ydXb
53uL/k1dRwp8EdpUbDk99IL7SGT9Uha9bTofzme+1pa/+QnqzaRKFxN+yj1Nyu1/
pcah97SMnzuWa43V1KO7cM86h8N2NVwksVHbsGi7kfO43pA2wm6bx7TiUkRRCGDx
g7HovPBdkiTLj7ORYnZLX7/VWboUVfR3wmTNGWiFGIRfHhfURU6u3NnPazoCwpCg
qwfeL7gpp15MdnG3iK7Jgu0r7Udc1uaSyiMChK+/KHxb2rkeZLn/jnTBohSbpCub
GqQH3uDbxpUVGwUZ9mm+h3istqeOj4aj9OFmLWPEWOiTgHSgCOaJYZFFdzLNL2RM
hyY/AIRCAGT0orD5EDLXK06H/TtiaG2KB1zdlCdE0t7VImGHV/qOYRobv/EqxAPg
T8c6ATX3lx4wokF9S32wUOgwc6WuRJxXY6iDrFmO83qRTNT9zkrbwoFXpqQr3JoY
5FTbWm2q2zZ0wvEHg1e2ubxi8JCt+P+2ja5FvJwwFJ0CicAFuXNKUSlUn2xXFmlO
0I87Zc+zFFr4IXZzkpE+JGhuSx3hZ2mE2xWRvo39xsv1p+qeivyk2ww5yhWxzDIl
X7YWV2lEUdgFAUORHTn8K2UfdBa4aWn+m5EqQ8y4fa0VI3dFeR3rlfksPGm88BJI
fhPmePcC2ArxEpbzjpkss8G4hkE/yJHVon3ktfqjseOTLujyoPDx9Mb5iedLKWYm
24uBs9Ya4W8LDtxUl2G/qRwrlWAwpUbWhzDm3Jg9Ci60VAmNMyUpb6qPZAPrUtp5
I5GGPemEuJ37xPsUAXNKD8mYGm1OqreQMpaAjnc1k3JWiCkEKJMfU+j3hohO3iq4
X/nUJEeHxfnFUOWb1aCiaJ9vd+431koj1CpSsIQmzrWwVAsWN+0mGdpaA7Q+0HRc
ttmwCPLFdso66p2dq1aMiOgpbbR48+V6V/5FBrRMZaMtX6rL7QU/s26LvWrb23hP
EBI3I1ZNwx/tCsYx/raII1saTP6ITQiy7e6+Gor5wm4dCO9eXqCIcw3T8s1pU0t4
WQs1ROs8lID4WwEyRbF2Loeqm2XU53pRlrECroPg59ObrrGpkJU6bb1B5jWn+DTN
/j6xa8/qSw3UbAtl4uIT4A8Z5yqR8Z3VbVZIiJxeYmmP4I96o42+kYrAl3sZOZ+i
bFq1pcI2ToDa6WpaEparXiIESaBY5V6LeeZwvVUyFg5Jw+UbuwQodeojrCkqP3Kh
3bTn4njPsmTI7trxVqntjuQP9J/rtO4uQ2eUfp+Dnyk9swVQzT43hVo8fPmPOSU9
Q4wy1FKWWySKlZRtRa5T7HkbwHtlmEN0UWcgBzFA1RYh6DX6DcNgkr1/hSIfH4OD
byo13/WucWJRBzVDmjUkvtb1nQ7fR5bGn9kcR/VtCzzKzTPxy2Mbdh9U8N8hayYa
EUFAj4bHTomlkRrkSEGOWdl+y/iRQRxTEgbv3quEabEIOMYF6qedbPelWaoxTg1V
rCcxAvrnCZjWB0h8J5GXgPVDP72ImAtMQGoWz2mwEb2P5WbwJTWyU/aHLWgrJ0c2
TtOt9U0PHyC2Hymqu3gZDPVkn2BcD9GNMvMtdFKSLw1vfOXqCpYVGImvNB4UIWl4
jstW0Dw8aZfMgb7wPfrBp+JuHnV9nda8pyDvL3gt90qC7DsobLCP2Llw2GQFMfI7
F6foyUd5oAtzrYMSga4ZZ3ae1dpVOkqf6Ebr2gPNBcuHDz8LqF/ejUIsbcMW69Rv
lmS4ewma45qXFILvJPslq5jNtuvL9PbPbIoqVrX3y6nu5+xjDU7z3owBZNQ3tZTs
3xK97cF4gjs+BiWgEyCEDnjffJtqnF6C3GxonfoQxlNKGE/wNLLTBiC/Y+QdKg5S
CLSbptJ7YAk/BMxwZCgSrhcGVbCEfZT/QgORAnhDQZ3jd9bq6xXHwNSOSl7NL1QO
4uo8Zv7cUJRuqIyVsIHm2MDqgjsB5jZ6G+V+093UuQXaymaqrKa4W4aevwQC55b6
hr8oJO/QbzoX+4ByT3jiu7ZeGYNBxMipGSTou5T8gWW/crsroh0bTw7wFU/uhpI3
nPZwtJesHKIrYnRfQkZ0gq7ccMrkkGfgZ0JDKckO2L6R+en3muawgekh3oqdVuNe
MMrt+DQLMFOkpCS3zGXzjyBVZO8+nTLQNeAmuWwlsNlGzXPudJ8fH3LLxnIGIidU
Q0bcTEkbHGEle7yCqZNDobQdL1n3281leD1NchmdsOgobgGh1na1y5neSsb8D/iV
7e51x7dHZhgztCjO6yHmEpMxRPpaSVpjeytN4Sz89WFs2uISZtmdaugE15qKBPng
dF/KAop1iFgtHmgo0mkgPIzugehXVJpf+3NRkVSjWjFcx5kAY9mqmF4phezIqAsU
L0XizMs6uZIPLWXRJzl+z1e0MxWsqVXJTjxegFpeQmSnhnk9Z0Rk5E7Kzgo5uaSu
Pw6SKNtaZgzgkOfRI2NQBUWUpZh7ks2V4Jrx69VkHCqmZpP840CYgq4yRPT63OF0
se5TsdEOXulPhStPJhiEORLro/umlvzL0zbDKrpX+ujiuyZSq3bTADvl0pHn9AST
aJA59fUGAsQtsBbbDa6VibU3ilNZQempfc6z9JUjr5QUM5Fo2fvjcQ7bJkkCw1YK
mmao42btPtLq98It4Eyvq7apetruQX5x4I5xAL489KhG87dkCyNzbg8FbcQOEwZC
PG/+GiiqC/kIdJxmr/4WW5L3yOys2q7Dp4szhinyfhwz3JJdEdop6j39eCD3kVrO
YQYn3ZpP0B50CCRPf3+a5KZX1dktOPWfO0Z5kK0Fa4jDwOLy61bCe4XMsUrm0zoo
EsWo3jQVSYFGCm5OYqzcj4U8+2uIS5Zf3A0qQNjnx/LG9X5x3evS4kSwgXc0Ixpu
Fchqx7aJ/Z5WiAFy8Wp/KQH0b6I4CPQyVoCNZlUgQOHQ0wwXLQiaYQgcwUrF+Wmw
eTCzUXAUvTOC+oOE8mUtzPdwMMADT9weLMcAoMzKbbeem864KXIY8wQ5k/Fhnx+E
22mg8YQ2Oc52hjlbhnIxeTXtigcz2JT9e1amsXkQyjvv6BbFrtPVZxZuED43Pf0f
U44I2BwCscvspFjq2dVRIf3jVZ04Fw/nbBu+rz98w2Rk6rsyqTcYkUZPRy2n1c8Z
TJcqrqJwv07sWyLs0E5B8aRFm553YLkEdjQyVgFDwtpvgYIFP4OQ7xPRSeKP4lZe
5dGpwLjRg2pN8tGLQbxQhCUNoYfiOxjQv8EqoXQ1PPRt/1jGgcs0/GV3KgaFAhQg
nK8RXwiG0ekvN+Nud6XYTXtpbg1EtC2sgPu4r7jNuGd0WosXQD06T8KuJfmrYUEp
5Z+quuL1LgE3l/KKh+kblTtpG280iQaW6ynrAkJYIrNzu5XZLAmFigUwSnYMXgOH
Kqsjzf8IDry+jL037gstY3YsDuXN8iDnFOn/a+p4tTRPYDZIYTR+HHQ4tzgvNTdZ
FiqkzvRlUCvApQBXu5Bt1vP0RVI9fkbIyhDw0CTm7bcKwqygK1Ho635+cIcTAOtd
s6X5tMzm+xmIfF3v19Cxu5PuFe1tQRXwGOoi/6VsxiLGM5atCG25FikUBZOu5AmF
4cZZ3OyQq2ZEyMvOc98XYlObGI1pZPaokVBZeZSHcmBJ9h82JmRfGI9uXGgE7Hwh
iMpPah07WT+bHoP1PxjFeBPsdGr1pcUk4QZ7aoW2rRuxE/DIiUU/LULDk5r1Cixp
uTBlHE1rB8WlOtWmlffXTLQ7srKgfkYYkjyWcFv47WuCL2epI0j/qwdRDuG4TMTm
WrUWIcCZ8buTzegdddUqqBIkf9ib4WveC+a6tX1fukXS8RQ2vMS7+qNO/HrUF9l8
McTel1vWvYkGlOdVS3nVyEwijhinvkVU2LiCw+jxedHh+zv18SiegSskEF14Qy60
T1LkZZlCmQlSWdIljEtK4lVgTGCbG5/PvNkw/tWB69ijq1q6Mtj/aVZAG10s6xUg
CDPqlqvGG/srR2etW46oxb8SDA53ZHQELDGp5G08njm5BFMq1KEbLk63ljkGUXJT
I9QfpUzZDSUYNX1wV9p/BPicODaHHMQ0mRgjLSvy7xY8xKNjrHeGdvRXFCw4KJKO
3hPPHdc2w8RF5PBqEkw4Wm68ghDsI8vNr/Ij9MYY/d+OhKh/zCTlj48pyWZJ046b
yJ2JXmGh+858aADZWhuyaooKxfxe0LUGmXp1q9m2qDvP/6r7qXwFVMFmMd/nYJ7Y
r0w2PFLe9ZzVJmvSQdNc2w76pluJlPSzZDHVbKcnm2zscd+91Svx2U/tZu1yHlW/
a4SglIQFphrto3Ciexw03XG+1gmFnFt/MueW4HHkoq+hcdfHmCLxVFw/MtatfrKF
sjg4ZpstPw9XHgk9oOH5MJql41UEWtv5lljVDRQbI2UPmYrOUlWXfLCXuwUiwrjO
FkN8ctF+b4V0ZPfuAUKCIbPyNGUcYEZCByoAUT6CSWFW1pipk1v1GzsefNzYz5hB
b97y0xL1qp/wPuCUKUEBwaWQbGD/vgTDOL5wnq+hfLhUwmb1PznXnwyctD/rxdEF
vAC9nYoFZC0Wcm9/ktXKTf4dx/saDAa90mLO5aS0T1s0uZ55PLJyhStnyYwJWjFy
seXnX/DoC90p/OY/5Ppd0kKfKCgDvP9dk7eqBXrgKoZ4XOXwvBCJAjtCT9jr6Cyq
A1cscQy7VZvFFxr/9H+S5/zrvtJdYCfv1x3BzlfAE947qvEaO79WvsebFY0f7o3K
Q0hhN2DToI92LKsMKQFT2iQ0qyl639oMonH5E9UNeDDBTPTo4hGZp1orhPTh2i4L
cZaYf57J8d1jbOFSK1jWXXVewJWfGxCDhMRmaSYfkRTkC8QgfomhvKZdfma/2JVB
2YDxGdhR3b9lhmtiIs7CLI3T9O/+BH7cdidqF4XXPwg1d5YmF5I8dlboQHm6exPq
GHhniTf0TUTvelTAK03EDhUa9zemFpIs9vjFUpG0fnIGba300A7bVlbhrq8c8KcW
owssQedGvzkk8v2445/mllSYtrZEN5BC0jVoxXCdmNSVKox0zgdbFgCzognWA3Ps
oa1Un7JIMAWCU3hU2CGAngMdUTtFZb6y0p5KLcD6gSEs3fdxlGF1B/oWMgB93Vp2
9b3jr1tUqn2uYVnKxcEO7dOIXOYyKBzcpBHS/Gt6hhi4Fgnx8z5RdtQW6jKhd18G
SIOno6i4WU1ZgLw2OJ9fnDz1JuozRWUWv8GvLKLWEAoOhmngzncfJ0HNbmZ4EQqG
kC6126XyDQSjLi+YsXvYlMvj7BEibMZ3TqB7hqnProX1sBdcmPCnm/WR3TgTZuMM
Zj+8MrPZa+VUroTovUYHT+9Mo/L+5ujzTjb1459JVsBjzVoO8uICkgbxYmoT0Pyx
ADJGWuqlE2CVnxUwTFmC4mkQakHqBHD3Sv5mnofR7uLRU6nOX2Gw952X58RdW3Ox
IeqpoXU10pMuzhjQVKkA4aJiKUxrh5Z8JeJFmxh8now00u4QKX8Ccgd1tNU6xj46
aPQLoiFgmkcYAPiHJPnQp2fQpN2MKt/AboGGCfEbXEpO29j8d7sFbtEAXfhPtQ76
gQJhq7WnyTpH6VS5j2lrOyLO+XtXENyqTzqs0kK1KHuNaWw38sqzu9UnPiVTwYhR
scrnr/fdls8SMXeQaLny2eKEISlmMNhjHoKdhoglas2Ek0wt8FEtqpq2iBCbYcBo
suS6vdD7Gn18sB8n+toia2LMP6WLUeq+lT6SLS7PnMf+rpI6QoT2ZzcQifk4A1Ij
URIlHalIzk3awlQnosWuvAer9lwvANCjJVFGVIRuOdN5Q2n0WpY36FS9Q+R2Pwff
6LZ5+hx6q5oIPoMG3Xt33mF/q8XyCAvIDLu7xCIqZ1xoKzjDtMJkSuq509zs+LVz
FNQDTEqQbkkF4/WDtHWhO2gX3IjNueVIz3llArzgNywfM3nFsHfffvC4m707xTrG
D4NieZIlxlrsgczUmZPuc1Czk8LYgp/byWHJbof3ieUn5hjAj4J922emdPJJG+G8
xZyhyuXQA7DOkyEi+QNgLm0SrcVc/TS/CRELFtoLRsb28VOAloWD3x4IU+VQBIcN
O4QDxeCbHUoyzQlc5B6pU21SzkAJNzIDOBBvH2ZAX+QwNbmqbz59wBzqx5PMpKdU
oQll7sVZl3EetpvsZTIrPdX9/U7e7azTghvhRvhgiV1PDeLOc+Jy44ZBUmciKQvu
M8F4YbRj+VOlLaEHmO7TNA/qULsZdD4dveyZ2pafeHYwfIqJaa4CwYM6hnT+SMid
QhkJ3btoSnIv5u9uH2lLifi98xhC6jnVfegRqzkaWF+5/uGJIC6H1i96NSwcd2Hb
Z3V6X2Gq9C0Yg+4mo330S9lS9QhVQ8vYX67dliD7iVtHnTrQeBceNREl94vHuOlx
S+O2BmAsbPPASzjLhdxZXqU5HosCT0oKHxmPa3CiYIJZnoaDRbfwGhAzwC6MnZ97
vvmGCdrh+SPAAVQUPipc93vKRjKTK5ePzzBhFiqhul5AWk9mQwKlOdateLTUdqYN
ee8gS9zjrFV5tKZLT9rTxQjO2I/rItk7AvgtF4HWCHmzKzRX1n/nyXh1vWWEtxGq
fJAG49XS1IeJ/yvAA1gREWtcho1i9FL9QcY1vprRWB3OH0+UpEm7Ubq1Aibej9fA
axNcHzLQ1TBZLhd3h4WOG0XGa729DXWgfHO6xnCs1hopIj3fcuqmhm9rjQ4HPla2
HRK9+LuXnDzgTezV3eWYBHavD/UF7ezutkm88hh4b9Ak0PrFgMFPgq2HgEy4vvYu
E8R9b3/yyymQEHAdWPUO7rV8PXPYrNuAyJNRN3ffu8FJNLJtPUrxyNT2d41FWx3l
HnEQFZnzvGlvWgYMXJ/oyiKW/2hYWVjcfoE+OMgX2fXmY7UkHuXp1PBdA3Dtb96k
DO6lGtqmzv3wiWtAw4/Mh1khUVKv/2yM8UjFz5fSCRcEq7SN5uIjDwXyzQwAQ85m
sJLLeXLDVSofi6S1RidpqHEarQo/71/hZKbdYcXBMTEgigmUXzPY+5LGrGUMswxQ
VdtZbcOiVEJ8+l3RGSrJLm5egJsMH4LT2WSYtF260Qdah1myqDlsQWBBLZqac62y
lTxzHMbj4Uuc5lb3V0aweggGLUI6DVa5fjzyHLgv+4V1O1xfo0pOTBCMozLPg3tU
jofRvk4o7DbDe+7BGqV/j2xD7/eZPjz2ETxupTUGUQYZp3xVRL0AhiHKHFWqeYp3
XtzpyodxydbEkmdMQZEEUUVJDsGbfsk3SM+0GLBAKcmTtMnZq8loVW1F4IE/HN3t
bg9XiFvRJwYwY/aasth0f+j3jPwZo//BYFUGgo1BXNmj3mVdICJFme6uEfJtPTlv
Go27naO/0om+jzNLAdrYxGu3VuS875d5tPa3Bcbjnk7gGslapaCWlsrb00Kjzh4q
inBtsu67ZjnxwkjV1P0yCs9U1u1leZm7uELi8ElmVuxEUGMCUAPEgIQXP6LPwkVR
/oXkVGCU7PLVqggbUvfypAgNDpSUBi45rfYv1S9Y6mGXmOoja6WpIAlIMthGobvm
dkKLGdPSRWUokVR4wjQ3szx5nO0iViwCvV/xWDE/k7ybry3wFWFKKqDd2H4vkhxl
BBRfXZyNzdJi5VDJ4j9Yx+FdW2ddgmFoqGYGQRUfZ1AXLGCodZKrTx5OJK3WAp6K
FMfr9FQlEK7DU6+4Urw8g+OxTUA+q7TrwsJX9Wxoo9fiyXuV1Zx89qzBKUOe+BAd
DHc6TAfIgPFUwcjsiX9vfpxcdUH0djoVObz9qLScTM7VdbDS0lfant3KTxqxkvT0
JHk7gSrJQyFZu/EKgAtHAZPc7aq6WhQT7lJ41W3xBm2RV/fLFFJ/T8pHUz0YNASO
o+0ggyFCUPKRHxerim89BkTWV9uYbHWcnZqyNIlc094A4mFbKV4QaZaFEpJ7keaa
z4dtB8fUj5K5W0kmotWMgTDboxAHPs0WykBz0hHHjt5lHFQ4POrbYjUe3LOhvR96
43JYC/0uRv+qyoaloaf2y9+aIsrEwG71tEj/q8Dsgc4NMUvN5fpZTYnuM6t4NE2k
KNk4vT220tV8ZrTT8LjevNUT9BWFuHjgaYeLNPG40ev15yqRdXss0awV3iPhD6Aq
QG35aynp4eESmYonrUrkYcfdJvQapvMt7nzsJZJctgEu38+KB9DJsDOrOym6X4Kr
1fhaOmlnLrwxjL/pD9xOombvsL3RkJg7+pAMWv8XGZaLBSZ4wt9Kasn5zsDsvaRa
Rlnz5fRVfM6S/1n+GRaMz7Q9ZlvauXZCKLqFsiyxQvCyBernWZnxZz7O/m0kPo6u
/K1vcabWoiGC2qXa0P5eLhXah6xIrGMpcowM6/mVpJj+gVhCptEGmwp9vQRgLAya
a+JXP5Jf5Sx5PKgA5kUjmcmE/fhKzYNmwZ8WuExFefn59Grdj8ZHF+RCyWiOg3Ci
j7zF1pmyCN7ooAWXJ8CAi0QJ/EHLyH7HU9KNb2WHgjjtKUhhPUOMLNTvA5bIU/+G
0WS0roCgw3Rnh+kwfpOv92jVFuQpoi5v4q432O1n9ihehzE/PDJPhiqYPQmznG4N
0+Rv9OMz6+gJjVRCXZ/vUGLPfrLe7YkItO2HREQu4n92lNTFzro7El3NfSMvyWqe
bAOqD6juU8hAaNh+ngx0ec3usH3V+OeyR67+UYcUGzM0f2Uz80+H/z+m7gcY1pkd
I9viJutGIPZ+J8fiYeOxAnOWkNBzi1rB7LxhHCpMpqX0YhCmZsTvGydD0FSUYJrL
El+DLrm8wibswRU/e56YET7egNkD3h4ltaFJ3wv5sXLIlcaqjm0WWAx/7RLJ7SQt
sify2FtVwAU6u7+DMxQ8ABnivHr742uXlFn7LKZxk7AFwPCrBLtiBOEm/hpgJ4B8
EybZN1Q2c4Hqxk+nBkM0IC+EQyDbRly6pBT6gW4jcMbaWYU7jmLr7UTGQaZMHNe0
fHo597IqWLZhhSHguXM3S53O2TuVrFkTaDlFNPnXonOoPyxwqS+mISxkjoZjpDlq
R6pAV4TBAp52Fsw8u9hSY81Ji9zxj4OvLMezRgaD/1Ty9wonorbIhl3C8qHyYT7/
G0d2xa7LW+akAXuahJJs+bpnAC4yyxgutpr7BMuPFFGHsZjm8t0cBHQq3Y5Dpjnp
MDXUoE1qHFux+r2YwYV0I2h11AmBjv51o8+4AxxuBd1ia7tGqSs2/Lnwws8Z758P
dUfOWrDfm54fCRzT5gjeivN0G9kPEu8a96ethBE/zGffShi+CnqhoMRd0h1eITqm
HMsep+Rj89K6nx43VmYOo9xn1xzauUp7kwb0NyWYMPiKjLT6kt6d0eNt5R4yrxyU
ZaxNP+ZHMCTve62zidxT2wPtfQcSIXLe4dlJByfGei0n6DzERQ69GtLvrID2OzEK
WUW0SMR70cOK5/kJMvuG9s/dO2Rvm6WLPvS7an/kweNp/MvAv91r8fNhVQulweKh
82YgLnDay+8VzwS8iDJibnL229q7iMgDW8xMR2sGVoZ5qHTcLlTFETEXu0ShVLuy
KfOTMVRximsTRWQ5NFdeHhLOtTsz3fSzWmcy+1qhSTNFClNZaPQn5EU4xLLO0B9m
JPDIwhuTjsDuE6GqCzP6Yn0K+yoo77bYRQFgW/YK0fc4rOfT5vHsZoBS1+Y34heY
rbcZmSR5wmJM4XDNCKBHbsPeU5Zkuw8ZZfE0lAre1svo3qSyHxZVHMHyjSLN7lZt
zcVu7TUkwPyK95rUjtaFBj+mcTd/k00euKHJQeykm63mvJdv4EnPhcWBX2tMg89F
9tCJN+pGS/SBpu2z1f9xfnOnqqrwjzVBTTXUdzZMt5bLi1zjML7eaaSIUMFUsfZb
MdzjVsv2/G+xkaZomHk9Jc9sAuNPSLoJh5qRLl66v9jhZWgXFyZwr458OcsKMWms
bCrOfsl0CCnr8cVmjhZyFgsHCe6wLqW8eOS4DjsQArrWWzpb5NrSRr5jSK89GDq1
dEqjyDv2vP228U7JUfuT0J8dtQEz37ddFdYijwnm5qFEjzVpY47qjVNyNeuqlZ/j
1F9EgHmhVgisSRmjJhFhyynO67EjVnnwBzd9MSomZpJsMJm+G+rUCZohuyH156iO
qhPqFqWRcyxyuMRaruInOLJm9rSUCvYLKmw8fJC2HSvKJjz6KABcok10y3JfUT40
9Rk5SWpEXRCV3D40zN6HFqfADe0z2tbamdZHDNojKsqFcXEXaje3t5POPCvz24KC
K5R9j9BswMisEBtnrxK15x3KrP0F8pVvviuLWRn0YGNauK0tNPaEVrm1MQNOB9kB
KqjzHW52NS2yOkhKE5OjKqsX46ET2rIi7XEqL4DsL730wfI8Mn/h67BjfSWhxnEb
bCHHJ6N7aZ1Tg1aUASzJr+hieiIlktqBYIE+xXzTmGj9G92R0bEJBZYr1YZMscKW
NObtFkTgeyZ5B6cMKVUHMW3ubLJbdbOJ2yIYuyerGm7mEhjaY+Gru0fsKn+nAcIN
GyKYNTe0HDP+hjMup08dPDRIgwil8lKvESiMPTAwOm7SQetY0AWuDnap18818GLO
1IvwZiF/uHJVIxdgWP8DYQzbv9CGY3oLyQVmiGaeD5OlGOSv0kNOexblAWKTLePn
zSJ8EpeObCV9uks7GbAedmI/aiygBApyaB06UPi2+uG9iXnvdQH52mPV/k4NxY/B
7xBCxeVVUMxJ5rG8A2UBqNz+MUzoN2zqjAc1d9ag3+oGIyV7zpSYvAx2XYc/HnRS
00kWuRlZGSKs6m5zFfuItJjx7d5/uIpGgROmFjBdZh7SAX0zqwhx8TQjcZuYxGOY
12/0CcAbMAvahG62TNc9N9wkFkCUcm2KMH780SjCRDa8f8jNSFTLmhJru/LloXaJ
mCgHQALSI5C16OMfRxI/M8mtfeUYiBqTgjxbO8nkOZm4U658zuPnHPjd0ezzbi5k
FDKfe0aY+7f6sPb5WLy2SeMjWFOpi0Fpslf3CvTxsPMhvni3NDM7fw886oeveG+M
ZmRDIfkoRjGCLwiX96H/PGcOTlcZqB6Jj4tDYanmGCX7XYAi6+qeQ7f4RLCZRh9O
EvjZ74cuQ0tm0Dvf8iCjF9qHv9rc/mMfgU6ohIqQzAfrmHk5AUxQdz/scCm4VCGp
22/U7tr8JCol+PjasE3vhRo7GSBOZIvYZwHh1cRQO3mM9L2IROSdgxQovGXIiTmn
jADBdfLElFFljwCfml6QBmb+2+me1VV1PCOwoc2qmDGpbBR+uSlzD8lPml8chdTA
/vq3iJkXgqZGOZqPl6O7gcyMBaZJfVHb10q/bVrVuJP63f59CgtC9K5n5InLubNw
uPOMgR6TdKuUyT4D+nu0JAtEUle3LBmGSz+4n/ord/UyMRhf7PFdEC+MDnFDUTB0
BxBiy0vk11FIaXTbnToxn8roa2gV72pQU+rWGK391Z0gm75AfUeMr0rOhiYoG4fZ
WFxSxfKr9qw0okbWUMmoiXF3RCURsUVZqV0bYYofFtijJkJTelS0/dY0TL4LiSFb
iBzOwOiMqVMwYhOgcDBasySfOauv+7S/JSMP4PtJmRI6hDlXQOnq3YVAfUEXZ2Qo
E0Vbkk+XYHekp4Kh0bca8HrxUesA55VKSeywlXQfIqEgJsNA5vxNrO1ZK/mlxDaM
9cJqp4Z3jOv/Qs64p8uwHzgnGaYQiNFnabt+fjPu3S+GvoHeV5Gvu5PmOD6Z1eyT
P/845siy4B9vLntTyO6Tb3cljg555eVVgkUx3IVPxsTpu78+g5RCJ+qw8Znk0+PP
0LBDTcNL8ULhWX5s81cMCst96QhABm2oz+4Po6IVMOmFIK8Hs/ET7n9IFV8QpmP7
vDU7GEofJKinTDncsZ2wxV1IziFHwc4hNrrY9t5pjDV/f1bOR4xNBmzhnkPSspdN
ZM7owbAiteo/ta8Hnv42+b0Qp1wP7ucoPvsS0xNhuzXOaojJojp90pUdSq4ImrYB
DEAZ8YEyh6ZXdj9Caunks4MLpDWXMdLraXBpEcYPxic9ccsHz+icmt+Ud89+6dYU
r7KH6H+hCyt66OWr3MzXsptgU6kUrERkhNLMkLfQnwpy1VXB54xPX9WdULw1RjyO
FyvPhndj5mI8/1WVBjeFnoqfTJZBEoAkDX6aAmsd3eht74vZg/4JtSxN8QsY1Ics
McvT39vCME8TtoQH2bM9/slpHTGMERXM29M5r6AYpKHTOglItmjineiWrCFayeg5
2kVdskiaVSvTxZ6AahVvjYEP+QGo5qMQEhKD0TLySmHxpRMJfBv83Z1DOeoD5JWG
k6Re96qliq70DQE00ocIeqCwwQyyt6WFRgWLUit+bbyLWkF8oUUFhi8LWMA8nCrg
wzoYBHP2s+bjVFGX1A1hSz09ubrEd0tVrOlaFfJTE1MqF/itUWdFU6aeInu7Vz/S
XvsSAKcVR7E46+ZICvldj9AKbrN7NjqDfX4j8c9DgvuNMOVxrafqVAXeRq4jnpbf
vSmX4L4fFMvEUmd2M7UuApG4AEZIT6lS7Qg85Ps9PgJDYeK/35BEcY5ApuBsrBiO
bT+LYRqwaMaKcCjrmYsEMhZngKM52JpiHgh2wTGQJnOJGwq+TNlGi5ucDm+AgeLY
nYr57u6PvWWzp4bybYMIMCk9q9RatTNK1la4ifabSWzHjrCigxmsugs0FVCoICXK
dIt09V5LGPnoCIDHGBvXhIT8YOwqFlSkLUDhATIqzZ1V2u870Ajz58tD76lOWLzo
LIBrfmEy1Y+b6cBfnwb+rFAf9iXFy3JBXlDbeMOadaWmrTnQFo12+sBRfQSUkEpY
CDfh+ouY7K3EnO4CBfLHcTq0XZixbKeaQOW7VoZpkolilp0SwJH1fLPup4NHOn0p
QZHu8tm3mm7i+MWsEYmOeOJfDD8siPcKUYZWZLxxhaTqYOIrgaY+URml7mBXKYHz
EvFcqMFUjC/M5QTSmG9mxoX4d4MQ2oBwrvwIa/NnSwoqLEjrzeYuXjZPY05/x/2m
JgGBHcEXQLQhejg3359KDlzjPK6AKVM0CwRRTES/OmRP24/eCaAwlg5I/qIAziNM
g9LUD+gH+ZEsRrUWm7JggD/9rEw/UXOO6UcG2wGTTeZ/HsXxE8yOhuD5ffozdnXS
erQPbZWScdX35hbBQ5Da/7iAork87u1a22Lk89yaD+GEcmCo/RrtbMiA/2zxruKx
tJMZ1A+sfpH9iYM5/qQCkYvzY8rSn4mG1CMVXBBSV4ynP29Bh6l273XGu9kL2ym3
XJKsPWXT9bXmYZi42bS3UseAblSFiB7nIQuCsLyJhg+tPUik22I/IO8ehv7xYN0L
hGxdGum2I5MItcU6HiKjKerlVJBBakLrbuioM3mN0QFhMjJYByY8WOADzyEgYOuY
ytZpozjKYe0+ojvos7lIuB9BLKTxxjUszqtS/dPDggLPYyWcsLy4Auw/V6Kx87cG
nc8wp6RsT/j9dFcL0oFiTqo+a1cbj42JU/0cAO8p4vrQfyvskuUJp/nvO51BNytn
VZT75d/pwBA/lwglb1jGj2xJzpJuY9nIQzCEyiy4y0gJ1lVjEpjtR1UiJg7CclJi
v+P0AVjgVlCenCSLuaZBuHZanxOE9oECq8uWU+zDCIP4e3tdUERqfGwsfnNDGXGN
WMQrB3a6bcXBX2GJk8sXfKlMmlIxjp1VBiURyFUE5WBL0FQqTb6XTbFnLXk+4mM1
Y+q5KHuOsiUygtzS8b7tBs4xGaPE8odO9Z/IP/fmdJrsHSsQ++PhV5I/FTBi5fbI
ZQEHZnVivkYR0j0c9a0/s13svUJY5sgZNFx9IWkFA+nqbZenkSi7Mw1yNgW0hO5X
CaNfavWE9G3dCkqmYglgmftGUSzKHUZinZhn41VC8BLjMwPSHexLqoVLzmwOLEO8
pnoh2AGCtM45W8zlsZeR/n2PyOwNnnmIZrZhh06IF7mc148X+Q2/mQrPuKMKXHhL
T72rikI6uO6DohtZowQydy5eO6+8vJIsypFSPyKjdLE1AaBJ66Z2ZMwKgspkSFq8
Cb7npkuO46lBPu6idSGN2dm57bhcdxy2voQCCBZBNJMfFbdbd1UChm+OKDyPZKX+
jSFriWvrLoZlrcPFUSi9vE17Dr6exj9D9+fCz9FJJxCvnhned93a325oPsGVhLEF
tdp59hNu4Iz5zDRE/3Xh2/tbVEBW7IyDNuPdrgzrmUCxNMlho1MoXilRNYAyjnz0
sGOpv2JrobjOCsNk+uf50wcQRbEOTprtF1NAdW0QUsSEq/rY/IPk7Xa4Y8kMACkA
cd3zRJwL5BOzolC3a2nOBUD5Q83EugIkHb6Gf5QYO1+LVJKbuvi+vQhiglMdBISF
sF0HM8B2N2OwhCL3b8hcOZeViYXKFaQZjgpCIbMWAO3//xkshJfhdRWiHl1wtEDM
t3sC2OEPjuEAkmUOALoLAw9gbcZxLQ9izAMzJq4Ioqr4B19KfrlNvrhFBAg+hjt3
x81Gs7/7zHzuEx1uIVe/DWJnakc/0UCJ6CV4B0PAbGF//BpYJ7vJ7bNzWerE10DM
R21Mrow8MG+m+tTYqpo27dKFvymCiW+HOdrbbWpTbWpEN2qJ+Z5itCa12xx8UPOd
F7fwDXuyXQh9FWMaTjRoSPMXGGSvQZhv/IaMGOSBebap0vZ50mQYApHIRQ8r0GAd
OvVDPND4fKZyrQBl+FvmkpU6jMJONumLJTn6UHaoRgy0i3GWe8QIqAqKw5TB3mIS
Ji0Kk8c6LRSbVFF9d/WRD3J05MhgRCsVv2Rykvms2B6+PIHa6s6FqxT5/WaZoPLY
xJ3JxIrEpi0cd1jb+JmME+e5Ie3v1x/4T1+Hn1DIjV/IGxiUywyDP9tqNFpcFK5m
xipDBMJCV51FzCIJ7OlgbxroDDnhPqn7NMxYbyT+yXu8VNJIDo+iI5JfL3u6uqpL
TiJArPplzwPBfuerNZjQof4OeNYbI2yUI4yeIEMWTV/SBdGJFLWSJ+vll3vDjEjP
YIQ69nAjo7NGVxmwbnVgDjDiGH7K8tqH9o4AOharg1BGi2IoU3YsLAnvCJ62dEpX
K3ZkkgrUxhMZoM/uTw+bcj0tzpul4e7UAbdx4xXzcHdWXSwbc2wWd2LwYQJIq3JA
6zYwNpc5oLOpZsRbLPUsY0trQWW5vYaliGsW5MKa0r46QevrxyW5s3Psg+vK2ahV
l5TwdkeI1cXyOfokF0WK416+ip0QhCEBUewzV94yg5ltlAXYb4MUphvLbDMW+PDW
gEoY6LmAVGcylY6gD+axICiivknBYNMjw/RO3zsQG6HHMXSEUaz7hadXliUXpTLh
ovSLVXcNIsn2fUKpgbc/kTU4i551jZpVw1JyyEETmmtuu3KQSU8XwM+Vwjr7oVlv
gJs+dkgrOYl5m30jWjBaXyLxGM1S6K5VC6CR3PfAPEI99S8N9ryI7S5DWOFJbJLg
5HPogN9recym2ENlENx/YMOv4VZI9nieTA4KJ+FQI/JljEs8VlUl+Tziey86kdB1
4Lg785nGvPMKp/uJgzb2BR+qGBYfjiLn1lmGJTP/Tn0FfUVvCYveILuqxRBswaJa
hgpUDqehTOjB32K4SsuEcPkeE9ONYFM4AAsK1bW3TJpYQyQ+ioHuOTJoAvbgWQYH
tl2TQFrSouDDaCdASn+uQ+8xsb6j9WuSWScrjC8VnNOFZ2MF8K4Ym7S6Q4X28GKB
xlCoxBH4ss1hyB+AH3sYa99rqYUI2HThiBMFeJThJSv36uDohF5Mp1OdJoPe4yzY
yPJouYU+ah1NNKnnRP9gu+xab7hul5maL2JPTzmer7ZCVhZWq4Wh+2g1BAfPzK0+
zEhYfxhpopbwosKDiXDqAgojnSJqlNvMqGAY+OKRzgTdqST9bcql4bTOqYnvjlgb
HPiOVTjOn9dh2bbwVBi7iZo9LA5EEVjOrGwyRTjAUEmeB8utKasS0WVNGjP987uY
+z5DbUYiNCeSUo7D3L+3Qr5TQ/gmKvizWvIJiZtnnzGP6GE9vvQyFSP2w/UxIJjZ
XYqz+Yp2cbtYsKfAHc6QGIC10OYjWpVqmYb8GMUe7Mdzq/vE5imtiwFTWN4xRcbQ
HNt49BGn2d9dswbv37gMhj+citwzTSqjLSLef6BOThe9b9CeqSuhLwnFmqTsbqAd
jx5NiRtQwz3FXtK1AZvtA22Hh36MMr/LBJ6+l/e0+3QCKxE1lzq20Lg7tzxONiJ/
dZwhMFA2HIQVHqvwWIu31Ml3ontIzhtxfm6vePa8tgrcWANW3CWkKwn7PqTdzo38
gHBRRIoxMTw1JVNfb0dRv80mmgU0geJjIDcoCHRpEOYn5EKg7yUJDcsyyI+IlTI3
5HpBcHVIYTYQ626gOinl8OpFPI8Q68ZKrnlLYw1syQGFo3jtRa9RMJ0tM2nY3u2q
CcKjUcSmcwd5pULr4/8k1KXiZ+rMMqAPJMqnSSWzrZlosiPncbqLGRXMwb4hZcMc
olOOorTWmAfs5Hfvcz/idfJVOEj9lE2+nQCVxIJavCu8t4TMBUp7/c7r701SDpGW
sDXrJwIBh7HyE+QtsElfmtWih7rlcUFVnWLXXTItAaoXJAbnaMvcrZgqGo4MlQVv
30524uGt5uMaN6M04KtjesZ8wYULqTiSYPZfwtkqvMdemCMisEtzPsyBcVw9V+Qs
3Heo8+PIZASA7Y7osbK4q2m+L5waE/IMbKudALBJTuM62v/Tz5AtZdMLL6hqWuCU
4YkK+yy2dDSKSIQ7SHDE8iu3xn/dyLa24Ic8DB7vceRAIWyP0h8Tb+4+qZzJSmVS
ZsP7neeSA3oThPPw0KUP8T2x8xCEbIilitzyO7ypWEtspQhpr9/zCZ/pA4d8YfKq
ioADvuPyGEYFSivbTKCnD+SmRpIxz89FTU1o37npRM47r4xpQGn9/H2lYQAGUfSH
D7Epr/n2iXLI5qB7P3jPmCovq2MMwdTidue0D82nUy9FGmRd/3nC28qKgeAWtMH1
G8OVfLRDmWiKhw0VAkAbq3r+z1W65duCcrLDTIyFmGHmwWcPi1nRzg1UPmHpsZQW
0QQD+NN01/pExHnB0eIU8VUOOJXk7pydS6RTHCpvcU3iLE6wKJ2qXjeLOBqR1mib
WvHNcmrK3o+Mw8ZIZ7nb8A2ebquL9SKSx+JvNASOdUP4ddCyuY8wkOnU3fbVnF3s
KCUfB3FnqBNudqvg3YTQM0E4wjyIxYvVt8z1uKk1G8uIFZPrHo6kry4EOmiqBxtb
OVQRq1XbUCxJCZ8AXhUbFrCJRG2qFQhWvIGIrqu6YOdm4Q4btkRzuopH2qb0issw
PY5ZZ7A3WX8uUtMT5nbMuPFNLUySQtznH6u3ajXHFBMci0K4g2vQEK1aULNYpwQx
M9eBs5p1woxAuitGAbfQ3DLdvc99Z2svlZe2npL7xzpbdlQizpO1uqEvCto3/ifb
fWg+6vZfkxAiT4FgQPyU348F1lO9L7v7nKuA3pzgWZueAQgB0z3JXMsAw+3f4my5
qk2P+vPVLlayqOuVQB/Q4B+PcCeFj6sLzz8ydkQeOHxgfr09X2bqtKfBLe3HyDMm
/sguxD7jAOvNOPhDir42WnV9F7aPxLDCpGexs27VNUkR+TxLVay2O6CJq26jppLo
VaRJAY06mjeaPLkVshC/PX0sAnOuPJrW1Nwb53ruOrbZME5uR4lHDSr5fp2OuvGu
/RiIrz+oRmPBRmDA/OC3+9WPLMF1UA6Ih2FIQI/E36fhAPDxei+4KkeG+1FcjASq
j6bgzx/5WZ9SEe4LSHrXTwUwgP5tSiifNWZtuphmfd86xYylzgWyhU4OnAcgqRPF
bSA6Z98S59GjIAFy4QqIxTZkWKV2Q8yceRPLyNdRPwzWhj4I1rMvWMFNPY9yiM25
O3eJ4ZeqqOvmkG0H/0IHrM1KEpZuVTR2qnZ3/rNdv0jbhXNU0BefQ/3WG8dXP2lA
X1hIKUh2yo/PC1epwfccbqc2yuYcHUwrs9zEa1r+eF5y9gYXGWC42Fe+KNUtTIy2
FohzeFmCagf6/6uCfS/Qa/06ojl3y33uWcyWca+rIph8mPyaOc+u6qdvJgQNJb3B
SFd6KXo0HsmqwjGvA2VDvirYq/ar7E9llJGW8B3iVcJddf+4Z+KRfH2VYVxM3uK9
kycx2JE0vAsNCsGIT5rS4JnaTYfcINWeI/jhIZkygbbm9Jjd1CZWdarxxGv0Xgi2
TQHPLLXq+7Ubs9FfqkVOT1eqjmwDknMu0KlhFSgGM/axU4OT9eqKCRZuSLD/rZOm
h9iE/5XvpG+sAbOl+e+v7wx+tZFHU2d/18EPpyk9Z//JghRiER2IpFr6xbP9faVp
7BbsS4P5v2/uG7SWqyTQajLInU291rWtr2zelGNKE9kk3EnGlJ5X9QeLDHeZ32hB
mo62KyFKr8MN2GuEOTEBY2bcs7AiB+rWG3g0VhOnWAN8iA2mgnH9t1Tfrl9iH5xl
ZHBozCwKvh8GWEYZli9EhV/2SwEtYRVB5QsY6Tc8Lmi/IXW/v090+bcBA1HSWww9
JR9S6QirlapiAoaWC7EgqpkKZQN5C8Ja5iTxzTsdkX+MenE6tQYd9GfQC3WCE1L5
rrJYrYMc/if4HKcI0kIK40obCcLu1CGQV8nQCH55DkStH4ygS8vxKRatKrOw3Vux
YItmiTGrDQ0FIxtlT9kzf38qOZpoIMCAPbLnpYa9gbOE9FCKuWqA/GFtp7KyRTVq
8GRqf6bFmUDGKyxR2FIMq02zEaUfMD0vNYO5jurYBqZOuRdiz1UykgQkMSaJ4+HW
v2he9WsrDvwUspESNxlI+OoJVasTjXYZ5gE5t4pLzhPQ4jtkzTcy/vZPs26u/FRW
5lz+DFTD+qumbsAXvYDfFEtL08T4Gasqd88HrQtcnOQx3uM1z6yo/Y1007eHXft+
9B1mxPXTW3Mg8u2T7/DVf6jV1M0oxMiREt2L3V9WiecyQzYgqgSNoEn9iKJqwVZz
qlzEwG2gMaSzGOPrsr1Ml7qfWJEgSAGAHB4n4J6Cf85SLwxzEmAT+S0AGLwYVpKQ
IF4T4aT/EXLcyI6ysTzlC0bNPO7KkydIsACisejOnPKv7A1oQS5WWKCZ8/FDOJf3
SqubX4sBR6rjcTwdkFEgTLyVB86JxO6EOwyrav+JTIEfsx5djRmWuFIwxXIcj0R3
cfq4xzTsdsdWMIr00UOraVpAkbqXkXKE7IGT7BD0n5DkMsDtlsJlKf30PNFvlTt2
pLy/UIAJeY+r5q4yKir1QoYSayTws799ZtZC9+oGvdO0W8fEozDpU0uN8460FDwF
bTfmKY8I/Y2ItUgRINfTTcP5K5fHREJ9M7tLi3JWhhzowS2fdwZVIfcZ6Y5axIas
g2Oy9YUNUXbJXpdA+KXMdCYibjsZH8ElhBk9rRKytUHUtfdEKuO1ru6bc0w//sh5
kiEWFLC5xL3U5FbX6EKAUPqQUK1fuPEbpNgGt2DU6YwBxQ7lpQCJ0sHHlej0qH2T
GgNhTklz5/TVP0ZJTofTCaaGqYXI/MR+Tg1lj3th8Sbodzeeg8zJUTSrE0yGG7mK
/Dnv/5F98w5P/ZjBpUKur0HYIS9K/dkuQbba0Yy0Op7qkdcQVLpQ8d6Y7WbzKSFH
fASvpbKRgr6YXgZd4XQBKQlqf79iMaVDYAK3wgnuIFE8pSL8NQXbQwZ5pj3N+hjZ
nQTPFWnefut9PQ/chFvFh2nQcdZR95oj8oPVukqunREBGPAtNsVZ39CUL08tqyNE
AJTraPyqr8ppcIynlTNFHLyMDxn+Ut3rmuApVd9jyuwZAHaumihh92PiQFEPREDF
rkDx+jmP4CDJBJ5ZXTx3rjpMILLw//yp1AfdijXXDc7O6VqnXSvHLmIbajq/oZbj
yrsHr5ESE61BQozTc/5hZ88LrJw3N4OK71B24N9vfFq/E8uLW5RcKVEIwq8iesCU
Z0rBAoT55cJAccvdlb6s835NTPUT+ClHms9BR1GWLdtGOKhkTbPdqYoEHKKVoEXC
MwLx+Wac1ghqqegX+RnZUmdvhrvi4vf6M9BMRZ8PykwbenNH/APywYhD38G0V18I
AO2qQadQHk4L7IzcVAnvNy5FqZa7zSWzGKLgcEFKRquTmAx1H41G6iG6GL4se6Sp
UlcMaOca62VrCiiu9MeZCee2MmAcpLqzLySQdOdr2pt63YliBVg8kzkLCVE6mE8I
I42q0f8sXPsDIgCxyJgwag1fo1B2oU3BlcYenv08QgscFGuo6zBbEu8bTWiSsblZ
jvIPdAmU2OEtNRQmy2olbcBSEKEDCDsaZGJEF9T6YyiiatqVNTQQoMJJGvTpxuHz
AOmte7G3nLJPyH175WweMBsWcIiKqRYAE1zfvGOCsfFpL9cnHV9uR4BOyeHJjxGG
DCMlAuSdJ6Xpjy2HsEX5VMc6N8//LEVnWb1Jdevw81MO9afr620lKw5Baej8iDcw
iXksDx2w2AX6B8neKaldgASmC8GB1z5Monqa2FeBoA2IFeFcLHzZ40IstsP4oBK2
35je3iWIOMomZadTdb7c+c5hhDKbpFz74bIayKZN9k27kOqYuIaYpm5YY+EzkTXl
AUS15UGaOQbMGh7AZcrKg/lnbruFY4yzghkZVESpBUbVoW8f2lgXlYSTQXidSxqx
Frnt49a7lhtWWtYFUIeA0f9MBPxZG4lztGrpDwsfHB+F423fv+41G32kCSvAWoXh
12ruEgPXxQsi4RBQZ6GAprjofh9PqV+DXYYio4OCd+8g702scSXMnMl+oOL/hK6t
3PD8Vy4s1y7bodNtTBXXC8tmSBdjL+cZs7XiUJuhRDm/fa4FARqCuT0sBmd0/e9D
aDgVBPKHGd4uuNlSc9T4RbHQn5NNwQu30miI6PlgOMEhVOqsRYlBrUeE2V9qEWlI
yzwruWXEX+S5QvirTdGEd+b3lvLQpIxLk8xCHsHkMy+dZALfdRdE5BhwlSTJ5Shs
FS4EC5DvYmUKU+gUNMPB+0DDbGiw+8WHe8EXklgSpmGrSmRN8P7zxD6lD9ztPtk8
Kwtx0Y8/E/1JTLn575WR/XBbPyZQN4BjttqK+WvAXXnXBvvzuEmMYVBswEIspA0q
Rxk/TMzzlpU03UlxlJddiZRPF9SWvdWdx9Y9syPaXhrDeTyIOg/pd6R4+s+s+NfF
+BgyISbdjoQlvvgKnDpw0Ft7qH5VaFmj9ewS6//7iOZ3SvTcN2ETt5W4zoLF+mcG
Bx9MH8ctjQVu4oUl+EXk6OH0goJB3sggvt9jPAiCtn6SIiQOgl0sJEYpiG+/HIMH
A+OOevsDlTB39qNeRX30S30TJ5wsGCUdLT/8oJjvUBc55j8zDHxVx3IpC/OO1IxQ
z47SfG81aOVs12UA+uxi9lPPbCOXxYsUcGSn6Uonj0Tezpsovz1/hHwRlHVuLcwj
VnE38YhuPkD1bA2L7rutPiPi86lSp51bNmYX1eAUegK4BOhAKDkoXGm/6UsY+zLb
McY+lfwId4rsClewPE9lLHCTUAD7XwQf/UFO1fzqFjR0mKgdkiBIAVc1PsKn1KvD
PULt+48jQBQu5JLsM2X+7oQG69Q+dPSuE0Ifj0VmumcApNw+H19OJRUhdYZyrUSm
4yWZkx7h3K2nz1JAtc854FIgDVwYmsvUjPxiwRrH8zgqXz9nAKwiXCB0CUU/6UnT
yspTJHYR20LiobyxYeaVUH7I4xr84rY2cF/SWzrSd5ReCiPTPk9LiN2t96C7eJS5
bk+cW4uKffC2Te7Ms4RbWwVx9p8EL49m8pSpzaNe6OE4ziuYrnRiPfwdYC40v9do
JHSz8tFJL/5eAbMGsasJ9pHBHbLgEAouFvfN1A3cmDZ1ChB0+wIvohLndDBfEq/3
+rryuGMmCGBzZps2KVayK+MnRZzjeWiDer+dKIB31FSoh2dEIceu3+LY2R69xxx2
KhqijbO6qBJij52LVs3Etw5a2IbbZUGgw4AZCkkta3s0PnjmkHWouj6+0anJbhWH
U8SvOPUR84wAJB3wRE8eIvHGMUWnXxP/3ahGjH4R32Gc3/a0Are31fpHU3E0ur0W
z/TDISIKL2sf7Y+LoCSWML2zME2JBlBHqr4U5LKhf7Y2rzpLzFca4DceKwnnm8Mk
pimlYJncFzzaozF168Fyyb7DjyiSILttE0W6q7SXaLnEcyTgi/HN0wITGkanua94
fnhopHa6eqY++3VRAJ0kuVhiYhGuO4GGpwG7SuUDT8JkIQp40qiY3evFWzoU4lTG
CLh3nJvV5RDay0EFokVTx1CbHsMtu3tZS5A0WO77ahKMuHVjpDrwaIYyS039v+yh
UqiuKS1U7zQOyL+PTsRyNbCvBwjmb83lPizk5x/vPucxXQZtc3gEoUtuiz7l8oX2
hq0CRzkTtshWsdaRP3gaE32+Sn3M3Umm54o//zk8jv/iI4Q59CAAkaJwbBXt6QMq
rW4Hp2lBaI8ctb5XOx11DN/Quu7B/PJKBOR+1l8ia+8ZMvfZWs5tz6+KQMDY1Dxn
SzJOezEOhrtjv7hN/OMa3A/gEob5X0PkNFTBvPJAbn/DFa3+D+70snqyZ/wiYamZ
o7p1COvBRtwWqWAdIagYI9/B/YSSvSOaIE4XdPPoBrVnKA4YeSIhDvEKFn1jVxgf
sZ2xgTFz5WdmesPwBo8CTaTA9UGymm11NoCs4GzDGqKzYtSXKSivJss8czjo1hgy
EWRAgsjuQ6uFIdkhLw6T7dLoZvv3gcf4lwx42Ppyy1Vjjm1oPQvFqMJH34olM30K
ex2ckR8jHIaX6fgbkhAUd4JjxfTWxnzNW9fXuBWti8FQDGO7kO8XH/u7ZxV4WwI2
hylIqA1pTws5+ptPf39fB82bSu2Jz35zD1KxDpbdpzKYNEXwrdwfBYLh5dPqZHRY
IH4BkNC9Lj4O2tf7CMOxSB9/jrecU+ewI8VVPHCAuKq9v9KodLj9zGfPLO1AqeYp
Q+1/BfempyVgVaNPSjrk0N+xGQQ8xjVcO+FNJyL+WJEEv5EkhoCFUibZnS/Xi1z6
gp5UjvDp7CRDgIB4u/VGMKoVt+DeCi6EaNNU0ra0aAGyXgDLCQmMMdzrIcsP6L/J
qs7xpe/n75JIz8W1kw9flmaFC51yB1MbenxOahIrEbGl4lgnwC+WIVaQnj7K7xQK
IFsiHvlYzEVFqdM7rhoW5Q3fucV97ow6XsO6gs8P/2j1heWnVu3x1iJcXoK+ZTVo
NSQBdSMGXqWGMeAyOtHQ+75NHKWCZtkuQoKFvq31nKAoAUVM1P6oiQ8/+caRx7il
GfSZmY+Y3BUk+C+QGnJFAGNdcULnkhCauh1BwAQvalHlyRWnIPctGHs/0ifsQqPM
kRi657+kY5BMh87YMStn6hjC9rjw5CSJsrU64afpRWZ32i4w+h0CnwTzDXblZ/vm
QTtzAr8Ipz1nUJwWB8YwD3oJkKlQ1y/BX+7/PCTrGTThJ/4mJIURZPwsnW9Z8ogc
c1LZpiNUkNAOtFd7ebjSmysvpcJdDQOiXn7mOGu8OexFASw6dMqMEgrxNXxgxPPy
SnhKrgOSWMemuv38/lgozu6/1gmnaxewjOLAXHf1DbwDNlX5LEzuKfC5GhFzwNi6
vDTFdaelWBTlojU3rK26S9jsFq4C9Kywc8F3T64s4hfcWssxsVqwN907FDBqsnV1
kB+rKBgGf0JdRbOVuH2mIZwup3lSmJJyj/ltCGRFb4jTTUi2FMCjZIFIkkC8wPAu
mEe1IqI6Vb5eIgtvh5WcNgWFtwByGE2Uik4GKe103bu/uWU1zpmqmuPcgr3V1zi7
sdaJP75fBQ1gVXL/oIu9iNREFGbEWjklaPwZI4uz6WNeb+5Y8MemINxxFsjKGyVw
WFkaHuVdAqfGFRa13YZ3SDcl+hPLdf5mpZYzgM8bnX+k2sslrCCYVzUeacAgY6hx
acCP5iwFEIcuWSJqX5hpwfPh+Z0Vgpw7KKRTaMg1Or2HQgbTGB1yFScxGJnp0GG9
ysQKoBAmtOO48w6g0/EjDrMdBlkF7T5EJUxj30aKhyU6s5LOBaR14ABytKC6JPtO
8exAm2/jjwB32riBm+lPOALAJGgvprgj/7bNaL0mM2i85ACQ0lKPA0dkmqVzlyM8
cP1ZRoKNgkj/uBH9i+IHD2sN5UDQEJTC63i3P/m1HOG3XcNIKfpHoxP8fVL83o/K
Xach/vXd0IVHUb/TByt/ioSwEf9wvUjXJH/yJco1zY/Gh6zdU46tRQIRCYCOr93y
0AnCyz4QGmdNUhaPhAMwsYkivPi9EBH7tFxBVmBN3y3jp6Vh/SX6BTkxliyjMzYX
LHR2V3Gm0LZ/ELkMU7FLIR8o6Ssq1yVSK7HtJnH1MjNT0YApux0ah8I598QBrHIz
TH8nDKftZeFu3q+z4a16P/WzGygHzCS10EXDqas6rTVtcQuSe5JRlbnc00aVTcI7
iLSaKP1qPVYtYVUg6PJLTaTDkcstICHcD6mbeLE9txWodqz+zrrOHIA7F0K4Wa1L
XkfsbKpmxnqQRbpYcjpz40rHpSnK+B6/dvnuOV9wtIOL3o9ZHTW5GObkRHOljefQ
8fPkN4Qq42+0pWn678eZ+6X/BXRs87VFy8lGmJRdX+7nbL8Tr1itQfFMD7PhtJ2o
fppepRycCLYtkOi6gpssWKgWPsc6hiO+fY+wUAM4hGQF8xtfibsa2OsCN7u1oFOr
rS8vtU6lGPExyhR5StCoxU/x4hkjE0m5I4PpSdv8Yi+mwR8Qf6D5zCso5c4lOtGP
3nrBsFD4NXemHixAzNy68zFJtOkQcfof8miV7S6cpbiVNd6U770/uUI1567Gd/ZX
3XxSdl2dw+8c4aL5sgG/gguaQZPc17erYPCU5g4ZdTcS8bYz5kxjWClySCuBf6xq
vT5DGhi7ON0UjyEnpD4NuUzCNq6ma0UMl6eayNIKmuvcxbIvyriMLJus+TAmgO0f
7X1o0i/bNVz3x1lfPLP6TE/1gpbiXWuZZYlNpqw6hu1Ed/7+o+evJM+BjUKMPTUt
6D1u+jUuoyxv24TciSfT03NKFRfSp06xwYT6lNaFBIa6S2BVncarjVI+KoFelnyw
lsGM9nazwlnHme8/kQcLyhrg/UyqHTrDiCO+lu6VlwvYH0fQljDS0rkmZdCCb+9p
iYaAB9+SnFlT/cfKgXS3822hvlPO5+3chPiJ9yL0Q5aIiks1RrNujbG+XgScD33C
vQIxmEtuHH4UWzlhpPvHeWfEY6v358E79Ed7ADEfliG5VgTDyR4vINlEU16vxjEZ
bZUomFkbXwuWvlCXJVT53RJsU/WBWU57fEjlQbKa89XMhAompFgj81qbYy13wac9
DmfnHRP8L1rJCMuDhuz08ZQ8jyv15hW55ZNXR7ye6ET1BwYqd700/Yp+UUc3/uxZ
HfJjphdSwQr9Od0UgZRyLqefgBBkTQVbF1kFc4MQHXQMRKwt9hnPwxf9IgYu+H8j
XBdMPi+yUxlXQ9qgwOueVw1f2R3fbKSmGfHwPujtFWhQ8DWK6WNL5RrkPUrSnOi9
krwakCRa3ZIBNLYHtvOY7oJarvgEp/oBcDmkFuONvlwmvvNG6+6HFbodQY2pyPON
tf0WRrnhjP5YvOKzci37l1yGb+CXF5x7XteMs2T9oJj1WqJ1/Q/BDo+Pk0ealJyE
8EcMzjH3g37hGkULriMxHedrXUzOsuYSYttzyfitnsJj1YvwYa7O7du/Z5UOTZ+j
N3jWxeUMrKmpJHSAYP+j+Hg05WW0p/XUDOLIxef2ubWnEn6xQRP1IvFShA+uichl
+thPoMkeQ59ZSv2jNzUfJBlEADld0SGYb1qReozbIqbn/l0ON7qagsS1HbgbAm33
zGbinbyU2vBmoQikLmOoN4KnyhtIdbJMFYChf9gmn4ZOvqvbleFzHyWfgZhKy3DD
yOoA3AaN5rbXxZSUOL71eqJQAsTgz2iqWVbmjaZqZ3LLXG+oLtHCBwaDC5D3elz8
Iy6W6kv/qYBMyCn1n2YgDn6miua7kp41DKNpcnA576AEZQmmz3YzopA55pPdNNB9
TcjgNPPDQ64yjKlkvOKo0md3w4fTh5hMJIe+TmhCnRrDh1rmj93BhbmGBgH8iQ1W
6oV2dzsklydunIKE8EzEdxb36wnOeV/EoMYZInsQRusrlzhZzoymyiZRuENPutZR
2PCGwZOhNeIw6s/HwAAUk8OEztshl4Nq7CclrlN5F/CKqbM8oqECL8NImL263Yqc
HBBC2oPqs/o8eDCWn4zYxsMHV124Ecykn9h3kg0JPHjcyYMSU4uKfcXxaX3zRS2L
PQiTSxYTzcKZQ2bAL0XN2WNwsfIFPPB+TWjj09s8sFkyrfvmGcnp+xc4teJX2+Cq
BCEsCc/o1/nNq9fpPbYM1M+nNCfIVQO7uUSVUtRNSd0FkVRUmoTx5LZmjZq+PY8S
E4MoYhlOX0u+6kpgihkd/A1s0ZrtHdgxUvInewOd7R19WRdQj2vdtZmIl88mUKzh
ypl41wEUWcxqCAs+01gkPGX0CUnkq3fKKpUTrUPNnJBy58P0bn/IZvwT3E3g1Zxa
AZk3smWKa4uHcAPOuf9/sDWrFbVFZJN35hQnO1vLbznv8Bu4TimsSChJEOgAMvaj
qtISL86xs246Peh+qq753nzK7jut5Ui3dSIJ7UgNoPWmpsdrBcegEJO1fWrMnISO
o58LX1c3VojY1kWYIAMLajlj1Re7fmgXpmVfI9BDWUN4QuP37STFjucFIJRMx9oy
fBMueh24tOr0SlQuNnW9AQIn9FAy0zfp24OCZIVpqH9HtBdESctG1n8/bE0nuLJU
Vk+4kpxAPQkzS49sg+TvRg362GevG0u128OITg+ZPoUJMrY3QJuE2h+ivXLanTtT
ytAuz4WNo8z6z7snNC9v+GpTKyY0XohbMfj9zxWOlwmLJ7GqZUASa9asj9Q19NyR
Nu0J3ajYdXi8SgmFqpol7do61usv3GglAjIGXHWcgfXLmAj/UrtmImEop1mZmkKv
WydhOs1iwZFZVj+evOULVLqzJkr+ivl5OjJzLrmghKNKqdcxsKhtD2eSML/jS2oJ
GVdqqPc2+PmJVFNmvkvZAHdNCwzdQKMI7LtruQRjN2DyM3ie7cvNAQO9MfUvvJAr
BtJuv00JkjbsKCnXMYK1w2gJydkIezhOw7o6Tn+i2iU7+0/zij/M+TGeUMua9W6W
WBUD7t2EceVVRzjP6h4ecqoBJUvRYE3gNP3XOEPJbXihefVwih4ZzzfuxYe4WWS1
WC8PClcQC9+RfQgki8r82PpIau/wWVb7jxxM7RvARN+IKBWvxQMZAqxfaiDFstej
0PTlRY7AzvhR/KDGuDE6pjr0jApJjZT66GRXtpp8dUUU0K8bEYhRksObHeo/rUoV
fCfBZKcnGnAr5GcJDWRhvD66qkf+RWHmMWG4QCb+HphNCQoxoBTl/BVBEtQEpF0H
FbHrodSVqn3utMPy8CMjVa39xuOMa00lVs/4OCsj+OUI0w27nG8PyEM873nyiQLV
7DbgbybwLExAkRapnrmj3dA4UylWLM8Dt2pU4EysY5BUO7flUYTLc8skmqISQZNH
zN26c8l3P9WpUL6NGFfYQj+r5uW+//jkWSmDLopYu9d2jscxkZ1NndIENFXDE15a
+BiJnAILYsgxq1IcqhV7O0Na2nAXaQmAbxRMWdLAm4S5P++HXKdBaMIoNiQesFcf
tmvTKqRHuIbFgninjee72+qjOrqXYHDzD/OwHXl85a5g74VKFOYMmq5fR97YAHp8
IFUbsHSVuxksjcF+wtPk0SluC3o80DwPcEGEpheYPRWipL/00i4ZLooBYCDC0Rs6
Z/MRU0C+H3hQe44xbjqf6FmXal676/x4lb9902VEqibwSb9Nr3lFIrOS0PMZloI6
4ED8AXhOl7HSBPX6wTo340wDT5aBgItv4jB7uVpMfhSQeUHt9Uq4nRuEMs59LKj1
aLbejVUs0GhwxxYTpQWP3r1XRmQBT0w/Ttjk11L6ED5CZ5aeIeEdhPALFkayQN+9
/W88FjABlvhnccPLbbPp/hfzO5bqPR/SB6mMPXmk9lm97HpICEB67LN6PTBoncaL
88SOOtue9JPXfzlaJibBiRcGFnCp6hVBWZSLRnMG/CiEeioXirQsbuYIl88GRWwB
O0zlmBRohmwr48m6+qaVOZKIGsEqcmD5+h8aNZdonGpMV4yqI4JnPXfnr8VrklA1
5m43ZQznGuSBQLJQeuLhhUUPS60/NXs2VuOUrB049wmtdsQoz7Gu9m6Y60cA4rK3
jVCMMkggbhyVhS5tJw/H8yFOCJoSwtCcLcsQBeNh3QerXsoiZTyMa71KgGPOmtHP
M0zvoIXGv/yjRpy0cKEC7hC0JlrfnHKYFOQL0YtPUuYsDuhkW940KtDdmtGtdQO+
RTndavsvOpZO49gwaIvz+r4CsuDny0f6h1tUE7x4GNSWafgD5/Q5vX5pjir6XXDG
b7uogpr5yjXoPicfCkv2zwBDHUrzk7Dt+PCU0ev+IXwdjyqtJWoOCi23r0eTJBLI
GsTh45PD+HHUT4sak7rsDD5X7Lt5eriz6TFJ1Ch/jsKi5IpT82rddjZKBKOLCyNp
Z52e+QMTFeIZOtVq3ZP2UUu2e70//gSCNtCFgv8L5lmyljtYZRFLK8xOrtP1gYsa
Ti6PXrlU57Mx17SNQMtJCH3uffOLZi/IweN4ymU+czxedoQY5pLDjBnv/Zhmd2tL
FElBuXxc6snM71x3A0+XF59j2kDo3IdZSrm4TDUnBfASe7M4P4zu9S+fxbMniUGh
w0qn977vIigh7CRYA1yElszz09lSKrLoyPHLl1vQ2xYj7tPGUJmn9HH5LY51cElR
/uwxytBes9PoHBNCKn2lKAB7I61LHUbjuJROrmRUCLBLd04F3dxX6EkaXPCvgJHE
BQd8YYU571LI0h9WZfZlVk8fb4zzCaEgNNfpskgyUzAUq7+3ucYhBjHW6f72iAYr
futWyx7jkTgiY7u98wiS2y4BH0RV0qLGb7cWUNd+NPQl2/buii/nJ/hQJOnc98Fr
7EWRT2dWgmnHX4Cp5eWs1wPMUAL8AiVjiaAz3hLLOWSx0B93NCBmVc43jlWw1i1o
oHpqP5yQLCPLcFHhHWOADuNRzBopHLrKJY/tvkNr1htsPMpLP+AHKAfUzXovH0LZ
K8NDFTbkQuMAMeBfEdxTLbqriYnfEUo106eMLUbm/CBowhAU1BHR25jAPj94X+SA
R8FJeR+9ipxQAEuzQM3czynpAaSGQkzcyNobfSufRbq1qiyiDAtwmkKOH2YEO1JT
rdxXHSMT9S1VeXHW0ROMfQtUCci6SrmUJEHSJSXtPuGTrTO2i5D+CWOlPwkcX6ze
Beq1h8rY6kenN/Lav2w6GBUkxbevvORYtkTvcosbFVU0Rl5Wba/6yD0q1clfwV84
gDJpK6gxe28QNGIPyT03s+VxnzRBbRVMm9OlW4A94ZWDnsalKp2MuoLR9hP1qIDj
mVRbgrqtiuWkm/vEfVB1Php08psOpzATT1qR7EFz134pLhIBCOy/2nxGrvnr6y4d
N9IxLkkSazhE/+WXah/Ys30hOtlSVRst6osEhQYoTvoLhbVcFLSB+pnErGcV6iSw
yw8ejPZc41kMDn9yxf1CTgcIwGF4WtuWURe6tdggLUfkbM2wMC4JTycpmAEeUNvD
MLKTla/7Z2lqyicp8kb0FUts3r/Z3r20TSb3f4XfLnkG/4TtcLGLiUSWDKKUEl+S
gSQH5K26xBw9Lk6bIPxar+WTpKSzC8ykNBowe1t5o4OHaYjXijJLdZYHKQBQYfUr
Au7E+rjS7ujj7Za7lGIVXZeah8JSx372ReFOKM0cmNnw4Uxd7Bfc2TRyt9+HYH/A
j8HwbF56DhpVgjNlc9bxDwr2vLv2SaVW+m07qDQhDYtSTGr+JRxo9ULcLn39aoON
XbhRmBnUNSRGpxK7X3CkCOreTRCUi2slSBUmdN8waqA3FcNJAhnJ4kndHTvkxZkj
MKR6llCQYHYh3icvWeVmHGYqgrTIYUyByRLlYlIywSUfH2qyworUX6mpyWFn84Vq
PeOuZIoR8JJNOuusAld8OQJawsa0kX10htpSFT/7nh4px7uOHRcEB6fa7+cYqlET
uoaCLn/C4kX9yobz7VkhAKmBgTIRsUp5TSdKdsWkP5lYELH9t4ehGqytbvjKusXz
CzvciyDB2ot9W5goYuT2lgr9SnbEhIDjPYB3iPg7ZAH8n2raqAXKaJ45LXwlM4cd
TIRNT0ZNWT2rHNX9I7U/14ykrvc7hIGTFNqnmidVVm7auOnFkoJFEceE8wr3swLY
SA6B8990/VQVHJCzxXGm1Y5SbQl8LWLCKlq97pnrnPOrStlAFmuyuSqWq0o/ohDE
WzFOLdixTqMjtbJAcwfOflVUUvqjd0N/D6j26C18oG5pCAeTCB95J2Dqp00/Svt+
Prmr92bbSpE+JyVBi2AeT3eXcyLcUA9BwdZi33WZI1loYkP7By4DY7mbz50d5/qS
MCtoqZ/LN1G0FYB9qk/bJuA7jt5u/Pm4ZNCRxzxAZERDEHXIgO1A0jmdd0ahh1YI
GNpPIzTGJPFTGN09U4CMKKBF+D84zrv0yUh3H2yvyzpl7qIPHsSuaTKa5Mxwi8Yb
Vqo9vEPgKTLVuo6d2WU1X4/Gz22NQ1E/h5GAqwjnum1p5np9Lm5dur7a5TLHz2Yv
x5RAbI6vAd4gxOYc/qM2Szm9zC+YzpemduAbegzzUSHqK6od7OWR68sqqYa4bW1C
JF+98VZJ1mCQex+cc53VYU8fooAv/0V8bcKej0rEvdJneMTvDDw1VHaDEcLI90KK
7osjCvDCwZdmvJlzFTm7sxYv+uzmgEk7sFY6Fs7JRSiDg5J75xC3pdHOD9KVxqA+
4iRrbftLc0yCb0/mnwQD+uPCTUDjzTxwsp7CsrtVsZGxXMbeRdOPXRMash0k75Q0
yECLqlQXiZl0NT5m0uYlRUXVnXxH8JHPkKscwPgkNAV/giIRCMrUvEvHgu5OzUfY
ZSf485qa73j+fE/VWfJogBO04YUDZD704ZT5367rXEUyv5C/ZtsIVE5xx+moxSYp
Mw4AjDCQUezepzY/rKVhE4Bt8Wz9cSHsCmiJtbEu0KqLXgm48xEmAU4P4aypyDjw
5v3bxlVdKdX6+sMXs8KB8fwHgGw/UgT7Bk9KrcgWx9KAczXDP6DtynPN0n9+EdiN
5GuMc2Yt66ALp3Z4shTVluo6A81zYqQ71j/j93kvMGDbfx0COtGq+fU3g/qQFDsU
yY1gwoL0Hi0SYU9au5czLFUWD+/BjOdW7oTeixJTYK0dlIMWes2bHfRcw0mv6KS1
PgRSjsvI3KWLPyZupFFoeI0Kg/wnlH4zJZbullHPWR5lGeg7EnqYTI4xCRcngE3Q
1ksgNgjKXoxqbpVrtxRkb7l3INuXulI4XQ+dz5z9yb9aE+g+W8xomIqGkPQmT+Z5
0vlaeZtAWyfObQb3Ol05CIlqGps4AFQWoeUb1KXDkvsI6TnR4jeRFKD7R1iAHG10
H45gvwsX8O28ehaNPjydEFqkyB8oZFOcOuDVtLLI7Bvank4S1Iud7MpbiBa5Urhp
KIIKyWTCYaA9tz88Up+r8j6Flmxz6E1zjLyECba/AojzuW7po3LgEDn7Y95F9eyq
y5sAEt0u5kA9sAl9vahvMNrd2djdf/13Wg1hU1nWki77WJjdc/zAuRNqteJvY/jI
8y459wyBNNtX/QTdXw6mOSMlhDuoUXz6kTRxyMqExhB/LvGu8OgYj76YOhBdiiiN
o2CMiV30hlVE/BSTwiuo0BQl39OPrXpayDPiHP2BXr/IeVzM6CD/iTEXkz6pns5d
z7xR9EB7eep7KDvGal5pNYTWjPeSR36AINgUwG8+9vVOcfmE7h6/Ra5g/jypGhe+
Iz37evVRy35g/WPUSl/BdEIJh29oZ6thAhRYSq7RYZzr0bBqx/BcnFx7JzlwwL/e
p9wx7wf+lBtRaebkWThK34MKjoRvufego5FTpoVxfSNOqaDKofmUhbMHPR/cd2g+
z6axkHXlD6Ba6rsmCxkx+cWSMSWMx9EbxDVs0vEiY/OryK6AaDg5YtbpK6VA4vFL
uBh1JJk/a6hpPLsDqpJLQvNrzyPuQCBbkVqoGIC80A3vV7WxR+XcnVzIW4nVAA1u
le0Is98WY/VybkGP1/qLVVzrhMxv/GbByY/3XhoThcI5vKZ68m/zGXdrIhARtgsJ
uQ+VFoz+jdEsAM57Kspy3GmhU0iQN/ExcYQjvf97gpLvtSkWO1/HXNAOutK+KoCJ
hBDPG6ve52MW1MrhL7x7B2iWuVA3WmYDcsakXyEeyVSdXU60oO0qtt23C3cqRuv7
lhKUSeyJ6/nQWaiDw0eE7d4OFL6cLccomcU+lc1Vj5jX0//TL3JosWrt1i7IJPMG
9BVUQUUR5K1eQLSIi0g9DE//fwyI4x5wH1hehGr68aNWjGk/R5SyRjk9WXEbBNz4
UeFUhxH3xMlPPgcB6qi5QmfD9P94J2P93qhGIdS0F+lXgv1v+/mNAn1k0KtMAjwP
bJIkxcraf6tlKABctj8wwsxCHXOq3LhFWH1mUYSUcx9kOVkaWAuodWS+sY9LHgBe
uKBddTWS7AkbGxsRUVA5w8kgwsFKf9x+zREMdBlW1Xnt8LZmSV9yc4kqCDTCgh2j
5P5YcGyF3ycv24uAgm0UFd8E7Q6uNUj1dQ3em3lpwgH44Pj2Xx9Bofdu7vjCJlar
HOABp7tbtk7hPrX8K/mmhpI3mhWpm6Xe9sjHrUrQDCyjQPDtJJKKJx3NiPz74Oyq
FcqfjXR9Vb0nvm4wK3NfuqstNSqUicOTdipOBEzJONEiQK8ywQvaAynHp8y7WrQ/
yK7MU6Z/EpDVKetp9MFWiM6F9r66I0bveQy+uvc3V9mkKf5aBwRQrZA84V2NED4J
XQA2UBe3bNzPvhtbGBlExU3edMxSPn0QFmacyc7T6jG/ztapRDzlrE8XVadUF5wI
WtGHp79hOe39cEVLhbrai6P476aDf8QJzJAxHyZdcYotrBrUIuReJjl4ABv7rjTj
sLB3x/nVT5ODqkq5/6IMXJhrRWwh2kD8apJRgyDL7z57nf1SsXD3hTPi3hYwjPb/
8FM2EDdX5G2a+nzBzm5+ajERkFhYL80bZiZ+P5zPVksShPonI0mPGnjYh9oHw9U8
bELkVVilTO5qA1oD1rTIQ7nQnLE4uQUFgtZBGniJ4bLXVOryVDD4JIFZTgD6aAzu
Fo8/9oMmlWL1tCNsdwvSpxLXFAjKItPlMHTVrHC+kfi2kMWQ/78kRZNDIC48xm40
7qvR5uDHoluyGsNcmWtWJmbgt71UC2Vf2kgb4owwWgIYdYsXYn5bebTi9IyT3W7V
FKv9tY0qP3dA7+CltFbJnKC9Vh0U9fAi3sooA0vvHui/xTX4vKlNRZMFg2GnEab5
l1W8XNOs1gIyjh83SB9kujV2JFZfOdeSmOC6nZskLj5k2md0Oh4dRuZzBUfgPdeN
euCOyyzScV3ZgkEVfMxkzTHKQkTgcicQAXt70cZWPX1/R++uokxH7djPnpVSFaRn
uL46THXDWjAYCvzE2egsosBfl96hwgdKcUoU0TFnbcqTmkRAIRD6inzB51pvKToQ
xtaS6x+5YNg89dfz25iCbtfROWP0oxDDYCB35zDot9NGeAbnZlvOnZ53C+KxTRo8
Di0KlvPIrcZuIh7VbXe/udbzv2EvQtlEWCTEiNh3Oy6irLYo2S7zABNSYc590p6I
elimS1KeYS13E3MQWjKn7JBM8bpvGAD0vhncL1VcXfb5/7MhxNkSWsAsuSFEj2F6
Xxxca/d+4k6iJQqqkoUDy9jl6qZzBqokz5NHYzUDtG81hp1R8daL2SKQy/E5Aknu
bYju4xyym9GyY55XOFrhUwx1vq2a8ho00opH3dMtOjsby3jGSkSy/XcNYqF0Ht53
g3+Zr/LFAHkzCe1QR4fd8lClLNRTU4x5LhAP7IK+iREeH5mBMvu9VxdGvqfsbfaU
vjZWN0qW2WxDHaq+rV97Xxg1QHCeGTpMhbCzhmR/ump9O2VODRSSF8xiyrt9Nj4m
bb7N3DUB1VnOppZL40UQhtrN0nlOWdQR7Jc1RABjHmJ6ljJdLOsnGnwT8o2anREc
Z8QCXISnlVzKuogLX2MpTEJ9WFw+NqBa9G8SauPxVMxRYZM2dpsAflaze29p67hC
1dt33ULuRMbgFJifdoYyJkvocKIRgOP4L4WGDrf1tx30FJAWL2IzwP7tuDDzVhjh
DiUS905Pz7oDF+JqDUEKlFqzvpZOuC/z5kgQDTnXkvLvyIoMj0D8cAS5WJSsprdt
3l9F6oJx2tfP3pqVQfNd2lcl+V+SNOsBpOtprVdyW9NdOLdqGmCXIdwgmFtGqrPM
db9FR/25rqyQi0YqVV3XpgthX7UOJpICFQ9k8RY1b0DlAQAGWkHL2ueOOrEruXkn
tl++FCKfpKeDnOFhvTGh4f59m4Pt0ztjqkWPaFBb3t0XgQ30Qe9+dgoPdWoCXDSS
DR3hPMaf5XwEkWOdsNp4YG3w/9/8cCYifiXHM4rAKVZJIHoNdnYR2iCWIVZS/XqJ
Gb9dqhxgRzw9kWhgHdVfy9T+aBgjbVMj7KRk+PKI97qi+nzLjnmvYlbNsXJi9eII
wUfyRW9AyFKCHqTTZAUhedYozhMh5VliVgBOJmvi/KGUP7R/rg+bc6Ijoz+TQwXg
Seg7U4wjlnDglfDz+Zd3Si30GPF7pqHFXqwI36ckRrUiLr39nn0M6pxIpliARg/r
ARQPW3STtIDVlfwLsIISUbIeE25PeecSUmGyUChlhGcfVoAKw5HLjBOj33RZKN2U
5+2ykWo7u/1tG7tsDFe6WOO3+wHYK0Lkchvm3adEbuqaj+RGLVtO2y8Sec884CtG
eLXzK/LlnjR/gXJjq2t2PU5CJWyGn02kmc3KftITFWkXd/1lYxQMxLyAylK8vp4Q
M/hGHSevPXLYoGO/svQlGdVOGS6Mxa3utKsP7KuK25vmxvaCCrbKWYUBkl9t9016
vnqHhKuVHEQio3ujFkLBkAKdu2w9C3Ilhujny6doqNkyVGyK3yavyiEcRDUWwGeK
Fq5MmRmw1/HAeBskf4fa1Kw07uWZipVriEeIE0nB8auRH3i9vhnTMVSnVNU1GJG9
cI4TzhH81d7U7gERNAUOialvLYTSvcY/JN2yURFj9TDPQrH/dCVh+r2fbV6p72n7
2OedMaNt+e/s+Ecd6k1Mj9VK7SiD9UFb+W/bYGQ5XIK6yJwqd7wJ9Z7llf7Q5NrH
aMcjOw1CVLV9tJmbSgex1EMXmgMds8FSolbOzCJdeL7FAeXHgk3t6hgRoiGHdJ6u
3UBJRjtxQrS3DWYbDQVzDyN42hlhhJnfww4gIx1hkCRv1opjwr2OETCGjN4iPYn5
FVABloiRo8X+Eh4zpU2sUY3EY3pnAb3HgbsVLl2EVIabqokmCD+Cb2uTZm/lJt21
IDJei6Vq48elhW5QhTmHkDDFXanjE8ziKL3RNSffQXmz+QkcslROiFhPayu4c/Gn
HywDecbf2ZdbwMwlartXeC5dImWSd31BNQq2FKGh/9gEtIZoOzDB+C1weEq7gnEK
+AyaHqK4+q9OuZJUY7FEjUeBI6l56qI8qY/pUsHtoX3eylgakrMpW/FZgeMIVZw4
8YWIrNg2z4pd+U5SntVjFQ66PPzsTaazg8rqgjxrDVeHNmsb0Z3ueCH8DC8LMIKw
d4bj09J/mTu/tGfAjnjNhCSHnbKh8iU/gephqx8cWEuj724Rgk+cnzYnMAFa19Cy
FAi4CTgQv3cNFiGMnj48avbOxrqf19Dq0tsYwQJsQEEM1IOpJeP5y3VitdPESN2r
31VuuM7YiYxQyvTw9cMpph4ot/qoMCeBLj+LG7Mw0+t/uPGJkclshf70ZeibPV5q
zZ8QNP64e+8N5v1bP4/JlWJEnar5CvGehWJoU0ysc23LwZyQCGYiIm07d4yVv7md
5au2fe8j31huSvv5BE7R/3U1lJsOoY8ms3f+M5j41eiclupzXe4pp2nr+MRdaL8U
QdqHkiyxW4I0BJp5MM67pPo3J+++vLYbhGJDiNKni6CTMWyYN1oGggbXz3CzYVmA
mxSobNuN/Cimi3anSu+i2O7ckCofhFTwiIMNoxYkDZ9kyFn/097G104LdZOxGKgf
HZKGaJYIsKcjd4UUAc997kD0vME417OmrBVKxVVmcrblL4RMa3ffFMqqcE36AtUk
BAw6nv1IEHBXN3f28l7ldcJpK5Ktz4aK0zsVF1l87IwCjQEq+6himaZkPsMFEJJG
2gd7tIvviBMOHucpcPzIV4Rs/APIrFGLh/RvC7c+WFFmxa7ivHLMqf5u97nsJBGI
gWVJgshdNvrX6yWXzk1t1E0VtyjBHsWPyJoS8vPvQMknDSyGY/9IhgWBnpnLFw7U
ZBbknGdJI4SEgQ+9qgDtc3wLVONNEL47xhU9bjGtIMZ0DjDUabFYMwQ0FVLm64rT
5R18uQtJcP5Ed775IX5mwXwZGqI4GxejFpna5V8lEsuJ3OsQIoMVPumsdnQS8Lom
zsGDJE6hkcQoCCePVyEsX8JjtVzFhICeSHWzaF/9KWQNtEWnzO4ouAEhVPQkeOz2
sM0tvg8OqQ4ZqO6kjaB58yfN1Cjvk6nIOjicsG9uj/i/mNeSFybJe5G1N7o9R3wH
vsUIHbp67YRyEf49MY0oeQYpnJ/QpPv7FFuHsbuSU7ys1nmLvp1MrrTPP5qwe3vr
lUx696z9dlWVydOVFVMzrl38O8lythvMBTocFHyoGKeI5adpdzKQ/DLSZON6eJDy
qcVoMSipgB1OqUqOGD/IVJBRXaMnr11aRrfZPBFh7oTzehKFJRVlWhlMPH4FPHHQ
N+LCxBFIsqzta27IFM4xPvHFTT3rJV5K3Ci5CUnDIv6rE3txrMCm0GouwDYT6hwB
Y5lyCEV8Dg3aIo4y1YysVJFnwDLsmQHYKKGvdpbyEew2ggQW1OzwAxlAEHQL4kS2
41/ljuicVphjJOuz8zEEEZbVNrg3ubqsEuk1XVw23KGcg3EeiDgwjcJpZvHRf38+
dv87f74wXWJWH7GhM4OymtTk1IOhiRkZFJ9tPGsYEFZOXg2SMODIfZiiGIYphaGc
i2g/hHcn8+Z06EWK0WO3/YqHWNDJJPAbtQsePFunTNQt2zv51oWcpEPBzzZe6g5E
kWSiS/LQOElJ8VqpM1bW1OAEJ7kOMTZ16+k20Paa9uQMrz7JZTOSWVTGaqcf7oc/
RyYoTxxWTGoxtsoiZxH/PitagMtk4OyZO5o2767APDEp7BaeoluadeE9kbBLG/Fn
cs0jL7ylO/sQV2BZn5jrpd8PpuyXH2kR2VilUS3ci9Ip3cGggxMtzf2Pn9BI0Vu9
HvTm9DfcqXOEThZ/rWEzlhKw/82PvN+uUkIs/GrioyAudsOI/5tKB0hRPTCnujrc
rWbzmk08Mf0/QLrY83zzZTTUQHYST+xr7ZIMwwEidWpB+3nzJ26O7j5/4/QR1lt7
1HeHmyVqkSerxV9nFkFU0CoBtOfJrbR5bEXoM9WxV2VVMoBXI1FUXRp54Y1YmFLu
dcZnALncsWsuxFyOUyDM5zc2sWv7DzvWmavTdfRVzal0DZKKnezYzXjOTC1rAi4y
yx3HTBdlcyJqSuwyZnigob+29xBPAakix6iPgHLXnfVdFjSvkxgCrkx4dXE53c73
eaWrlHcktn0Z3xii365BfVjsyfwdocflmQqXx+Y843yqWN9IrGRGCUOSB5GrYOmp
Oi0Fpho8N1o9ss/QBeu758mcLPx9tL5aqVQY4eaaMZrkJwxCGuM6mkAp59WR7yRd
c3G3tU0nl2wq1q8gp7P11HrkaybxB12hq12cl0qAhRHvOxxF+i/JJRp5A3dVdOWp
f0zK5UtWIFh4+jHLuFIElgAL07zaULfK07t3MF/8I/kh8Dznj2tW/rdCDVWlKZ7C
dWMsRVwMS9bXjrfq+kSmddLiulmzWFoffICt5C/dLwVdarJ7bl4ynSCHFFDHMnk1
+aS0TNr4/D8zxBlR2k0SbAOJp6YBaI4yu8OctJTD1OeZEH+YwGSrgwBeXoIKAsIP
VaM4euTFpKhR9R6GU+QwdM+MUqIhOkIj7WCLqH9eofeHZEGCQynttAjFFzz8tOce
Viem/eqd9PskasOf3zcUOsQGWoSrgoNeq6sPpOlNmwa0LvHSTHN0Aoc2+7BJlHOu
1CiyA4qmx9r9Rmlo0CPx+9deU2Y+5k6tuB+iWGu1lnM6N9U+zZVno6EXyBwGEPcF
CC97TsP1/L/+TS8TDvqaxPNElUgIPpVMMK6lBJ0ptnkf0n3TM+m/l8FjRPCBw/YE
Y1+Ydgl8yd+tRlgaZllo1V9uX5RPwi99/fB5WOiGXF/M7zYvh6XfS5g9rVtIsBCo
JaqzCVYzgW/pOF34fxgYGGCPf33eaLePjN4vXmuTnNQH6h4eFf9m3E83dsF4JKMJ
xFSY70orCkBEJ8Coa8uR+RuQvgQLcurehBMHWBvPyrjnX7Ft2eKjOe6JK+jig5g8
EoLyDUb9CzMJgH6jVyPDMcCOeHJkr4aKvqN2GByelARx2rqPC+HyBu4KXTh2kjtO
8abTEqN2ovkEV+xisOLgoXP2k9fNOlDQbP0bCE5UAUHB+Mna3ljfqXxmNprxGRj5
7nr6fncxQgY2vjBUXb8mKo89SIIgcMGX2JYvYCvCnzqdlyD8HxttGbmuU4vgfIPs
o5UaE5axsHlcotWqiAuAVNcEyuf6Bret7XmH3/1PGcsiw5mK1LtNY8jD7hbrZrzk
bl6n6ubtOEUcbQwvTn/RVzMlrlBeau4KeKSHSoPe/hnU2cdd+b+atlk6aL1NrIC9
Ms04JtpRfU6TXZrLC16TVfCcVVxDw2FPVEEalW99erIZ8658iCIMu4OQH1wh1ASq
cKOJ0l9891ad6eTzyiwHJ1TtIz01Nm1pH+Pyf6N0/O1ky2D7TFRIgfa2kF2JKXTl
4xCz0E78HeNDDpw2+lw+NAcsfPHeSGrU1pSpGQB8Qa5LuNo6jYIl31UIDXJUbSUj
I8jYm6oO3bgfvC+4iqrTaK9/gVDZkIuRlc33ITpN3RO522oL2P74ApO3KF6cBQSF
HGq8Xv0iW/u8cSQ9NStuw2IwoY2ZYGp/k/rYRM/E/kpiIl5VHCOT0sTHR92TwiyM
r1HoeBe4MnHg3Be5RPVlBhc0EM0t2ZFQ04KBZLcOY11K7OPTF01x1AOPLpxiCURT
qjz3GzyY+TNCJcEOhEysZg2rLbvDB5hj4EGb0JnUK9EOe4nAIDWrogDZASFVHuH5
sl4UUpt4cS6WwI1zlgvv+PYvteMYnqIK6KsXp/0fu+t5tlpHGbiCIDGlYDYJ31Jc
92DxPsAxfFTZGTr+5F0oGzHqFzpt0mc+P28mvQFBp6LlqkYUbEpn3Zusq+eb1MuA
nFZc0bGb60QiAThbz4qXAm+ka1aXwqhBdrag6md2uGjixG59MpyxYKjJsXkQcJfC
yNwECtc59kktnCyHzZCae6BK0zcR5t6eRwY9yDXxH+Lk/6DVJ2evN4azCq+96XsB
8M9J08gcIxT3juxLMAofV2Q60A0PMa9vqWmg3KbfPVxprzvK3oE1pF3TlfPfnHPM
jyuHfHcanhprJMux5kNIdk5BEUxxc+AaOnXfU5m30LjUjqX167CMr6rYDeADgW0r
tIIdZnRVhYs1WAnuUH6DaNWo31dHsCn2fO8ZmZqXgY7ODfgbCmdjNPffc1OJXlx1
0bAWd0ugQU7jIelBv5eWdX2GrdcJm6p5uXw08K2KmQkYhAH7OCD7UVm4gmLw4BvM
Ig2CmHZoR5C+P7keC1d/991a9lX8dZ8/h/Jdn5e6P+MLaS4qxGkifsnUz5DQGf59
K29gPj0LU3nrR57OUucmkr84Jn+yAQ7FRpubv8NjofY6zmoP+usSgifkNrLxmMx4
Bqvqsu6RAHVUZpUW6lgyYdB/Yef+e3yi8CqmoK+3xUzAR7UktvhPMQUuuhmbhvFs
zLSZQ3lBW7Pl9Rz5YB+SPFkCUe7OvRsZyJ9WLAX2n7qi+AaQBvTzMX6TDqSt824N
YCRvJYn+5v8pE0BDCIgcB1TK3XTe89SKTdynMBSN9KIuhrd1zy01MsXkFEVJPl01
YGcTjrxgCBrI3GeqUnWQzVWx66hkPNjI/vC2qTH/HUl0jjDKEJSKMhyha9Su9A70
5S6/1WCBCa2d87+JOLXexkbeRP7fr5ZuRHRAWJFe0Z6g5pZyJkSU+gePsmFJHrrq
ELHqVbNm8Wd1WPK5c5cAbZm9FKCjoaTObvaLSt4jvShKOpHY1MY+dqLfMZPD0Qcr
9JUAjCH9Ft0qnWBtJ8aqxhxbaqfd6C1UOzc0hdhLdwPJ2RqcgwWOQ7AVEL/1LqJ0
TXK8S3a+LzIR46X/PXHy+ejp4EVF90jyZ1Ed3bdjn8GSpcvt4dBWMtoTBBpB2+/Z
DIJCNkjJIcZIJvgRAqvFQAku/slPGlc+oNkucJKNYRs2m2bwOUyNL/L93OuLB0tY
vC0Cbnv65AUfuOBD4oULGqyrUTtE0xA4E82k4StkoSqApKHgILjnf+scixnGUVFp
aWoW4tUq0dMbLF6JdALb0WQmAFJ18HEJLL6eY92C8taLiK5SPLqYKupJ8png2ecb
m8tFmgKiNnvEawWhJOQ0JXHIdNOXw6SNwSXSUuF5e9WXO5Z0EVXjh56S7siUJtaS
2lxWNyRA37x4yYVHGdeJg8k0wlUvRlOvhcVNpFIDOxD3Kjtg4Yek0ZM/OeFsGV84
tkcn/EodmQUln41w3rAPRhV2YMDvsRJvGZUEEBkB08UvAr47W5YjosfJ9peb38QH
eVSy9E6BxXvaOydT/0WzjUi3Rueh4XmcDIjyVddRXoMUrhZXJKm3qMKGczhZ2VBM
zT0Lku8SYG83KfhL6BT/ebbwyttAysvyfCp2nkpuTO2cp0LBL49HAtdMBIihaQqy
L83O/xBLgGyQPpSreKEcNlbI77DRipP+8eZvh9Q4QgSBKy9/GDPZR9VMnV4A0kDy
as/NA+GIpjbBJ7mQ9H/1mjdvNyGuZJwh/T5g+g9lp+CfnGKQmQo6KeO2hZ+i6AlN
bIYiGCRAgzeVwlwc7DjaPhAI5A0fWDyeXaG/VIwCbn2ttfXKwRbqxkskajCba47Y
r2lwNK14KkSLTa4YTvODzNJBmiAO/ncpeo3EQgbrgphpLbZ7dLz56cqAnWBLawnZ
TCaDu89Vmo4zIrD5E3gRgR7hJUbyGO349366nj9Thzbma3y3YJ08yXAlQSfQqbET
De6oEOQW2Q26kLFnW9FrigxUalTNOGm1KSb/V0mc+0HKhAJ5Bv+UC6EJN6rEjGp/
qpOwjGINOxgDsrGjgYyEFK0N3NIPaxpBhOKZBefpdcCaar2fR1/tf0N8b4HQxIyx
y/DXXGSrVYYUnVUuAWNiiQ2MxxkEY+Xpovd8TVoUn/smNmx1c22v6cQQCwhVOqVy
PdhfcGCJCLt4xSQoWXUGEjtb1m7BKfr2JtlPvrF0ylgJBIyfxl7D6tMOhMqOkp8I
nYfS8XHGDiuIspjufvpsJGtv0N4M5ymdoyhCaEU+oLUdJjzw+iafmPbmJdYNpGNF
/cMUL5HL+36H7cieSszFAqJTL4gEEzNtocTqo8729gRCLheMzLr1LTGzsr4rvk6Q
WxGIxgSgXZCSXcpHfsQdQrQhlVv4hwE5i2/+Jbmzv0pDEkL0t643zqOIdvCGNs07
r0uEGLgiLE0QJkFFLb6rGjJ112ONnVYdSn0LUKon35KIwmiEhDqxJgqHX/waByzl
HsFcay5zcvIdYEuOELzJTKn9CLtrlqjBekkiR8krAS51fLfQp7nJ0wUtJXVIQw+Y
vVMq1wsTzX0d6BZNu8+i5Eto1Tl5YDTvBA610q8hYWCZEcd1EGjBvbDWQft5CNgY
QUnoECiyR8FaLpL0mdqpCjv+LnzctfkT+xcxebEL2efcGhjhJzrwfZCnZlrJB//l
ejYHLxYwBLHkMgmHGp7CyRzFJiAoNcn8Hw+UlMxUz9uDyM+gK/otD3JoEZCLZz09
FI37jWZjQuYWfwqbkEYMKQwlHCN8TjBM/kkt9g0k+ksMbqMEh5GBv0M+Km6D6wO4
U4FY6r2mt9axX5o0+w1Fig7OcYZ6rBhvfyVwoO0lr0qlPyix1SBzhiAPpEm7+6xo
PpvbJYURRfsJonMHv3yE3Xhp6R+K3WMNM7ckxLpFUU/itSNM9wnCIG40GF7C5Ur1
QvUbom6srxSyFGaKcd65Mb1DcgJR675aCQ8cKYLKZj0mG1S+b+1wY/by1LC8NJ5W
WFd/Hg03sxYFwgbfsBAN6od93BXqVTQMbSPH8Tfll1S3UMqLsqH7KBbLok1BgALX
fWdfBocRV2jhRAU4oDr1nV5+QMx2dwFn7x49HnTilEVlbgeEBWQJ/NXK06jcQoiy
cO+3koMyEEPaHoT4wYYSoL1zbhqV2jgTGxdRRYwaW0+origbosikxayMAY0krlk/
5ThJPHPN0cDNpWX99RI7haBGhPOqkMnQjeu6yNu20YriqSilmV4FjcBLl7IHw7hm
lGvGX/ta3rkljUcRJy9ge0C+AnBTkGmbx+491Fg/W5DanYFeUfHjNMIf7Ymsaqy9
K4jyTQgkOSo0+XsV6AvqBMrh7iB1CVkf7UeOhHfqT8Bt2zDSkgbtYDNSvQcMPvKX
dwxtWH1rWSuDuvuF7gb9IiP3uuc8JGrRA6cQHqSJLQenfYP9blPe+MSa1jon/Sa6
mocPObNa1iVU4K1hm+i71wTz0KKUfhzXZjf2ySx5uZqKoHYseVWgAnqaycjCKrH7
3md/KgbE+GnKdUxVuIuHPQWRZVUGQQY8uAJoZToBwd/JN7A8a+qgEWqP92uReMAh
l8bZla+PJE+U/1fG4j2aXP4bv/sPfa0UstNtFZaIQh47k7bHsGPt6d3xLuYI1mDf
kQZ0zwo0ZZ/IFz+GUG6ltqb2cE4eICwN+3LekIA8MOyoqmC52baDaeQdVZomBdTY
imFjozG3NFIlpp7mc1f+iPIJi1cYvwlHNiK5vwOMfKFrTUMA0jY89zgZTzT/rsM6
QYT2AqVovrFFftf7XaT1JnS0I7RgSVBNvMnL+joii2xRZFFSMFr/WcSDj8NFI+EC
2WzVo3VVVox2BrpApWuLviLAcnsahAnR4Y6etevRJTX4WsawrOH2F9bn0m3zmf5N
c+gJNlEE5+UbivVL+vQ7CYG8GCLbt+uiz4NiV8lk1nuJFZlf/XGjY6BafovYrdY9
CGqgpbwRE8ktkTJc0E4nuUPm734I58c9+3cQC5ttyOASa13dKi+1oxg0vYukSS1Z
D9ndibIf5EucSL+KQhLvXxaJt15w/QxsP/Yn572xZQCFgC7HrLea9EqG+PAUQMqn
J+Q0K8leSjNP7mvqPPgtPuLsfLvHklyyZinwzVq2NBWuvvA9ZusRyRt8/R10u5NG
EUz9cQ5z7n7WbGsrNM4JOXH9AGOqAcr6qqSyFu8Hg7wDdkVUwg6wUueoan2+HwO1
kWdllKbY2wGTBCzl2hsV0rXrEoPBJBJiUKttqj0+X1ZfPK6AkdHEW9r9AjwDyWlI
M0XbRu9FVriNjbjoBZ9ZudjVsuKFvG7kMq3tNgikoPVUVoxuz1KphZoPErdKFTde
RHyexnLzie2QFKyiSVOo91/JsNmL+2BkwRYmqBUVIDTG8yKQFwClwVQZ7GJwn3ei
gUHnnWU9CzB7QoLuyFRXcp9qq+zsIhw+UvkGMfXpzZgaR4e/fbtreYw+AiqY0wUa
vmwRlYavM0bY4nkMVK0/VUZaG53QSzvzpYi+o+P2sUEEIELnZ13r6YbwlYGYYOZ7
j/Rnt7E1w6hqk3Ge/OkCCxUEf9u/aCUVugGZYX3EGsjq/2+2EhpN4zGDj2xNg90y
PCl7+SkbTz6T5Sz4KhsCXCSjx3qqD2aHKnIFUrEW8lDXYSLZpZNEy8N/7sM9lX9e
lZBpQmgTrJj3XKjioC5y2FqqVXn7lOw+N9JqDiuWlvwJYiMgWWR3lKEbBJ0lD4a8
AER/U4Ij8lm8FeQQGf7QpLwBuq7hVBlhWKbTtrPVq+Nx2jRu4BjXZfNQ9v5k5CHh
ZlsUZ7ngfZOdJx93x2FymdBtsDVa5+NRG3bcN7tavmkUWpQq1udwk5Mq3LonI0+j
cnjF+aNxU+kvNXk30USh/eHKXIrMBlvkD3CDac4cvG/1T41U4J7Q55RmBsFoYFe6
cLEDFAp48tfwcr6n/Hfk7ru/eVdjHMaPyx14CcqMQ7mYqbpoFqdFoxF6XwyjrdOs
q2oqlwInlAnGTBSAIbI40Iowz++9dLA6pSShFDEvXeyx9EkIJQ49nT66iI0LA/7t
sJjSYuj8DBWtGeuEmf13LJovja3ZclYIUL0M4jhjoLUYcLCyzuf1h+l1rIfwgJkX
5zAdE2dXK7VDsIMkLNeZnUTpKNXkogZEIzUl5bkbXCT/CGCrEH8DkgYqz0SBN7us
FvNPZH8iFwyjYMErTiSD8VfkIloG3PPxp4pPuxYdnoE9L5P2ol0sQr8kj1AtZLXt
6DP8QMRN9GDLRqtevVPmVg7B60iO7Ybs1OYMPT5ikMQR1x6uKeELMicQ1lv0x+zx
Gp9uVQSj9MZbUwMDruiquqRowaFXSM0BtM21+ehEfeRpwSTph1dszGvh+Xe6XtE1
RwG9x7bNubbzbQm2LY5vwsG1YRzBkoIC/O8DShGzsnFVrYkwiqwhfBK1NNoJklue
YqsEl98tGHWG0Dh61Bk61ynhwNkLjz/jZtofjIOP64cp3QEUPUO5jdZ69buDoldL
WyOuwtbY3BdlAsYlnhSNAspmVhQwaAOjG8QQVEjM1IfBw7T2Tub6EqfO+M3I9hNs
53WqnrSIsQ/ZZOZEp9ghfwRFcoUZ1E8XTgho5UM4fdzGuXf/psE6abvTHuzJK4VB
oNKoo8ugEJoWrmjokuKQmZ6oigGmj64m4K7jSkkJonOHwCQ+Hg9JMdhTPtgIXhyU
S7SghDmKvrAee84zanqGozN0WZKgrWMsJo2VE0JAAM35GCithHtlIyGKbif/twEc
790PUMSo+Xo/HUFHp25MJo1LAuViuZdVL4c0qjmNTLIB5igSeZ5rMVPlg2jJO08V
0612WEPrFJ0Opo9DDBnKOnzmrUjbf4sK6fv/FHui6kAUgdOPOF0w0zuHg27HJy1i
CVJ9PsQ4myzXVmRx6h/sMa1mGAx03Zji2Rg2FWLzI26zzwAjqi+8tU+Yqcg7RB9V
G0UULqu9OjzXqIvV+vQIZxf2Lkk6GxEvBQV0/7wDnwUX4KhjqRU2g3yj7I51MkHm
nv/Lnw25NvymX51aczD+acacASAtCiUfSl0flwFr2fUO2rL2/RptpuGTndrVa3c4
DlP08rq+cPtD+Lcqya7HpwMxoAt8tU/eP0LDhFoQIe6gAr8yNx+MCBKBJhn9QXju
ztzPA+5VKbm3rbejGmHFrbBY6k7vlxrQCSppGeUApJ1UIPTdKfZ4yKR1zQQAsqIc
MLcVbWHhA/O1hvmDTuBkc6uuecWsKAkW8otG+BVAdeCPb9ZfbYu4WFT4DdVpdgiO
p/VZ+CvBTjsZwuFjBZpr5x2lI/oePvRkw8IEkRQstARWhA/gi+pi/Q/8e8kL7WCy
TvZPzq47kKYalo+0e6+DrQZjxQ3bD25LnCoLaXsG21052immGX5TA+e1fqep9a4z
mAhSLiQrNSeznsnvWXBYcZDqYNBN+eR/linMazHaGIt+aE9A2xjopfNb6ZIP/QAY
oB5o+898YglfUtK+lnrswlceZIlU/gWhfSC6sn29jMc5LZTiIMlbqHsET09ws6CI
qvzCSnS/KfHnAic5uQ4HGmOSzuWeXMKmP7vwXmC1fyxcexuVFDewkUdfN5WaFefg
EqbaPUb3Ejm7wvqaKWNcxGLoveA9rMKOb0dhfKWCFJrT5tcq3ULfsiznA2aTgbmt
HLH+U3yLhZ94Oh4O1taPzdvsPluL/JPPD0780j/ksDcfXdd7L6WS6aDsHE8SvuZy
p8tli+yWSUcj6vLusmk6F+fEMBdxTiTXGl3U4OQxtRTTklASPGJrwQZyYUfTVf/I
i9UiEPAi1yyHsF28CxnvHj0Aq498qJMhNE5aLtGjZ6/iEFbaX+Y30NPwjIE5WsTd
bkG4POOOnRnRK/nHuKfMEo7yrzeAQS7HeYx2x/Td7LOcS+q0gNVxVsUuUoGZWWny
yf6f4heby+jPAW7TbIE2XAn7Z5eJAR2Q2OpsvsGy4Vq84MTSk/d8gqIosZ6p6ljq
59m4NXz3FURQWdL1pcPoodjtQ1w0F1dxm1lK5wXGAbV+LwOOwS99Ifd10mbq+BgV
xc+7KDNGMn/+RATag7INEgbGt7AUHmIewKYg9FM/cAE3Oh6zO9tpEgpqzRiMRd1e
7duvOwatzTzWO+9IRXkhyXt701c2sZ8WAg4JLR57i8GjpwirbMB+hNrrfIxeTPsu
NgKuTRLtwoe1TcTWuBae3h6QahZLE/BWO9eZxt587YJEUrtmb6n8guvcx8E0vFEj
7B918b7Y7gfE9G0oKT1/fouRtPwUEbKa+Cxd2v3ffMQZ8T/FXOqNXIPEBUhrFNCU
q3z5vkQIUdPThrktugEgmlVnVfW/e0ChpVfSEU/jmGcSmV8U/nzB9AXufcDX4KcY
53AstzjBdI1x1G5Y+/1/nLvCs6w/QoNIFwIKVee8f7F6+rtodzHh6n/P1C2Jzwrl
iUEM5Yk/t/9jnOBQIDSR2ly3FhIvB7GRV5IfWsgk555Aal6UA1cULXcaCamQAFLq
dURgGinAfrGBNpKkOf24FIiPK4eFmKGGvOeh+5y4cx8UxekODIeMJKfoEqZOwTcW
KIzdd1hxLr6M1Eo69xFwJamOhJS05iT3W2F2EAFyMWrkZY9+1+DlHIUjO0qCUBk/
UXsHfANBXJxA7RXPtockEr13cg7CUt+a9YPpti6VpZeGjTeICLIvTumaXLX8WFFO
OpcAr9gBVvJYU/DV5gfXeh8OMkwXT0uUxrSzITo+0Uwc95psRCXQPxgY9REARYFg
ee4SNbu2+vofyo2CIvJxEiKYLcLIwlZge0Q+hpfWCzkmE+FW5M/Wicxm3x0z3AHH
GA/fODZSq/Jxpsq8XOj2fgciH3Mz0CHVRyt9q4Bl5LRznJWedwEy8KDgPo4krXUe
s9ggO7Xsz8D+j54h0c/uHOf8HqR1iLUVUnFBb8Q3u7bIQm0Ov5M92EZQYli4TrXa
tsNtAJ0U46aO2cLXKT34Qjkog3ZLHRXdGOH7RoV4GEFYDMOc6EaOctOKhRmW2P2b
cWSgOgoL5Sljjgtf7O+iMZY4QmVgpOKC/VYnPfqrJKlH44azCqGDVk8JorZJM3s/
bj6ljXJc6Ip5SMM1Bf7Ymd5dCHTCayou2k0kDE8nthNXAWErNCd6/Bcy9V/TSVWr
vP5EXLpO3yAN+Srba7VfTLl8COMPKTyq+4VWwdS2jjLMSt8pIyLxTlux+LlVJIOb
fcauwNHlVAc1bN6CZpYp+uMX8efsENWAJqoZ03fN5B/nw9wwYJ6bcMAQxlNSwJlw
TqnrsaIb+r4xazH5mkQXf9xe4by4dHjQPjP1CqanHLHoNOulCxbySnJgdFf7g+9K
w8Pc6d2Mxumv9JvOoge5Ptbk/oZigSL6XEegUgPmfJxfSDVANkCDJtCZTzpDQRqB
AaH1cD+HLfCEVNZNIyreBE+pJdjyPBJu6aBkUwA5Vn5Quvr1I4/uUArN0xmC29qL
cWbW9+RL0ZNWGLwMS1AsUa72WlzKlizlo9LtztSFYVBdsPWNGuhjCO/WWM9TzHSC
rwYNiy2N4DrtygMqKZAGfkrnJB2DJKXD32VgGqSAv00u5/bY1V3zmPf9twtw+UdL
vQmvvQ2T0W7E9JZ78/XiWMValB/7jUD9BUm0tI/RMljziyWmMnHaYTmJAjITnhyI
87LwRqgDylEBbE8gxTqUhC/X4sX519F/tryf+mgwsxoVaiherTVKsvOZBJkrYCDO
UjIKQyCsphgUEC3Xjjbp13WhHw0cHSyrJ3Vx6/Y3FdspIhdlnu3j7J9eFmiEqidK
dGTeUZCTxACHLi5QmtOsRJSpwkKjDmnL+gg1ZrxrK85/Wxj4kAAfjsgXrHRklcE1
yN61sxwUUAUmeAW6/A5Zc5FHv0FmygERn3lCbeGaVuy8hoqC1SVFRd6nV7s41J9W
UpdcKhCQrWXdJV7xGWjiyhd60e02oEXOlYZLT+tMHgDAHO+VNfdCIhNU5k2gvAxI
tKqf/Bc86KN6X2bqcjUA7DzfJsXi+mmiV0kV2zVQoVtsTjAscHabnLmU8ZCj6p9h
yti/1XnwQkrOjKunxbIWxMj6TvtU05QIAt4WbugMh0Bq2bo7Bh8PrYXVVh9DsFIE
0+NUiq5XlErzpqRvzbqhEONCKd//+//hcIM6tfU//D5aaUbFOLlkXklEPlvA5Y8g
tHj6bvoVl1I+dY3455TqadoRPkd3gsnCMjDvJD9gZLWklxGKXaZ2uP7SPAHjnnGK
Xlbxl05f+BVyXesDk6tiq5jTv5UAEVk8+1gURp6rV7IPzvK1z+EYGJ9m1NX/OGcr
gpeck9QMlefUKbN9DQDpaFNMnlgQ82SjOt4nW0NZubuf5PEnbn1ZeDKbDcNUyTvo
q16O+EH67za/gliwcZTQNrW/xiWxgn20PAXgL871FU4RSi2CValecYtVY9y1pikc
RJuSWunHgergU+iPmlY+zOd7wCeA9Kpu6ez5ExB9aEYjA61HmArR/1r4GTzYvqR7
vIZ1ZCwmqKt7he05EXoPlQHsOrVK3Gr/1f7Gaw9is5dkDZlmI+72yxKOsVge/Yy9
zT+TjTMbwvkdGaNFVGwZeO/9LHg18def377enD8thCcDASbxoBFClJeQ55q3dZmq
hlYsGbdBswLJgmrPqQeTZ/QOXD+CrRuq3wJSph5VELCFLU5SUZviEzWB6qwpRcnp
9DbuwJcnDOOeIjmZGkkMkWvRDQLW16JHvpk0lH+Ex8QmENrcSaUrZpb+0AQNeCQ+
a9yFHCqcT2fGORPcmzKC6GoRa9SFVWQsEV/5mKv/+wOiCJ26aIbUEQfFH/I/U20b
Qkxz62r+uKfqmsu8LdYl00QPDea1DHncVRdCtYIXDZfWgitJRQISo5uTeADhh7kY
THE+AANGUjlPnUTfWnedVN8XG1RNmhQT+pF1T5FJgp9kEaAgrgLWod+9SviFsJna
IYBiKd5uFhANeegMKfJlPlhpJebHYbpcoDenf7J+rKfozQIx3TuO4UTytiGAgpNV
3N/Wz5//rqIF0kmKW7BAFYmoiD+CnnPvGNppCAhTBSve6imKfiXhFfpYMk8GAFfh
d1yOj5aWQ9mxUuggxgo+Ah+DLiPYW7cSdDeeNFvqtCl7Qjvk4bniG58Bq+VdFg+8
PbcIsi4guzd5UfTASUk9bdxDUys5pf9zImu3xiXZxV3e5mV2sCd/3klT/5NCNeek
PSXbTvggXGxuBzYWz2qvaIcQkcfyMOos7wJlgytEei5YK0Oquh7gGzzg3W9HaQ1v
RlS7Et0AA5J1bJfK1IUoN7VzvodaFgc+U5j7IJUEqk+JCmbjzy/G2u02jftsYsM6
OQxPxyxIwVTHuvubRJtLAfc+LB96RNbdd4LBHyiC9mLhAi0OMKjWrsb+CJA3wmC3
LkEcSNnw7KYVuODTIZL9wbO1QOXnER1hwXsWHj1+AXVcvcbUkl/9QkRQrciDVNsS
gJIUCLTjlCHbDp03XQk0zOrCxfUNEpGtJ8s6Ioxvar5DWzdsMMhCrCIgR61q2UQ0
pFIorfB+tWwl4MydrWgayrI7kgw5N+nv97erY6tsMwDHmVfhaLCrO6w7wpPIiFsU
hb7t7TO+5F/oPpirnQKg4ZvmVm/Erse7/FYR4AVubGwIEpq/VEvBdq97P09CsvR9
Btc2cTdSHMk6dgPMGW3v7M+lxIljFPHIiNXxa5P80WfkUyBBE1xE+5P24lwvK2x7
aYkukwmJ+nZuDSbkLjWeQ4xfdHZXaeF3mJ51adRzAySohBOTl0+XE1Tnb51vJYMJ
zqlv7ND0gHy/EYhSH5r6G3zIdkWe7K+MO8VbI2PbfS1fSFrzjQNJ99JKVU5/+EpA
D9kzjPnPp1t7uK97tH7YGMdH2RjSIIpEKVPf62Dgmk845vouSjniM5gOocn9oKdF
UnSz9GOSPgxs4MN2FGPbSH9HPTnnWSK7QMGG6httVebLX6uPIpNpCQbJHGOvdr2l
OXArAsD9OwRHBEJNHcQrxMn6xZ7JMs7jIFWoMZaQ0qBeWGMX9BjsqSiUnJrSouqu
HTabO2OBdJX4nA8HW/niE68wgg/DfCmgIxOYpaRh6xD/b9+zBAtAw7i/kvJJz43E
/aE2I8ak4dDyGx3d031XYYq3AOc6BCmPmSJZp5YnzX4mAR5e/47l9Qn8C3PyanP1
n53B7cvuuxUeqx9lgvppP0FKl/gV4SNwjijHc++X92kzW6s4zbgOH7hEcMWISfm4
kekm9Pd5l0ZKIK6o8czoIP8DwBBLJw/2gEkaFL8qP5kwkOCao6sys44DFtHmpkP1
4m85oGL/0dbAy+em3X52ffSJt68NP1BzMHVQ8DpK6ZySzVqtOC1OmUWFMo3/xH3G
oZQWxDul0uP6jCFsFU6HxrwcFdW444L5Pe8NKyyjxiIEwkBOW09/4iIS3V8AVhUu
0byZkyTnENINdIwvcoEPg6AKP+Iq/bR1pBr2IsqnYkGuHkTdkrCn4i7oFGH8VOL6
IHFFkXH282XaKoQ7c6dbWviOX1sEcuBCkPcoi4b3+39Ivra2fLwptZUl21c0bKvE
AjCHO1Q1CI2FQD3KNBwtCNAdomyeUcDPZfEpspl9K3BrRVCkbxrRrIh1iEUPOabI
F8PmGvDyJGZSkR9QHJbLisBR94OS9R48jzO8pA6DNZzH4PzhBUHNE56gw7TBt0JE
CXW+W+uj65CI0reV4kWLWwdSb6VpX3jCWCyzeRQDksiLcmVIM5ujB34op+YGcAtO
0aZzfVeL7td0sM/UN/0Bmq46whwYiIjaAMfW919YfGv/6ssDNT+AZr1HQFnnvBQd
s/b+CbjSe018bfIBjRA8ojOpvXomu7tjjY+Dyw4CqSG00WTn5WYMZ2M4IqC7nl38
HPASrSk8Dn+jdM++FwRJUi//1xqyOmLJqbNMQCLUNK0scEX40Ge1iECLW8EyGCNz
C8vfhVMQVWFXb5bJ975VraRoP5lQ6ZbISWgAC0V31ZfHKtZMHQOzceRez70mix4f
MJ1pG/d5nic1R5aU4yiFryJxdlqEMYRjTasrFr0uvdsAAvbvFMWe+20qxxiZJcul
yHnifOUazVVELPW8SkB7Dam9fNGA4AsZmazTkyDnVasrgV/C1quYZDFJCxbq0Mxf
JbwfpT5I8UJnxx8Jyp4pH0sdcB7DriNex73Te/2+qJz48c4N/6DVUErU2i/HScSH
+ogzA3TNAPIeQVBDNFJ9MqLVt4ypvk4y9do647RChJILFByPzXSOZYdN2Q8Juf3F
Rek2w7v5ywfGSj06+wdRTzUp2tIJ6ganWi2glJxYHJbJAR9hEgJSeLIpUUKixPxw
PT8Yfd9dmJh0zSTH//H+6+vcpDdQpb1WK34rz0YGufDVHdyGa4k0XWbeNt5P4p7a
acrSrgFfAn+DKwESPYD4deJnzFUZWNTaIh4KtgCIrTWScuPgR8dsCTG+Ezbeuyri
z7gn/XtykB0Qka5ja7lugWPJzXZcQfWCSIl/H1jUMqwcIyfL3dU8qFdpHwBmq/6G
IlHVFC3o2vHL6EYMb3eBRIonFWRD0Ue5MqeOu5+WEnSQyGJm02VPI5JM5i0Xkg+l
vZsmY1mT+v4F0M4lRO4ZvbpP/rWeGaxnOQyutkmESLjYRirSEpLrMG4ig7U/gmbT
52PAavTnZjh7WWkaxIREJdi2Up9YCjUBEppUMRafwAFkKd8Fa5coYo6Hjf63X21o
voMu8+sFj5chgaVkhaStxD75SMcIDFY/uqYTyO8MFXe3uSjapnwTxR7/7Dns3LX5
Od3ueJTUzjMtE6eJTFTaoNDI7kbrVlZlp86JwJGCkfO4fzSPPDSg0sOSssXtOzON
DVZheFKhgFchOaXAequwuEzSbJ2vJMLfDS5i4wuOk9jXPfxRp9PVYxEoR/2Fk0nQ
VY3ZFdOdqdp449qpY+KuaMZ0predq1Faa8OUDUvOXD/vdBLTtleB2Pov978to5JW
JuQn5mQVh61DuC8RuyErMuhSECXkV1fQQ+NbaGRYCwP5VO91LLNu0qCkA7ENmCx5
/E87IWrLOlzZW2T7jUZrPp+YM7I2gu/9f2JseZ7j+O5aadC2ZL3lrHDk1m+woGGE
HM0ENSnRntjSpua2mWjeHw+3WM2crWwF6NLaPuG+PxAf4XaDxFtClKliCbWL0stp
vuh+dnVJat5xB9PYWI0+f+qi4Z3Mw1ymTZdP+XEaZ28gH7jVjNl7kkR4cYoUovbe
SF8vtzGI4x9iiESjVRM3X7Yh4fgF4wIWq4GVwQkyBZD1XejNP8UwXwV7FvY5WROv
UMIUwW3uOOhqtmO1CJjQ+7pO/9JnJqHdewkBKojagRhKV0MgzTQ8+lMhGjzHQ0rQ
a1+LHehGQpCRmoMQF6pPnrI+ifNF/XOedrbrVcEZa/dEejAU01HjLUY/YM/V1aMt
77+SU34hKAzUE0/6j5U/E/mjH9+1untPGBjgePYubDHEFN8NqI6dvVe35PkLJezl
Y7qKAjvSsznmr5JEZ5LDIBCwI3SAdXLABnsn9NRzDWadB5zfi/MCNr2y1jSeSEWD
b+3xmXUctv+8CLQ7Q/itkt7Jbag6ygZQmgNfi/g16vjFkQqf+0sUFBJbkWThusig
0eljwluS48iGeGsS4cnqk2xDV+XSO6nblTqWR/Qmtn+Ewawik13CTiel7WQv3hdM
izQl81PXFu6wxPG+cYbparw0j7EPDf/7CYaOiZvFxdFUhxxgpl7q5RHsK32GywFN
vAX2SN51xXz4sT3MhzW2gMjK8puRZOz4GSFPVYq07oXS2yYx3Fi4BPZHHx1kH6jL
uTtp+hp2iA6gxhU/KqrA4c9Zdy8razrPT2qAPMkKONivLpB4qB4+GgL9z2u6JwSJ
snn12YlwgqWDOO1zGO+rQS+qjZRpuHXz0xo4Er1qnw0cenFbSp9vAycARhSZ9Nfu
AXz9eXOqcbH+02r4q7g9mtRWqFAokYgbVtuNjrbNrKek0aDDL6YW8QqR8E2zbUza
GoortbUcHOY9j6XM7FxCCbheczqJdhZxuxHltY9HAWWXvVoB0iZg6hEqbv7ZoGmL
w9YpBui4ruLzqZY8bQfOMZfkOtvVnU35H0uf5cDEmVtANbbhPoylPv7xDU4gXD1s
G3BINt25lK2FrHbmGIe5eOPb8jHrJ8V+HVT6pXruveGJnLc5YNtQ96do5nCN7vig
Z0HUsND3bB36FAFobY4OQ/a3Evawd8q4caa/2pXfso/YnNuRwfKDMPJyqziGOWLc
0CgRDjSOuldd4IOsSmQUekoOBackhitxhHRpnESHqlStWm11Odl1SsmqYte8wAZ6
rOIZtTaOAxwHCnfLL7MU8C4qb1bYfGqkecZ3OqU3mQ1EAeKkKdgyq0AhBtP4Gwbj
/D449PiNRGT28IylnP6+f5708TpYFDtAKAVT/4F0SJNfCzHSNsnoexhDd5+V/cVs
GFN0hyiYsczhMXfGDFf3xrr99iihqr3Uy+TtiKf7HK662sIpIRYladu9CTiLifM1
pj9eDXST7CncU3HiANS+RqEb93AWVgrrNJ8Ea7nfMcebJO9E67ejCa7fXHzfW+ME
15+dptcScuLBiEqHiGpYW31Nvkvq+HQ+Tbl/YDoqxxYKqa0/eIx3tnWo0ixmIi8c
vu67/+TgKsqAxYkS0UeG71Xf1gi9fpv+1HFcQIV2sdfjV4t4pfHvxgSY5JNDL7iy
/yN15J8fCCHeGwz6COZfbnWpK6BdZXPslm8MLHPZ65G75PJJrYytokdMtDxqWVWF
54ghgK3b7NlmBRDciCDtdO5Snxb5Fb4TFaACymHNvS4XEHpRHv6P1Gp5En11d1yJ
dRq0/D5Q1uu3DKYEcLwzRIR1WwbM0210EzGLJfByhEwGGFYDcFaLC+nL1txHWoOg
oO3aeNs8Dpyc5JUvouRUAzggHP7bPv6iKqdGG7U5HtDMiCYcuDVspwnUwE8AGHaI
Sr5BLKfCpvLn93l6lhCDYrOXEI0kUus3VL+S1STS1ijP47lDjHu3GZv7RUIlii3J
QPp3CfbyRZ5c7gnXZ3J1d6h5j4HwQ9jxW276QngkspLkwRqqddjM2K4XMHrT3EQI
bt2XQFoUDnFdINRxQyP1k8dekTYeKB71WLnlL+/WgQwaC2oj7QALtKV/q9cVwamJ
iDNaJ1y/pVTGZCYJ4/Ycz/J31/8HTjdO5vU5HiBp68L7mYKSjnmoAzu7w7OXkJnJ
/y80WGJwY0AuwMZsKd7qPkpf4Ck8/kYe/aW1fBdCZ3XV+6TH8kl32fArS656pv82
O9Btq/Y6qSeqVTKhLLzwfYXjQc9ScfAhW1cCdEX8A8aHBmfa3BXd1zpf6K6zfuGY
ZC8GrlrcVNutboWtIuIdCgvqxWYivEQoSsONKDGb8YBIczrXAzm3lWJCmlIOgZb5
jiWwDfZttSNfkXae5qj+GaRL+W/mmFwBTZB3qJQuCooLBGy9MLSKLDiAgF+6qlC2
L+2a7hRZUrng9WPoR5KRHUeLs8BYKlGYK5wktc9KCpK4dIR6Jbl5wT0U71OYh921
ZEcpWabC+GIzwXM97FKq6wssfTqixgmtbH18D0g0u2UGNZGoowNn9xjVEm8HV+JW
hWhqEv2ZQP2Luggm8Qo9CBSsyDKtc08htFAMfbfy2+Wgswv3tqgfDftPME2877Pu
OUJbvVtgiARLx3h7vRdt2dQ3l3KIeb1z6ptA0GrVKEv+xAVNbwaylfQ/3lMs95m+
Ee+acrn4FFbpRGCpQVd2jtXRZ8h/ZfFw2NgFttd3XW2HLUmfwjYztRGkE3O5UaiW
I0xslr81ZXdRSQVonGvGwIQLou5zez4ADsTVdV+m+9PNRuU9buF0ly2rIXO7bbDN
jFEMaJuHhmSyuCQEo/RGDfBzTftA4sjYt9eakwOApVW/9QzmJWur88KPvNfYaAY4
7mUYwmIJHANq3xd9CSiaonj2YSjn/3rnBSNwuXsczVAqC+TUgGM8p0bViyt+0Wxt
3Ex8E9WODvSieEExsZQaJVuWWQc6tXipSsEe/MV2QBp3QROz00cz4I5AXCUpbqDA
TYmV7wZo3O4jDFGJ/22nNm8qX3t8Bz071FDgYMje/cb2RE7YYAZl0U4hQpBP9upU
3ZszNK0CGOhV72o+gQ3rwk/gEGkClMx7nWB72bwC2f2qNKGMgg1kEM83yjHEscLQ
Q8g2ddM8NkdbkP54pf87bmnSusFjFI17xfWwrSNRRliKG6eU5tteyxYoAJ2XfBlB
+plwZoYElfqYB4CxoxcNzKoBq3ZR5+nYnd8YtScHDXfPh6oxRbHSutJeQ5LfVqXy
BxS7S0pjIytVG2CEaBneC4ieIY/OztCesydPHYGlrpZ7Iw0QVftl9GicgsFYgnr9
JYO8vYSBIiaOGNogDqLSPWQRtnK/vG+GdxwzWIT6DLnqXE8/x7y+4smX5SrXKsam
NkLf/CPPVBcFhfTyosdvkgu7bhtvlyl6qeV9I0u8PMLgCOaOFFtew3RoWQNrbviH
uSOhNrePFgfCCrKHVs57FA6kD9O+3ivdXJ98DFvfhJ4=
//pragma protect end_data_block
//pragma protect digest_block
800UDRli6ObcAvq6bCFy7EE4+Dw=
//pragma protect end_digest_block
//pragma protect end_protected

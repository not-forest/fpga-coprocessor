`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
g15LKjf/5x986XpJ4JauOFjW74R81FC+8KZwsSUFYg8cV3j0qqs5HpsuD88fgjLE
M0aXUKcEgFaoG91HMO7/RqXr1crWxEf1hdOOHJsJrLVc2RsqHi6yQlEEgdKK1v9p
VHieTZVX8fQbgUfBGq0ohWM6Tv1lSUF2+jE8jQDpWJQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4240)
uReG7Ea3a0e4kmsATC6TIJULgIxhxeQUdCPVfwlex4TLEWwgDsM5LkOUC2DDZqCi
bVdVjIhQDhRR9XNTV9q6UpUZzu3E5kVKfTuXaXsie2sRdHtdR9r3K+3iKfiGOKd0
wgVDI6+wH3Uj5z0MotUup+lXvTj3kdJM9k4/Lbv/SlcT5EviUT/bPPNE7LDNRmEg
B4/CKRxRjscpKIJvY5gHRMG0V1J+iaN3j/mUsW0Fx5+5Pzf2SqhYgynKTZMzv88m
+4F+Pq1RV60T6tQPkSYHOQGB3R8pxh33HCcpELpiu/pp+xSAX6pTyp63KyddDTYh
L07V7GQlgsxX33wVgt/BRgPCXBaWcY5OUmK/49lwEDXvysn+ugawafbYlCwcmv3i
Qw2XfPOudH32nrjaWjyqKq67KjYnqsttYLGnaOJwtHUjLJgdisHHzifXP6JtZe7z
WXolVldHhPztAqPILmrfwOjG42CWn7QZ7/2P3lET3WyRbnzP64cOr4HUxoN9BXKI
lJG7+E16axnHgCalVYhJhYRN6jNk85KFREfQR1oTVnnCOxGbm3qhmQNijnIvvwfw
kuIK+EfPkVo778L5WtgW87lTs/ALY4t6pYWaYwDystl1377dTBsJYG9euw0h6/K0
ndr1M4iGiXiKkmNOyMNtmR+YxB4PTVltTWWh1xjjszj7/Uk+mr4FfifCvORvIhvH
pXaEq2SAx3+5tgEH96YTSRLHxK629Hvdl701Rq+kJ5fbKjTe9y7CLocb3SWQxcjb
vcdiHPB5PsifQUychGC+MLqOK3XvJI5nPmsi4UC4Q8MIW7Xv6GzmJYi98q2nWTm0
Mag933eS5eRSm9HT9SGgA0gc+5WO/JN92GeLYrQvmtC0Da5Lq0qhODmzSdgu5Pah
vjiL619CLSCiWmHIiJDbk3LC9sbWGkGBceusGOwEwLr/G1QKM+8YnptumSBai4Qh
FirMz7vbKVt7h093Tk+jWvk5ts5fZQcdThnjdx8gqAAXSqrNYQm5HAubuZRmZKf3
Im75FHYI3GZoIjQ39rjHjjTUO/XjP+TK5YigCMQRspqytOd8LSxp05Yc4iTxtlIp
BdfiWkBkDC1YcFffU7XQDDnHjfTKh4jCDmJcacq5iRrD+yZ1lysDHh2x11x5VlTT
NhYeiuf+Um88s9RaQrPAw9iVMNxczabL9xp4v9C0OUXeovj1+8/OqGywE48HLsgg
5+QLQ8HcUES9OkFuV1ymVqpbYoxjlqXgM5YVANllVlYU2PKqpg57j/sApI6pEJab
2uAnIjKKHA/o9+kPUwFGuDbsF/ZKb+T5lXLP7SyJz7b7ZnH/ctmLGHp9VQmyzZPn
/Pc9SJT9kBmYhh7SjPQG1zyU9DNXa1OcxgXwRKKDdyW9XxS8jt4YaO1nSV8DZFp5
H4QsONc7i8IY6Uu3HMZ5nvAhsW6Vn6NBP8wlzbL/vWFvOqzQZlTEqJnxtieMnqdq
US6abJZgbV8a0kfMdlkCd+NBvPgsu7PvihqIMKTRUzn/x3ki3g15lm97UW0r9cPR
Lgt/b75/315XueC8UVjJTnkkBWLsMltLGJVmewvYBHy2n90NqSpUdTvQW/IEW5xU
Px6JWlGflGbyOslirxjkLzRw0CkXjH93fI5SBl8XyVM74kjaW5mY3RdueainjuWz
oBmMxxnefXwp8+J3rKyYQeswReL8MN999qnVruRiG+rXS6M1DZ7Kf3HZR6uKyZVc
4ksEhA0sihZnl/oD2CTa25cVhn8rCcM29or1nytDjNIJt8Y9YsVAKRJUZN32TB9h
bHrwAP/4DoIKpHQl8XZHGGRWVi4pqHWH1ibxE3ZLsspWQihMQrTOtZlMNEAwGgGK
iZ+gf0DO9vz6H2nWcjwRBnZULqSN/1KYv+juxo1ezwZIq72hRo+QTe5SXy3ftSrK
FvknTEVjLH3/DrH6s4UdSntFMNGhH18zoBSDBxhb03Y7fxcC21FCY2oXv9baS3wX
70xhOslbwzjQQbaXGzZoOUtLabpyRrnPQR/Ma+d+3r6dEaawlRaYfrmtvZEfsiUS
3v+s4JIVL0+MOcFwUS1wl/6N7pcIaYLrdmYnbBac4fh17XVHnbjlKAD9oNDwcHa/
23tizbgnoPpCV5vTcGYILo5niG5BoHj9zXOfpmOEbDpR4+Q6rN2yDutdng6594yF
esk0T/fXLiKu/bVQPxH64LpUlikIltmsuRvwP66gt10v3bHPTWryaUv1e5OmVrd+
4/Pk6Resxp3CmSreMxQM+d0yyCFxF8B4fv4gqQy7aLGqGXHZEEaEHGSJKBtc9grS
DVqO/C+4gf+zRLTIAlZfqkW6bKq+b7icPL9KZYsW2g2NTiOC/z58ZXfgNQnxkTsB
2qaqivlHWu8JW3+Rkn1wo+KRtXMXedqDz5apHclu/zDZ/QE8Z+UejzYOiEZmfZ28
bdC3H/2YtygWwPqpU6FjFg1be06/ilPHe86h0GHuFEzso6eyoFQVbK12epMIwjmG
J3GSnO2bJy0Qylf9jtmGljrjX5EwotPhYG47B2AXbEYuMinH8+cjcx4mfucc3jy0
nDdk13CPjOjRO7FCCKyrrTRfNckTpyspq/t/VxfQ0nbDXZgwZ68qtCNG8kNqEE4f
KUKShjqhjcWWxY9fy8QGDkhSEUJroP7Qmmi6FpLBoq12TAbgVdxEb09SXEp8EZbG
V/9YV8g6ciex97r+M+yhiiab5HE3R5UCwljWiKKQv5i9MdpMY5w5i+XBlj31gjkN
wWMznlFKG1KObZuVOO3TYPKJYsfJ0UqIQaOU0PyOHFQ0jYh2oNIyaG1S0HiBkjOr
U6hbsbmMbLK90aTSCBpGaXrn7ygDSrOm94+3lssmeIUFjbtO//nDZaaKxiH0udsd
nScssQWR//eYdEwDjiuHmkLgtr1jgXDQx1dvb2HvbWsQ5KYdU/pMyZMXaQo7yHHX
EJq22W0GBuvOOR99n/BlFgoy+oLT8NLvzg8yiaLApP2fJ0MTWicG1MSFTjUM66Yd
ODswL1z/bHtSOV4Vq+7nUi3oDBZdpiqgVIpmKqqpfhINtjfIxGLk4yZsf7swHFQs
/51/F4f9zwxfZBxidmpkzmkRkvpiUpi3L1VTaoP0Suhri9KaHDT5Ei87JwLJTv0I
1QGrnIfcmX/ieOK8nY8Igb8KUt63I1EwkqYwn4liknfoJGfdop9YmJUPAuU1BEkx
yEDDSx2XkTtGIBMJUMsbDMHutq6egWDVRWi1nZbmpkthxtkuh0HhfL+V5Do6ZktZ
pP2vRKWkfTPBoQM/vwqGu0dVdZhmIPUWd2EkA3XjDcMclUUKu/aordID0+Ek91IN
Pw8RtwHf18VrDAc0CKE1uhQcLZLtexGbgJM8HgPSU2XzBQddn5h61wtfXBtvBSvg
ptjR9uVjUWiNVawEDx8EafzWYZvi9FpC171LAknVTHtsRCjDnfEXMv1te+YBdDJa
fnVT+A55IwXAXVzi+yBxTTyDiPO4lvCmQji9oErD/IFSRvowS1WLJ2dcvaa7ggnG
KFZcIAG5bm7yg4Zfn78ZBzvv2qenNAOBRZ4ydvxCMIfq6UNwezk989tjOJjtzIOK
kDFS5srYIJOo3/eLKXmKMbbVf9KR1YcFwKaA1ZV7B00Cc8dGWeTCcZ5QMUUoRsZA
gKFfRVXo3OSzamtAWfImx+nuGDIniXAG5KjNjf/F+NpQ1dxgk2fvVovE9T6FrJIm
eeWxTsjWMrIG232joQX9UeeNq4mFMSqIDZDbxGnK96aGlerXX3zrmUNaU8zuXEiL
STEeSY0Dl+MSsXK1fl7USzgk4HLyb94J/W0lWPRgmB46XjFG0XHSMktq4hZ6G3Kp
6tMOMyGBSrEteyp+/D0uF6+lIF8QXjOuztNe0DNoPjKUBKKBiTe+qJtSkdXCWDaZ
O2VxxxAsqE594cEKS36iidRXqQT66Uc7hgg+g8H2gfjJD9UdUoFZ5wsr1lmd+AHn
0vv00syicp1qiiVjJl7hhzy2kNXF02ADRNlBL/7cGngU8nxU4iqlUPNnB8PLHOhV
aScd5laSplUM624g0/yjhi+ExSsUsr56IpUwUMiGNiN8wI0ZmhWiJofV7skwt07f
mUN3XBBW8niTPyNrBu+3IVC78JG0iy7KFNgTWyovg55kiFcq+UpvVjJ/JgMo3NMk
ocxFULG6RrrGEbGSsgWwlSCbDEJoJ3fG2NudZFW1GDOOhuxx5KzCp+YlQSIGcnAY
oPztMHqAk2ZOBz+GYRzZcAL39KvJxtNukRzTWzpRptPHKwFf9uxLaTtLoy8zTkKx
2RatXfEznBAPG7LTc4JwyXYOJ6P6l3nnTHoN/Evso/9j0KBHc0FxOs4wCyFbxa21
/fPzKwkS7yEW72IObgY6TlKBw5f0G7fyi/bDgr7hme+8rikDx2DeO/au2w7lebhQ
olIFvL5S149HZpfJsoi5L/zXGHyDZgFTqP6YH1fIv0CQf6N5Jdt3MpRWvuaiErlC
n9kTRkOxpcPnMFW1LY0Isr5dm745yY6BT8omZPiDkd0+GLQlwLdRnW8SGzuD+DLf
Ru7TuXiiLVK8NnSQFz93ifmWyua1Grnw7A6ot5RXa7zrKO+tjOdv5LRSFF884Vee
6H8MoaBWMhgiVxlQj+f12VahDrjjmUEL1Wbpw5RI4X9BPcposf+hAUGOOZfFe8+l
dYzBvPtXB3mzot3P+vVjFFFHhr95t8OW2JW0WRLCfnNKSqdSaAa08tiWPFWCGF++
R3VPV0CZKcGntzaf7H8TFd+dPVUGNeo/RnrjSWqZExfQu+GE5qnroIKSGQY6/FBW
8esCpvo4MpfEg+WAuA1D3HNzb5Z3rwVKLIyO+zHvw4FdAMSid+ihOqeb45MszVT/
ee1HBcmqvA29FUrLvPvodixibeHOcjXnZO08kFo7grHVvSTHH4TYsenfKPScXjdS
XM8lBx+1HoRbvtD1h35RdG1CD0S+xTMlVnGOf5shgjRipUsYQvwmhFlgdCvAVluB
ZSoc/SzkLn2iuHEaaNlnIqz7WsypHadrfeWxMEiR1yi/hd6/ifEYjIl0Begkduqr
UVFCAtceItGkkLQ0CLvBzTVem40j+HQ9SYo0ap7JcEhKLxdJ0Z6ZTY/viGUNOxxR
KCXtJXxTFJcXpkGHYDG0uNJnD1MK/yaEK+aW9EnZUHgfRTmU8zOI1WuRar6o8h/x
rEOzIOj146+t0uc9qjOkps1aMwCpsP+1Y5gN70EoRZu3r8SXya67Ie3McVMBlmor
knFL83NUAMShi6/3IGKFCcTdEdhxHLhL+6xMC6QW3/Hi2o6Ymn4LFgNzHIgNThXa
LOfFzUuR+RRQOaUd6+7+Iq3U/3Q7cKDys1JOc5VW1Kj/QWGSi4HhgvsYz9MjHlAJ
R9JoeXy4dROCsCMxeWG82yfcGX0LKslV3X3elj9yw0kVD3jI4V3Ovbb2yJX8Kw+w
TF5PtqqRLXva7nGVPcYAEHNnrykyytmfjONwsUW2IP+uTrH2OVMDu4+CwNPujKU2
XRtBA+Og4esPwomWLKRLHsmirX1Hw7hWiZ0rbIKfdEfp4eALE/KfHyn6s87TU/UH
c7g4Tg8607k1KawCrnD2RwNo2SNw9Me7L+NS7yaLb7D7A8bV2juVa1gX3hGnMwNT
KGe9kcYzrF2wvRqCsSczzA==
`pragma protect end_protected

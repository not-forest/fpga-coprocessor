// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
GvbMMLj1x6jikUXRqqt6itB+GNR0+ifsJGSF1f/U0hY4Z5umQtmv6TjJjYQHupKh
blBFkPLnlbUQbxijMNX5mBJ/eYTjo4cMZ/I5ONg1jKKenv0E8NLMwqehfmyEn94F
tmrLw/UIJSFP+9irgI5cfVr2fnRNrminojkXs2CLL6s=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 13632 )
`pragma protect data_block
0fFFDw/0/1xPTYSstLG0zRal/O85cW39B9hYqNSx55DVEZAm8dyrfv44bU7nN7a/
PPAH1RiZfHDdyMA/sNTEaItvOfVPTfQExt593CDvjMrCLZ5GsYrf0yKHvUKmhWT2
YzwcRqM3FYlC6uck0MjHC1F8HNILsvN+TnQOqEoGT6AwW6AIvvB241ps2HlkBBvY
t+5oQdCAd1Yn7VOrNngb18dBnN7psmAMqpISgyvInmYf5isqmzgZ95gwAx6HVcPA
iKTxjGrMtnuu2YaL8+5xstUUIrLvAa3Bt/3XEjbPOEbKe1nTGGaTx2ovGUXKd/La
BUYnrp9CSYVlogV07SNGAUCTpfXmUKLXM0zUt4HINEpixPWvn6gwhnJoknF5nn1y
ls9pLEaMrX54sOMdo8X3DkIXVs0VRcD2duW7tYdZ6+RxKGf54Ju116Kh896KUWbQ
/XghhdD3lOA9PSrNVA8t1Xd7ew239IBqzKfPipVfWBz3msl8BJreeEI+qvApLlH5
f2V+tjP7okQzJ1NMNCrKa/1LZBHIAAUT2BmofttoFQMzN/+JFoIk9Tv7sJ/qZPZE
WDy3HnChdNd0ZH7dSnZrnE0oT0HbgThnhITk18CB7yRMKgY1zj+4r7K3ZPbCcMK1
PuVuT0q70bwzed4cul0GMfbBJwRwJfdrtBBw55C2FT7GghFGriOpKLjIM5crvnTJ
/lclqkaF+WINy5Ump3cuE/WXYMHzKWscKQcrMvjJHl6D/VaBB0nSUB5OoJWFutm5
78yYleND6rSlvN5sCLrGM7WkRoZADPkMucrdnHLJ9PfRnPSmEqgQCNNQYVeIdJ6p
RpBEZCE7E90SXXxIqemEjUYoex6rmitY+kpPVaPGzRu2GuonHyBzYgIyT6b5lP5Q
T+Qvec0PjsWyFnHqL5tiAbhtUq5sMP24pwNVr9oG3DbFSXNrZP3gG7ER98MpQwIo
O+Sf+EgXeAkow1FgTHYF69XAyXBk+PLZA70IaWgne9Tgb1gv0Okade316h+vYpde
BX36lulG+gru/XqLSd8JaimKduZ7CJaTcKr8KUECbfkDOb58+BcOoSUP4yjsAkSl
K8cXSEenJCrgEytCO90Q29WPwP9jpEwSjP39DSE1FP8nd9KWzHKLKxX7b1EsEeO1
d++rNWEPnOuhpQ1b9qderjlBpo1ozJbIx8P4457jhWUxqJPLDbJFLKZRIFNjek8L
SqrFP8mg65rrURBaNL3qoEQJd7E+nU1kra4JZv6WJlSf5PyTUZQ4NRP00+UhFyLH
pepPML6EFyAezDx7gs8s1rXtGFdzJpchBdhm1OyKjFR/tlFgGO+j0elSmwbBHdwe
YCOGnFcG8hqasbj9IZ8JcHtwzqiT+clrsV/zoB3IQYSesQxHNQ1uUjpJi4qtjHWO
L2BSXCTx0bUsnUovRgsEGAglglN3sqLOdyahfuLqKiB26GY58E5Ov6lBYdz1enq1
69ds2BM2oAY13+7YEQd5SCITS+Wie73cOWxXhS9wJ9QgCZ4SyD0rN3QIFCav8R5L
TBtHW0nwGiTPnTyYLYEuBayc3RX20784ZeJylsBFrotMrkpR1srp5tnunMFIE4Ki
dnHFLNp/UfFSlVAgQhsz9iH4hUyS2s5g21zHjuOFUrYb8+NWqSOH0Oh1wYjaQyLt
BQtHrnvZCZasdJlEuLGYV77FQ7CDNs2rj7u2LVXNMSaE5SOvsc8VMo4UNMIvoMNZ
M2DX/+C2HxYowlMD09iytSt6YNAhyH4d1+yK/e9EUt3D9EOfXu406tDFvLbbaeXi
ZG4NgVOfoW/uWci136A5NN3vC9mDK8sNNC/u5LoDD/iT+V4bzTpmHO4zO/sEdXoQ
wOCQS6UQkOfUVdPMd4/YZ60BJrqQ38TB4X5HtKgjPdysOqyqpY6uSBBuqyE0eJCj
SVESJ+dApegIc3e2qDusX9EdT9ETHLEdj1W/+wldEfcJglNffe0lDWpR4Rodf5a4
aIWuFBqT3LwULJy0i6xaZE3CeEkOpfpm04rJXcwrMWE4E8kfxYIScUNg/ukrJpfB
MNVU7Eztk19Khn4E4kOXK29jQyMrZITywUoM3DYcGGBeMCemBaVhooZPbpOXrKPN
B8kUY6S6KRUF1CSOf3F9Hq4Mg5wAbtcMQjghgeEiguDFhPTd9keY0HvkSSpZO5U9
q5tCoCLoVViaHkxrhWSkqL8qqQm/Uw9ceok+JT023242mgYQDcYaK2b5mOpY/Axp
ijY99mQV9+Cf5niFLo8Wgv3oMC6I1A8ZcBLrEZ7xlLsdf8vofls/bva+aSnvxe7q
kqf8vvSuTv1za2+3K7w28cRK6xHkpHw62LbLTu8pD6WU5yZlKrkJmBdn3STDD9PE
C+OTHKyztXMLVsXeNvHqUjdvK7we7kEoz29Dmfb3lefq9jqdBnx9ksWJdcB1k+fi
RO2/1GKEssD6A5dIxCbpKDIOQNiTlvZzLrenZq5lud/3gGCdgxXQDrBgoUHNmfgY
7CFKDJWfO/iN4r5edCaVDNkaJ+uO3sSpPMFhFrGzwo/F83LQMoyM679O+XjTliLs
K8FrvGAzZBp3YcOJS5v+tHsh554Rwr/MVfwFj9w4PpMn+U7JFSI0ztMXgzlGcZhT
cwYHUUGwPZbziKG00BGsXQL+G2B3uN1ffaEmN1U/Y/bay5U832sGVSw4yPKc+4Sr
3MgTDswxw2uAKz5lKcVGbCVOdUERZAjbkTPB/oM24kGMHBXew3w6ySXCbn4C3D3W
kBYyGnBzmG92Jj/7G1aXly9qxqxPSmWx+AUL1MZrTu8hVwtOrW2JQXpUoT3o7ykM
DtQC4EgPZmcRhb9912hqtkkKrt8WRCcebsXaCoF1//KOEFROquZlRlyaO5+eYLbD
HibijwFDZnOHktUYUOrjy6k3vAscJJ3mUy3VA5oR+rtJLLWjDaLTvM0X3ASFjC6i
u/pmVW7Cxrn9Rrwcb+xefJEze/5EUPBJeCChoYp028DriNrlKT/q0pLrzWd5HMdH
FbLTmbgLWoc7L7A9g1WteKDh15bDB03Yjhx0mGaDM0nz/iGJ5L7+UTG3sZT8ZbSC
CYrH6Przz2FijaSBVzjJj8aqCFbqLdl6y/WGkiKJL7fuhZAu7RX+CCY0m6GqE+xd
c48HJY3h/ClfKXYbbjVu2HG910qyQCVlVgw8kXbDzIgec6B/ajYJsZ5G1phEABNL
K9YkAiZKY99Qax2OysvMNS+GCGwL7RmIdn0nvvw3GJMTZSy7z2qRDecBLxzK9hjk
X0nHViv2r0SHFLRFp6jbCCA/dZL1gMYrVkWGySliqfo4ZS7e/EoaxKOFF1kxC2+S
lcecqXpWrCWwVsEl0UCV+v8rCaGv/05G5CiuR/jkylYNGsGjJrPTrW1ls5BgKKhK
HBPm22k5Dk2RbkzXItIEXRFuIDtDN6CP6X98da7UPwZ2jtknjjSC7Qo2IQYKL7uw
wVWDCRL9a5HxKHFduatEbJVxymIsZCz5ha+/NYK6nb0ZCk4osM2SavAkmsFei5OK
BxDTRK7NOmd0YcuxTjjVrfejhcv0MNWm6a+sS1a3hjU9Sa4f13n95H6GKBeaE2Fc
N7HrMZevEJnY8zoNUqerARStlS/taA73A1E1d5k1fX4uHmCxDd4/o/FwekNu7Clr
RaGrBms9oJsa7uQIe3KrmA6cF8EMYpZJvM9323MVnJaicir87YMEIaEQuRDDlGAe
KjdxyR9zzO9KHuks0EeTXDpz5TN9XANRF62SgCMr08VdB27WQb+iWwrM1E2oK+na
RgGcNrsAAHOECQVc8daHwmajUCD5UiUY4K5F+FMqT06CEhxsMZTz6WeOe39jXb7w
EgQr/M+PClbD8FSwXJt9dwOxbnFBw/c7zB5TXM66KYgVthzE+gWAEPDa9WuxHhn8
JBa2+u75bZC63+vq+FpxEUdS7rYui10fLDePOUR3owFqOLGoaPXbs66Dy/T86xRH
sqiOEb4ULB6T4TUBUuIuo53AY/8MHBUuV800FRUxa5VLjaFjwNGcegv5SQZNHQVK
JyZ1wCBx6pU2cmUiULVzDMNxyRVYnE0qcXUB6Y1f/AK1YAcRy7EbRGiT1ooPXI2/
DZDPYQ27bQ1uYZ17j48/EWGMZLRU7b4S1MxswP4+WsG47V3pb5Tvh/TqEHh9L3L4
OusHfFA5waop6bVAv+ghtHNLqKT3EHgahkTOFjlB9zmtCnSvDGzCzCeULLlmEJeE
dmP4NufMi5KALCS80mXld4xApUrpboRLAh+WH4KXMSxDHhVWVn1UfJSFU6QItB7H
Uv9p+HdwbZgLGRKrIaGpygGo8dLo119EY4gZiwQ5eJD2e6NnxHBTSSAKnbW9wRh0
HaqMFzwRFLcM1yo003To+6JKTZLCtg32QjjZr7dhcYOAp8rRiWp0tApaHBXnI7MI
anXrhXSat2+SIP/MF4wNZwfHtZMskVaD2xNRHxdz7NX3ksHcMcHHYFL2QpH8HahP
71NFap8OG6UHoTweAFbB9Vt1lR1BqKA9nr7GgUvRMQcZyN9+21p8UMwrGu3sQdIH
dRJVhZmUVvoSc5qmH+R34E4flxlCnUiiCW2eARJcKT91BNNP3V9IWNpeWBWW8nS0
EtPX2aMlzMtVs1A+3ZsxDfi6JrOYNAD3Hy30EpragWMSUpAnk0ZgqrctiLPjGER0
hAYOr2MZkj3xJAfkoW6CafiAYqFUtPABvyz4oRQ+r7ryi7fz0gy8WTgprSOt+H5S
Q9iXMczLTOQp8iB+pss+0897qhAd0jYqgDXFYvXIXwAS60ahPZoAghSaJqh48UGR
FTzz2eZqeypTSA2iyMycQo88JPvX6FIAQt7IvsFWeSe0aOxN91Yh44le/2b47VKO
XgG0XpfGfJpmmTBv5OC+NpRjbbC2WRmSvM8ubTU2m2hsf/5BOPU7WggK2xRtCVMI
AZrrUYH1+bqxit0YNYRX45l4lZgOeuQGjlj/cv2Rrm6E6SXkHfW6I/QRaNY0MG82
uJhif3HXJjTT2qE5hYxIN6FwPRn9/ohDa2WSohiGzPSAAA0RnJPrTrDcUz/9KzDn
92lK1M4kqOQcqj+OjULjGsIK4LIxy49AK40fv1wwsEHoi33zIj3SBv6lg0F8pA/E
aSMcrHoNpckdEFWBcwhHscY2yosscF2pDv4sbvNyVIcmVMBmdZbYm4GYF55tdGBm
Plbl17jP/HuqWTiRwuIr8Wb838U5Btf+4Q3AU4mxFGQG+X6iL2gIwJ8lVDLtDWBB
Nmf0AxSlv12+M90jIIBWZkE2SGd27Ct3AWgELRDw7j2XOA59BNc8SH+pWooh0h22
gOCdJ1Kwzki+axeZWOarZ4YUbmkLPb+svvb3TsKGAe7JF77cvTtvxG0QftilMXkG
zngWKWNTXKzIQ1ATq+W0HTnq/RVnORElx34jijJOAKMQ1Ot4F78d90z5GhlRli5H
A5bHY1kFmaWBzHXN6DHpC1ZbISOF/lZXzGE7Q7CQOr/jj6HxjOA/r1Yu7kf4DsaD
XLP8b1+NcIVteOmCaFXg/PNkQdoatwxcUBxKn9moM6CFVwXa1OFU5Ofic7V+ghga
pWNDVF86WnZ1rhY1XXrRRrNMbdTs97w4cWIgVhIyMayUTQDXSJ7d98EoEViAKPxf
Ctt58pM1uHRUk+9XygqrcDdCByejDBmyN+dTEpwS6AJD5zmfdyZVlGLwGiN++awo
+Dxjt7whRXHv0g80vpyfnqKLWHa+5G/OdvcZcdA1Sd61KYD3f1Wd8qxrI4Tkb3+U
QZyS4jLeAchza8gCxzZNjRgDgLk3QKLsHXjN/YxLufRSu+ali8jF/xH27EaBn+vK
WQQMKU99wQtHuk3F5rXf/h8hJN1GCs1hsiU7Pgb3W8qKvkZG6S1J/ZbPXB3awX1U
cPCXZHiDAy1fV6ifJmjFG8XxYs8Zoe62nR4odvEJ+qD5wp0C51KtKBA1z+HRIV1Y
OqyE8iiRFUV0CQZF9JYNbcho6R/OmTY93jZmuYFGGeXT8LsRKOeQTvr1sc/ZimkU
a0J8ahxM+tssVkXyuhbSYb94ul03H8FVKA4KP9/fqDa/nuSVlvoRU+nIEqjhqEfF
RxojFycGn4kGx0+wljgDe/tTEMfJE1c7ijdbUNXsWckl/ypGfe0/yJtIIKFmcmTU
HrDVlRRoVs1LzOlVRCoyZI+tKpvBuz/Gt9wxoEhf+EjFxlrFHhDfEOxn1lDH53SH
bONkE/a5tgZahGIZZoEI2PyCNoGxoT7a2XiqsQF6blIr2YVDKggPvWg8fU+lXmKh
ms9HjWrDi/pPXWbZuMFrq/1LjCx+US262CdYr0tojChExbmSurgAcQ8+zSSyboty
D/vSl1hUGHGfeRZ5rYpuKsfO1ZnwmxpSQE1oaz6JienhfZV6xUSmDW/fpZhY9G9g
2EtHDQ6hJudLSrAi78IoloRnIRUnyPM9gm9j9u9a/cehEnXTSOzSVugao7NISEa/
k9fzelf43tte0wuR8jzDApLJfMSCycO3qIA9NYTZnN4e3/+d2dEcCPxWsYHAgg2k
/U9X9BdwVBi72YjtcrWbs1MIJNH5TkZmUPcVgqD4cD3sBp5Fzl26DBQoZNuFEw31
EaCM/fhyok7t7O+1kGai6zRETAbDYG/qJKFiqcldrVLw/Nv+85l8d7PLtINwFJH/
cIjti9JkyCZdCZSDN4BaMuAgBqtjhaQX4AkGP9+Ft/M8YLJ1xzxtPqT38pgAUlva
xWumpPe74M2d5IDBGhdqMhM7L34pMWRCw86VsLme0YDUlC7cfEnNjkxcOy+eTRY2
0rZoJQ9GXEzHZcz8DVNbS0eWMZRoTNYfnFboYBvh+DcggguMTTeBdXvPlrMMoAi4
8xjn46yAbIfocBa3B4lMADmja3Exh9dDlVoPIZ7C0N0TIAM85ZVpe971D+jfw6kD
epyNLZMfvoE323h5EzRJz++LrLZE8dW6ioEb1wcpVZc/dTszWvKGGQWH/fzZQUOK
F9Jnf1JaD8YF0p6k/DFm2x5bFVjxpAUZr1UZmCcR6x0ohc81ljGd4gjhbXw8ruhg
cko8/Kirv83Se7GvalsoksaFVxXyYOxaNALRUxNRljWcr0XPnk0E0LJ+PA8BRMwo
6lAf5PaBBLcGiLsOo/ep4BjHiy7uRk+TWyUm2WwCSSnhjed+J63ZzHdnkhjeD4Hq
ZtsP9lVf/9hJm+IZnxTTKrrxkDJGNd/XEnORURWhjfg2xFiMtix5dMBsFUHjnfT/
OR8DTdtflQYZMfuaiqAnsPZ9lEsdDs9/3mhBZ1oMXg96WN9K6nQiuW77Pa4AZOap
6VtIazho1+/WNZbwz0o2wyLpjIXT/byfsbj1O5ecok7nP1PLhcz4NJVd582P3Qi2
xmYaeEpPK7w9XdYKRpebXYQGgB9I0aPSD+VOzcxXg5F4efJcrSD8j/6bJjnlN7Bd
Jnr1TZjtePqncEUtkS+Nm8T65zOPI0H9VDsfB/yZCizaunysB2aPRJDE6tCwiRXD
3Q9b7MJibSjJ8EjGR1P4QtM9J+DQWqlTbOgoUj6O7W4j2dbum5ze3hT/R589u5JX
JcXUzmM9MiXatjPev72gmy/SFf9q32JbHGRpSBiHLcOOsBDK11NaNudLS/7WDxRc
uKxchrIamKUFDJjx8FOQUIDMARNIc3b7eyUSN8bnaJY8HJ3/5DWdSJ160U0aHNeE
+o3KtawnU5vpHNv6lpaKpykjqR8LKCWxH1A5sB23+/hvolBqbv08Dh9hWk+TLpzg
IYNZS57qGD2sVhlOBUAjMFY8PtDtDPPZ6HyJHd/UVeMB34ZX+H5fUCFrPhQTDA1o
OGtTgirMSey8rSc5rhiNOS02G8N8yI6LhY1Hqsqj/6ZxIlsZLBqlsEj7tl8Aa79i
f/0cVjkRlVImITCF8JSK3DcH4TlvsIvRTlGClNXh+3bvp66fQLIP1e3rDLvWClEv
qjAlwmuFAxIDtmhmRy7qWNBSzske6J5UUb9nYUZUjxnRU1kXPnUPr/UG+/qAo0Aj
GTk7QMsL3F6Nw+vkssxRIgFE6ldEYBww6Y1cyBOSVTQtVeHSoonF08uTV2xMnK4I
Tx1JbJQZ7ww4HlMPpWe3H5SRuP83MrlBLy9mfCbklZOZq/i3Z5IypZz4k1040+bA
ETSaXEuKzQQKX6+wtHuLykOeiAYeFLAlHtiAemxa7dZyH8xCd/xXWhiOJPmR/C+t
l9bZ6LR0/YRL5sfKSlaXM1WltczFdCt1dx3glScNqpsh6eMz9UXQuTHa2c6mPvGD
3vYYMIdN+STrpkmXAc/FI3b/Q7+zo7l2+Ed3afPN/umzJ5ofp4XYqUwl1RV27Jqc
TMG9Uyu7BL3bRAX7NhB9joAlxiN7xUTS4LfrLNDC/cPhNvak396W1pG59/WuP5BD
Digf8NPEP1nIUFTQUVdsjXIzCV1fKCV2jWpMQkTMOd/3FRFEdzm/MMUNCYdAu6P0
v04xHArPCwaF60FgMEqcYpHQEhiw7rzJc/Xc4SXm+bnrVs9V+cA76/rqboMWmLt5
XFsiCO8xcY1MLPqgfjc/mV+sydkdS0K1JpG6/SZOZv6kx+2Mfv1kAatMxfIBJS72
B31wPSE9CLNGLrSSXjGq5N23MkEbxcsqEdtgh32tCFhsriEDb6VVZqCULeCaiWK9
wQBiATSMAMEwpf3k2VcZPOwwu/wnWl/zPnQeb1cUJpykv4ZeG4Mgc2OgNabfiyLu
9/r9Y7qHqGv042i1sn9FU2AumUNvtDHY/z1Rxg1n42472l0hW9TgMlu4LL4eUy14
ceAaSHr2OJB1YLWYoQI0iWI333qfW3XPe5R2CTs0corwXkd9IEUPQQxgRkQo+Fi0
Nx68QiNtc8A1P0X0rHJE0DfeqJArdDepWQlpzxAUaMCxU0QA5iQqu0SbmZL4NEUR
Xn9pgRDIoeld3iYNVqdqh8lT/pf0r1MfD8h1NHc2XtQ0+j2bKCyuVt1AR8u7Cf58
wDLMe2L9BSLN4WzKKPVGziyzLReUXIOzKHRqQYl5LaJVlR6cirALJPF+RYilStmn
+4+1xedfYAm0oxKpbrUBMxKku/wIEVeNsXNAByQ4fn2lwWUjq+57djUImxbvo6/C
RCqlwK5ubpDRFEtZY2TZTsrwTuoADDdikMOXtbv6LeBRfS80ZDPuVPVF+Qrz7pJ5
IuJCX3ZUvO1piaf/sqwN8O4uQ4WnZ3OR+1Ett2kms8mxCfpRvVrdERUZFJ5ouBCg
cu+Ji5po/G2wVLnwc5SxVqUH8sNhyETkLlxCFz+ck/2/Er6H2dk9TpNgHHDTG/ZW
gmHIaLPnY/yDzy3S+vmFgSHdDsY0XxYXDHuADFYEzu4oLyjEP5f9fK5YPtLTFpXd
3KZNatv6c9BaUQGN/X1R0u8y844trXlVaJ3+GsJh3i840nhbg5VXgl7EEx/oyQnM
7NBhb+Cd6uuf/j9mMd9G8vJyZUeh6To19OYKI0FBtxUpHUXSe1UrPe6e+8qGi7TG
ikgqimoFe8pbC3UqMoiNOrlqVz0VmfwPV1SacF0ujt6Dq/i6IrwoJ2fWUFWMAhGt
ZZ6pSvGyrtsByebwLHX6L7iFuz4Jtrz65aqMdBPceTv5Sexf5HBPLpi76N/avMQv
lVvczMYNe1TcyvXketyKh9A+DWqEF+8Qz7WKekpghmSq2eXvsH8GopXiTgcZtNUu
Uo8vMqAsqhaKZLrn4G2lH+z9vN0zyye8udj6L5tdYaWGwoIV7+T6pQ3GykR9orbD
2bjR1WGwBYRGeYW2jzTdoV1+iUwqSlbmhSN5B/Ywiyrc2ST7/PnTaGMWl6XiKANG
UnDaw76hxNhJXDHDZffklxE2c7Yy0P6rJoljk8R6mHUzqpEsE9ofBM2mzyrfkFkC
ROLS42sQh385UhoGegAlFzHnxmdhBktJrAm4bLcXHjz08mH524zRF6gdPoePd2vJ
2vdVlvIuKKRCw5fYPN3TN41YMmmfJ76UtvcqiccdkHadAvkjYOHDR3JKaMczxaS5
bunwLZUANrGjo/+YSj6F5rB432OHrKd1/o6NMhQDu5dkgQSlDPjId+vP6dVCO961
fzHwSHooyRl3Eke1BcTI0LLYnlk3aceY5QEg4fKea2hGBcHkjp/sCKwVlXW669/X
XX9UqeNNvvJf+tSad3ENXqybUsQdZjolEcAG1xUct2aBqYVzp5ZS0uAS6Dr2nBPG
nlz3eeVt1NYS2E5e+oc1HdafJOdU/5xGaQKvX/tqERjEUQv3ohA1avr6AOa3NEU9
lx68pQrHFzvtf8/lQXsrW0bvGxttKqQzWzv3ZKKqcaHJlRPg3Pe/3TC4ySmONohm
9v+FQf4L6uBp9EQsG070E7MOsfynbBGyqyIIo+PDthMWMs5HnOs4fLl7vmOG6yEA
QNHMRNybhVIbOXevKKJhBXsS4OvO4BnBJ9UwvLCry8ccXrxvUCM2lYq/B3h8F+AY
B8oObKIjiG/Dj05aZBwP/G3gUjyPqW2qhXbORdWMLN8zW3xc3/I2+mReE6+pIgEW
1l1elg8STmlKFfF7rV8C7bSOGHczZuWLWbZDhAAaH1gCkYn6DeEAPT/UtCl1xrYo
1wNMTtmgtVXZ37Ky7kkFzCxrM6kHzkm4h0649g+Rg4dRic9O+RPsJ/6Rk8IVWSrg
2+8kTS+Rv2KoRagBeZlMHxHS1IBIbCNkcv0WYhn5ohpafcDJIAzp1Z8irvm0UaTR
/KQ2Edrvv0SP6sWU8fhGumqlWaOA66mjNdpXvqCIeJOhEDxzJSKefTeVknXSe/qB
rnKUNygma3tKhjWWakzPxqPTLtZIKL3dqYPYzr2Bv9Uu8i0I6KDlm20xHILTbcqN
7iziK6smd5eybXyOXfqHicQUmtAZLEhEnF1oJLrvnQND7dUAMf2SxCZCE6k02UO4
Qq9kPWd+gS2f1mCaq/V0zhGqucEtkyhs1IVdks92cpPbCh+7o2puD2wosFTih2/g
PWfEJyINUWYxAKlGkGt8D7doqvX8aC88zFmGSlvkXLC6vwrUbUO/PqO+rU4KJxBT
d04FvkNloYLbdHr/0i0ep+qaHrru1WEzAFDa8uiuh6+oJjLTeGw3B2NeNPvol4Li
B8rsv+H7m9THkSy8mM9tUb5KLf9LkwjJO538aWVQ6LiP7RHLHetIDSs64qotwBex
01u+AzNIMttzQywVzjt1I7723Bc0Bd6S1zGIn14AAdlOd2HETe1gOHzmoMKUJdg+
D8F8m2a0ybgsFgihSxJgAUP3DPVyw4n0DikQb3OyELciamxgn0N2BnYPe8/Aq0Z6
xRZDymWpr3nMJ6cWE7rLb/9zKSDSEKA5PAEcXkAjKFcMtUol77otFgxR8KEWMI1R
uxyZwmRzUaQQyOOePznBK1NVqT7n3mux+c0MFGyylJOqSOfTQUO/cGMVkeklB8Q6
FeG0tzOQ6MjLXy+Xa/meefyD2+ad2Oe/X7qBTwcq2ofvOqLlaapc4uLsdS9QttuM
V7yQd9cTeZBH7PLd6Hw/hQ9K1e0/UmKoCZ0mcyjYINb623kSQc4QsTyPkJMGLxwt
+WqTVDLDz9R+tF6BnL6vcfYHAlesi8jpwMwsxyG9RsWgseqqUsLdYJzSpToeG5Wb
ZzZAIzZOOcv/A+pOFkTq86CnO4c6A8bRoubusuqKR0KMZN4Aw5pkn2FqIE++v3l7
ixw0Pkf/qzQh/cuaJEkqa/wfMPFBPaxP8RHtLcEGNR9YX14moa5BRc0yNzIjGJ5v
kGcf+WJYl5yK0H/lsHOlc22azzeXztBHOBgtC0WDnoAqV8meKJ5rMC4UUHc9YbDE
oiHhZFqIxKdY892DlbjVTo2iUY4WiLtUrZHkOaNsorQB5P8kf+SlJlSvfIrfBdWw
xWHstmFzuuxJ2A88abcX5+RUiOdmTUAuf4KIal+QUDvks5nEXgXFyKj+QfT8nBn+
Boq5gtsylb1HCjXz7KHX2AM4Ud09jFLtVjzMKNcDdbQgqLoBRJ3kZ19fOaz23eU3
1yL9aYNszq7g8qRa1as9Ib1RxTHl7Myni6TDhPrm8WFYAMv4QoOCMAOwCjjh6bCG
v7QcAPNeWTopCK7+WGHSJ6p7n0DYioEKdMCY6zwdYtlN+xuJQunfidSknYSCIPn6
4fRhQk8Y6QSpYfMFh20s6dbSGHZQzjYI8IT6e8Li5JSnChCC0H3bvfL4fUNb21a0
XIyRx0J/izfrBWFoXhkdr3z8OJ1viZLHmJJzdSssED8DiGeE9cdad0AWMFV0vH9v
OInImnWSbRq6ewvffckk7/IpbYK38Lsbr544jJ62fdQZVxfMl0Jdc2jZJyRE4qvc
4VMkrRfuoo3TeGaT7dweGE5yp36+dN9RuKO0JvUzJYGi2GKRTVcp0O2+rw4sFRpW
doa8itouFkS26wX6CUXPmlhcKlZEIJyJQ/NazipByNjihdYGj+ZYD5rqFjsFDX5s
GHeHi8RxJM6wYLhoUm4Xh0GtlIi8NkQrVWToMzQpHS4WYjJtmUbGMCBBc+4tWhB1
PlsAihkXffEXZE6M8VYlh8q0CFnGLNwzQIs42xaD15OsmgET4euDy1hzrThhwpr6
AyGa1VMxX5CzPGhPu0WEToO+9mel6gqhXBuVh5Fst+1LhtDW/H7+wyaqPo4Dus9Y
k7p7Lb+PkEeBs6aeD5VAEU01twO7v1ThKe7qmyi7PVFkUudWqWRTdzYG19x1329S
5D2PvFD66QHMnFM695RT5CImwOOU0XMeXOZ252oDHfZVKY4VUMhYEMtOcD5mjLR3
B8Y/mSfFjzS1Q9Y6yySajzjkLWOYZPejA7iur+st4Kt+DxGaN9jA8N0eBLQ1hc2q
M0Yol7OwDjTEjIGdBD8fMceIlxcWXqLGiO0/QE98HqrIs0XJf7BPy7RPTTft10Z9
sucgpIHa1zVVpmNZTHZm5L9S3l4bR7IgdvfxtpLi2WWKz/m7O2ZkFBxMcejoeO3z
YoS8w6+OHhR3XCqb6+0NPlfp8unj1xfr9zCsDtYS0+ah9jfYLKxyyfy4CduYNKC+
4mIculIfPM5fKpCnhu+OpEgaAb6CIixvn84zYX/0ti9wjte+3Qg2x7fptBiTDvPS
XY1cqhZiX7Em4gcL3psCRHYDxrnxFD4fPWnUheDt7fCAVmn1MDxwpq7joA636j63
MDlGcKwqn4ZElAyZklRt/2Lg/aV27FUuROvYGF3P2kleBZMIal8i6AqVHFE+fvA6
XDytCWBDt1+CguQnuvWw6Sdpwg8/DTrdb1AQMNbPhEQBRCoe25OiCkvNmPlLuBNS
osoK01Tqai41RWLCDZAFuULPxFluHDNHT9qGh456zRrlmcAfOcXtCE3qC/eUzB3Q
R8dqFBsIE7RN4ILg88+UMMCReq0qv35GS4BbaO++9FVzOTzYuXw/ySrah5tb/CiS
KSm0gnG5/kk5i81l9FLrWi46Ep2xrBgx5zCp0xekM0/sRy/4ihbjSZOEfEZrP62x
bICQTkFt3Xwl938Xoz3yyytvSasKgDyUP1jAd46rDQWsOKml+7mHIYIXtqWxy5rE
0XUUI9liSDgEI6gUzGYR+b+tOGORJeho1SzJjrlJ1Ng/37+NkhUKujehCYJ63CdB
NnwdmIlM5Ycfw3lGlp/hoK18WhHp3DAOA9gqfvA1tkFbB+i8QrcrrmWdOb912205
cJwvO0dwe4q6p/7HQimiI9kZOf3CP0Wft2+8ay2sOgt7+ropo2IHbe2RD6oj8Kf7
6gJJiJ+GesvqE4hG+WSnMfcDofAVt2nVRQp6LxDBU8EJaS/hQLq6/UwD8Uisxg6m
2D0Ygz6g6x3QrKouoCFB5JC3P5gphqMhwlrcxHU6/GFFz9zfL/s/egttiHzzNy9q
T5Bsg6zVm5bC6l8rxFPWh0Ulw3JVwdVGtRLmACsmXHBxOqBwfTL4G9OgH37Ph4wr
g8sI4GNASmjbPyQb2B9+Lh9W5WgSvg7D/sQ5AXoGIvbRuKuwe9DKZhwcDQEZQGj1
Rqigg15pGOwP3t3xevzdNheu6+Jx2J1YiJAx6nsQJi+1sQp5jR29w1L7NICVTcgg
zKKugKne/MfvA72IT+etYK1FKReZC8SmaLnqLY8laRtYkb0PmiHQTH1GXdLq0Lye
DxMmnnRWik2UUf0g+v7ZBV7Td/AzxpksXOLimrHT9oySUOVZy1fA4mmEniEoYrFe
u2ZuG3S/sFa8Txg23ZQRWDqGXyCLqime1wk0CGU+6h9QwwU3bZiuW5OSWzbfl6y9
JiISTlMqaZJzF+Q57KcprTW1W6CwM/xK/VdqPVCM8c8vkjMX5T90Rmkkz++V+HJj
WIJMEPWCeP+n/EUjwyJ3kQtTQaXiShmDXYIGuc+/3sN6eHhm1wwR/4UeWpgOKosn
85QQvxG/WepvXZMa4COEPWLZ9zJfYNqYpmec2M8PHSSIppCir8sM+OgIi/YUjy2R
EXW/QxiOAhIBfKPzL1F1M8Vs23qAwmeWNAMTKqIQ1bUCrDd4JcKVd7hU5Au2/52K
yXLyeMbWpMbgoq3zlqr8YFE/CJ3LWbDeC9FqK230t1EuKI5iqQRfTFe9SpKV9IGo
7h6WNy77S+AQl7pexAI3NoSqoln8bLYV7cwa7k22Cy/5ApuK3rXa01enuT7kYEkh
Gup6nyJs4UDstqTyTH12z/v9cM///EpwWNLZTI0myEbrqurJSPls46dZ/p6BOXsz
pkUJmXMcNCH+3I2e+efj3BH0vAfyPsdIgaEHYLU2wMCJqjPD/WtjorVuLLqXPA3r
rYE2bZeOEwIWV49MCYPeb7Xkfkbkw8NalnUAU2DYxoiREVfqVEgCUDlEe7pOTH24
MTw9SnAjrgwMYUMOA/76+CFjMFdgvvhvifUi3OllwjEf+k6rRo5m1ueCayDG5BG4
cAFyAeZNqn/6OlzZCBvsfbtkIF7jtyJ1pJqkY+5s3QDWGJid8yzaB9dsFJ+FMAD5
f+hzXDOic3R1oUKl3IxEsMnI8U/MXuyzkLxXhT3D/qsBQn7ELJmvPWANNxwg8xgN
LsJFY8VRKlUHqYFIkA0T15mr5lRoKWIqy4jCQEUkYcfLYmRJ4RiDiXyPYTft6aVj
dtrc6/RKWyLSOp5IMHYVNX9no2ktmODGs/Tm7misVtrvv6d/gkGclEoVaVQcDE92
WSQEAmgbM/puQJbXbDO6oafGgltLWr73FaTrg8An3jMJC32jtmYtYgpxM/K0jxpA
XYSyv/KJVgfA1nU2G7ACi74iW45WgRLzFj7yNX9fGllX3LE81IYp4NXnR77FPROD
EwA612K69Nt/HG4tH44KZk8mxwT1X8y60XJTDUPdlM8mZjJOFLamRNVLdmq52tCI
pGsI5yxmZ7b1R85gkNbxTUGJvybUJec4u/syFYRrHxcL/DM0sxJ/GaXa9Fb9eZXb
nhwZUxzuoQMk4UwsAgtmH1YwMLbiXXfbh7yxr4UO2vJUahS8QX/GmVUvbHoYCJHb
l+LWtlQQb6Tt3UZbEoR3B/1ETYZ/CWxIZGbHhQg533hVGEHQ13Bd3UVQ+xMAAr51
aKrDUxwP7Y+TdljA3rbybYsiGGW5jscKXq+zQBtymMFVuymHAIr7tYL9njI8Qddw
1sPY4bjSzuZCXNvWi/ioehbD7CDllGGjBS1xa4Sr9UCpf8mHRcQ1FQmFCrgX+WiH
Jr0S2EcguSXyUz43tSba3THbXMx/E2AKGI/gobEIi/vxsjWSKNiD9/hcxjed8iC6
ssRTZwk0xKMfckvSBCYU5e2sIBaOv61Nr90WqJgTfdbWR6gI8EnDLDBX3Xbi+5v4
6/UpSG1eHLUyQgAncZcojNQZLuisl3gxv6cfaMFSd8890k40WDXEaVAr+odcE19f
0XhRWoa41F0SJ0lEG6ASWNRSsMTTAl0zMTODn9EYQmkpyK1RGJa5W6VR6J0aqsC7
+in4l4znsH956hUsCo3zjiFOpd8GY9hDI4xP4Mmwr1hv6qPgxniTp+0yCDDDfUZB
WmTc8VhYHZTCHRelyWSJw7S2Hia5SWa5MgfEWB4rV13kgYpqMe30lQXRb5ES0rBQ
fAaMBly53vDVM0b/CIEK3a/W9/LZZW8J5l0tLmTLYMLO/v4jCy9DE4IqIdonbmIT
d0ImZnxuzcrUexixAlH+L9+SgD6QlkwYXWlKzucnYkHNfzFrOFAHC5i+NgzMF7f7
+zEZAFQeOTlZSXY9Oh8m6N2ykhwxF1+VCD5mD6fEkLZIACA6aGV5BgtUAViRgGzb
hMhYKh1fPZJvtO0lRBkrsgKyvJ/VSbXDne19ViEzfLmjwbcSLTZDdgx5tLzQ1dRa
AjyJL4ewdvAail3IQsOhsXqf1xKTOE7THxdhW025M39Ps8a8i6oeWZI2ZTnw7E0A
YayivMyVNfMMqOwjY13JX7bTqmVi/hli/Wnm0ECSI8upL3W0tZZ1qFGPE9WWm40y
JyP0N0syFy/0NZlVtZTryDYlJy7X5dHW70FbxihC2q6iTjLMMwpdHZi+eq3ofbnU
+CTzBadIixYaxDbMygAqv12iqGpqUHE4lutChfy0BDf4E4ckh0uvoSVAXB9wKZOa
Quc4ApTEAYjRZZs4xu1eKT1FQZZt0uIOM/8yuIATWVeHG+29YCfnq7EuERb5/XZ0
50CxD5egiE5YXKWeDlnfMdqzTJ5q2+WMVdIZwvWFUXEbkRg6r6IJtNQLB1+oS6gU
Vq4h5+HbeNHhnlHPzODucrmMaVPHYZcW9sBzkjRGBYMEr+ttFndTIpKVktkWhwMs
5F06Nwjzg/ILOH2CeGiVeRZf6uP3sHyRBGWMU3QFSJR/XetQsZATiDL8e2X2886B
PEMmv9Rse4vyhy+Tiuz4EnMeujIYojyt3yBTZS34GwL5JDbpP9LnISn2kyWlFIll
fC2p6LmLaDvD5OR+Mh+86ZrYZG48Wdy+zaEU+fQYzlYGP+ppWPNgfUq8368hLSbt
pnbRLSvlRDry95PWwFp/nhnyaW1eZ6LE+jAyt6LDmcqTMAPMDWgcxb0UB4Iqg+93
NeHlYSB4Dbd/ckU4hWsoxAbPtAbHmCo+9KSkkVzmT7QeDVJ9qVPMLjFEJo4Wo1KL
503zGwvi3CRSCWAbo+bODOybt+sfTj555pC12WQpArwKDUPNDojT9VvfovD8GHgc
vFZtywgA/LsAnif+qb2266We8QAYLU0NbuExqR6XBbp20DoHkZHhbdPGEvNZ0/p0
HziK2LocfDYeQGKPbK9bs8pwsAXaTHTRxgiscsxoIHm7PWxNea+qoCCctAtPAs/i
8T4BnQSWG2ANJHzUUUqVzQOmzYKNz4/UyAHpH+SPRFszd+sHXyId1/0Lm8hDIJae
EoJ7/W1+FR91B1vGrg0PEycdCn3fkoF9lL5NDdJsfXEuG4XAdg95xeLqnbJRw01Q
dF+dCRCsb9o6vgJWoKJRM5tqEalDGGEM0Q4mS+N4wMw5tjQxWjVJZyHFg+KFfEv3
7GeOXYZWu0xGbEwfkhaWU9+XPE8ytYnYusUAmAPq2bqK1Dw9vChnE80vRzDoCfY+
a3g2CbTw5NpYlwa0HtUEODSsIZcuRyIto5wWJv788Ll9rYKfEnCQj+mtjWgqjqme
V5f+Oh2Xl6/QmqTG6OqsY6jvGELpN5BCQjCcmjb+V90MirLJrZJv0HXBLHpBjoa0
j6OPk8Bt7O2qyanQPxVI/dKcx9hup1bI/SFhf2Hql4SWJ8Hd5TP8i7SM4jy5AyiT
KVM0bF5J92RK4lMrPKma9P5m56dR/Zqlzl2xbxRY9u1Ips3crM2oIa1j+jSvbXIn
vrxiB5GcDDnu5VpuzYjLXeYaF3UcDyuuXLOeOct8dDSzHYbKKH8FSBGBx5Jjk+He
8oBWJhQCNq6LA6vIFS7yffnj+yHin8hZwHg81TLAOwPmoNt2llIDw8edeLkQXd3w
njosMwHnYL0pZ9H44A95yhfJdoOfAfmnC8J8ZKlBZvyrHKzfOkyg2pFjv2Czbkyq
0kw7Z9OEp8acJMZ120F71KK4M68HlY/LbAHZJTFSZZhFR0AiqY4ZC/eolHY+rBmL
LrvU3eN7PzUOqux56kKU3M+4kXG2MSHSsmXUsiJuYpWGXLQcbAUpUwqLvN3CM+gG
qsBq6AmUxwapTebCfK6OIYTJFlSB0xRPeNIn3nZW7T49v4f1IS5wPig9Y9ULKI75
bmFU6TIPHGvEm25Flamt19gaHCZV3WqKPWsaYwGRcLw5vtgMTTWlXg2sNMt0matU

`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
OwP2XHgXrTLzUT2eWa8LDH7DeKF4EEJLuyIUIYQVo3tp4KegHMcV/kcGEvdnu5eV
K6qdRMLCLma+CUJSTueRYi2Ia+rEy1O96fy/+VZQBkKeGzh1fpZImQADrN6C7vGN
cULdks9WdfHvcgWsf+QG2rzhfgUT+7LGkZUsXIOCZgQ=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 8736 )
`pragma protect data_block
0xbf2xqlh/LV9KcxFlZiw+UZtdUFlQkGQPz0qeQtVbuh23YX6Aik9JtTcZ8melNP
R7E9nV2EAfrY+fCWn0TlGu1+lI49mJnHP8laHzQYsJr/gD6PilhSlBoJNFjGV4CK
vmHp5kzNBNkcTfCbaemYROHm1syh+xvvxUQDGrbSEJfKxfKMghgSFfuIQe0E8s25
f81Wkwam+n9hdwN2IT6iMUrjaDRAHCEnh/VHID9QekDQA8jgoGKds/1sm+0Bw0oR
Cdpey8fn3NyT8IWdgycoIfcb1PtouVyaIEs1AiYNRcS7O+jamiW8TAD0LLfhDDU4
HbhsBwVFcH9ft4FfZ4oH66VA7R+dprMKRsfOgY4ZWxGJZbGNOtJInnTB2qMNK08P
hrNzd7Kz7unaKfh375tkhXGneQYVv2ftp4g7zVv09EPhmjKHz7YJEWa+pBaTUiRN
hAKdSaS8b3NwmC66jcmHNdRuTnbaLlfK1KYl/fBDIrGCqV6pnOTO1cnu8v4x1C/B
cjhPjhjkQOBjQDDmf8hJsrLuKleuaQUP7FbSUe4g12cQa16N+572tjfEqXNUdILf
/CKboGbH9e8pL2b01lTtAa3FzdK3Xp+ZLzCCeELsQKAPXV+fFnuwwgye37h+SE8t
srCuCrNdcIci214k5Hrwh/WBOC4kL3T+tI3PFUvUoo+rMieYIQGwihMWd9owBrRv
D9GWN8HydtaGFs2i4vOpiaGrbRojl3ip+mxBpkYBOhUU1+ZPe9jDNeNw9Wc4qElQ
v9dEk5/wXVyL0XZpuAnKAVsTQ/vRHs+hinLX1TcFdg/JOq8jiFYGKSVTiH/0QGMl
8iy1YRtElAyTmwed60R4FFVIy5xBYm+jA4rIs54qiXo5kaeyFummi5N+sCrM7+Jw
L+4Xb9G5bOSTuAyP/aLL9O0xrZjUS+jn3lfXWFlZN+v/0J4oIRWlUOgcxohVv8b0
TONXiXiicy9dzDcnyzmZ7eoDlNv24SYDmM3HgrPE8DdEiy/PFkiNXaYDDXmUn2/z
zfCiq6PUJvmKgExx4mI5L8UP1+34itt/AJFs0ym6plQCu2reO42bZIBJcGzrBZSB
cPNdu0iXTE0VRD7dTCXj9iAvhxqiVe9q6DYw5ox4nkWbXosvhYQi/4ZENL8YFWyD
3dTF8ZyRmvdIV3iSGWGslVGApv3QE+OYvKuUXWtaW6FZoc0A1SXxmi/dDTileV2z
b0SyvF2nIeUejv8cRLZK6cSAHUQrAeOBo/9N2BA9AtYIp2vqRW9yKg7O5tD6YnWi
s95adfRkCvXmIksoPF6/nTBueWxTyGYrWRVOi5KD6YiiovyP+6L98OPiUHcDMcXD
gzYmD+BSt5EHqYSlAOCwzraoFPtXtbKwd2CFp6CnFKchm9UU82H+x7nDZDBqwbEs
WT21+WAh6qCp9WgnpDVbCVzDndoujITy7sLwvq+9574J/CZTmlceJ+8gVJ6F+mfM
Uusylzn2MEAo+73cXIV9jQ+/8zhSEILqsM96jfZATnU8mYds0zszv2bPUJXk+4jL
iX0Hzoocq68eA/Fw9876q8gIKTv3MVaTFPX8AyH+K2Si9FaA2rfQkOB37FRmxWG2
O+KOOWx2iwzUNeV73AG+rWXMQiMa3C4JDtf0V8T8OFDwSJhFhgITCKEbJEmmbQ0q
jyggT7bZxdA6dst/egwboitBXLhkqIwo4B6lO19VMG4v1TjoW01uv62tywWIgQ6/
oyJVzVrwv2hraO+03ao7SiJGp3ZS0YZ1QXnu4BcXpiI72P0yT0kIF8Pg2p9iz5IQ
rN31hgM/c73yfCm1Sa7cV62Fic9V8LZJLAhMmP111cc8IOXKYusqmDLAnNPxnw88
8phi6lefywONeMc77uuFwdPbACVOkXH1j3eVOWCd7QJLCa8I/VoFlbUULQbeucwW
VhEoN/ybkT6bZ9O3xwyH3gJFzZ8SMS3id7lvUb7DYi7Hqpvw8sMtesyTfIn0wasp
7i1Yx3EczwC4YdMELdmNv+mcbpmg4/TUXB7gqRNbXA8s16gxOaF8ineFRkwP0NDm
FuoFquuvZP+uWFbXXjGNmc2o1ZHqKdePMl4h2+B0ydAiXd5BcnrIBU3dNfgq1Anj
o5KvVgQvknMqMwoQv+VwuyUxzVvZfXPjPFnmx6+fdkZPGZkSH1Z9xGBxTguPJBGb
5nKd6JUiZoHhHF1qyRU+mfyN19Df3WJitjA7fZK44ZRvc8FDv6Q6wa2cJURiMck/
WGXpooYKmkvFWHQR7mga/oxg5lF6tAxNQ9bFs60T/b7aCVarTnzVCdz9jbfC5Ozm
O1tvfNlj3qucFjy3KTKf9qYm1oe7EgJPtji9O3NUhwwt6xQyCEfVUFrWujEeRTFB
6M9vNWsNk58o6jvtr8rZKn5gSf32aN5GOfdgrAWTg3nCFpc8bxWvS9e+wVIBjBxu
mt/ejpsCGxRWy4TadtidBWwj8DCu1W5ulL0seQp0tzvCsIGXRxPeaCzqWW2Pu872
q/odsRLMx6mDEn8XoHS2XEGcMeyoyEr+vxoxWVuZwOupnWiek4kThw9UsGgQsxpa
uZVIzsagzlG4BiBO3gHxZGhaTaktWqR1WQC6qT7yAw2FP19CImsVMj9XkLUUjqYP
i6EDVs4SmvvQgJAu97OIOyGocjhpWMcUN/xZXAkquTm9cII8e0EujDYkU4jAoxgs
lYF8zKJ76eBmG6ValsT7eUP+YQz8p377yYyIQlNCXJR0XY9qG3mPX9uiJyvKgoJl
GoYGF0BZAEQ/AGgcQBy7Jltz46e7bHYYZ6THBjgGhfPpt7WwEJg5IEQf/eWA2YKs
bErYE5cr7Q+rjqY4Gi+H1Hf+ZpLXk0A1WUQrvEWWiWms+F5RNLPBiZ7/BpKqwOBV
p0dBKjlxyKHblYfdtUw4KfBlR1CZQceV9Z/j35QMN9eDyfWt872n0u9Vb13TgD6w
ryqBXetc6uvX8v3WSoB5sQmcc1duuODq7c4UJrXKaL0mo2u0SG/FoOLMspjrk12s
G+k96LU8Ge7ZgkRuHyQaHRhPdcUWtE+LSECofhUY3SNsGZmHQoebzWbIxupRpJqM
bbbJmFL/XWe9pX/i38R1cKGXSRjDXvE95VueDqx3gxnaMGFZbMIkcNQK4GsXv/47
8bAWh7p7DGOv69Wp15piyKTkJShvRuyBdaKuykcDsp4UH1B4p0DSxNkaNGnnXt0J
Vc37jamo6pqX8LJh1YlgyYe260M0z1FDhPvyioPKo8Yp8CXN9Id13u0EAHuFWz2C
qFpjkgXX9X3qcyFg5lYlczjvse2/umW6ZSPS5dUlesfeO5bjgw15Gf2gTr1L9ag+
w3D2HbpYYxDdsV3chSsU1h8hJJKpnGcrD/IlsqUMHRTqy8QkZgiP7wtxfj38HH4U
JKVSdWr23kGNzhF3rFqwWtqRR2kZ7Mgpom/MJgud19FAABx48tBqPI9VhTAQqtrU
747MVGd/0QYUgXDsmq8vMKCQl7HPqZ5UiWQF/5xnILjOQ1rhxHTT1ozLaRHsAqQw
SqEAiatJAO7KYG4SykYgeagIBMdiuvwKBJwZGWq4sme6gW4gcsOFI+1/og28GAwr
03YluokpVaEwMeMtWUoPP+WeS+GZ3MnvADJeqC/8g2KyZUaQpE1NjvBe5NOOmUi0
0fbznA6xNd7X8uJg9bH/pYPofLTB8jHnG06Lkd41Oz01ibkLLNkTHsWCvVY/cXzG
XSwlxJw2xeSf55SIMXh7iFlTXEkvxmfXyQdmLJ1VF9n+edwSyVkIgD2TuhYiIg1y
n2Sj6djz5zsXcPBqK3fGdU1rCyaPB4v/FpGYgHTRqBxwsluei13DebeLy0J+Yu+T
R1S9+SpqVNUgLcqfOTqN/7p7dNU3UKmLyeHXgdVaPMgo/S8j9qQOlBUh99dylIFO
REZ1+mb4VMLJIFf/H1fyg+geEqXiLW+gjcTCivgcdvjVJcnw7VtccN5vBqXguyHS
cLHdMpQh7dQ2Z3SKDC03tZBFPPIfQA3c3sEDGrXw96IKMaF2CBjgHAUmnr9amIel
xCVqYJkrmfZdaTo+nK9MxHrnPfz+iq4PuJUsxZmsLs5I3Mgr8ChXCCIwJoZZvBmm
gg6aogbl7sTEd/dk6qVOMbVKCfQ6gR4BS9TDc8HPxgKJu/YiqaCFba5UPrUaaWNE
VEVUL0VYN2S0QWg+9pjuW9Xc0y97p1piOzqc+Hflr6qbZytfPN1BocSs+tBIj1MP
6sIIrIyyrEDMReUTPzdU1WsKZW7cclWlZPSjpb/gn0qbao6dFuFt1Mdi0UkjABfk
5rtIYbq0clRqP3Pmaaf3jM8aSiOCgCOYS5Kqw5EpizuV9JtdUBa1v5Bi9jPde/dT
RPWEiIriQs6KK4MVGvBVYDFq9CY7UL0AcOU1Ri4QI0sbWWup0In/katAVfYFTfII
7JAQjH1CRNCOsnikIe/sTnnaKjKKKYLhK2U+v9aLYOFMmIVaSljfc5a7J9oX9fE0
mWCSqLMHTkHytmP/cNGJZ4geAwP/Z1AFdmOx4RHSmOJUqRtN//8Xjj40PBl1580v
YdcGYuMPe3f3wjZDk86xoTxyiU5CgxaJucTf6F4GUvdjVSFN6mRHlhtvt0HxHVQG
ltajo9pvhRnCVktdUuBNs+ULx//6kaMSJcZCHDHtpCw0O1Lz72FSaDCLMyccAgT2
h04gmhfaKzNxXfgKuta34H+oBVg9KQkc2AxuDWCWkflTkQcdMc3i9zTc9AofkFu8
fRK6FKiJ7t187OI/eNd8mNkrQID48HwyzGTVskl0qBNOU0fbnj7hb7Rj73shi/6d
IUpMISX7IiKfQ6od1QPE5CPA8ibJrA6gwezGv94FZAsXV56cVTjCs06tKrW2AIeG
FS4dsLkYdlkm0zJNN/2ky6OCrYIBE1B/0SasGdiARMvr/ihtRKWhJP5N3dW4ZKkh
zhVli1s8TYfLw/H6MYPd825laoff4ufONqUcyO+FPNJWVPA4DtdbQdiWyew+vcYw
3Cu0mdRv50OtHB+QcNteSdW7BDvB7Rie4ynij/nR+9crEQIUf0tK46nHPb775vIV
uNLw06nBLXISVer1nY2rKHVyFvIBYh9zXKplY5LuLT+h3OgqpaT1RRh0QRMRXGSy
jbhsh5Puqp6cHfLR1nMibmSKr5dWu+z/xYdvSxjNMQFiNpknK74ar3oYU2EVQj8y
aT3mBx+fUlgC9mEfHD81r3MVzxAGRVknixDTJk5a/zUC7ZAgMaOq07BtKWSOHKaq
bjzzyzzkwIJCqQ6I8q92Pea1jVB17NVsKVMRb8SEtqCcTovj/EPizi5p46Gb/1Mj
hJEmLdz8eYNybnJtdv3AkTjmXxSXDCykCM4OvOBwRRskrOTbutuIEDss+NRUCAcM
9zr7L4f32ujay3MXnOe4Dx4z5jmvwsxpCS1p73zU/4wwUI0tkySgXkiedyTpLSmF
cLY/dreRfmhi620jhxOPoPHXiay/ISsn5lLpJr10ILYdjp3mrXHWgb9zWAWPVrEc
Y22icsF6hLw72Ai9sdZq6S5B1RYah671mrvbLiYYxAfSCHI6Cga/PRSmWSLcgWHP
s9EmzNnqlOzQWuOvgAyBVGOU6HPnqRNIZZdqX7LArRGv/K4SAPeRLZLEPH3pDIXn
0Ezc0fxEuO9j8Hh4N1TeVGN9Fm/Hsf5+KptiB9FPGmoJX0uaThUEUvHibkI7A0Av
/w+HnfMvfqCpBUMvA8H1qJ+7ijUqf/9Zxa+r4Z9fM93V6H7V04X5UUXr2HWNAoWm
JUz8g65tIDeMCerGEaYdGcsBdz9bU9Gtfo+CbhJdBEVgexkNaUqPS/t4XXRGRah3
Wdh3AHA2JCXgd5SfN+etOSIAA7WAKwfXp/oCehzpi/bTHTu26cXlCBktAASz3tIX
09shsc771rUwoe4zu9N1+NeA215IyEPOPj7Q2noF1jU1Url8u4z+aeVrBjZ5oymt
ijj4RhukhJ3jDmNQ2QlVisLjfVUWzjv9ql8sF+LooQY9DYybwbGGM4CsWOIP3Oqc
yflY46VVbXhosAAaQNueXRYxe/gAPcVFif+EhL3x8rGEZVDYg/29OFI3EXEglZwd
2+RvjEcZGYXZgZfv8Fp8qWvoUJcHdNd4cncdEtGYcH4UgWD2fFqJsOzl+p9rCPlH
DLdFP7fvtomw+YDOc+w2uo8SA99hE/A2EuVWF1gceH0v4pQfZNBk/hfHIjP0ZjSC
T5jyiGj6/U87u8dlaBdBHE1wIk+61xJG/6aKL7DRZthZVAiOCKrSqFY0/prRuyco
RnbiEjDPFvyJ/Fb3GjMDqgN9z8THWYq4ki/jMnABqytjBRpnxBFEcZpPrb/g0iVa
+Egz+5BvSxetsGkd6F20ZT4f41eNapirKP2BFgdI+ZUGqM40Ti2whGZBCelqRZ+/
EtMxO0DUH2jHMb3Qj8BjS8ksShLDdo4kga27I7LyQK+j9noeshKQpJ971ees98tJ
Vn2KmE8iWsxIVPkzCtrFUc+5MYwEd2za8FrZhnlnvR5PXPoUHp9/oIDPOFmiduS8
TpUFBx3MsbGTfag5Ur/z68vJwDazAgUYhbF7IKkPFRaj1cOHMGIoYGw6kNcDTcZw
FJka84mdvmFSdYylO7uErE1Km8D+3yDrIFqm21pLKwaKohFp+JwedNSUrb5qYjC+
KW6VG2kuU6IzsaKLGLCM5DeY/RNsd4AZ/zRa94TsnjszGutn0tnnFn7jLeC/bY7F
AZnhPS3/ejmtZgzqb9LtQHZaIAO7EfEKDkwDz4Q9VJk1qaW1Wnv09GaQBlO3t2Yt
qPo2/g0xwfjJkoeoGlAGQubHp2PcD5ttZKp+YI54bStIGFz4ejHChs1VC14CZFeZ
oZOSwQjpfmmnuRE7Su7/Eo5u1ntk+PuDoFahyXzKqbXF5roNit2ikIHckLsO5uxu
nWrXGj5glq3oUsqVO30j3SzPom8YRLYDA3apa5wxx0obyLbmge/cSDDCVed4Su8d
hc8s+HoOhsrCwH5IqGRj1N2R1r5kXVuZYlzOQFOLxIv7t2WCwGtjmdGH0rKn2sPt
pb2uhMe7jyleMHW+itOO6uAtojwFkYlVJYbM7mvic06/mB7IcB71LfjgeomXoxsj
4j2fHRKIjhrTaX1yV6wfJFBkBwVQLBKD23IzgftaqUymN2fQyyMrBYYutVTSpD8i
FayK1Ly3vm/+GluwfjjOb+myATmuY7ZVjd7nKeoDkO2X+fckkBx8DLXLBgKO9HVw
TZwU2CCwJatwgYOumfZ0CCt30J8ffWKNsmQK26MGSev1XW1nMGvrM9DYW9NbROcJ
J5xjtB3yicL63vnbIYmyzpWmVUccAmFoRZFgfkJjgEm9wkK2bk0bJtSNxqnjljPz
CFhC39gmBR67UhKlF72+7YPuXSw+BT8PvYVH1B8Y8O9VOMwENWDCPOwGbPqVpYKl
RtWX4LuZ3Sufualu8bLZmBPflyL0GCf2vRJtGD2h3nE/YLj6v9ey8y5FXzpzX5Hp
nxRNS7fBtjTMSXpoionuIAIaPKGgb6NtVqehe85JBneOL6lydRqH9MppKrSrb777
E9pPxs5KmAiK2cImRkpLbYSJUnaOoIvjvrsa0UcqXkTMnmi/9LpQXkYU2TMs2M3s
kSImRyXr5eIIe25O8CjvfZN2vXCF5kibOflIfLs+FMmzglzQGZzSeXsWu7KNfP2z
9SEWb+zBGiMua8QEPokCj79ooGtTyZH7dG6xTToC3StpRZfJbaaW7TQELryBuJrx
g8vBTxC4t85ZHQvuXRDxZqo//vSVXZ2h4V919iUwLcXqnS+D8kC8/+rMJZWyC7wD
FdVaucTRnCeWSNFaaeulg3bGY1eC4o0Zh7eZnYA/ZcnC27/c9O0EdOFuE5ZiOgb9
8ONpAR5/g1xfFlnoqIZMnX1cetv0sVrmN3X0sMh57knUmH6ONNjkSZDttq3sipzl
b5LZ8PbXuJAD0+Z/flYwkudV8mD8yamgiQ4dZJl0H3hpC3CsumftY2pVl00OraMI
D+s49bEWleQAlYDBFgpNGTVBxBVUtMwFUFY6wy2xbLm98c/aqMbHRJlIiyRlQdha
qSAI73438R+3T61Z4Bmt6XxEPi8jj3xDEx5P6gxT3WxcebAu4I6GVK5UTbM2s/Hx
0HOd13EoYaF7pJuGBqPXtWVaG3z7D4M2I0EDHx2rxGM66uuN8gaf8IyE3IyGr5u2
AmawK1c9oL/4Rou5GOpy7//46bgILBUdOzED04R+wPvSkq4roh8PSByGrG5Go+vA
rkvc6mcoS9zJRJy8CUAR+a7P+U4xdAIN6lWiFrBdb+jiv+j5bnzE7JwwKroSC/wD
EDo3cyyM8tgaEDGClxxtg41tf0aQoQWj98e0phXpG0NMeVVmpgmFX7XQdwY2m1GG
Mk43oC4RijANSCV+gLrL/LC3vd7rV+QqUuwfS9NI8jnSUQXld07sJfizB0huoQYq
momwxub70D3fiW0crgSOVqhHY7TvLh8yY0CSNxDaBPzWNmiyHh3la/oc+cLxGaMx
r5paLCiaI9nrBIlZmfhh/zgvwbM3k0tbj0I2uNLe8yC9b/nPro1WN8jWzFoW2LQU
qx4pXf99blo9angLsZaGR3APdjsXzzV3DIb645h433V5pJ9jVpX8fMejJnq1Vm/l
cLJfSVo1dnXBatNwUYO3iOlFXunng9nnWO+Y97krEvjhP7Gy8j9DevECFPmD/1Fs
d3Fe4NEw7662hv1X14T1d12bOdVhdCgCyVCVb/8x8dLMBSLazW7ZhTjXBcv1IW6A
OijDvIO5MDnUfG6ia3/C8MqNNXz4Fy4T1Hj/CgzdzkkykbbrQx+MOONxF42M9Dlq
5FR/d9NqqumkfHZMlC4iD/O50RoWo0vOzE5JMIueiMvZ5hdhqlWLJRpRK5EYi0mW
vQSp/rImq50LZ8FV27yTE7PSsNGHh3CeAgQ1w0A+morCS7Fnqdx5IfH9Be4BrHnd
AfHjAfuh+7OqUNU8pBJ7IqeVJ1q8zfNNlB4DxkuZd28IDWXM+dRAGMcQUUZ4tNeh
D1JBbjHPgwxniP9BvYUUSdXMAhTwIyR1BJWpBE9M3yR60IkU8EUE9RllHLEfIbXV
jhayG7asqzdtsOFgCa4xBb4hfzVRk/anYLTMM0JNyX9ZoC1fJ6Y1VWNJcbmx5hCJ
UGlaqJHMqoeg5BKY+VrnE8TBGgT5yXbhP/CTJ1J9SOcV6rU9Q0v79mQ/230VTHk9
6CTRCQrdbXmFcfrLQkjrPg4sy17PeotDueGoZxxlP32n3QrkTqo5/tLlo9lqvFGD
8azwD0uywrPBr5LfE0z8X2x4QGq4PmkuGKI8HjKPcwldOQ1bg0rTy67EWzTzvRbM
Cx+2poqOS2vpUJsmKHHLyojsyxOu771DExbDicQ/Zi2rBvsyIlMlFxD36Ibsyytv
2niJDDKEZy47dxYrn6QP8rcuiBEZVs1XCh/xPvfdj2/Wl47pJPf70bz9PCGJZvnR
lbwwe/W6BGL9RuVVGK6ynIg+eoB/ygtaGXKdjj1HXzaW9A0AFDljnZEl7WRnmZXq
exyH2KSSNs7AX0MEQrV8+GOM8CCuT8DaeslmIDiEvQ/ZoaiMFYxvmyhrzrP0T26A
K1Z9Xz451iuUH1EbDrThD5lYM7cw0nemZbZSESyPFrBLrl+REDHbH+cKAXlrvS8u
TuqFUBjvgXKm9uIOSuB35kLiZAVR0qIypK7X4yX3DKPTYpD5znPGdbRAs/+Kt72x
/JCM8eO6F6PB0V5xvRk4iBbgOdpwgg2l1e4LCPfHgFeKrNpp/rCQfhzyUyJE8HRA
0VWCGDFKTvnMHP2oSo5gjB8rCGn5R+PexKGZM7S3F36k8EhSZ4DacpxZEVwF5+ph
u2kCLYrn3s+r7bJVe1SJpb13d+d/UDH1aHL7Nk0ctGvDA3hx39xbYTW4x+aQ/Cqp
LJ3hIpq7BN899oorefEg8IiQiyrQhh+RXNe8mPByj+gz7PjMELIaMZtluJHBgpsR
dbGVQLVZYmf672CZjAhqOOADYr/skKC2/54z9z+lO/htfNeDbZVOGJZK9wydC7YT
LMhabSbfsoruliBlddqNjTGcWwfl0aGe+OLcddOCIeLyzZED/Ces8S80EfdaFZj1
qgLBK2hHu+fh08C6MFP7ONVHjBsYjrp9AdpCBI2IwAvoIlI9/HF/8dfWtUop8B7G
zeaN6Ukq6p0px8PWpIZ0/yKfCfUy8Roj9NRrfCAAudWIhlW8IYcZQuDqUAAIyuNC
VAuRZTTRCsMfnH4Pc/KyoTgjsUPd8AcWO6mBxT2veWZyzEJZozRcvyMBtX6e+kjy
Mr0ECCZ2OvLR4LPFQn5r+G5wlLgKEWebwPjMlypXEUDzgBy7qsABJ1iI23dpMkwk
dRX4gEMBItEAwHpeDe91VQln0xKXMftet6Zpwa6eTkJ2thF3BNrPhYyUaSn5sjWz
kWgGXR9A8zQSn/lHClTp4IkYgH33x2gYTZHhx0aSF+m6oHTcjn8ll7YdZPnBQAan
OZ6ApQi0D/hTIQO54Cy3DyIWNxYgFZ7VBC45r4rvlnaBOzMnLIncEclw9Rq1OmWR
6cCnefxDFkc8BYPYq/yo8GPgwM2uxlgKWaRzKjxks0yX3S+uHgMg+kMzZn0Gfl2U
AkD4mIG1CtkT9PyWBRVwSnpWd5cJ6ZX0ZGVAHAs742JG39+qQvRlDukNXC3gJwI2
F5hEAlFhiMd+HGRvv19BsVIKDCYI6twJCd9vIsC5AOf7w4gef8CakOwehLQaJO34
RFY284+/dOwBu0GvwsD8E1YVgNieUJcr5FhBoRZvfbcHQElEJZ0slqO5YlBb8B8s
exVbII+HNQtEKf74ujc+S4IXHqVhbNGbtjBlBESa36NKL0BSkSJJTOGusGM5Y1O2
YskdpMPRJxLzViTRuBKrPIYtqs945JMt+wT2OHmYv8MW3lbLpcWoVq529jJ18jKT
6ooaQPUa4eu2BM9PUjMhNcJYMmNnKxu6KlEHvnPGBcn55BtyL9cZr3uZ+ux+yuMo
XOfSb0NgiygcYf0ev7yMSQ20TQCsgHHg3oElFgSXn6/gNzghLAxyfOgdH5YFnLCF
VBHMi9ZU7haVG6GMjXIThDNLoL3EFNyLpr0yudpYTbYcmajwF2oA9DL59sMZvBpY
iLRSF4RJj5P1kBSsbLBcusZuakWWu1fV/HZO73YbIRmHQ7KBN7JQoqy+I/Xd1NaX
wYEtKLaWFRLLcXixbqSeF8BC8msyslrKHWKXqOEtGpQFB5F4h485iBjpDCE5f5Ln
AyblCH080L5RpLwWA/hL7EJ/UbtRutDr6Z4HhzvPna4O8vulf+SABxKI166DLZoG
krHm+Qs5HI6XyQGfxNB+gfXpt7zf3Uuo6DvkLcRd4DgLT2QB1WMe0+PY7XEooBEj
CJdx7p4LWljUx3pnHf8mXo0mdKIX25KGODrjnZegrDcfKSHng/twWyzOaBMEHuGc
E2Br11xI5zLyZYvmNtygxjxwSUTf5AEwlb965HSUZsYN/Mk6mTu6t7MQnXcozMCv
nFSiy4pBIpAIXYnwR7mSTqUV76+bH9pLyLJoXDJQprNsDxtAGBaNy+yegYotV+2M
c0t1TCwc5Eu2BBPq/DcqAzcHgUQHGMzReU1Nd2o/7QjOYNNZrGBkDTxkdBnnLtZJ

`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
EDZT7JL98PZtE8JVOrhpTav2abExKi06qi8o8EEfzSaGR59AbRqXRRFS+/eOQuB8fj12Bl3F9kOk
wZETWyHi7mB3t91zkUYRoWurL5UvV327yWzuoBXBLDheWQnmEjtV8SGCq93q/hnyEYPKAViCqh3B
91ZQ9s8sV2cIq/rIFTfpC4Tch0tkuMzZC3n95bjknNTcTRgv73GC4m9+UH5ulM/axaBVfmR0kUQR
RKkJNQAdlreRDSL2cHvr1LN0utF/l6Zw4qeJt6Tv+t0DY9lnEmEdzWuI9ZZeSUerlqCkTRnjx5eW
BydwCDfJIIcnLZGqgbcCQdKotpNp6q1q4gY8Xg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 13632)
lQ3Mn5phVTIiB+5LbdJbmfQBf5m1AKP1PuyqIB+IJCOOJ9TlgyNBe9fozjlSusXKYXGn8MKg0Ob3
UyYGSBxdh0ME2JM8Jbu0V7y284DA8Lf9WzqaUN3w4mdQ7Tx83wG3J23wnSf4sX5yppNoniVuLV9R
SoDKtqhABiCkW5VABL3uukqy8VsSkNHvB6oD/z8SmDDIYZYAI88a+5LSOMA2mbgHB8bt+sX4bbBX
jl/CeJ3KXKwwv7WmXshdTir6nzX3kFNfLAksQAZs2zIMIKZFYW+IcmVT2CzAkXvUQRviWBXpj/qU
AK3ZYj/TfIcKOaMVQQ2r3B6srQ2yEh56ROVzXlk56Al83vcgbS/DIJY/cGmdmc4M9vL4YlqINKLa
uGNwOefI048ab4slXVXD/zlezQe4v9kx1+9LxCfKYuTJckG5p7iI7S6pQdTWMdSCKPwECQU2E5MZ
N+VvA5cxPH7JkeXOuSvuSrRl/UozPctCEk8XPJ6bi5aKqElaAMyUh9PlI80GPp6dNBhLv7BYjEsQ
QXKKPThPgeYHNoK5f2YLohPqCxYKylsFKnFmkYHHA1Q6weuP2EvHhmWbdSiZXFHUZm9mQeYFXjYH
QZd2N3ijix3ws142EAI9wM/lqGDS1U/zjbGkzAM/3gWnBFuRJj9/enBgQBmc2Yn8iZtcmzoWatCj
oJ1sNevJzyzDzzu1Qk63HKsItMNA/WFRdwVMaXDrovYNg9iMo9OQWw32N11WVYotiuTpXaE7J35U
Z7CgjJsFECcGJpbtaSMwTqFlP6qOuGq31sVencLkMBAomUiV7XkzfHbcWToWf7sZ3X5r6gAX135+
C8ZcUI8aoXmDiIDCbT0Y/SV9tgTXx0lLvx51dnLBkCuC7z+ut2FyrWZahNzZxWlJV5d46wiVREsJ
VChltoh9Rk2ETfZiT/J+0QbB05aFUC/CYw8MIPQvk86adwL0jj0LCIxrEUd/6KFPM2Ok49opNgZr
Ye814HICZyYI6cRo19cHJKBKzYm4Q1OwpHapsI7HVi02YB6FO4LLKFABLs+tkKjKE17jvA79PKS+
CCmDRARO0Ym7PjcvVsDasLphXZC2rObkrttDyviVDX+OVr1mu1ui/hZ+5S/shn5J2Mv519Cs473M
vcVomFof+VZaN8OKbY/PiI1HvqUc0K8Bz3RQbOXdHQ3OlqnnYDoUSC25SiVdeJ8Z41p8CIcsQQtH
C5Qt2GlVnLuY5pWLloLsEhXprbfhDvySTqXN+8jRlAwC6Ot7MFj8ob9N16QQyILi9jLjhUWjCX5M
NHF21oG4IcrcIjEkQQ/E9kA0eKz+x94AIyv8mcGLouACG3Aoa89XrszU0zuh7fM+qt0ZkeclmbCt
sT0tVBcxeAiMOeM1j5xC4hos3CbWhsWhP/eec/8oIJuStFQ0MjzMvzLMEl3K5TzYecCw2Rm69f1V
JloXcvxUX5KJXk29eczd4Csbs6q3zcmggyArGLdFevDRaJkvaTlXXsUVY7QISQCTqLEjoTaN5mVT
1FRnVBHnNl5mLd7gUneZDzgW5OfTmoXiKC6VgUBtnBPoAb6/dxpLWsJiFLyIykv7QL7t5G+de3/t
g9oB0aCsk4+iAts4K0kaR3xO0c2FMhhU7dyn+PCh7H971vUVaGkO0Q8arY6ZuqaRhbIcEatI6R7q
FFLh7SVG5cQmIOXdCeLF+tqPLTfWEbhUaObEwl+wZJjtmjIbgqu4kKZjhsTjSl7KvLP57g0Z7O1Z
gEPI+gVcfHda/OQG64e/xF17bob3fpM9eqZTfUSyJu/4adV1NyNv5tn9uP/ZHRNHpnvrSurSEYN7
Bk3ITGmcOFJHiPNvjstgnALuRdSJY0D9b9+BfvRCMsLzUdpVxSXwbTjjJWq/zV2FepaAI1IWH6vc
Hy0eTQ0taL3LOVm86WeZ1Rl2l3CS1xMaoD+3+bhKE9pOgt1f1ls0q+f/XN9mdYZSpEDwrdb5OGJy
YitFnBr7ZX1hnimM6yBeyqzZvwOxxGsSs9FyzylQeGS/B2QlW+pnZCkv4e3k/WRGJRkrrcWzfEbJ
mkD7AFDGv6uRLGSBNn1rOaRlCSsjrRQrDtqU9SHgTu/P7lJMoTtrNqmkY8HczdNrcKMbWRymmgWZ
+8qZT21U97sESSElehQ3+M5junEcRnIm5I780QVFmDfYQMi+bb/q72tOW7pN41MzQBtmrjV28Cia
JurBWrGs29+p9tOF0ScXtsP6f7scFIzJ9d0spd4y39zEPLLhYORbTIH7gXAKqj0oIgHpJTOcL0Bj
QX5JE4tgSlCHvyNroryjizZRGWmZUK97YZvEE7FsGzJshDxQYlyW5KXkVcT42RaFNsT+0z5eDv3S
HRplvMlFZzeSweXEAL8SQCiC0iKB3uqxtsaAmK3TGobtyhhd9+/HRO1ovE/U4pQQ0ULiVENoAkT9
ng53EyE5X+f4UcwUzhmurA5x/2eKB0H9X+GnOxEm/nuQKss5ElG476KN/SyML6AllwcOyh4SG3hT
9XE0YWti4YAKOweay1OyghCmXW8XmfwsMd/Z9XP3ztWOz8qgf4lAKsgykp/bR/CmmVzMvcEH3Npo
71DI1toYKdRUK02/h5tc5iLocSXGBRIVwvEVz5nM6cr2MwjWA6ijpZ07BTz8NTWiMxSdt4b91u4w
CcpJ2Dztn8xykVpjfiAZ1lrTptDDEw/FQdShko4dDGExNEVarXsDOM8lExBGtCclmMzAGLOxKhez
7OXeyB9SAcJD/fclwoMuc+/hsW4ySFO6rDIkZj0pvW2uJ/+5HSKeJ5BikRKVLoH/GVv4RoBjCz+R
BnIhA5O/7TZdF336+u+eAvhoJTnu1ArVsgLEGgECkftOPUuQFlGJ1dEt/WrjDnV/3FO7/VO8gYh7
c03hqgjfzwG0c3idE6OWgIAjeSZvrfpRLnQKvth5VcI0EyrjcXdJN4dKIVvHnREzcEagfaAcyEiA
B7Q7BkBjljk3Iw2YCVmw6oE41BRu95Vcgff6nkNmYZksOGdF7Fb5LS6mljW8QV4MOAQrfHXOkaRs
xizkOVgdSJUbGaP7zNuvwPxM/ZsCnKQLVHP6Vup4wNKGEqUvtlbAqQAwN87yLAKUueIZi9Wl3imb
PZhZv8d5K3mjJE/AFKiCrt0wtR2C80RkGkZN2V0ZLpfq9NiqA5Pmyub6P9Ojry168drbQ8fwY27S
2MLxfcb0goSzPKLuD1Q69DvCwdDfsJRqqPriZLk5wR0jFtT9citUzBC1Fz/UaRwV8Jdy/9cj0Ore
WmSVUHbMBHCfx5vp2aGkwOGq/I7br/I2nXno+/FMy+Kip+El/5fxEh73mbqVWOeFF+VbYmKJiLZc
wndjumTYqvs+FLxHBcSQgxizTQvuNep5IoG2iNbgvMdgeisQ3z92iI5HbPGTKE4+UKDM0Zzrx3N8
y974/37aRCSG86hZpjQY17+D70wqjy9CPMX1nk1vrWTTm4A65tbED4Pz3R+7SVQf/R0io/WWf51z
jNS8JMSCeYqc/iygVhDl/ILjqSjdv3WYR63k9Nohtv1FSxCbSC8p8pJUQfM1YMACngUu9pryfmVv
dHB6+M+gJRTaWCwmTT0Kgnb+Y+WcNISCXyLYCIqLXJmslukoMN+Epv0QthSZ0LjFrowEUAybdxeC
j3wXdLWpRqi0cjPLpR0ulRXCizGUAd4p2w8/SedVHkoATVT93XSWbCjz9Q9h7Lyl0f6L66F6r5Lm
iheMCQ7NcLCOtls4aKR6rVh9iysAxXoZR5N4iV13ewKAfk7qy44xmOnEjUg9cSO2H6EGwDne7gZC
eSG2D18VbdLpG+jNgMjhPh775ZvGGJW05Sa4zkOzaLFfnKtCn2ymRNh5vz2IvxS9Ev11EAVXKyUF
giUHiWAfmUzht8exnf1C2mLKh/AZrkynLL9clbvLsICppMzAdRpUuZIY1/dHQ93DUCk55lee4egU
DsDEDT592bi2rGJ0zJHrNwhFeYb19JjdCDmQKz8Y8PL/W1K/DPWRrhrcNPPJrZoZgrY8QurWBNEl
R9FLaUgQyB7sQwrVVN6ll0MEKKI8VCsr5pXNi/ymcvLNKZxeDz5Zp49vWvdvbG3bmR99WYFdvcSy
JsJ8ZZ9EoRkH9b2Dd3OUIF+4LVe5FAwDIIesICUJTwG0IgNh3eDKsX75KRnZQes/TipZ9TeDDViQ
Sw28ys7FWoRG/v8H3MnxOxJPnkg0UjOkCzUKNw//Nq3iWuK76ZHZ4PkKUqsAxjOkusm53HzTi4tM
mGIDSBG0iZerB2N6mg/8deuOlTQteB/z3ho2zE+3qe1Y3IWLcyHUEfXEt7jxk8G3hK9u000uapCz
DV/DQnl2qJ9ra/8evzoEjYfSjnnJBtE2n72IbuaDuTkmo2zBsGSH9TZYGCSL4lactVwGP4KHQecp
n7km+p7YqWCP6anJEmdrpj/cL9mcm8CfQL8/vRaNeC2SGgg8/dGi9GDiSNsaHUREcGl6EudD6qmf
raj7ZSPNVpHLceYTHv6Aq99Y5eYSdVggM30XJXc81b8xotSPes52Y/Ndvqie+J07MQf383ShC1UM
w53/W8yrrrzNbS2DdNvm+PbYM1aY8KXiApAJr3DlVpoNLktlpCK4qWd7TMwYzGNPmYrlbn6OKknG
PnLiQVUoqPwtU88sYG7Ihd0BV/luJkBT1evRcBI18+TZ1V2Iuu4BxonNK8VbnwOYnJpe/SHdEKpV
+Nc86muGBFme8iskJpQvYwT4s1CSl14QR33lpIgyW21N4ULO/AtIwz+ODi5Op6JThsb/5k6DsKhb
Ouhh1LPiJvfXwtAABVbcLu1A46TzZXRwG7Vp8PzG1sWR84p9Ph64msldj3+u+HVjs0QI9olLrj+y
YANWn9+uNCxAPRNBzY5whp60y7RNeXH004lR83BgBg8t7Vk5plDHsqe+Yolw5IOEb6rlLBs3YkSR
61saDt4XMU2gNNpkcFHF26zv1JeznLF4Ta0O8/iYWkOdYRrNA0T5ltOzf0tnN4Cp/R8JWZMQWHS3
cWNvLIzqDgAA/sqxQM7tuS+MOgZ8/Hl8FNQ/VltBS9cda1D4nP53EW+fwfniaKWnjFIlMpLzkRnA
OS85Icfb1agNJKwYJNME9i7OfO8ID9PAVwPYcA+1SQN6TsJBInRWNQNuUmxBsYu+vQdlwx3ZQPbg
S5thJonGLB7a3yZkpZ3CXVuM6beCpfLlD45NvTaolH3/ZvRO+nGlLLtXkgSqjXaXXKkZtVSl8/8n
Xij7ntG+I5vZuCpwHNWmyX/DAii5qiUV4MLJbwOjt10qFv/OcwKYMNuymkJR99epFwPxTLONa33l
w2DQS9Fk16Ms+D71ywE1E8rf0ZPnUqcS1PCkvqK4/g3xx3fsYF08Dn8lOKyotmy0lLuq1K6mn3wt
7KNMjExx51uBavG33dP8cN52N8nXvCYoF763hugZCzb2J9ayHuQ6k8CkWNjAo6iTazq6t0xooXtg
PWM3uz93Pwjli6UR1lqzdFxRNQRZAZ/YEd1pVf9dagLKJGIYFMecP6JpqYdJN6CLYpKsolDNbO3D
lJcI8lq4qsbGwHd9ZTiHxZA4UYEloDup0MDqwWdGGo7lf9AARbzBguxRki9dmemZ+kgTSKBjhZgk
3OlbcE0h3XSefhmqJsLEFoCpsLNdKEVnCApdwZQYiRjj9yaXusOS+rKhzZAcdRMB1IMszeKtyRYR
Qsa+OXzpWp4cW1exaZVUinfqo3E1HBML9vyJKWdexxkOcjzzFMnKoy+F/aeI6Au0W+/Y86VIXwIf
mVhhtpFSk8ZGhDBX6ckOlpJp2XODV8GeB5ma/rU5o1tk0w5u0BgA4TFcWLLEaU33CXhpk+F3tiMW
bN6si/Od9T0rbeSrXbCaKVjuC2qAN0iXDXKNneXpzbi10XcM0BL8xx2FGouPMzz+AvEGsxjCi5TO
9TmucULhdu8+CTM7ePEZPyjgNO9rZl939tCxxF5PzJevimpRqnkcyaCYq5hpKH8I8iNNfc0XKoJE
ymEgHlgwXjWY8DBz4lO1+6TWyUKmZ+JXqip1zpTWppA04go9TdwMUSFD7HAwe8JuSM8H+VbVNJIP
ih73uMJNSZx85+p71HsnqSxmAn+4/4Tv0Cnjg6QIN007mwZAw+Oeq2hL+f/m8cPxJl/f53+1Slfg
Uh2aukjU9Y9bCNiVXyvxG/Mj/qJYtzdW0R2bjt0MUXe2EZRTTnYIl8mXTPO1pYiFxwXm3WKCLsUD
JynPpfULniB4EPYCA3SNmDCjHozKW14nvhrfF+PpfXTFmRd5SVWDhdXWQ6ZkwcQ7hwNS9dAjjsc/
q6b6dbhMxEJR5d2f0DCxhIdK6WjqwgMFtZbcrWdJqp7q6cn+WRmg58pTGbV4Wd8BJPi1BnazRXsf
VPeGcjsUoHlf6eVjvk0hvbX+6Hus2tQhCDIhV7LxFH+NLWXuGoxKVSr7v+Qa2OXbBfcFrE+5+P+p
45wk68tI6VrH8LQjT1oziAGLVNdMP8swtRTfY1bwkxuHDKubMgkN8m0ZVQUA5M8m/SzclUMzg6tY
C8K9e+ne/wCRHpvjT2N1rxvZ7UmP8EZlto9gK+QXTXXyhq2wxs/RsSEvfHma4vILJZND/dLLA15Q
my4e6zPVVS+VyfLplZzZEtjYXNlEMuHBX80zkZfmx5mOeeRgXroZCchySL/O0BBp7NfrJhJyXQqq
i2IFlWyKMCIiBAW61qG+Trdi9ku+hIWiwWusJoN050DrekxQ9qrfAg+beDmjGGRWP9SPz2fic/5H
IFyrW65w4Ix8lKS3OtbaJZ4fpCaCT377pN0yPh7CmFPzm3F2OEqY6i1lPN3bUna+wlQ+dsSAjQ2e
qPkhoiDDh8lQuLFIicomdb5vCVfI6QM8x5yES+ZEyzBD7WQ7obDsoJV8PTvJSym7qP9e4JO/hgWV
RmgZo4JZgxdgpGOTNR7xJgTSxTv1RSlTJE3OBZ/8eWjR0KM9bJMTRmIQTwvfwYShHIdalDeecQkw
KjMqlHaNZB9qWovFSEwyhVOoQ5PV9zNCsd5uQIOS1+7tZL4siPt9rw1oDLsod3ZSdJnjHVeui6oc
+rZGly9j5hYt1RnvfvXaAsatkNIUC72R6rIXXztUpmKzJUoHhLGJTpGkI/aL4orSR1ffyX9F7Z1Y
Z/GLIG1w/9cJxSr1Kw+6fvlFNanIHlxkO2slpRKOoFkZW4n1UIe7/gRTouhluzR/grOxaZ+BDLcC
6xF1JY/lMJHRcbAVVJxR5QaJlK5insOYO6NQJeGDlcbKBHrBEW+u/5f0yTZeSloawLhKjfSLXQsT
OYfPMrMRZ7teRYkOOxiu7vMz3i+8fmf382XQsHmqRRoSWiLD2wjd8J+K33v2ks//c0sRwfTf9UDY
S5JuwRGEh3xtFYmBIIma+SqeLVqYYPH2P8j8/LgYlNs7kxJ/ZSyGW0gJjSJZI+6dSYw5Dw4E4mdI
PqC3PJSC3md6vXbwfewlvit95JdHNHhW6/TDL1BsQaMx5XTmspC85STmAP4ah1AdHI4ABLTIU4ic
MD1oWKtHtGXivEeuH4ODsKu+MFw934/yoMSEYu+R1NVqLn4ihLq5bGY3d31WG0xPcx09Xv0GA2Sp
Q0yanCbJc977WnJQ8B8ERZWNhWyd8jcCchWIuvl9/BIJ2qM/bZSU+AE53Mr2RShV7nMtvUPkOaC1
5x06F8fMbd6VPh8pOOfrT5omGiJ8VGgtGVjt1PhI2dJFb02oSaS4yzjDxqTBAh+pM1bwPp2KW0pa
CmLWibGWs/9CZj1EIf9tW1XoBS4vPYEBLy79gd+gBZFH+6X32gl3VlvoJmnPEZ+kknWJiJaGPn+Y
Dn/LBBvf9JkqHU2qu7SNTCBZceKiYmdsyS3arwMOmYgv1Dt3jH7ymckQkCfkwYz6LWOR8Pz8LmqA
fUy2CeQfMzNcJ6P7QOaOLFBZ+S+Or429bflLSgtBrc/T/6H45o5dQxg79d8JtSYlJLIvDWQZgr8m
Ex70vwc2JaQQziKdArewGbW7gHN/stQGz0SBZYd56ASnrcK2oK/13iPDCH61YatBxxb8n6iCgDqI
kGsWrNRcmkDh89RgYiVum4PrX8+Jh/AjqIV8spqNZdLTwfqRI/cwQvtqmPIlyJB9aSzU6KqcORRv
wb53d7KQ1t9k6CKoQrOBpuzHLG3qv99F+/5/7rd7lpksdWmQiMOV6TnF/6KoErynX136PGzpNK7U
Q3dQbiAv7TKQrH+Ht3rrEp4EaZrZ+XIIKr4xTcLewmAJxzL7ksAYs7OA6YYe4cDx3tO8QkH/TGQK
BQHeKS222uGJRwvhjrNz51H+mAHHDUm84n1A+dOhK5hMMnNCU0teUgVyMEywqc5Zg9IjzBxTJ/rv
hVozGvY/uZXDUYFSw4t6VfbSU+woDecKqTRCsYI3fx7Jxs4OnWPyXnAVyymMsVHEhQFV+e+8Pg9M
lGle696Y5DsKYRdmZbeWVqrJXYmg3J4ByYDNgaTFCBdTQXeifmqc7rxFcSV6FIHZcCfUCCFZIYU5
XgiCKJSfiXzIuy/4A0LtjCv3hKdpCbUts3xwwUm0oGzmfXcwHfC9xGDyE1ekDS8KvLPrsOenbNo2
R6tpAYhNUr6pthyBqm3L5CbCo6VoFbSyhodm+QQr9uGfyvCGbEj020zIwF+GfDzWR3rMuHO1LhNy
Yub+6EIhxa0mpDehIPuliG7jUPnBHja0iCHUw0s3oGsgbhg1+bVBQt5i0zTgZhlPLRM5p9vxDQAA
ZndPtX7Hss/UnI1imcM/V2gkkACsQ+AhMMmqgC3jvIGxBqGI3IXusb8hbaVIhq4/r+wGKYVDF854
FJQ3eIaUXveqQ3pS3SbG9wNPA2iMQBqDc+GFYBvQpDFfjvr3TlaeROjlhM4NMFdUnpQcTQVawPmR
sYTko4web36OOGmJp74uBQfKi77VPGRlWB+/ekNVzSZFCUodx+bRbu/+UanIN8lEaFX30PkghuxH
B5KO/k+Inp6pGOfucXBK+O5cwljVdiw8nDdqQ+W9bmhqlppwmmp64PbUoExXAvluwIWm/OJjHIUw
TMgxuu6LyPn0nzyZvArR7IZeS7IjNeoblcVxSLkPwwqeZ8t3O+JtneFd/Pl6usL5jB2iuWULyfQA
Mlz4bAZol+L5A/Ji8OVpQtrd+5XBGRexL8dLVHPBhro7DmRemR+FPHeH54ToxG8qAAnWpPiER3kn
7q/wuAIuRTYgKoGGqKCh4ikdpvahFZnO9azEM26HkNPEBk/l2xAVbt6W2P0JrQmNC3CdQWzRiOdu
drMgUQ7bfGAjRrE5PIyUCoe7obeuX3X7XtzVVN/XTlUtEjwgUMSNho5+bREFS7RtnvQIGzU3dsYo
5B4AWK/ue9+ulPboLAzSWARGg4EaKYuTmnaI5OsR1Vs2uh1l/ekXnCpYAPowqyuX9rvt9da/nmFy
0UDolGBx0KPJeNKejjQeqExFoCjxP5sPavmYnoYYohuXfPYcj0ddEo8oJoymGa2KKfoDKE/H8Aij
28jvAnU5QWZGFZc7tQEfgLU2yc0juR3LXw+OZGMbRGz50AQclRUPnTaBq816J57jOjQQvB9nl9CY
AwyYjvdKJvsTfBkOv32trU8bVtrE5ohk2o3SEGuzr5GEIZQdFA4rja72/QbDu1iMzlHYIl6zJgcj
kz9n5lkiEo18rMIeK2K/8B5BQEn0DUBL9GrcvUm2Nr2srd9QO+04r1Sue/x2tfFX7Ts3D/IwoZKB
rUvLrQayaXzhpxVfYq6OfwG3QpJrUonDRoGj/15mT9UntWob+wIm5KK9alsc3UxLcXExYCMh+1KK
NtrURawmYwY6kpx7HVIrxy5cvRzNOeZN/WgoZfF3ZC8qZtp+d9SC9u5rTyMisppx2/kRuh6QNglg
aVur/wCWWiw36EJg//i1mbRZzKRUkj4k5fLIZmbWLVoM3xkadbaNj0ztXDurFDHYLMwq+aise6iT
AQ/yGRerF2jVjJPnrHYBlnQtLcpAvfH3/qie0/HBTd08bcP3j2Ik7cviXeZM36vAiKIXglxP46MR
lVk9gEOtveWL/+2feczDh34gLiumzNd+r7XKAOiK0gDF2vyX4jb3L3I04WzzgpF3jutCqKDUcrrr
yWjmOrIch4Ziezxr9SLp6HUFLTuYuuMcYPmj5akvNAKHxUAipqf9nhrK6s42HgeJ3giQF1eQ/lzm
O+laG2t7BZj862FwQdzYglrjB55jns6Mvm0ubTiXvhAO0R301WHtQjsP2WrfPcBALvYGgjb+3Cjq
gM+RFNl7iTSHMWl+DumKKVGLBLh0XmC+XDbZZorz/1ybSdCFi3UF7nbp/n8A5IQ8IivgYEutKkbW
KmaKQN0Tat4j/rBXCa3xxDd0aWuqF+rx+ALnY9segv0usvtv+a3W1ndoANTGGSTFxvW7UCkhm8so
9lJ94tg4hdfrrZxv0Ec4MD9Ryys/7NGReaZm1htJmY33DQb6IJFkKeC8EExkY7CXGNIa8TGKXjrR
NJEYazPb0G5cmNswPOQTW+7eH1vFd44lR7Nz4Z7VIp9pSgm8SbEp2/FmM9MBVr1GvqPdUz1CnWPa
RIHGo03LeZCW2CUB97kY2GGASn83z+fdPay0uLhxa0nixRJ1a2Z0KqykWhS2ZgkLWdRybeodkpW/
iW6lflBsoxTK5c6fvdiaUlAxaCtd4cLDgQlMkR7DYBwVX+mYqoqeMu8XJ7QEZK8mLSkVgkqHhsvj
lMCuspvNMBp+aSn78GDEaO65W3I738UQPihgPz/eP8Mzg4NAeIDItVqI3hRlSUSL1RuezmRdtMmt
HdckKGR6xrs70S6gcXvvfn1LC9MSdCL7J+yjNGpQ/Mu548tZYvnQiG/N/P2MZvc2FFY4icCbmTr/
ynxoTfctaOZn1mkEG3bSbrUMipuVy/jBPwPBJAiztgFuR7rawBNjVt7jYQfL/QeaNYjT5wlwQRIO
FQePM4qodS3a3pW0Bl2p88SfUV6qvBKnQz3ERsbuPCcsy4eFUEOL5Zebu9VK9cUHeFKAscHVlgZy
UuVGcHstDKjrOc1LLeQptzpHP8hFYtnfZ1gzCRNb1g3hQcfLMX3rFetKQzqxB8SjK72RuaiMH873
DDsPGbgfWKdrW47bg8xXDWBidlDBllBvw42dpmD5ThrZjiI8AYLICVaIWJ1UiUgr5pGYEJN1G90B
5Ba02cKoI1pHzGIEPDeAv96prfqOwH/nwEoXZrvnrqqtNDIz9zrptSzQ10wRDtXbHoJ4O01fQEN7
P4jU6qtZ5sQsONpHJtyaK5zWt8MJnD4N/MMut4B7frc5peXYmGgaux7tYdc5BookMirpktFGHEkr
fr8HuoJmz0UWjIYh6UpcwU2Cd7UF1+uQtNLHTKI1Rm60Qq9CoGSq7QRRYJHPSvpiqVsQ6xd5sn2d
Ypvp2K8wxWR1icSIMmu5lwviYK7LXgQaCffTCKHeG+PQGNt2P0ahZ3G/3w4iOzMvreJwMMVnVXKe
ngX3E7kfhpyflf8ofe/kWFv7M41Ijwsu6cUlNyJNmNcCp6C7nqaTidJA6nXxGG+RvaCm8F7yIQdM
Ik4O63ZI9TK5IEigCGf5zV9sqQtOqSbBkREiNdWrH2g2GjmZ/529aprREcmJjyQ+EUZuS0fTYOzP
EbwI+zXR0NrrAStYdIWA7uN/qCmLdQ9qdX+DZAtk3aj3mMRxMN4d8KCQlt+SBJSKIKVV5Rjpp24O
i62cLuTZOFa4fxoj5r/nRwNF02lofrSSS997ogyJhrrrkdbnzrwQTu0kIFJD+HZJT2nAsRpAH1jN
jDj8XV71Ck2yA2/hM5yVUUO6Z0iG8l6xnw3YVsc9jbqbA91dnJ0k2/Q7pnIxL9bML7C1I2oUcBBS
WHnaFiKOK7GUtAdhlA6qeRhbZpoyeqsMkloo6CgFbtwOWMMC71V0kdRrEY6+NqEKJaGYvxIpfnUJ
6CGdYkZTVBpWz1qWvD/F9y6dCFBHYAUhs+CnGkZ9smeH6UmTVkg/Xk0qvYHURa9kotagpXHC5nte
een3N4Hcik/pRw6VvVDh5QTHKUzLcBX4/NpGqvOpE40Es9+yEjebmg5uiCTEutfHgxvBHV6ifJRF
2h+NX9yRNm2v6SlXKfUWWKg6NaCpytoGdyHTVRt0EB4T5FSJaR9b9phwP7swt0rzRBxoh/LOMXfF
Ua19YuX9yl/ZFigrRTHRFZI8EmHiQd4u1Z0NOKQHcy85Y/ZBLsggx6UqZK7swgK6a8f2edg61SOt
10E0dizGc8KCPK4uyrOEOHzhYzZLGJjjX6PrscpY8BsUOXu+1D4k2vTQJCKv12C3xir0HJmfVqH8
4vu1cIG3slyExjkOX7doIIFpo+m/K6mW9iUaPRs4CMdOrXBW1h3KbZ3Bp1yv6nyeS8emCC0sBDot
xCwHqafOUSpGwvLTMNlqLRk9vUgvxxZjVk2tQyChrk1pTxj/wcSsMwpXERZs9q3CE0qRhYGLfQGB
Ku/fFf2eKze2DtIfJmdF1HLbeCWxG5fu9aw5sNWBzAq7Z7snKeMXC2j4qIlibn6xucfjGQdRNdTM
EJlh5T2J3m5J7w3z7NY4E/p3d6jmikHSruIVLNPQHlTSWzHG42gWCERjgwVyDPSDxcarjXweQDwF
6LCQ4Oha+re4XwjL1tiDwpzUzKv9yl4cdJtJIAFEDupxWN5O2ogUkuKlcrikZ/aUVvRKJMH36eZm
UHM8D3csLYUJpskdCCUJ6kfD4CBJBU8a+VGsZ912RLJ7c8UwVkYLtpVqfdSd8cpRkuLG0qbiAte7
OB2qvx6dErnW8kILPzVpEdPZSNcc2QXjhdruqUTu6F6zsdQ93qwJGChHurv6wLwF6we4xJTEVmUJ
u4HZnpkWxUEo+1+lFWtQP3l5VE62l27ZKwWa/6mx5jfZHZCV2s8h2S/vxQqubiDGv+sShqiBPxqD
ipJ6afVX3bpkVu1T1K+hiKPUf30TAjR6PrkdYgfhWFo9w9pN9mizLEv9xVsJMRHC/HioBd8x2s4H
rKPx8Fs8DaRp3evuvvlkqEYygn4R6a/PKDNczCJLwW9fk4TBDsgW6h2Uz47uVIu7X9GvI9bV/fOT
MI8LPgedKi0v2zjRhWPcr5hduhJZ6MKdSAy5K3QhkQf5r1VNv/YjyL2hVSO9moPZmtSCnhX9jUFO
rq/DC8V0El8d2ckGTLk8y0z0te+8DX8f45Zf5MD+Lqxp/gWWQI5XdIwpB8bmal9wTyvSDM0SPZuc
3UEcT/rQ58AowcsGtgiDkiwqC7bNmMqX4Ix+iZRS4tbmEDxvDeMSGENXqjcnO1AMUia1uv+VoT1l
6D+TyBNUFkvMO18Ih/x52jgvP+JT4cLYgl4TzTB32R2hdJ4MWnAar2ri2Ht21C65mQtBkL16mphD
D0lzC5JUEnAoF2VOVA7K+b4kDyCgkQIMioC3ip5+S2mgro680uUg9W+1NpMwk6z4KMFvLINKgBYz
piaLQhOioF6aC1eW/ugXKxssFRGxgniA1Acz6Uq6XVHEo08Yh0hzc5t8EQih6sKDA4TFMM2wFCdF
DaQz+pA22o+rsf2fMr2YbKjhvmNBeaHYfrhUi5IbiEHHihX8FtFO8HhZjoDHpqcoiHqJWDzfNGtx
ArUAHHajyCbDUoYoBAqyL0mdMi76dhPb34qbuZOd5UsKL3Wm89oiQnTfR8udIokvwzsDshKo1ZWZ
dHuUTrWuX053li2N4HQfKTzHx4F80KjXDtkeMuVrlrCIWauUitW5qETvwXdXxg84MDslSBLS8De8
5h3hLL2+j/W8g3uuVI9x+D1d5ZBXLtrZGu5ZnwjxSFDt9WreNU0HtDv17heXYpBPMomUtJ38daEN
DvrAVmqWAoAmCrftRz2HABQfLHqzLJUrG2UxAiv9AJ2kQ/oK9jlFX6+O7s8dMg9M3mxvPC9Ey45S
JfQiAh1YR2Zs7++0kD9N1SSryOKAhy+cY+zVRJkbAsO6+MM2PbQ9z44nbOTPPgNtIos7XxqKu5hT
jx5TLrkcuE/L0zV/tMVZqBbNuKBnTEUy9FyT0cqW1pxCqZt7sG+qti1Whfddmr+0EX7ZUtMEPQzR
xSQRxwWF3g3fufYY6zapxamxkTl8Vq1sLFja43KDuL+eJrQXWtjghpnh/JE5VpMgagNlZYZc39Cm
IchbccneQ2uin4mJ3QUX9SFqikN7xscLAbhBtMHvNk9oLzfnCvpojkb/7eCSVsjsCyP4veYQH1rl
YQ0WqV8XhG5sWJfgnJkV6qP5Ev1JHgYZnOxSyIVUwdmtzQbSx2PKIX3YYM2AGKvsDqwT/aDwKCeD
yHhn/wqvTRafN8gn65B4pCKfloVwJUeS8CoBtSsI0+/0U+YSHpw9oKwOhwnWBEeFxeDN6qObLTS8
VDWdSBHRUbpwMoBBMGrx1uiYswQbCFKmXa+Xybc3PfsPS0LV9vMQJrR2evNy5tF4epqszGKg54Fq
CQg/USV4fsael5n9ywnFHcCEUhE30I837nIWXm0TEvP89F4vbaJJnGalZ7+Di12viHk/ENIEy44h
CaV9/Te5AsQsDbhpHwzKYCb2kfUxoEv1cHLQeC75KzaZErYon/5i/4jsQvUhHIl+cdqKGFGUVQQa
znCc6h/rhZ72su8jv0tARwswqDkbZ5ftKyuZ30jhGc5mNgbjVnhbSSYGJo3nTjcBN6xB+RUKzM04
TBLJtupUrMeoz/90lEJZrbYLWUynsUG3pIpsfPz7uSJ4222aP6x3RLjnSGnmLL1nbPzZph2MhByu
t3e9h26PEKrypOog0ElhNj4W0DLW+mNdd+qFCABTphEwgQ3t1EDSOC+2jGm0BwlKVXzqnFhaWlvt
S6gEvBAJ95rzaeFJ4JGao6TEeRWOawmZo1CEc7SU5+8bDV6J6yRy3Zw/6bjIOVAlOacvGgywdO/x
wby8xTRSe2ORRQYY2KnsSpZmqMXktfXd8Cps+FaCPUb19g5EDGlVeZozgiawU+OMC99NKUikQL7b
6hkboR/VGWM/nKC1+2Tc/cM2LlYovOWu4pN88ahLpqxTLbsZfrd2CsoR2OwwxEkMQfaokMcW+FHI
NjUMVHyzeoO7UdhuT2/GokY9wOZOUpa9mRZ2CE/J2wDKyzN+XgCCXrIffxdBH+Ccv0N0sCgUf4Kf
qY7DPTC3vjMeH9aNNAJ+iHsB252x1sNABUetvxHTeBHwpzhpH0K7BUrI+WHxg/nfru1ZBpjCVVKk
Dl7xlzbSqYyT06nS/3YwcJBQTNGSyn/K7U9Ya11tJBmY5QsHSqI/CPO809UBIEodEdmkm1maE+uo
e4guM/uA440aHsojQ+4op33kqW8e6uotTLBOqxNEaAu2HGN5fX/P/G9T8luQSvjkXtrAdHjD1uWF
nB3Dj1GkO+AKwRzmiVE43u/TwGwDD9hO4vCafpFPBnmhi0nZr0ONaqnNg6JFUPlCCv+iUHm16IBl
s49SrpiBirRWxJ1vE+oOgrltLeE+Lnm5dfcUdPWs/8kwWUsXc61kWfdnS/acuFw5If4bpyhXLhtC
dJP2f/IOkdM+6aSOtHYJpMz9gzgmyp/Up3kCUglieDRiVFf99YLgEgjc1+koBDsDha8TwBJyGD0A
0WfwVihDcc5bI7oTmY7VOuxJ/e3874flGEwhiWj6Qp31/T+1/GP13nwVX3fcwolvYHaaN+17+pgP
BFrizmVddBamp7EhghxGt3kxmMPU0e/9KHrQBjs5/Eokzcnx1S5ImYFORTarY7pW7u4GKwk8JJf3
TCYOjB7g/OxRePBFPTOJ28uJa8/yLMeJq1Yt08dAPBYR8kKvgAF0xNne9i5xm220VzMZt2jRI0A6
EXcAlrsOLHQR6jiIPYKBzXFZfRpN1vlgC1rQDCBeoS+YTwHnFpO5v6HxrlpTM/rBr5iQ7UdUGBRH
k6IQuHDVhYfLIrrP+JcGZG3mB2E1k8gBV9qxYcbTF9NhBGRu7kTCv24A1rpsbZf+JUaYldeo6EEt
s2g7OCjRmW+0uRllDE9G2dsmtufbVH/YTDFwFCqgtNSO4DjpNd2lm82UsSK+vKvDTY5AZwP1jIQC
Dyy59rkX6MGrR38VK52TLGHNS57eGDxCFfSXittvHg2plUnJIOeMtqYEkwf7P/d5K1S4UL7/TdAO
Qxtl9Ve5myeygqxJc8Q67kicTCjCsitc+3A+F9Apa2efetzuUlFRk2HBLK1UDk62vxECy7R6OCJG
Z5x045wh3/IqAb1ntpf9D9KMGJMSUl568kGETUu6AgyAagal9P36Gbwaya4bRUnThi9c9nOUtt0K
2QbJJZO6VD6JafBXcp96YteDERGAaVr/h0/0PLjOhbH2hX4KHTIhIKXBD+qP3rHuEEJWU4ZU6nH6
SQTkHhjiSzaMKaqi5+FjWFri3m6uGhkg5LqfOeF730yP7f1zhnlMkMjdyJM2+JYEqGfYKzIL8D30
AN9L6EXXsFfOgy9BMulDCwb7DwKZpJSYZXZLdczzzbvzltJd7cnugK7mlDVsV3KxRfkC7suUuNwL
gYf9JELerqw1L7Go6q+2G4JuU7A8jVl37UrbGLmYE/Pr4dH9Mz3av6OAorpWC5hQiAiDM+LnOfu9
ZEJdI47N5cH2OTLYYONHO5G4ArOhjQbLrwgDeH2Gy5tEPxdf8c8KoGoznxx6o8p8J9muTiCwITz8
L8m1XiQY2sekRvESYoB2Nmng0ECWvl7F07toDLEKx2NpKwECfZTd0JZzxrE+lZBvyAM+mKhoOemI
ZQSDTuna5hsGSHUVWLR0unnODeSTIsv/9tazhOHBe0/A9qCHMGE3Mhgh4XS5H+ouGOCdhVev0qqO
Ze3vVL+qkGqWKzFT5CRGahaXRYEHmrnp8tb5E83ozKoK94qxtdTnVYQtb36rxxaZXISCMkuLeKEL
PYS+NazOrNyXb2dn+HdIRDPTufd5v25Z0c8j76AiS3JXmWkQvEyo4rYI8aex23EMCgjPlCOjeB2e
oUdAh9AMHn6nImfkpoiuDaaWe4EQ9dsgwuSW6SDc3sUmUOlZc4aEY0XvkSitAI4Zc3TGmJRtWO8M
5becFIkhYcROLc7XGPzZRK0G0R2UGMFWSNWvZnuhybLIJ8vzsEs8QMI5ZbATeXs7ERjdkhYKeMtl
wvEScYQTDWeHgfuv1ogDhlLZqmZx52OCYk6YaYPIPC8VXHoqH5rTWytzeMAduh4Kd19NpvV8lLPx
Ts10RKxwwAoN+NLIuc/zumYpX4sgVqlPZQld+4mT0yQFt3QIV0yTIriHTKwlJ/7ZoT08eObpqlF7
OzwtjBf7aLAWO+JRL/jAfbcYWfWrbjNLdSBfXFU12TQG0FESs12AuEto8WTg6zuShSFKPnfhYIrw
kJq+emge0UVJKCwTtWDlOCeuzVm0xBX2rOeWEg188JKsnAYbSnR57uPqZngZ6GtJzyfZvdHYsLIQ
pDtUKOKhildJNNoZhRzi3yqYGKgaP6Pi6twzvakc8D53suekS6tcx45CbMb+0UwrRd47GmgpyMsp
kZp4kcqFF6CkimQpMbNysbM0FYLZXgwhw1kXK1bvi0vfH13Ffyzt0lw+mBnw2iwMrwqVIWXjNq/x
15ygwBqtZBFrnX/VXAi5eCOJHtVKDMSmVBPV30YzyCS9fC5OKavN3shfcmaKkg6VSQ7RAB8uIZPV
4AbGwUuTqGDvn0zEZkjkq551LTX1DsyOxCykSDfueG4FjGwQJQOT/C6XEVit5lbt9TuObciW+xcb
FbvQwgcT8qfLVfQOi+1/RpYalWk/mIy8ZkXHPgxe9/4rTUlXDq7kCuDo7mDWZrOtBolUNVFXW8gE
nub/R35DUEBLu0MZji/yeaNNCb/+DC+4mo4oJUel3wTpd1uy8VBlwVsP8z/Ow7PD4JDjDWA4Siwh
dwRCalWeapVeFy3zUmBguaYrnrXZ7e/spBuH117+fD7PRr5LX/WbQgh1Zp7I6s80tj2NpggpKhDQ
VRbTF8FbIGPxqx14uKkKaI7dfNo9fWDA6KEddOD7wViuAsmK0BOfWl+gZ7DVwa9/dAOkOJPDA99G
F8x9BrZwfZDR4TuRAtqWpzafHfyRVSR22cBPgQ81HYnwrjONMp8JSCkbmgdixZOn80xT0WX5puPd
/DUBtSXqZyfdXRaC3hAzG11Qi7VhJn1i73kMm7gUscmAFFveqYlC3+ARyu2ofgkdYtg42yRCwrkr
CUikfgDiNWXs
`pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gb0PVdjs8ceew1zNMMFDynFmO7Nryu5D2IMVeIlyVQWuiXG1eT4cmyfjpoguoC7n
i1+A3Ui2+r7t+njeBztMN1cxyrnlpDEaKzAWxjLglIkAqF04hTWqDLuXvdw4a/PV
2iJUsPU7hyEv/FFvLHD0RrICyS8MPWwaQSwObqGDLr0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9296)
QzjTG7AHK3vXrv4gDmMYzDz4RbhbUjeFALHd2ViSqrhfI8GMhSu/PUl4Ekeu8s7g
FyohmhWR6wYq0G1IVbMqdwzHcOf8G8AJGob3HqwyEiB5OQW6Xdmp2Ko+rbCKAoqM
406Yp7DIctIxhR3TlyKj2fsw/2Du4bxwaB2IvxBqJnvsiiUICkNo7OFwnQNJieQY
Ffpzf9rAdqdqbf5A7LO/xQLdqLsKlvvjufDejfJJgv8rw8IYXXHzHVi7d96TI+8a
7+35o+fY0DQpdfRbom1lvcibZW5gShyx+ZpbRa0WGKbH27ruaxpKMHfcJ2g/kEj5
t5GPtFMQDqeGMFvBH+zcDwecwi2XMZ8ESHVGirxX34+mxrEnPm2vop0GRyhcmI//
EGh/MNDfz0PCtzmHY1qALo8iwNbEBt9UL+lKMOl1t2okSWbP4flVxsNW1IuYczsj
wAy0/bBGPBusQUmSukhZSkWVcAk+uPU42E6n8HjThBSHakv3UAom32poxSxjD7nH
//+2VPqc5iW/Wi8L5X7Ua53wi4mFfrKKS4JmVQWs7vi9VFdxPM6RAZcyFDgr+pOi
KLOmAd4fO/CpVYlx4+fHRHk5c+tVRRBRfzNtBUTOhh2pSbXFoiIXxAAVIUXvkhp+
JOTT9ItOFUfknp4RxtBW6WmzUiKL6QHZ0wK32ej6MrEvZJ/7s+jWpwoSx8a6QP/7
jmHjJDSsmBF+wuSSayKq3zoIcAdKw9udysvSQQsytKINewqd4q3A++/V1y7tviYV
3Aw5ttvbZE0y9ZgZTAnoakDiWjAA+lW8EOYUsArXMxkhfoDZDTX/U2lNjbGHDNER
Lvspj9oP44bj7B6hFFw+2MqbO5IOThBoqezsmGrj8NF6AJmCIOlA5cDmYHsz1AH0
ce5l97UtSGvBy30nCzPD7aWOi5K+4qaa8CeaCIyW6npcc+z4B/dHOG5LsPgRoDBJ
gjjgmOTb1r6ftNc7FFjjKoR0qmB85QJh9movBM3e1LN5NDtKgF+qowfsbjS0SLAw
bt0EJKRLpt5eyZIhqOi6O7XfB0aTaSbYBOUVZzOqxmM5hMZwslsBZ3nip+mQI91X
3FoupAkUCrcrMl/9ffnwfvbpC+H1eERgYXVThHxID2uH6BR5eNgqOG9bMLAG8Jbl
P8MLRkakkfk5P5Jjfl3kNJkVmRXAdLphNN58wOswLd1OLSVsWcteXa1gruzvhQ27
0Bw+QvZpBic+5cIHOohk0+YwsI4E0G/J8czNgTT5Xr6bAat9dxUL1BBscuWdmZMQ
NRF9mt8M0yNvkkb2QoqaNNN2ijCBwO6HXITCJiJRmB962Fqa1QCtI7r4cDjFVc+3
DJ5tTaW04wocpHJFpCGlf/NW/EssflAD9wxYKyKAcSJF4V7nVdL1s4FHl6BZrJug
SiVlbPNAKosUM1LWwq7fImzdLV/VSXaD3rmFmJ3hFbncP3Cuo4JKMSKeKRZlbr2G
zo8XBC8nGBEnEF/z8+MwHfEamqLNeplh1sNrnfMQLhl1yCdrShqxofraq62Em30x
tjvs2CS/DYWoyOYhiT+h6l7ABBplcNgwIE1Iz4lH+ddIt5B2sDxf70Dmh82+r5bl
2/YCEvJu66pSjCeLm0M1/9eH6tLCS2a0CL4LPMA5SYFicY9IEYbZz6oaLXoFYId4
x+26XLsXcOL79dvh9MX0AkCp/HCqtmQ8qpBblR4sneV5KxLTTqOoODrRgmXjE/II
UBJ569STLNwAD7LglZU+z8M63NYW+dnsrgo0wqmYhmT5QMGfCUCXaXWhUDGo2sl9
bKP1zMR/UmXC7+Gx+25YJsjfzQth7f7V8rGFMa/AMqC7XxHk0J58I0U7fh9JAmPd
NCvYu2iYbrT0/Xy8+AI9mOgATLJW/mL9ZOznn1CTjl1Ft/c530SsTG2OdszcKoAP
Jpius/AUBHxS8o2w2vUseWCt75wqUnAfBa8+crdtSRyWpE9L532r7lCz6IEBVvjr
EmRsCGrA3kNzLEjdN8Pk1dtCr+DNkaIRSLeR2GMZtPiT/YhvocBMNOi2E55bICQr
Z/lYjMlCWGTmHrdOUeEAEjZ6ncNC43UD2yJdUwvdQc1qTo0mzh/LV9j4bQsCTBbm
tBhzdvDcsF4mWPj+JL0DtqbVXYaQljkzNLdRHNym/o5lUEDPdX3K8NKRuzFZmC2J
/c0ywnyUzxkfdXZ/s9GrHAhGoqISGOjCiyiUCQlnWjI4VLd+xCc6pOsLZHZH0BM9
vSKgJ32ivBL0ph7K5B1++ywfLEV0eVnOYITJaknGE31UIpT91HEWWvO2MECWaYab
nbMCAc4ejePWJlFjz0IxFev/6oXHSYyDsYNkE90hMYgQycPQg6BupUA+wbxLz5R3
AOIY3YT6TPuxHvF2XRoe2DoQIR3h4+vP9I4DDx/74rA+ZedfWLmCiZsqcE2fakUs
P7sQ027kWOQ0X/FkX8JPBwC/dE/lF8zTRZI3degMNWVw0hWivnwpPGja5XIdhGnM
/AO93ZwHSRk3Jt2gBOWmJEy2FYaatXLNK6G7JKXqje1aB9UEz3p2DxrK94MwIVEl
MIzw/BD634rjMeq55OtAns33OBsCy4p7IjBAZKhLm+a1Y2VqkIgDsSir9VJew5rJ
SvpBRZiKT3chM+tUJZ8sarAkM9MzfJKrFThLuHWK6ltTYqw5+e425iAuX0ycxzRv
JZu6Zh2vieSA4Ns5mtozaxvDn+9YIu1i0369PxdsF7yNLyJNf3cnFVdMS0jcbLtd
KdL4Nwx/g8Qe2EWVu/BPwdGXWgHVY95sDhjVtGOl7qZ9JcY6g1k/sa8RDNq+tPXb
h1yussZ9QDioRmFCnWc2wznWWLGUlzxM3sbcIoopS1qR8bD9sF8CMvK9ef7HtjNA
F1t88ryl9R6RySdzbTD2Hg/n03nu/g2IcKk02Mi/TmtCQMXByv6fJD7AQMI6Funt
TDU2CYCYEEGpAdxr4G3kh0xR3k/2YIcQO0i45GPTu7stdnFHaUht+QqJ+wu07t5M
LSB3/befARAA8tsJ6MU8dzJpczfBYrLqF14KfWF5KihL4Dyx4Ol0lHLfaJHblRe3
gKCquoeAPLPLPdnqIHlxYKstpt0f/UfcgoyOgbcnbTSQvjth9UxUtq4z9oT8OGNK
9aQ1CSVenzgLx8UEcI6gWMQAb0DwnwRPoY9ZzH2NFCbf8RyLpF0+w98rllX+H88k
LcJsUVT6n+sAFbIUpTBENmvIm7IEnSKyd8vZQQC9b7+2XIp61aHFgj8LHgO/LJNP
WXJas8FlwYDQZNFJ4HY2ktqHivfff6g0VheuFA8WHR5q+KtnZUEqpCWCYK6v09vm
zA4EeAz8yQGeO+2uUKMLTmIVXOTljcEQUqhNNcPKjlbwD6lTe4dF55PMtXDo4r3w
iP2Xuvz1+n4XhwfVJWewEh7Li9i5fOmFMKXyMYWaIvo5MPQmqjC6R36atJeUcFn2
AfA59vFQJQ6K2cwh8RmkFB1f//hX/hjNTlSvEXzTH3KLSMcxA3ObFVMLQKaadUlH
Eoqkp4d4NyZIGX8aUvYQ3wH5V+I6Ib8s4/bPvLnYc54yXIbIg3uhyut5y7jqcNJ4
zaXgZ86K7qSzrpHCg/5Du34xIEtMRN4wT6ZmY0eQbZX1ty0VRrYDGggoi4KjDu0T
8JXt6V3t1GQBENA69TwZy0w+dgjox10p4MUh9FozN+2FExpKFqEWeua4PB7ekMaN
NalrprzaIToMZyqzR52HST7U8fQyQJtPGSCzQv2qdMGE5UoSv0vQh4Pnswp0sn+e
P8I/HlAbt8pqcAxADnythVIkPWoOYyxdbXwrmsrffvDP3nWZFxsPeVByAFv704Ds
NjTBAvNaB57Kf48hDc50tzaz4ZyW6NNtFvUjF37rOHj2OndQDqe7BfpG04A2fYd1
5P+ILHZiVNbUO+W096oSvNGA8G+NsY0fysos2/FaQgskdfZcvCP3Mz+tQYauqQDr
ooJ6GPoSvNiqWCf1ewRrfFtPWrh9NqML2NSarfIQcspEVHtviqOiSSIoL6v9Z5CA
bmkPMvFsxWZRXC5ulrttNvELfzfzA0N1bMluwv/928SAM0or+TuKfUHpHQxXHnj1
007gaSaaxNcSvOfUdxPQZcONfFEfITmEK7RJhOzsEJGsXD/INfIqetEWr7klZXKj
nKc6suKy//UBRtH+TukHWg/mOufXUBSvBCPe1lKCAGeYkUOagtAbSMs7AIbA3ck7
Rs48YozFvJFSG99Uk6maiHAF3rLKJny2B1FtS3DGcOtNKPeCpcDG+SbDg1DJV30R
UfjVxC+t8Flsw8NGMegZF2iP18MuZmmNZZZFNragM9CE+t4fIGSvryJ/Yx/8nLWa
nfVpDpgvTI2RPwVC/hEbpdskoCNew2EuMxwY1rbMT9nLl4B/HOoF954tLQI9tdLs
U8yWnfhYQ3RL9eRigZcK+3vRhMMwBvu4MqpbmrN/ZogTTjFAfMTTSKkzdpq/XODI
t1mFBa9P8WG4582me4B2HgKiYpexPNfELad2aE0a1s0SFYuI85KtoCWyk5LSfuMs
xWCK6xk+z2Z04LZed53IWszxbO9v+ypDlxMeHAuooD9TsKFOF7Zz1ljtepoIZJV1
m5vo3lnQlRa7fv36fvFhygtXV+St/CtYjtCWo+qEIWwOJUQPWYylbTX8/pgsAYcG
lOsQXNgjKmSG8jJn9Uj65Si5MKILzscoay0DT5UsqUXIiMdIZ7qqtGFewgyDQMin
JW57Qpwfv/dIwW6u/rSkdMc4sayMlHG0kLB05d7J0DURaRJHVZrez3gGlblea+Pi
LF3Xt78qX5vqwQ88t8nuLLg8R8Cxr/ww1wlpoRJhR2sHP20zQ6BinOeoTkFtf5y6
z7lcnRDlwXSEe3FfHY8EJoRMxpdmlYW0y9NrO/YDkzx+a1+Wb3QAs2Luhu+ZQbc0
n1mA+Ojz5vwhd2FXG+EDEDY2bSp/kC24axiEUIJFc3KwWKIL0N5BN0ZjOXukdTSP
k89leVVKMkX4WL4588FysDB061eyFODT3RHdH0+b9UzO3XWLFoZlVTB1YPYtF1R3
Kvl96AQjYbMlfGR34uiiIj0/jfQHfu3PuoUK7ECrW+6M1nAbiuTwsX2eYyo3go5J
qxFb5MJehsG31pVWU5lxwG2ElmuFziTUsp0Yxm6w5olCGDrqB+hjHm8lfRWDletu
c9KcjoGsjjFxv6CSXuBes0MTmWoMqmkuOyO3IyY41oxk99MdKeCoANirh8C6BmwG
6fF/U+rBeVnw1osXR/MMhXcaCoVOSpHCD93kLqS930F02lg3/1IEGVUVo/4WL6kR
yyW7231Flo7mgTUXJa9PWnc7U642IZsCcS1Vu9uXFdybSLhuk2GG1qU9i264gz8D
mwwrQObqOXu6z0SX/g4fOEG8AObA7Nz5xHnPUE/5tbA1bJWMI6APmaoTYKg+tBwz
kJX3SP2QLHx1pDmMY3v5dQLLlbSDseQDea8bX9GxAReNe+CzEbtb2jAmkPFm1eDE
U474QyfDun7lkSydyg7Ib9hZJXGC83ob/5qI1Imghm3BGJQmPLC//2cupIS096QB
CIw8Lcmo0NjHbfhqAIDjB7S3u+sK8hv0oTBoYDI0Sexm2kzD9X0t0lkhsk38m+in
0BRKZpQsqIMVboF3PggwVwVZyqWzjxdivCqITu4+GRhTdktN4i7rda45bZF+BjxE
ridGTbDnR7Ho0SZ3vwo/nDF5Qm/S6xGKP3gD22UEIsFdgJL3qvzsMf01SIEwgtPI
RkmE2E8TI/1vM/n4zGTQhg3f4tCfD4FjOcOstk03semgg8LZDfUrvcaDWpNxZiHY
sqSDpnfja5dYEYQU3jpvHvXpm82ijpVGEZC20IAkLKItbKm6nUAFZxTkwjo+1YDf
Jm5nPU7BoTr4HWp98afft5l0qgM9BPTAC4CJJAYXXvVxZPXuxH98xA39ESH1PPFy
kF12tK/Ph91ElWTJ9sHAxosiuGgNXR8ubfdn+6dVnTmTfyOeeNAa8oNJYTSzP13l
m+O1QEXbtwgXihhnLjTgpg8wrHgYr0jF+N9A2SPVN8pq47x9muWvDyaa0nFTd8uq
4qfgWKu0Ri8FFKxNeaahjGimqbHtbeiIcVJ6LyCv+op3kLmGlE1jZuPatXdIIl+C
HLwcvVwXuvHULxV8i1W9M91eR+2LmRhzNG6vzRfDUbtBhyMfWhN8I9Tp5/oOvDsl
BQl+u6zdceLEEkLdH/3XLFFG9NYUr7oJ2A9LCoUlIHAvK+Qe2a/j35m8c9NV8R02
wjc1A5LmhExgicqsKQb/cjfzIMSrwQ3Wytjfk5s0bz6LfgantyMb55wrLW28ROMg
N9thxE6rfEsCvPyVATuAL9YIfPAN5mdT+GQyUKFAedyjndSQnrWE5A9Vi1SlFPhu
9g91NGoY9zqyrbgm4LgiZEcEFK6ISeSDUrK8KbHE7vqwAhBzgcTtcK6xZ4ZujUj7
/2QzZLOAa873iY/uAfWnsadZ2DHxVB29TdJtFDBeok/MxRWrgIfR0Jh291Pj1M1D
TjYWQmPWhSFS4F/JmM051Wqy7Mi/g4KnU9BsLWRspGQFLQV+pLNM9rF5zBN9Sn1U
6RkhfP2OAPXyRiW8znIklj2APR2VImd1yGjZs/YGICXXZ3lwpaUtU7Tvy0UeF4Ul
n5CjJWtYOrjXqgitH/rq9vajh1WxC7SW9oCMty4Zs816o8bcvvu8W6L+olYekpkL
KttiIWM2kDO1p8BHlMvYIVqE4URbG6oQXA8yRXArGdBt2D9M0pGxOR/iJlMm253d
w+Kk0Jd4ZOb060zMX89z5tOIHGqo85hxJ5tF9VL3CWkBJxzoWgN2RJ99tiDKmZyE
XCnhy3GZrzNr4HmaRIBWPt+Mntwi5A4s5FYM7fXA+1kRulM3zl35KfC/MM5GYyIz
shtIlYZ5cO0akaKgJAh3EK53JGBkmgaKC9IN0c/SIVoRnZbq+xdBpeNicU6dQJfr
yC7kZYNW5isYw3WppAuXxTt/sNv+Nn2mkN2u7FEkZztZFc8y7epFfa6yRxfBi3TZ
uV07EfY2t+uD6yK8aJ8+AQPxwmwvaI+k+W4T87R7ouXo7NDLQDp5HTHDfOYJ1VTt
HZYWOkeAkOuhFVD33MSW1pLMCPhNI9dPk44nn1DTGjzuv8mWLITjZSKfj83LtCtF
L6SP4J2wvBRXFOc0evQT3e+lbCIYruXxpn0ts91j2UsfRwCFi9OuGT1cvShnD8rx
oYBTVUKKt64YUfqaZeSPmRYT3idxtOfWo3nRMbLoSBGKQxoNZmIT0qltP9IrFL2h
fZoDOgxan82krktW/G+uIqmrWJkRQi65SfrebcZOk/BzaOwzA0P93JOxweSH08Tr
Mr+TqU32YOXdNCuajA5rHJFY/lHedeUGHMRl3ETG5EMQwSk324JwntCoDgUDJnPH
gBfTChIrpTkNK/hhmC7b9RcnK3w3vrhFTepkvZskOBtJf2Vw5k633cPYgP/MBbJX
PbL9njddmy24gZDP3j0XDDyZj5MRexUJLdShpxTt9dAqiOIcU1JUOJ9JTW/BlbL5
xublNrYPyqu10dgRJbImDuQDqjjsG5YGhj4Bcr+F+dmVhnVkN7GNTUVoJ+B42Jl9
SUXNYp1AqOKvkjv17GvP8ofzdGC2pstvGb3wyiScXlAAWexF9pJqQAJtHt5m0U0y
N/RPYHCC8FTiD2s7poOohEVWWTAM0v9xRcIAsRI3CR2B3frgxZjXunZlcBlW/4Gp
K/dHZMexq6C3Gvo+j5L4vISGF/npbtI2RFQEFXvdEzKwrU4Z35FqprcvyqW4fBUy
XkkVZzeemiAD8j5sXUGkYXvRYM4y7uUcuRq79k1A1wPip3XSRs1DdxkcyGtaQceH
fjrdpK24g7OGqjxe4oI7HS97zXRrgem1lg8H8yj3OxI8GCLN3SnsPccNkDo6AV7K
f4dNctJUoVG9zQjcjMRC+kK+/8UfeTimTom/LtXU1Fk70ecZq6juKSjoU1fby5VK
FyKNxUP9/zLDHsYFp4ZJul9dJDJbLpzbleCnrgtbtm+RJoFW5lbi0KKDfsbYhZ+1
5j4EjNdwHQ1kRrtUYhqrBDIznaRPsb+nHnLXoi8Lr4afZ0goz4/yOM8j7iGW09yd
Vyoq0Tbssd/xkz2+tsnFAQlgisyCl5TT6zT66ItWCrOL08v7mJv9izEM7b3HRyXF
Ntvs3wKhXeFnw0L/2kw3LUWK8I7ErNhVh/Fd1775RynJ665vU+RSh6wMj2Dqx0Ip
7lFXTybUfeftZUNWwepfWJABDcdwZodj3vSEhId3zoZuB4wxYM0TP+Dfor5NCrak
CIWlM4b5OtpAeDQhASdiMiG69Ej+Nd/vNS0CZXoeTXmHR9ZNvKJdCLQQ/bYt/ojr
h4Zke4FK9RsSBQsr7+giTlj1PSPBDZwtgTMBZ8IinGL5tOh2fbCAFpforBwP+ofF
aP2NSfIjhSradh6BfpQN44jvg3ovFw48PP1CmD8RvRpx5GxiROGhkLlw+gk6zpMN
g1sWykYWvgLW7YzJofH2LngCYa5hnnt9Wsu6XPSRyDjeHRhom6Kp9VE+oBzIrw6B
7sWlM+aXatj1MESxthfEwAEn4Ook1BR5zopVBAjL3SozX2sQwC/cCxNz4Eoqk/FV
rc660ud7/SDN8uHjRZqZjdL8hn8pJDhXTBDoz9wuJRYZHJt2+08YucVoL50xzK16
n7jqoMmh8sP8OYItWieYER5UXw3kqg3I6k5Ict4K0tHod6IkCybHbrgPKDpa3PRl
FOJdRQH9wZt++Tp7lyaEtAzJjdkKjwlDB7SEREh1GSrW5cfcavrraG5ZQmMbd3mt
dBBuAvcpir1S/YmcYAZ46z09BySTYzoO38cAKAxzjCQsoSiZBR2yPv6xh56f2jgy
tDYJEoNN7xbUMAOep1mxxuAHJpOissxMvcixNpQMr5k2nnEnUgG1f5+XYjntMku5
QzBf4XcpnzMmam9bTYNvDYUUKAOyoFcr1SAVmzrR8joeUtZ7dFK3/zo8zGJ+PTh0
EK8U5URKSb1Q4+qCvy3WIM/IH+S5DBOSyaghfQZz6dJKHfmgauHL3+Vr4ivJaXBL
Ejjq+V3+K4T8RdiJ2u9MJoQXf3EqSm37czJkDXVd8YZzcGyt9/IFqlwR2Xrx9kW+
unId0rpZZgnV74STfkYeM8T9TqqNa61WO3U+ZZTI2eLDIrre8Pz5FRf5kViWZCy5
CHlTg5yX608Iy3JatYYPZ8+2ip5vgHpATbAFopRnQ+DJkBwmegmrDxzXEir8xHcT
RwySZoHecu2bnA4scOBtPRHgweENqbfekzm/rMCrmnxl6Jq5/CJ+AKlmHr1TgCfg
3TLdN8LGKf8SCXPnevKRwLiFmS/1rOd9NCsPjbFY+Jx1G2RIKOZQj/16p0mwqM2H
1uVpgTirps166RenfFRTL2B+kqCv2l5FbDOB/PyENSymGv5RWApRTy3IQhPCfuez
CoNBwGB2LMpHWEwn2KDjIa4r03goHnoDQe8tBlo1IesLRrzd0mDCLti6qnMZcIsL
bxhUbnhLGi5FLkZeRKL6AM3aU7ktpsJK+eAaekOzAOclYoBrM43vj2zqQBoVQx4Y
zvLlpXcFYca/pnwDhFiAx1GMycS0Y6rT1TYdreSvC/DJvE3iTzF5eawI8aXzOQ3+
ErXIrlnS6yYOfkgyxGM9C6qeS40xWO9G/7D4tgupb4JAm1iFXxE6HV371s3FDJdQ
pc1uNLsCgvHzfAYm29ko/b2kOajHZifX+4QIuzkYxE5x4BI/Hs0zRZWM4BauNVGY
oHRlZAEJpKBna0RDIuuT9ZF0itr26xbp7Iy7elHpqb31Uow6QCkaDAWg6Sth/l5b
YTwyk3jZy9RqW1FQJhpW61zqLR+NdGvZ7jIwGbDdT1/xgSep+I8tF3aIRS0QQFj9
4LtdDR3NdfjpnVdSEXj+n1vVG4nfyqmDh/n/jIODWrhXG30QNeV6L7v0gSVuW4ix
bHgkZZw+/ZS93rRhf4gfLRjDb8GMMlYIHYgxtv+bmqDp4KnJtUTsfVAJfc6j0uUE
LNK03dX/A+ezrCxPQRjMsZJ0UjqSPJXBxlZ1TeYJjuL4bGtuFDZDJo6FdXSZo2+i
Vue7gXjm6XCh+N0+0C9eNWLfqf0oIn/jOR7aB3kS8skHYRjTt0H7Kzw8hpBQc1v2
N5KoVD5k0SyVPpUCMmw6yYv5728NlNVHc58jnxOBnZ1OH4CI5UCuQi0VxsHHHonz
WsEkRsWvc+X18FgcO/02VgXjyCUBW5kQG2PBCvdH9eQ/z4d1nQuwLmBPE0EXdHTS
K+s8+OlXUwY0ZtOKYQx8gMBnWk7M4Ddiou7HO9178pGoeFgRvEQNdLkQ5MY8acTy
GjFH64XVpeeeZ7OCH2yH9yLibnPGrjA/orfZj/0vIwh2klqcWd628Vx4J8rYpOER
hcUVkYbQcU3uyc6kFz9i4+4sk5fmymLZbqaJNe90qCBQtODpyx2gCfcmDwCdIKY/
WZBsH7AbDAGK2BB9iU9mxxlBZqe3YzmYJqXEqSIGpww9lLADxzVup+72nPQhlvWF
6LiVO/zLJH4W4X6Jgrd05/e061oy/6yUjsF1DJRmnh8iA+3cnZ9WJAC9C4CXJPwY
w09GJnGH5nCxfjSuyxityDTB6xzQeuqIbIK8BYFgZbZDmvd0lGs4hT0sG39Lfzyg
rBN7j+uKiAbqvgjy7O088NKtf6ydXw+kiOvQiGeIf82J6wvrFqefL/vvL60C6SOz
5tH+iZcN4JCpSKIA/bLguEErBnizaeN4dm/Euiy5hCZcRhaNdH5ftuC1mO2UVHLz
A9ZpeE5pV44QH7wWFRAGOYI5YlbQMah3+WmYqkylS1XAxt87uRmzUGkvGLvVgY6n
WIPPqC6XERfdCBxQmGU8O684MSEcueS9ON11lI33wgxCuJODpSCFv/lpkjUxLG3o
7+JksRw1s08Neio6dgL5F2bM6Zs10lCNrvPt+8Kf9h0KUTiv469QjtELBaYLxNxH
q25WRXf9YlwWYPLKwqs32oyCDipkbDd8SskzRYAsUPYZ/VIbBdOELHq6uBkAZdBQ
tNUFkl4KEtdHxxv0qOyblTWhwT3+vadG1EZbMxbOjUe5np6K4u2O0MNdQ6jMiQFB
aWmssN1wPr+tC/xabUPAjWYoa2h+bwMqS5IQTg/ZkHFszvt+lk6V190nO+Po7W+I
2B6PsjKKkx89NetJ+R5xxljBEIhSxY7VPPFfwGxNMlY3gXa1GewtAy5wr79248NL
hISc3tRCwReCXir91qBxAT4xQDBsAR6Cs+zgmiE2y5Kf74TFDzqM/w4bHsq1Lw7O
/KE6uVA+W6bUGvVgMnetL2COh3NshqikvqrUMjqOx6Yv+n8AF7wk2XLFONUxctVx
LQm+PkuCQjnfiIBfGKc/38tZHC5HabSBXv6dnUj2+8EBW6jhdGZyNxF8tyrSVKV5
Mho7EzliZ2wy2hPbLwzb07PKqttzHewXA0uPYeMbe7qrfts8smyQRIhGihPUelrI
zUepJnBYBTHOD5RRGkJwAFJW7Kb0lgbHSAH8Eo5iKjALbLWaCS7/ZHh8ck4m/fxE
d2eVXylZyUV991f12uSvHRxskWPFAA9a9zTD4cj+gZyCg6rTx30cv1MANyILY04B
Ijrpm57q7qALUplr/qSSP+5+0law+lIkM7i6uGrxgEfhHWxBTljxFce/mVF3z8jl
chZNuUSpMNIptHdNUvzuKC1UOzC2pCahx1v9T7BWvtZobz+ebDEvI83n2Ybe8eAL
K45ep0aDwp6Gc2NtFq+8cp5lzEtRM2u1xqaC07v7SgdSCus1vLQCnp9Vrv2+DrbT
Hqlusi9tV/iQE0uIFtusBS2+gQFNLLrGUM24X+fK4NgP/UVmWD2n67SN4L7Pftb6
s+uS3szRyTyiBQKd+UUT/EfzPBdlN3/uWQWgrOLvwsHqt/FSt9bpv8eRYkpoQjJU
XnE/8KIHQgbJCcXmPJJbEY/F+Yxza+OarLOOt2wy2EMOMchYNorWQ0kMZ6guv+tW
YqjQbyIZWaj8LkuC3Tic8VF4+xlXrYZ98UzCKcscVzPw9poWth4baV0Vi+mBxEoT
rwmd+jUaKuDj2kA24XH19k3j4lktl9nt8rt+iR+rUdSHfUtvvZsQKmB3kgD7yVZX
Bm4BzNR2DxrbyeVSKn5H+r26GTuJxDyNRThgA+w1gKLflT8pLywXABKMKhuHAh6H
J0rQdw3CviqLGuoEDwUmRKoX8V/dwnOwjIfd5BQPjhuRBuT6KdqI68W6mF1lQHVc
jUV3ylXz1xjW9I3bdd9nImsDSQQAyNJqeIIUkybMYpHZp6xlL0iXG+WB18Wpe9Qs
YN6XommQxaqksa8FU5DXOYoU7CDT4f7qwK7c6bnR84Y=
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
ZSz6WlXvokuSMQdsvKNPxvgZi/JbKoTYnGkZx6fildcM8vfphh8t7I+Mqozk5D4sfk/aQkiWAIXI
3SlTIpu9eQBUNwl2goPm/K6m375iE8i5obdBefRPU6JIrxcMmxGbkMlAsjpgIQhBvYZ1ChDDp/oB
n4kFOdVLdhYLXlrhobvSYTqwP8ZHSdkB7nKobJ0KHqVZyOHhRWvhKAbg9gJ0qwyRIJ62l/6nstq0
c2xYfrKljjns/SHqHMHPL1kqLNCDyie3K6Yw4t84gdIUy7sOAmRq4fXEMSYhahzkfxqf3+i2nuiQ
75yHQXZ6gCmSJNkvWRC8u4PDC2VQv6MzVqDsPA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 12048)
Mg8sYzdmett3GIQUdpo0wAijpvhuoPh/kZPItO0kQZu9s5lSUfSUxD+KGWgge/7GLo7AO8VOOUnZ
p8fDksJxw1cJ4Lh1q+HRTjBmpBNidEHzrPLCo1YciKaz/fJx9/rzsZ4eLEz6XKkRywdj/RXpeCBj
owl5OZlE1lww9pMyn2akBEgD9D3EKf15IljLyWBgRlO5wEbS4joNZW3tMRcFHeEyIMMCZnusBV6Y
L5fvLrYtY4hhKn83Q4sKnQKpUlPb78V+SSm63uqSTNkDVrSDj7045Vvbh1xjip5upXIybcs+7nod
QyQsAmyBqvjqofGtnruLavX0NeLWC1aCvPqPwn5n4kBxFhKN7EpP3SwPeqoKWWgFy/C7SVa4yoxF
PMRJxW/rdC7+iXh1R0xN/ZvEcwgB04P0AsXIKfv8eMgFEdyTj7og5WVcZtSvKOuR5Zd4MJ0TjDGo
FSynPvx9PRpYbKcl5f6OJAl+Kvl+RBkn4cn4KuagBHHchwW2M6U6m8NAdi4d69XgfkRCOtMgUyV8
gzU9vD3QiQdc1kyFW7FaV21IwcZ3bws83WtG2GijQucuyCFiEp+WXzlJsY4Mv66fgn5H0pjd3/Sc
Oth3DeQ/k1Vzy10gJXFuZguWoOboOFHAwJ60pBDDdKpVNUWNhdVNgj+3KXL4ZGJ0cGFFblljmIcH
XFJHjFnHZJHtC124fOUNF6fsGKob55FeZzSh25IF8Xc2YLEWVGc5ueTO0U7s3wNa1Bpg78w/1CeD
zK+5LIXj7RG0MdVX1PTk43KWj48Pop2/XEzVrpEColJ1xZBatskK7s2DUrctFQXiPDKMAfO99hUY
CI3RdQvYSnPMnGWEzGUyJOgIw2ozr9s5Ytkn24VXbFAATFW4oi8XV6MkZuVFsuNk1ocjrLTWD6BI
hLM7YyTU6kjXpF5t2brwhPj/GhsTG/cwSLTcwFfraBVfQCPjinWMMb+l/v6Yu5vlcrZUaD6mTL+Z
WOVQfk7ujZoB8QbYAr3IzsLbdiVLAa8QEUHhF6+IlAnnWIZoODJZwPFBQNNZt3UhLgpXhRXdKU+w
cJcVlTrZM82vXXR+EHUueWKX/eVlNoGtk5Zr3s6ZslP5eepPodN6c1hlUyLIYUsb2UOCxLKTAPgp
FhBq2fKatvZ0cGS920FXYAysbN1gDvugOx2rOjFmG3zHT5WWHkYDVrnbuCJxs/BAwqBwqsriqqBz
Aet4jTIBAYnI8k+DY7chhyoLK82bwKn+8Mn/fbsjZDjeaorl1o6viM0wlS6iI1R9VTKbQkTbzHMl
ppsjGibryn2LWRiplGaM+naA5ypRXsnjmkiuk8Gm9jJZRrG6Myhv85yTs5JadPR96C92f/R++Yfv
sCLq+sdMFG3cI3dX9JIxXCfi/no8x6G/rJb2UU3MP44L7F4jfpTOctTCUTHmtSfc2JTO4/z5808+
1lfY0lHIiF9j2BqpkT2nRk6fFTcxF6XG9JEtGaehFrGN5E6TaXAj+bG8uGDet8wjd3P4nWpu6poT
h/2fp5UW2M0C3Jr86VlE64b8Pq8zhCuncdIkxypfMoIwi5ovI9Of9151HL9W2v1mmiY2NH/eei+e
+IntorR8DnuiZxVWQ4xDx+5ZS20RTFIf1TXn01wp9VT5X2MhuL5v1aGVLLtpc2YqP46or7tVKmFj
Y5+UJMeSat++UqD2iwA8h6Yx96KMGYSo9+TgT49NedAVDgoZ/IiAkpcextGVihFjSPjmwccyjmvO
owdQGK76tFVB9UvMDkN5iUXCkM5NJFvNAMXuEZKH0VxN2F6vzCVYRUdldlIlsHx0/CaeyL2CNzHN
2+i5k6Y9fcvUJVkTWMecgjN7GvZ8PaDYWV+5tdA056pBXMsnFOjlS7zM9HS9WBtvjDlEPVLSATeo
3sDnvUEHYQky19F38dRyGNbVGvM5PLfUaTQA07RwSpVbM7dDCmAn0kbpwkHTD6XkNnSzML0/3AQd
zL6sBRWotJ89tRFndXMfRrB4OcQTBZbwAb9dhBg9kb0rYuXs0Dl/5r8Sq3jAGd7es+2Kx9JoDGMi
EBRJYe7rSxP34WbjQWjGnw6SKlBm1NHhg39nwuw0NunwyClv29ZAxGfruq0vWPqAfxuIQjSPWVkz
ulbmpSMlwCPrQagre2jllLM6CYw40skyLc3TuGqO+acRN5MGSyRIVHp5+AaU/KAFBrtO5tn/YaSc
vZwNqF22BjgMal2O4DbaBGAJWmkfAr0LHRyw68wVpxBAs9H5/cD0ef3C9Da21UlpLnxaHa5ge8lU
U2DwCbw6u7kZfqdM6r6Ocku+R+TZ7dDBrIVMjnD2r7gxpo7AMUNdH63kmZrnScAjiM3Hee7uhJfX
+7G9bhNC+4dZT3WujkfnfgLEjuVSL1PchL1UVF1jvjCjGfvehYoWWVo2dRFQz18rnmA55LIiKOx6
/9qMnpEDQaIN33+V1uxpmT6pwmIKXPORC91cKkYQgU9yv9XTdgKrx23yVT6mdpNaUucHix2wXJmH
uHHtER5gvIQ/dQ48kwfAQvEemymGKhrfVw892zzZ4ACDTEkjeY60I0ekrRChYRX6P4hzidqx9NaB
GHe3xJRberJ5OXBHGAt8DqVy0fBL0VXNUd/o0EDH1tCTSbKjBrKP1TA6IJc5mRXH4bFs2iouZomC
hrhn38uPSQy3431pkLAnWyf+dw+IgWHOpTDwlTblGGo1xetRaRhwVpWCEzI202uxsYyv0rAAWECw
AYCYejNL2n9uUN5sVvyLXG35TlAP6HSQPO6PP75DRM/rCG7z0T4cLjPACpDUso5KvRnpduIWVa+U
WBXF78q1OvkTgpfxpxevKdIJRt0xTFejcLW9kgW6Dgt/rldw57N6/6913VnXwyrUE44mYpI7XUSI
Pq+Bt7F7T1MEa4Lp5wm11Vez1Px7LCXk4k6n2MuJ/PGPyTK+T6YHTBkz8Zdcc8lebOqC+DGbm5c4
000SnefwFAWh/qQrFbZtzLDUL6KLBAgRkTpbMHVaC2jDp+E3sz4qVuwwlRTddBXkoc3TKDlN103N
eGaW8Qm6Ad+E59KM/ccn9tXjOYCXwxfMRPcNAcdpBSjxlvffjl9f5PJHHALWRSpJJGY3PK7P7oFc
PQCwZMKBgKopV38ebxSrcDQDZ9cSmZegtI37otQJ9eQF8vQCPZd40mZcX2J69CHhXrHPWlu9zZlm
p5vtqou4zoWLNNj3qsXSzD2Q2Ur0J7xiOqpyXNRhBfaS8aXGrT1I1t70SQ+f/IbH4OAESGHNyz8a
JpRccMTaQLzQjsKKHDtGxpT3JadVEd6Cwxz4ebTIdrJgRtmLFR40C0aBl6e+r48mRoc6gzM3dJaX
cGEIoXIeWUwLBovRvidqrt8JoNr2PPQAZvvjCZVMXcsKpVU4+SZpNvmBafjTsl3xD1VM0o4UsUTO
JurCIz4D4WQz7o6If/WDrj9r2MhRBfx/eKKngkBQqFBtE8VerRPhACCXXSHPF4qP6kFV386IEpDI
Z106EebzDkzrRnH09pc1L4utCPGIsUAbnR0rc4u+xObUrIVcHNbx7+wJ8KrQdD4IqULh8/Peg2Um
BxViSiS/n2QFaq2FcU32jrmZmKtB9UA3b4ZWyBsKNauSzFMdxUPC4x99kI8cSaaRMApTelvlzSae
kf05HpYDV26bFb83ZKAUXuw0XWMXkWBSzaRZLglISTg1hqUawqM8v9rAb+NrSvrkg4wMGt14cMbC
LISQkAN6HruaPFdKG+8ninw47ZWQ8NGj6b5QeHyn5kQcFPYfdELzjibdoKexZVih9GOST0WKQ7v2
UCJqLbBgXMkTYQkv5WaReVayjR9bSmbl9byF/Of9UxDwBqhye2MZGLfyZAoN6xYwrpCIdLGHe0Mp
0PREx3fKRz3BFsM5YI6IQL59Dr1/HV2GslVXQ2kH5ze/ziwS1vKoirYIOVxHBarw1IBt3li4HEU0
ZLr6pv1zA328zRGvXG3jkjG0j/ce2f6nl7XKPr7mCSCMSajBh1xR6l4T6XmYt3+KZhQ4XxugM/bN
2p9DEPDdYFQX7twMt/qxQh1+QAyclCZ78QatG+D5Bj1bdqf99aCvr4DR4ngRAgXfWFKTA2M9XxVc
rC7rOkChRUeUhNgupitaB8/m7+xmdhs23JuHDhm9lubzKXH35sGPGb3kJTJmgb2hUOaEDyYeBGkP
MBANh9pmB+1+KGR8PBEFuq4iJ+TDBQvT+g69ul686ZLozVFxDLiRdDOspem4eO+eEkVAX5BwZaLW
2O0uiA7xTtURVc/wS8hileJK+Syt7BaCOTDF09Uy8kKoMRKaJ1RRS7wNxQpnSS7PkRooLyTHji1E
trZr0AMKBeP0LDnJ7QC3HdAme0eWjIV3zZ5qMFTTpPBMPrJwja/RQ2B4vQNM0lttiYljdqpz8ryV
ckXWLn8IfG9jo4SbCpIVri2RNMfgTK1aEn0yVPYHXmkOwUf7fUSNiu+mnqnYX6P9F4Z6wb4jNYeF
r9plgbCryotTavfXUEvcxdFVJBMRweDkBKOIc5E5K+FaFIanNpCsM/pttKOyspNFk1HeVOi1UfcN
a+azTA13VMrfWvdrWFgo4MPFvRHAR4CL0siugVT0Ob4rVNgqTGFkWeuAmXC2o2MePYyBLdSeCnKJ
YWBxJ6RR3b7QetJAPTQHpkBL1OHT7F9DeEEeU8sqcBCHEWh9PpDy7y6NlGN2FRtEaNK8In+0vc/i
5j0YFXrph4rDqMNDeBprVNi6QY8FV+chDY8rcvzIWO6Dz73x2+IKvz9IFK7JBc/1zYYgbwaYCOrH
Hee48Qkn8IzdOH3eMEt3d0BOBVR2UJ/OY/PoX+/6ot5KM0fft10JGLUf1iugzgSFib4ixo5IrkQM
ntkovf6MSbxdJHqpCh9CiF0ZxmcaSrkg95pYfTbrmESK3F8IwKovzpuZuudiVv325sgaDZCuo/3q
hqi9kXuah1gfdBe4rqqYHEvJyh0UaHSTD17KH2VvRPDJfeuO633qmhYWEPxUyrxNAlMZfVvZGPYc
umSkzS/HHCfFq39Qb3C/T8f074hS87BZhGFxag6jammpX9/NlG+vZ+YVZ9Bg+YkrtEbT6A2KigQi
XXPb9Jf4YuYsysoEChkwwbi+6scMAbSSeGpEMu6PAd+F/Q8gMkS6f+VvCf0dZUrbV+WddpsLr5cD
wm6UwZbIv2ZZmpmMruBHcF+NQU012xyCeex2qHlevAaJKTMbhWoleh3GTsTy8Ieftj1ymugSKi0m
Bv/WfGi28Kl+/Ja5ngjKKSLCwQdg6FFDavoy9sn7gMRBbJJAe6+VIZabipc3O7SHo70d2OzSr5lR
GJAWjyilgSEElItDnmBYwHFMtoumsWMuYB23c8S1vVtMDWDedPDzzcWWEAqu2CCipM9y6TBuDPxg
bQzd0OrYrhTKWWBoFdzJ9gezLC6aAjhyrd+BLLYSQn6RY4VFvIVx+XC/4VOGtXpRq4vcfl6xXAH+
azRewqW0Ov9cUQhtM4eSafqOGn5Qli+/UCvQNv1bh+b3urx3L6xorcRhn6nKurdiCb6pnOSjdoBQ
OpiiBLC7aIcwRu/myTwALzVSuGUz9+VpgU3xFlFMyyixqK0++N9tI4Cjyf7vRnUXNPgrD8FIidOh
3yTPQQ/ECN0FYLDcyLZQiY7fa/bZh9gTXtHLFU6L41HWdP/aMIM9rkZJl1JtfvHFKjzASxqbSsQD
IjpoclevZQ74DO8QbmoNO3T58gajYRbMYFkEzPUFlBybw3iw/snl2tRjJrdYvJCEeeefyp209LPt
DpH/8aDFFxUdZvqDex4nhYGZOzYuoxMrv9YlzGW2DT/lH+FZZNh54F2HxJpyUTsYMPbKIonqSnBO
rVWt4aSye9QBiOnYTdXM8LbXG7uhZvobNVKI/FBlm9VAJaZJxzsBhr83QV3N9fuB9g6uqgR+g8fd
HdVp6Pe4pIuDfb9EGcIrJSSeohXL5f25YfO03vLBxUlO6Un3/f1psLtZtcexqkUQ59xpWe2c4Upa
rw4O3tHXeW/XcAufwUYlRrg3Z5xTzB7D2lzgOSv1g82y+1+Q7orSDmm9pM0z2CvTVPBEXQSjHwr7
9bvS7yiGftpNDhnOHMb53s3Y3z0EGpTk2ITCKVp6Ah+A2V9q8YRC4r7MNDWxkZgsMJLzHG3i3rFr
zsV1UA5b2WrwUp/nDxRK+YCQqWVVYY+RLES1MyWYAKHx/rqul6o9VRPgwUuG9DOs2RKzaDCEWBBR
oyGUDSGP193nrSj/kn/x4VbHr+iU9mWuOECvovR7m5xH4u3nvYX58SG3njIqQtvLUHKLEnWza79n
1iHD7B4b+kvW7ZjfxVWup1jXa9KP1mQCcrWmJ6LH+yga5PjHiCG7XfhmxFYMo9QB+nkIgBkdasYV
WIRsbF5B4WhNgyK5VB8qIg4Ee89EVMsr00Ojmo4BFZqQxSPPVy113Khju7Tdu9hKfqaaeFu0VKOc
4fQ9icEmoCDADKMvtyHlckUG8P3HneH1Vec8dt/HCG+W/e2GDVtjsjfptrFdiTDy4KakmX3wlVd8
W4wRQTmsjQ62NAScWx7kQx4qyDl8CgrnNn1r98oSllMXXzLmpAtfa0P8W/c19wq1whKqG/jJlivd
iVZHbxzbso3HIekIyhF5UhyKA6wTeLexqACL1YCkERqRQl5hZcEOfE1gCZGzf58A7vGYE1XwT+N4
E37ipvfOJYhV1LUA3czEKR6Fl16uUkpp5TfnrBFLbZajivMzJaoPdHOU37GmMK0vdVQGXD+CvLiG
Do8raAzwZrbVgyL850bwihnQ+709CEDy5MXd2pdDtcqU+ZHJZ+YyHVUKd7Miqz6qQ22sn0JBaySc
xA5AehN4ATZmyWGAv7Q7sGUH8DevjAgNqO41NTIgNNZ0jGHXLlYOOViQPE9rsDHwclEhwv/TKOSs
CdHGfjw917BXlZeuACsp4TmQRVrllZH+O0HjJeMME/3GlJm/EGsAG5zqtq1sHMw2af9HdbXqi+Sy
o+ex5NNCUTKkd/tuod4DvGlZE5EONcvzDzuLCA5SHa9vIFMb07E3jnPIIrNEFHQxvshCWOOvGqAa
HaM9YbzfTh7k92mS1qQjK2Gsk2EWaWlOKY/FhezRKQkSUrulLOrfQaqt9ZW8vZjJIQme/Qjy5a2z
LHIGvSkBQcEgP+v7/pB6TY+lxR1xsJg6RUwUh5dVPrVho4YvSxOoW94tD5RbCjjjaYjaQjVwAnQp
tDY6m8txPRX1Dx+aJYtiXSTxuxmYDk7ED8jyejmSlImQXUAJ5OA6mrSh+LtZ4ghtU8fbShCpFoCj
T7/HDZDSCouMXFLFGbE26AkzpES44WWV/V0yXyomRNO1hHnMkYFVTM+VPqT/QgwUrHYNHW4QCJQk
gLd0BG9Y4balBRt5SRDZu+MSZe/+EKn/1y5HeLPMR2xtUZY+lV7Sroyn+5mSSwe7Q9qumJ/tJ2CX
mAJRv16PFyn4+k4kRJF/EKQQAzlLTuCvkJobdR778pl3A92qDvetHhgWy+1ucuc42xaM8p3jPnT3
s4GXXYkG06c3n1KwMRDc6o45Ci/0plJUkIOtBZCp9fgKInJwFWNUiUxelMnwet2hNqQ650yIV5qV
LbPTz10U7OMSuZbk6n+HWI7uez8+qa2At+EhDOyogfk0JenZ6xI20s4Q1EE0JZ0CL+70iFcxLX3U
D7CJUzG+y01dBAhAr+P7RbPU+vwfB5L+mORabOr6XfWlFmNmrDYoV2vmbssDfDGTTfAUlJB4qeZF
s+qucrlTKJkhJKciXTBMRwC3T8fAsU3fJrijwWyxZ8bURhA0il7ae1DJX2MSrb/5xg75AGEj8fxM
7pYjoO704e3LLOnkwEWHHfGHBmf1jHhArMfJRcYSrCT079Rm6Rnd9GFwKuHPO/ADt1jmTGvRgR9W
FghcWDaK4u7AChu1Pf/IKph93rxYcObydbQlHtzqQl5nry+CfYNFg0xDiXAc6s0XjkzV4V74n3ay
MKif6jAMrg/wyodW4HnW8QAqRxSXx0K3dUcubWJLPQEmShNxTm75zfZhJgbdwdf/0LJT2kZXnrbv
kqGqhSk/2hoa2UWhLv7II7HEBlLcObiqu9nQbGDE1d3B9NMbywUhLzuDc2vt74WG0mfAl1mkNGd3
ur9z5cUNf8IM0hZb0AcG1c8Oq8tqXO3I00sDFv//xzbnV6290zJ8anoH+X0y1JZ49PWuxLtha64N
0tbQB4MvI0tWoEUUcunrALzm5OlLMzUp5eN0qAUcZjdKsCIxUq6BFoDoaRyaBsboys7KZEJWz1K9
nnPKtnNtz0PA0wCnXjrdJiTpgvSTMnqPyKHDQtqyZ1EtiGUR1EN8PpJ63H0g5He6GhmpKkhLix+j
170AhZEF93nA96HCmp3rrsh32t5GtHaVA7g9JUArxQjUYRXSdBmrSDcGhTlYpzpz3rq39JlQw/Nt
z0dSEa0qKH8ykJeEnpN1MviMKn/gWhPcshjNIKPkDpeiPz5fWkOZOkIzcicd8AYNmgO/vlRsr/54
AuHcKGGbY+CDV8mFGSbkXfPgy8rSGPXsC9HxXkEDmmyeV/u233Xa+A3FUsqAiwUyU4yKHVlkXSxg
mCkI0MVoFQEOF9uaigFj+gsBQhHpCoC8K/QIgwfmdtUDHtvmGDGJe1fEQWwrSPISFmPetYdO6g4b
SSrDysHK7r0K4zKBXMuAan7IqAqubYxWNl/ukb9LLml1xr7g/AwKLkBl7qHVs3gOU1n7mSL6KEGB
PkjALgvYX+jaklAF8DCB6LU0nL5gpqB/Y+fZfl7B98Gijhg5D8FDUivF46/l5B74WZoSOIp5Lz8f
uyc1eyTv4l9j6oIMrVm4tkq1gwcM1pn/Bcg3PIaml367uHKnojLtJjTNB6LS0XvR4yz0JM/dRT+j
HQQyWQ9balXhBNa8WjH8miLnGz0WH7zP8sWwndmJJW65lvn9nfrgqS4CySEcxad27ytfeNaHf/AB
bnwdqyvVX0Tbn1T7ZLpfIiAdkJy9fYi3mdw6Otr0uJaNDwpKsPSoji9Z0wml7zU+xoYoJcZYLKUK
oAGFGd4ZWpIFzkflr+sMi/9cT5gxVSfDp3pzy04g80MpIP3j/xiaMJ79Jt5xWCy+vWiUdQFeFDAT
M5ytgxlIShEIvHZS/fujGqqeZurn6b12TdwrwNsmukP2qHQeRTCIy3J42f033hfzJnRvWh0zz7nd
x1wsnEzQzpwug+AyfyVOYgyytw3o2l0Yf1BahEccFyICPEm1EtRvoKqEYrxlw4+2OEwFbcYPxw+Y
B4u3vqjOBqueZXqLLDyVdqdHh5bCHvIcAI9IHxuTqCZo/tUCEcJf3+WpKb6ACnwCBZ6bua99aba8
14/uKiUpd+xSVi0DOcqPK8rik1dGLjcQlXik+MoWfYzf4bQy5stIk2aIWPkQ98YRxiolH9hffeMq
B++WaP4ZQWjeTFU7MnnTUUtiIx0hcJtNbxihyCRmw8hNPNRN9YXNyCxFUJqwBHIQIZMqXUQa1ILU
c+/7JZZTxaGhWmu5t0tEomYSErMUKZlkE+Biy5IRf+DYXdPi8tEqo9tG2V4eFcSNJVw7Ht5pIBl9
iKm3EAPhYnE6jY6lhA1AzoOGJIUzmssLWs7VtNzfp9xIW/TwvZSFjY3NIkbU6StAvuK/+CKaRNoJ
SGSyviC0WiJ37HIJ0PbfcfndT5/hv0UDiNSgucPbzeSq76QqaDbTSBtES6jWwBmDiu0n73Jv5ehX
TVSIKyX3v2czoNX2Ql0goWNxoD0IzkVdw9XYhqMsQJ0xoDmee2puujOndlc3mFA+/6CxfjCL8FyZ
fn2RL3IYCCsQJb3rKvDt5/TJ4Ncr89jW87Nt+QvcO3SZsP2iGrBS1sOYfEyubs69LRmh6DwkEINp
odnBrQU70d+dSqKNW9RENSxUna/7fJgj+u/618r6XkrEaGGeKH8U9RyGRN/FLrBLsi/GqgCPIV1L
yPE4VeoqtGNnTQzN9tVkysO/a75D4fCR93BrG5Qvx2bl+Pf2d/TR5tdnxsWIACjt1xDIjUOs1J0G
nCb90azJ/b23wprLYMyFbrValvZiDButBF5FnOYDeKoDAL6zCm2g1jpx6uo4OVBRbSQoLBoF899z
URF57mAICtSjPtQhnDxASpxopO9TR3HRNpZYzNZrwnJNRC0OMtw8bJUht4c2osbpneQp5ruLh08H
QCZERgFJdz6xWvyxhe+ZWSmBP848kD9tyuDcOoln81r0zc8xTKJ1ApssDJjW/RvwHYWbo1wFUQqK
fcmHpEs5sFjdeOtIZFUdN6GZAby957Jy8jhX5AtbnhRUL87QXqljoX3YNvOtszLw/vQhESrqczDa
sNEcEsS0Ya5k4od8I9r8ob9tLaM48OKX8D4mJF9QDJ3YjMB8b8A1j5VUFKkk+InbDflvSm/oUaA3
Sw5zP56Mr4JmX3CXI8cMa4WngkBQ7HxCF0a0B5/Q6nS8HzH8fzzSdew7YzsHJ9rXid+ZiwqBMHLf
dLH0btLrv7eZyQeuDa3lDie/RGPSELtyX+l9Jkz3T97zwwFxWLzyQ/VhwnrVGXiRrYZilDyV/M1H
Hoo2Nh5ynGnD0ErN9h0vLcIfVWJRfqnRk0TTfmEUvy1JyRcM+x0UXT0MUy7Nd1YXC6wecMLRAH2r
25j16lPCNvm9BE9UTl4N7qb+shkFEJshJHYH5kjuNLPmS5BbayTw+28VsBdtAjy6e3qQZHPAZdQj
o2LxhC4JYj2lfAStiF6NNXAgH1VWWlOj9xQh/AKrK0m1g2HeSDtPUWHQcb0yVlPwL3BWWN0jikr/
1ivGplp/7zOit3f8Lqk3FMEq8BMGsHU75oFI21M/lqzHDJDF67e8Xyga2KHv5BksA2UvOrMvCdV6
d08TWBZ4/KxwgNoZ7iMVQahigwedig6Dxt9PsxXJApF3WlXHtTTgrCMLNYOZlEc1IjtP1gonC7re
Rn56yInxvuV5vvUwq/wjom67nqcuNqvsEZFbAiW4+gZQgH1yBJY0vdZH+oEHfkBR4rW9+n047RkJ
A/e4qkV6V1V2GBIN44wBqnFX97+nztEtg1WRMK2kaWCMH+aQzDeuLVfoTqae+sCtFzlgE+1qQLOp
aEqGDLFGq4H4Msv8c5Ks+FrzDYn+NYAdYADnrD0yjelftPjITYwcrmFF0J5K8NRKBCm6PnyLISEv
VsdozNiThlAYywD1aUTTWHwphFRja5e9G6EBYz9GqcaJrG4mPm0z8FAO+iV2BaBzeeX7PFDjHO5X
PHRwQ0oNumLEA1dOR7WCQocDRydNl6htcvZctuysz630tHTq39z1PyzjcvQyhnFJs0fPqDVDxBOB
WJGko0aR+41KSs8TY4CH06zpqblry5zYdSe+ZzPmnwxmuxzlBzf4I+QN1o6bQcA1BhnKsnxd/iJ7
vjkKCOIbQMoWylhMr/FuDL9TvB84B2ggBgU/DqaG/zlqrRl4ZoCd7p6fXI8Vh5Bg302/dp0pu/fJ
p2/Z0SfZ1VVLE2GUaNJB3ywil44OR/sVFljzVGyUyXgHOWobICL9dykSexYmhm3bbwj2Nga29n0m
eQrrh5D+QzcOLBj7TyHSUVq/GpLoVw/CmsJQvup1F/e/b7CVV9xg6OCUCFr3B4QSPKWHn52hqMqg
JqmsqEa9SOEeA+eFCzxiB8J0zjNdcShVcXBSbC8AzG4tbMDkpdxIDtHVlXA+JBml7r0B5W/7Jq5W
t2sQnxExeHtih0KKFtbT6Y1SN7Vr/aHkdMAzuvL16++k6cq8MLLrUrmuqY95MjBWRxpn9d1Fchhi
Rsdh+iTKZQcK/iaAbMJ7Qf6lh6ssdmgO3PLVM9loI2gQUxZmHxQDd3/cmMO7aRvGe4VDKEBQVFJ0
cIs43wIogveME2+obAZEd6/t9XIR5iZ363MQo9R84kncMFQni1ktlWvYp3+PUlmwbgISWPetAmhB
pHzBBbjFpU8qQUeN9WOYNUnJsD3dgm5f0RF4xEg0qFESgFznZJekGB8O8WVniaHH1BhT1c5oGFsb
Zl2rJGupC0QK2J8wExNgV1sv9SBmA2Zp+GLtQA40O8QyEr0u0oNL/hELxsv1OouqZv95LmZt5LSF
mwrx0AN9GjJy5z1C7NUL1tn3YAHMqgos2V4PF5FN6/G0uqykieO67xKhdXjo7vplOXgN1LeDLm+m
N4sIDsb8xDG7nNBda8TzAr/EE5p5pIBb6Rrik4mhbXzA2jdDfvbAv8B29NEjkbEcsDOc+LcZQVmz
2afWDulz89iCL0KmFqE9BouXyrJnLUhbDGKUQjUrPnMBHbwk6HS8XreX1kp6ADu6kGyu+moSW/QA
A0KauqmLFxHjZe13XiCCiDtUNnZgUuWfhmVTL2WfAQAlHiN35D4kCQsJ6a6o77o92YjmfEHY78L6
MV2jV8QOCos4i+X3ObRe4WuZ+tO469afZKfewfsakwJaghAv8jASX5yfGI1wR/6e+vbyQFtNS6aU
oY1SBXe7miZbn58ruXP+Nyh/xbY/35nyC/sYORXkscJOEMoVauCKTPCwwGJXyJrcuS1oToY7iMrW
xAHXWve9Nn7TgN/EM4EQZO4LKWYPLOeHF06c8xdZuQKMcP0oV25zwvq/fm3NLJIPvKSiPTEwVoJt
MyxVJm8SEnRj2pQJLPe9qncs+jqBL3Jw3h0s+0Y5EIZ2tn1VRmmkDDlu8ZtzZ0Zqkmm6m/5IHLIF
3ZWeCaCC77ivE2y5GXSqrw+ccd13PLU/9GcMQgPMQVx0a9f+Zc8tgsOUkTtvi+XaOrylzx37J556
MTJQYyKZSql8spmITeIsoUsk9qcRjUMngtFq+dSnTGfB97eAJRanVTUFw4b0N10pw0c1l52SbqEW
srg8ujRZQUdqmCQYCRjjKgMfssa283BNFRpkjk9O4RGpZgb5c8cWz4KSx4lMKCcCIEhKfwcWLcf6
4ap1I2VQjHSZyEKaIGakqp4XjvHzgp+Hg+5KZpYLRuPPaQ2Wj10fwaxNDRPPqNBWQjdRxlNmf0V9
GaXQD5advg8+O7Dz7NOs1YTgOUEksQXY0n3oe3Ng7tycPEnLuGzQipUWjbvBwpQfrMCJzcgvrajV
dDfSC7nn/34vM6bBtF3gE9X2cNraHfdCvnEcnyP9h6QzmPhxdH/VHGkZw9A4jDfx6QNiGVRkTkuW
6Ze3mlqlmjuCINTgvC4DOh6YixdC1+3HZ1pvWVP98MUiFqN4VLrC4LS3CkMIHvlZWS/BaQiIxWOE
XwznOsw+TqCuIIKUc0XCqIJ1Wi2t7aMmscRqDXW1twU5X920Gw+n8iyRWSBVPMqX+ikkjywimtBV
2543YN/+Pl7ssivLCNWJSmSaDX0s3u7tM2Zgd0Js1zWpGBtsHCeJa0X7DAAKr6wwUvf65sCI5BK+
2aanDCCyJ4BSHrdSh5fhjynD/0yBw18EuRazbVQfJ35k6s90DpUt4qyKvUI++/18wW5DnP5hBT5U
1k5TP2lHxk0sZGvIUtMf7WVFmKB7NZ8L6RMuBXMoG6e8nvU3VSU+uUnMPD5MU1GLz3GvRZfQOTho
BOoatT6DnpPldt6kOCG4O8OP5lpw6LEnYR3dSloBfy/zdnMA07f/WfwP6WG6VAoV32RdSDzyD9gt
4qjC28Rnm8xDrk0+qx9xa22h2sW4EH1j2SqaA8fSOb+gDeLdufV+c7h742o9F/TVQCo7us2nMQNo
nNauqyVhbHhzK+DT1TtIfUOzSPKiqrxReTXcvvP3VbCMmm+pgJY6Xv/OgXsQUlygN9ylNOTCHB4h
Dw88P4LVb4PUU7CPZe3JmJyVfIqJrDPZsOkPL3/tG5G+ExHp5/KJ3Cfs99rJX9rDV3v61VdUd7Ev
ozQHwFNp1+/65JOC6ACp2uOKq9ow3c6k//S1ECRC3+ODp3QBg7Hc+ugGbsK2nDyydAjZIl3AX44H
s5eMRxm+l9eDmI4/ldtbO5WnkwHRDAacbzfGW0HuDaH/aNi4nslwbPF4+RRjj9aL5uXo9hraa5mz
uF8U8RgvE5w5hY46yRwiVaToSkEsyq8YhRyEYH8FUPea13jiNRzNshS8LJOnz63fH/on1F9kJYN/
HzsFDYs3FCzp72QxXrcrK3O9aWGtHd7DAskc/29HIFXuar3osHhiQfTYGleCMIIrQnsJl2Y9LHjd
DtJqTWVadFLPIYNKQ1KVtPaGq54SauOfDeAFvmflswvFgQxE+n3748w61yIuJrj+YYSFRguerLMl
POseqSbP/xOJcvvSGTXht+OMMVLwbt8ZvsTgBZzQ8mnAOe635Urug+SKbDHiSp1FalxCPCboP8Cs
+R3L0FtLj6UyGnv8hwfb+EaBI5oSzXEq4hPsukbZoZWAK/TFBRbKYpZ1t4dV4xE5ifvWkl1/2HbK
eEIbjBr/jQukd6hODqnbctlZjJKJXaTTHCLMJuQeNnB/O0PqwQR8MD+KTcDCr5ALoNJl2CqerOco
esxkZyv9TWVD18uTCCZF7HcxTs7Zvrs6i9HUouiJmvuSNCi2JV0Q4P7vZmJjIfWk1fSx2oQOWuIN
Axmxd/MEKoHdEGN9joS7lyXuk4zpb4DgTjTA/olFF9ZO5wS7Wb9v7Rk4T0B/i6Kn+Kls4gRta9Q8
XCNBRAopN6pcJlnS+CxITEE9XG9uaBsqlP18eBUPTWaE6ChcP8KyjWr0UcCQXCZi8RTzGHShNT2X
00soBvVlZAPyq1tB0VkAnKpBvI3KJi921ZthgB58z8f/knFAQBFx7Tvfz1CrvT7J9ez4ovYlVHkV
xSeMxBhRy78QOvZ5+M0K1G/noWYAPEJjl4k9d/IueSBYAE30vdhSJwjW9svyuFtGHCKvOiPYSHDM
w1CmREUYuuUxRrbusYVrlsQ3ULqqoCXULGKSzXmwOhEVVmAowP0O8KLWt0tvB5tqQ6NdAljZagxA
Kg+u0tphiMUbPV5k3hF3wJuYAj6ZF+BTgZO0FrOI8I5hOuOE53SVTRqHD+uN56auyJj1XflHKttM
pvz4SBnRb1Yl6DrfUDPF/bZcDcHGBbN0P/0NRmy6KCT5UJgAmj6TsT6XVVjbyTnXtQLGhYQC6M+A
NPlFm0SXjTw0I37iBVKW5+qlHE3wxRjTIEKKuFfEcMNz24L3gS52MCcLm6yOs+7iFe9eIkrq/MeR
cD7RdPQyH109rlgSQUmWCTeXUXCf9MOhk4JWysKGaVnGOpbPqILRHepjkTtOPFdzaNiPNLcmBHFE
g4YCO9BeoGV0+keZP3MVNZ1vfatmGU8coyOoOJeY1EaMqDsGbN1QOg9SFr24EVbF+5zw0hqaXzs0
1fVcKEgJ+qp+TLZTV6ncqIJxp9emdfL32Xic8PABcFWaVrusCCloTDyrMj4a4RZvu0EBEs+ERKWr
Puu5bYZX7UlUGaCgWT41zh/6HY9PcNiUyPOek5Yt7vMx2/gzAxJSakkJj1pE1r5tyjtUge/A2nZb
fHC6gYntFOTQRzGbHL4NoaebDoxGq8LNiIhSHxGoHhgIFm+TY13qG4DLQTAeofUwhaSY+/Q9l02x
ZRb9Z5Uf1G6olTmaRlYtZEQcT+BU93jpW/potyk7P+Gewx8e67HwJdLpE4eXuRT5AHRz7kDfmDFA
zxDVO8k4+yX/wmROvVOGtuANO/pGjz4BpprG7AvKC4ynd3dLK2luKumDKDjOykDxNnCiup4l/hsE
6jZgHw84ByC0w3uI2ONBII3lUkFi+BtrK1B85yHPFToNXfZSJi0hroJn9y12JHt7J+ZCDZlDrpDn
UP/QpGQQJ1m0bqDCFCUAouw8kqj85DMmkeNDlxqAHGHOin6la+T9SxRVYXHnmDmq/+w3Zb3S9CFt
NabnUcs2Nc1p5Pt6kEK6u6Qm5zWnMe/9rV7UiBqrPL956N3pjTx+cwZS/bLsFTuTfeJuQQOr2UbE
Ew5unXH+oDbXl9yOIZcFuyh6uPZiZJQJNPUU1Xa5sYRGsHuxXUc6Y48XENWSBWrnl+6MLclhaeZ0
6p8POb3Sl9w8oPcGoNkV2z+msUfT1jPgoXhEnZIJrqWBP8Mj+QVWw8903/BBq/xZIHULmbnoAElP
+rzTd2o+Rr7+7e46eDKYAHBS+b/B
`pragma protect end_protected

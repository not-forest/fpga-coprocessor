`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ifuRooJxPH6qnRzNHXrpi/loCvqNJQETHHSXAdAL5jEX/jQKoxk0+bvGNRU2ABiC
2nYfwaaJQJ/rDpHJOBmBKbpiL8K9iSsdgkSuutyedqvW3jLgb9b3STeh2Mu6dCxF
LK8NTb/tkZzNLDpHMLgLibYcsiSjZ1cLwz3x4jnVWnI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14448)
RKYPUSKme2D2tUa8g29adOCFau/o8I3a5svwOnIQ3ZH8K2HOsx4rmQ8MF3VfPld1
47DCYS2/xFCTIbtt5d0CL2jIE1XdA4T4T6QMHreIRYSZrr4tMSAtBjQjQiHLQgzU
nFwaXpYllVU1CpZihJyuQtelr3I+m1hua1TjaiAsZ5djcdg/elLyd3j7PN1IaBpD
V1aexMqPImxMdLjMSXM6OcD9phsLEagvCG5nr6xgBbR+mW3DY8wa0fhjdUxOMFvj
Wprj2Jr0rtkz6WqaqhbDn05coUpiWDvVvNxDVOXhg+cpkO+2tc4fOEpCKXMPHRV8
BN9XAsqkQFqlUJVRFPE7Fnu2gzs1qQdXAgXDoGj+hMk9G0ZuSxYry0+xAGi5np6N
J8Z85mofcF/wTPPiou02e1kQp638axCE59xNqjybTXV7Gur3F2NXzQGKw2nYh2SI
skEPuJQ4TZhaJUl1PKRsPhOMgOTFvmQw82kW48wOEZAanwMnewTOV2pmTn4uyI0h
gaFDroLrt3DEh8/CRRkslkJD0rucpXSPiDkrb4Yd6mgu+o89h+FcE8TJjj6P8QVY
IrHsQBfPC/q4Q1O26GDPTVst/LFGqB1YNKGFmNsLJ2+lnmxEMtrfk1mzGml3WoBA
A9aoisbIuCMyARk3LbhlxPKtJk7ktFyA1eKxvbnAsrrmiwZZTC46tOVR7cp95Ibb
1srlaARdjW4tUk/Axme7orWjiwv2LKmhkyr6tcV38sFUyB8phC/ooGgck57BPl09
WJDDKJXcjkdytRl1Ea9Qx641SNOfsfuwOztrnoCz5s6bcyG2YJfSuri25e47frwY
stYZjnxQ45HVPH/6qhnOjNBwcstGYxwWKc8kGBuq88rM/6Ya5F4WTEKUPQ5psFgd
b7DbVqIRArpHuJD8uGvR6aHhMO9EWpyknJW5qmzrqyJwBcXvdkgDpLkY0CUNRLsm
f6ofP/kRcA13d1U9Z9U8/pSxe/oM8Z3g6bO4raLhQ/1Eu09vNmZiHsgMjhGdOj/+
7dSD4mi3LNT5M953fZebERQCt5QnnCJhF4ku+27Q/slcDRcwwkNCfiOwZaBuCA6L
tCfpHClqlt0Ke7J3OLOF6wmRjNtX94VbX4SKgcZ2OAHhMd2JjZGMQHDTPWA6v3gq
o1uOrK6EHRoJFFSdm/9gI6atn4f8giIZQLTm8wauVtJVJMFg7J4U+UTbH4Wbrd7M
UR0Qt14kXbrA0qUFVSavoW/5XJjo9zPQIqqIayIIODs6qa/Y3zo5macvL1JSbyu2
709eeSO4GQM6MtpYi9Peor6jGjTdecNzUGLzStjFk+gR9xp/Lhlu09lDgZPOJzhx
9zYpXwyvVRY1fJzNaJEaidMWoEPMb3VohNe0GM5+SS/uGhRzK3p7iLjQe64f3ifd
f+gKlRzcjZ87okQXSOUquh+w0KFAQ/M9qmNad487Qad7Gll+1i3N6plxEofKMzoO
DIZdybCVmbp1AfsfLQT5glwDfZOCXQYwKgNJxhWtA0eq7OEh2U2WFSQP5ud9kBzq
yMF5FCaJ02KjPHbyT8fUzOHRALzgV8LyPSDPJWKMu+FF1jbP/v3VseW+NL/OiYcb
xaoSN6rNRebiNxfA8bkes/5G7fOnpTdhJribVQltGFA1hGPUen2Pvbs5X9uldd6U
zRUmBsmon4Ojl7NEjFB98nzsFgbpSSrUmNbv3FV6DcbBdB7zmfOh5dcphMdLeJL6
IZzSkSvKTFbbP/yY7b3AMUO9OPk6S9Ft7YEaWfj2pJkvLgFnseVNTEGYLEVjstw8
5X1vU/kcHW10NcB3Pf97YtnwgJZsi5EfZvbiin7HFU07CNlUfZTo9VPzxCRRP1+S
oTvVwT8BhgJ4HEvRy9SPbtF1ZkbrpJsDRFSImw2qjp0D8x/cuy1Akw7Rhw5WSzIG
FgPR43HhL6GQlDS5EYlvXRb1h5vejhv1KbVtFhqwNZGgZXGjRBXoA5xEnoO3dyu8
jbXWnvLnlI3om1E/okiUfojZkxvpVK71Q0I3xDP6S0nRKudKubsvm9vo1yhV8nS/
Hvg/AW/CA4pXvryTxVlk/SuUuakCrSGuB/4L4THxERmg+rABcxEJJnQUQ69QnBHh
cHqvY2LgF+V2u6rHzlsle8ls6AlN2rQWKdmrLe6z7yk0HVWK3xzwF4IQ5SNKg/yw
Ym7JE9v/0mWmzTjYdd9Ml9MsSrEDXoUFpywmJ2svG9BvUAC9v7+8oAE/xowxWLrV
WM6dTb1cTy35aFpmXqlor1JHidvC4T4SxajGtE5v8YnYbdBF0zrj3+aYGszX7S0j
nAOcUb8voqoTximObpGcxePy+wxbjPovDHLmfWTxjJ0f3KEf2kTsh51nyAt+DWRE
2hkTuu+4Q7oy3O+Y8wD4H1HrmeZdkM+9grutkxFbKp8jmSuuyRvl1tMyyO1FKuwW
N6dUsZ5bKRzNjEPPYC8aNWSodRV+fUVENeaGw4gUy9ND8JarEdE10ckpLA6cXAQ+
6AdmPqiEFQdK018xvN07Jscz6x9qyYUnCaJE3E8Zq2Yp3CnnSwoxDLoxiVEwXYEW
chpAQTVSkLOgfTcyaNiYUGaJcUboV35ijQBVw9Mz21WSpaE3epE1uQon60HMMaZ/
FRpPwuLPxexRYcoDWyqm6QjscaHLNojml2jEbSTqHuvzAHVaas3tqKnMvhJy9DbN
egy+P4BcaN00wNDM7hKmSo93jyT2fu5TPCikd77ajgj3AlnPCSyni+JuwTPPMrjO
lRrX/nY/aPJ4Pe5LBUU482OccSBgD7OjcVscEsakv2DlneyOQN3nTVIKRJ/ID6lN
qOFdZNb4WxQ4BUxIwvUMvJlpxl2nSo5c9mXW6ZMuD7F2aQmoMzf3Tsh882E8m/SS
x6B30WiPiAroe5WH5FGGakTcEfy3RCKV+ey935WwjUvw66yY1GPkuPGcBi9oF3wD
8Y9wExavYa+Qfrak585q/msjrGUOfFFh0UvnFYysH7FTxzp4ZjlcMwlqb5sPizFW
4hPXx0qq4j7To3Qy9iYbSm38EVcWaKHpEFo57mxA4fHEF6DkqbaDBgfgd0V0UKRB
sZcfcn/kklvoQkXtwSiUiXTiAcDySyVyRUOWN4pdJkgEAm7dic2RaQDNiLkY8yMa
uc/bxmVwkW5znF5Zc/3bsK2l8Chu/Km6r4o7Inu1rbbyhY/zRbosYrqTbNAbFwaO
+sF0cffGa32dEqFKAsUOo0C7QtcdLQ7qldyItvs1/LnrkVXzZut77jo95duI3DT/
7NLTzaJa/eiWF8s/oPwO2HzpiYnrZCg7/YPgcnuh4AEbqrUMweg8jN5za7KQtbLw
Q7r3eQPKCZqSJIFEbPYpOHcg9tEq08ZkewcQxuPXGNFxi+pkDV9dPTSKXi54ftDt
nWJCjKRnpntU8m1ztVpl4+awY5ralZG/nIWgzXpZm0t9JMaVjTdApfZ6RiJr4g4N
YO6j9F/ejDT1FHPQ/6o4DNioAZ1B7bZMKXV4uA2rnop0WALHaRhr0p/+LDA+kTyz
ZeZB64GpPz8c9n41CpqIit4/bJSphMWtKvEOJEtmAP9eu0EAVWNWtEb6+OWklxs4
kO5JsI44U36uja04czU7Lvod4bYvzPOdGapuu6mBb7yoXgt5JgsvJKf7O6Z4aG4O
V6R3gJwZEoWtKUiR5NrqW87+YB0CV9BIE8UordKLl+kzgYYEHn7QsBOBX1Sya3H0
wLUl5fzFSh0pXCUh3cGNoJNHushTPrTAZBztUEA9KyNtt+TeVtvYRzaLVV9GfejM
aPkNH7Ai7ojSa1k+DtRMj5PTczrXs/K6MVNZeaPaDKz+sZqvGyUcP2Ke4bPWDp8Z
wDM79cS15a7xrizjkWas6ebdsBQeQHRaeq4aShxWi9mWoDc7Fi1MwrlpVBlIOeYZ
fzGDYL+jcsZSg8jhL7sBF1ZLm6Dx+6gs7B1RZ4tsnISj9lRT+m+oxN3nhnhnuFaS
UMvHzlV91i52r39QqNaXqUsHZJmJnECpAshcBaHZJ1X1DuZRkyN68e2LEBYbKVS1
k8Wlvqn/mocc4KweCGs3jIsCcJ8v3E0Flcj8MvwuI6URw6oqY0MiTmCFu5DPqy7z
BcQprn0e1AEHOGUqYpwb63mEpMnqCFiDc6AQS46kLh0KWtr0O+x79zJgk7el0MCB
m5B1mzE5mTFWxFsKMTi4y98cForBUGtuLEzTfv9ENev6l2KJNaHqF/DNl+o2T81N
aIpo2/2a8WZgjSUTqjw2aWch2SkJeTbDLJ3O6SLuVSKS6iov04E1uBobg+DWY1y/
hUMt+H/c2ohTt1fgz6WCSwa0ciRmNZP6ECv3tfpizcseRr/Yqu7TNCvnNw/Oxp5/
XyxonjOq7WEd7WbIWF60bB7r6CExUqD6mvjn+PgLDPMEPS2TbRW/yDtl59VcUSQg
8fUVEKVqJcJmeW7HosVRHYs0fNSSp57AzXq4Cc9eQ59RHRrYL8iTKBS1QNSLDHMF
vzkWICdCWaWV88YKSeVL0a6xd0mjWyNtkmXGRZEgXceNQmgeY/kYe5kVDjiTsgpg
wn+Re8YO5ZSoMMiKf4kCOK9ZZRreUPuveQO62iqTG5lqDX4MWC2O4B46aIR3bEpT
oFyqyssjm5XtB5w24TGu/E6lZ8F9SWLZs5SeZxOwOo58zbi+vvXAbida2wj98Q5s
RZBD6GE5GmGuWNKCMPh9pX7yVdNIHqrrnMT05x5a/kh/9nvfkw95doiCaVSRmjNt
beXc9qF9Glze4lOBYiMAZicgXK1zMgR4puAdHtActQEe94ylLiA5LWknOgKNenhC
j0pKn7vfT/hf721kCsn1NZ4+rAgiey8dF37jf9BJXz1lMhNRmEsheOwrdrU4vJ2d
C1NOG8eNuQXJmmTkICFDy3wLHDf9ULDicRnSP609vZOfvN340xu+yZUYzrUXKkQT
OVM+Za2CWJBqw3TCUWLJfic0cZQTJYPMH7FnMk9qFGFcPtH9yEbCapOUoq8eSlPz
kSUNI5SmudJ5pMvjKN0yHKd04ZnKiyLv9pgVFccDd7zkqlc8kFajF4Gl+hYw7WhL
A8tlGSTkKIaLidWHB8ZL96b0+wshOxhK3fil0YbqUrinnqU0TEmG0Sq5TsxU8/A0
ZbMike6TnvhVN3wlik89BovP4CPTQDvU1NIaGULvVZbs+eg348wxZ2IDXVJdGRvx
2MKTdFj81pRA3cHCEL6DaA923W7q1R/PkdugmaaswbEIhHD82UsoF9xq4xHyT3Rw
7Lp6iBeTiX48GHL1A8cbI8OikxdxsqGbg8jdKgg+Avw35KtGzyX5xDcvxw/LIP4s
z2PukC4qWCvh++IokCWQmplnW9gL3v3hyHwJTKegn9xPjMpoa91/y6LkmEjB8IVF
OsVkXhmTlxpma+nHX4YBg5OdH8sp6R/saOLgWugPTmXDNwpPRhU+WATsfDhUMyNb
YvmQNvZvpvOxmGPYd6PPha2RMWiPct8MzpIhddCqVwvaVr2k7WvIB336lyNNXopH
kEaa7vJ2+eTBhVPENzs9U7CNeM0AMbakrD16f0JBb6gsjmHxRJmonLrh0Sd2+7Rp
r1+5bTxLhAa9fKLU2Xo0tG14HYhV/ohGHf8o3yGQRrzqPzdniThRiuINYZpEcXB9
Oi0+HW9+D5lwccnXO27k1z9iK6EkisFwVV++Mb/YwrxtjtF+qJPUso4hu5rCHhjl
znAox23O8bvkoSR6CLmpQPq/Ju2UNFDyjnli+oFARMMFe7mISFTgTVXMX2c8DHRm
sbivcZ4x5NlmgSqqK2dWL0Yh6VdCmTwB6X/OIjqfoeGkqirlOotckc0kJiRTkGCa
zhACZGfcWCz2pLTvytIUAGAlRKRtVWcKmJ9AZ5+4F+BQIPkVhucUyIX/TZNZMgM4
H1ULeC4lSYWMa0NLV5wx8cFdG5KNJtuO0DvpImreoE3d7pLhYhSYIyWw0G2T+5ls
AKzHxTqKH3gVZ1a1GFg8NslN7GDp8/aVq2c8KD7QLCeWK8W9QC8DKemQ4OG/GFfm
HS0k/l5bgVk4JSMsxRVvwht9JqAYvNU/epJ0BiFpIjkbqO8mzA8MRGzd6dLgGzIT
hb8C1T+kxWGgqSbl/+gTUfH/DNRh016CzHSciTsK3LHkJYKiLg6WYTCFTDfqbCXc
yPHxX/C+S7wQK4pa2+7rDy7USWR/nrFbb143y/KXJmhOzEAsu8+B03fIPCZvl1Gz
G8DmS8QlYe7oxmwtQ7JdSNsbNxW37julL5XQaT9jsAc32yJsbWQYpU+BNClGXuTy
RZctZnHN33+GEWT9M2BTcnumLRiN6+SBw+v0W+c7+s3mory09MzFIRoENsT+u5ye
NCe+sdo+cTOceYj1/yR67MolsSnE0kRYYBQTIZMV7sjEK0hincKUhyMAraMXAHbB
FNMnM12lMnBcV9Y/A6xLliysURdl91q40xvqI4Is6KH+PLSPgi5QOM3DH3Qn2JPX
TZq5fZ3RvFnmURD+A3ZbuW4DjMS4HZ2Eb3hzmyrm6GJk1k+O/7aQzg1RwYmI4Q13
FLxKbxWUCWhwbwBwjJir/4dGkega5BnX6ZJl8dc37iUwfemLPxbaILQaHzjy1YnC
BPVc/eOeFDc4NuHoaqGJqMhrJc+v1Cs57620prx+jpF1s/xDijBriI3ItHSiBhuU
+nMzNzSI9WtIc3UKY62auuJ8rj1tYSJU5rrYUSLFuMy3t6yXBVw2ERAC9kICvsPY
sjehJWRDbMP0l1u94H94/owIpqhuvxmRYMwFY/Pj5NboQ5lk5dF4YSOJRGPDZQCa
8mTW0LhCaTYJeNpnb5KRpeO9w+NyLX6xJfHh+iJCzLfSLDNIkBe9+zdvKU9BaEZn
pZ1qw6wcwJj3rbgsufACH0RE3r+T8FsWITAo5DFIcgbStdubdG84YkqHSKOvr+GL
mCmI1IxFWHEL1u2dM39MmE8DeFt6bkMqQTtu+jFCxx837r2bMhWdS7UW3RKH3CqO
VGZMTOzUzWmzUeKLdcDyOyGO6kB53JoG1RPne/bDOkPBBLg4oPojqdCUsqv4QPHW
FmCf+UYUblHDOiwppaE0aH+0WgsN11OINawTBod7ZFBRLTvf06DQDxse3oB41fhO
ieAvLkvpZAmODX0z0+KNEHn55Zxxl2HqKtPHWrxZNTEqPXYuDXPUUHElwUfbMDkZ
lnS0Ci7OKkb6UUmAxz2+EnVTAj+sCA2GmGDs+nmAn6fjQHoSKFVEAJM9p6B2FgJx
usocePuyX+a26BKU8z7fYrdi5XttfQqXixrMOYMf53PonMe1CZUqlEOtOaqkajU1
xR3Dr0y9Pk+EWSEN8brLN/X1lixPv7m3FqIutpePu1m7a9qjXNGZjOX6TbecUjEC
ddEyxBWHpfCnd7oM0CM1FzzXevsgsiioT4/ED7cmp5DYgYIei+iiLReF7lBKoDVR
Ohn8S7hEeD7pOX2iLd05fx7uz7f4XNxcw1fC/QyENj/M3F4NH6zpgkw4FZWPzzxL
WU0ORj7cZ1ynRBrNoHfilB2XAkmt5ljTAUkUYaIbkf//Qmwe+W5UhkgGy6Lw53tT
i0QduCDq1FKzTElEs9urMc8vium3QzLq03rAq9r71vz8UOGGopFUexlSGvxw15dY
nfQZCLchHKzY3X2Ca7p83IqyQDsNL7IoVd1ikoPs8FMnggR++BL0za7x6YB2WdNk
rU4XQtBKAbvKjIP04nxTZhb1eok0+bVQVPekpgIWwRQ9+15b2tLqiTDbJNfTwlpi
sCSVvkAGIxGLCDNogX1T+PaIhq3vE/MbW0QKx32SRW7nsabQE3d5JHzouHelxs9e
lxo10WlHgf5Ev56J2z3BJqxvBTaICD/zqKMaOJar7IOoTkfyHoNhXu7LJk/rUGY9
44/SfS/I0PVYmPehM2N+Wk5156sFTaW1mxeXXXB22AFXlOaFAPlWnEM0sFK3m4as
9+C5irA1CJJBaLkv+TB8vfYejijQuqZ8LMaMGpYQKECpG/kirmVTxwaby4H/LLFZ
+H9RgPj50LqaRvuiP7YjgOwh2IVtyPWR6Wv4UntPKpOTazP4iwGulImZnWeF+8gU
IjpOCdMpSD9C6gQiEHG5UDz7SsZZURQ+BNXSTTTokvrcGXswoF0D/1cKN6GN7XNK
XGimWC6ewcuZAzKTvpnRhdQP6Dy5muI57/NmgX+EbKAnjiftbluhOfepvq23sK8w
FQOsdqjC+I7mZQXUaBigl8/kmV5/sdz6QmzgD7pC/kk2nSZgufI507qMKXs7e4MV
vAmP+2/VqAAiWX3RycUqPi7UftyZ8cvFGiQAihUkOIoWttNSViGzJ6addJB0/0p9
rrvIplrHSaPmrpyxkQ5//htnF988JgfNr18x52C/B/keOuqe/a16DoFaG6NE7yTj
OC5raROxmRHYG2uTGWVmwHv0Mh+HQoJgUe58c02HVP9PKph1DKllM5g7AJyfF4Or
vtscXiqJ39n64VskI3HyMjSHluz3wuOVCug8XbSa5jhS5xyzTnpRFprrcORJO32/
c8nchXscMAcjWft9CAK67EHx5loDpXPI8RSqizXGlF5DheFSuqfRbdUqxWrDr0J6
3NMqV4JUrzxozypuzZOJJCT5Uq/4ibyuYaPhzPLCOh+Bp4Aps+G2OQBNub/lOIrx
O8//bAQuCy/byPeY1ZvHnPFoguPeDpuv2mufUpUFz7JNSMaxOW1W+ENToC1Wb+52
xhlWs2QuB6KmjAFdPqBKAXDM8GLID67c7BUyR848c+k5ZPqvLUuMl2FbhyEPL9TH
CYT3CkI4gwREd3Sla/mytcINsCafjnW0REEqnaUbSRD2xPICtA1KM8WWHqPD4oZ0
6d2eW741kXH6IwLrT+8EWYyQijTIz1opt3zpbxoXhciK4O6RyfGYmtZ394Qu6QY/
nqoeyR7KybSJ5mCLIftTJc5wCTER7BTNVkc1EyRCFjpdI58U80mczbWxAqb9w26g
xrpC6sCGLdbQkcz7txb7HDc5FGe+RnE5a7fHsBQnBTtUJSPAJ/zqSYtK5uv/hncR
cS7BS2XD2PCoiHTpdF+KPJMR5XRRB2YHjHPwg06QMEwIxl65HlmAS3TfxIr1q5LJ
VXF/GVFJjOptULyDXuZVlUrN0O+YhffMGhkCJ5sR6TuYSkIeo1IV0Aiz9Vv2zk3q
1Z3WymQ2wFe8yC2l6ecvdkswSs0ETX+Bc4Hn7qpdTvMgb6f9CKV5FFGELlfF4bcg
S0A2NGs/dQDNOmYQs1AsWkiP8ikirRYi4I4yaVTj6Q2ZGOkLv9pwvfT1HqXQGy/c
OPeaIjKaCMbyo/8pV9RRkapGvhxNADi4GKhHDtXNsaD1/yaYavsBL3q7qYRkdlFp
scuekVbu5u/WJNjsGBxkUDxuktTHAx9Q0WDPbJvaZxEZNVErFDHpGEi/dSbQ73vo
aPB/5hN9TZXtfglej7wXxqNh+OS6PhhieiwWYj72A/XtNs2BKqRfvyfljurkd26X
jzT1nVh8wOESEKI05qS666FzYuLycHh0G8zhH7536mIQQNK9w9A+4XJsXqlKA27N
zkUmnlEFtjyLMTVApCgq3Pxq6dNUU6V3ARByoqWCGBBOwYjQS+axArFM2rOGKBAK
hzxncKCp1Vdjz/Yreu+Ea2tpXIQRhkxrU5w1v9lQi46762n37DRiezuQv8jv874j
gCC4oHQktjy05MHmobMFDsuNrXwrFLw0tGI2OWi3YtMLySrhIrXemu4ua1kZtDpC
re9U6aL25mXd3NZyBAQv3NFiXORwb4TBknDSFHLOe/m0QHEak92kMVjk5JYz2UUM
Wfla4j5ans7p/+11PV20WcQhqik4pKliEanA7bssnonE9NRrsu3tlWm0pZsLPFMF
vv4EVXHk8iP1/mWTwXgMrzDupdYcK6tvK5j3sOqOgR9tucMoQclZq1UpDee5YT16
qYHLuGzwsToPtk2UFACQkA0fC3oePPkvsywp4ElmEIwMIyKheITdIyETNbWVjZuC
FqI4+jyr6XBvOhKN75POtJRPFZSv8dx3zFqDhJ8fsOKnvrgx3Oo2gImbSfP7kh76
vflAkV6U4gZkWx6LuT0KzK4BdvuFF+RC5xoFMcF2mMHjZeSnv3LJ81fjvi6QUrN9
Y25riC7aBMQzTDYAvIPKcDzpv3C/pc2gQ97fxvqHcDXUBvqJNza9f4DTYnDzCMFn
wHVxHqSXGCFngNuTwpbzyONOWf116tiSFQ5CozZs24jAqeEtyXVt3BdAizL9o5z0
bNRMYL1l4v7lSRs4jmx8y8XgnUo5wOqQ+X4veguVr5EjJBbI4HQww6ykuGN1Clau
LHOndcxY9O/3q4OmjVtVB6A/kqW25O84LoirTA8jeB6ZjngBC0J/pzFoc6eQNo9v
/W0fzGF60fagCdchpM161NtczHz2mcs8RE2vcEdSkeQYm3dIiPtLStXMGJ3ZRyaJ
Z8pBJacZhD6MWTsyfIxI/cNGOqAc9ngb1hnba8N8GtJqSaIhrjHVKpuw2PpBov3S
prZ/V/2YGS+CMEeC74yHmLBEG+1/uiHIry4WIHOppxvL48xUCqzFIUscDpE2P5Gf
7q1ojQ6EDmLng/fvLGjFOqFSglziC8bQOBeo0L4bQ6GUro0f1Io2SfhvKxBVIURV
YPakEJYYb7QgB+jmGTiohZK3sJoGzf4bZlxfbvQZsp020oyEzRfc5thlzd9aSen+
ycIJP/58r6qZev0BphFA2lGSipxwRKYrEu063EQeL/ZIN+p2WCNZUxT9MCvreP3Q
lQvE5q32lQK/ojWpOO06rUwBvhS79uQohGy6tovJYeDTV90Ld08LObg9R8x5CT0E
AaPPbuoHmTTbD6zroWHMrTQw0ujTBkB8+ceNbGRgsSnTxZCrylpslwAMtkW8VzzZ
DOL+vTyR8YV0oXyZrrK+/w8GAaXWdQG2FB/1eLg43M3+9UhduUJQpd6HQftD1BEW
+G1qn+o30QyY8eAky2Em+Enx8Lhc+kqJVfyWNWIvw+1JLvOVkmtwiF8RBcBiK9KZ
hvlbBqBwDU83WKJFv9TyKuBLnbJ5mulusHAFADI3db+eoATFZoyaknbCZN38DXTi
4OViQC9NTCKHp0x2CXlvNv3VQ0M+lgZJmJ+DMHzhN+PbDrF6HO5z9Rldkhdy76sl
2w59koJx09XeiYCDRsZSGeS/ufA+MLX3EL0/fA1IstyF9TLgt9Z6UbPmKDonPazD
JmVoOkvGX4WOTp3l9Gwszh6OFOW4fR9KvEwnsWluTeaIqf6gIQqVm1oJ62CWLmdv
PvvhrMIjKxdT9ohbEC2/FFK0Y79y2tXy/q8Ff92j1hTg6dcXS9b64m6vV68vU4mr
bKGFkew16hauCdHqgTUXjXm/MIssp8hk1pySqtSR4lrp5RGacxBeF2ZEUbkVJ/PP
yfhPvEEQ3peQS7zmutAGvVCa0pG4EFSj+rtGdEWMUxdSB9yoj9KFUk74ZeDQcjjq
wJMcn65GZJQDmFotaH71X1rCAif8w7KUgUDZ0eWhbUQe+ktwmWWfH4ypaZgi32d7
0N4ATuZVuzqFcujMTQUC1e5Tk6J3U919YoB2t26XU+R69IPA4Tcqv8aIbxy+xzkM
vF53q1yqXwV5GH0GdakhPMWnYUzLM5GQczN4Gae0EWHDE6SZBUahxNpufBGdgAKm
f2z56gBDgueb7fmnpKjQ5lznEDBKcuh8rETk3cIHCH9uKAe+rthHgw9OuL2112ps
iZV6Y2GHUUrvebw6br5kGwccNqVj0NT/PK/ieNLSHSQVgLjYtSaoEKMFeyhQZuhq
jssJTZ9FMAk04OxM2eLZHIsuy3xDW9+F3rSIdPfxV3XMWtmt7l+DX6uXqDydkIk9
IW8/Bw57qktmHucpL/R6+O0Vr8EcwXHS3DfciRtcKLd1GTk2+7GTXHalIH3x3qE7
mPC9udTgTlai0UdsmSerH0gSEaueadFbmorDXxjdgxlBuwJmyEz2oVRRtuWM4bni
SPNDHC0XQKPNz24VuDT2bRqDJOJdJoHleh4dK7bAqtS/Itf1+GsPDsQ1lUS4U/ad
XQF14XfEG41VSNjzBVtKSQ4Fh4jIANdtz5ZdPBTI7YpZp2s8jpykQZymYaOldv+w
xUurJGY2BmJTDsIJWBGbj56rIgj9VtOhgv61QX7zTjeH7YN+thcQxUF+dxUPOdIb
Go5hCLg53F+1oqE1PorSIHPBc1eTyo+z0d8Ow/xddnRGUySWXHBVnKgYFNN+H2Rv
ElN1aj2cwGJfpFVDAgnp7BfQFWcgQ7Fs0Ge5XP50pUtkAYSPXVSuqz1fJyfVm1d6
Q9teRogalA1+O+1oN60BHFrRjS1fOkMEVEOy+p+Yt5VpRvLbBJn6Jo7X8SdU5Hw6
q2EBqj3qlpkH++i0VLM7dE/iYqSvfaMqX21T9jR4xYsy1yYL0RBgLRZXUMIKR0jF
wqQdBd4DZXk/BgPXiTuZZEPAKLM99jnJjVXZLrPQYR5zSdq66o88lrRjr0FwiG+N
918pH7TxaCvErnZfb7PsX7OIL7B9spClUNBxAoYNZguC8SXjMoT93Y/82CxRZHma
3DSmROAF5UF/T0aCGgifEcY/+4U3Y7cjVrH/Q7v1KjLxBjnsah07Za+zRagZY/8k
fTKRLay/ucuvC/vNyKEJKpG64+O/88yybOoTrzPSM3elWh102oPuVanLX6ojMpOl
LRJtmgsbS7ciVhIbPw6OEXQVeb9ER9V3liAx0GAZ6ooYFpbk+gHjspjRH5jmHMTc
kyEgirobfGpRUSsxXaP+FCZuBn/2Z3PWr/YfsN5o37U8LSznMT5/P8k9Z92xpidK
KemcYte90zmQZLZRftos9bQ5D+smmMbVwj38bKRB1ers/4u+AMNixD5TyWGqZYxt
T1Xs5MLiSgYncSqLVc3rSvcHTt9xS+EHKmDijsYiA7Nh6kPwQ14bkpZXD2RsgqdL
/0FAi6jr4TnkL1WlJSUYL7RgZV74yLilh3gI0waFgyAZwlRDkjmd0z9EeviFuwQu
WnmsPU7vCCqKa2R6vb7si2GtmU2jC6qDdcCAmh6J11G7RCWtfDNd8Yewyptxa3PX
Gwzhoua9IWqRagXYb9JbiuUNCF0jlFNSjNqcSeQooDA4TvHaQbLzT0t+B2x/3ifb
1et5UIlU3cqUhqi7UNgibwIFMy3jeYIulElRv9rpnURrdWZx1jcJywZw/lbs6kqw
AZEnudLBnH9IWkTtoeDzv4SYrVMsY99nikJgWhO+ugT1Vao6a2DP6QL6PJsF/l9V
3Bb1Gn1D+kuXOSt19oyaKHVU3vzxPQ+HmxbdelS0DQam3rLQYLVZ/JCwfRf0UXWf
7aeUPgNKt77pYw6HaN0Vbd1XUc9imPyxFPi3NzgHkQ8EWXbuOr17u265/3NCRlji
pjopSnaFHwZklb3+Pi3YB3gKG02MD+y4SHuuBrFrQyWLzAYdkuUVDiNhSlO/WqRZ
WxkVA7yY2YaodXMRFbvUtMDO2N1R6I8VKeFaRBwpNIpnb0IcAwKOvpCs/aOmMPA7
7QCRNBzr88f9kK210FumYSqENn/XITQZKZS3qhpMoNDwxcYPfDBcSIPztTvWaav3
twRebiQ+JZynb43gVAOE2VbdMonGUE3Jke3G5vE/dNbFBmXS8AlvZF0O05fUt5iX
JZFwhwtPb98qQb2FRZUhgE/FJePpWcN1/Eingx1qV4ogejT8oFjTu4HgJlsM1Scf
NJ4cMBIBCu/hAZt8KQPTgCpFjG4ER78jBJqrin2MGGevtD3bTz0xcUPj955ZGrFc
C5bxnTOtQ8Oc1A6m+puLrOcHPEP4bNOiU2PmjXI7oeL1d0CQPbGHd1IZ8AAGIOTh
8Zy97+2Ik7CKo/trXJEPyMUm2TtBfaOsscSCXAb1EjTaFfQ6qas0HN9RbDjeBayh
VUOaxwfkKB0SP7BZBMaiZcJZ+rcRuN+J7re1ebbLJf6PpVVwqo8rYR+9lTIu5fAf
8W9FfsIBDhtFmJApkJbALNEJevmFTRfj+T7a1mSFDYyPb5vEExG10ObKY93/HR4k
nTxXPH6+7a1lbf+54mJQFonlLJM/VXnmZ44oG9JHqcgsNh98Y+NLH+kwhBHLoM2t
/aXLBPD1V02XYvKJhar9/A6YQ9pBD0A8fUGyi2S2OiqJmKSnIqwoeP4svzzcz85e
s4At9vYr/7OkQsP8gNH0RWMI1Bd+uZ9RVZgEb13A1aHugJgTJVgpppK6wnMU8Vfv
siDnWR5IbC6ZiiV82Ofu79rcgikAjWBMa0//k5mFkjsCEM+6bUoxMrPGiXi4egxQ
bZhFWnkD1EblXF3KgRaK6vllTU/Yo5em/NIRio5/YgFjIDmsYQEZta9SFmGTHwxK
p9FBvHqtRia0vOI8sshzf6n8O5BgKUuQPFcXK1CeBEaqivz/gzi3Ci1sJ8RpSjkw
SDi0TMj0R2z/o/9ak3yWe8+QfzkmNCcY/vqQmtppeGiLjn7hNT1YWyeqqCqIko5X
w73Xtg7hXa7syITPLO1QwJXnDBWrGdpNymTmRrC+06qWziAuJq96lLpCZuVt+zWy
4TRTOLSLuHLM90M0iqEh3ZXEiVV6LTRuewGyK6AszcFeNGT8Z9wwK5kmSw+9vJ5u
heXh8srcTAVHt9FLsBvkbxu+v84ccXDszyQgy61EVxP+k2YTJeU4Tkid09ZAo3OK
JTRuNd5kZYzc/d4mSrEdZZl3PymBDjgRQSJxaP2i6wkXCVCBQ4+W9lPo2OktkHGl
hmybTlHOYjB7ALDFhGAgAdMDtUG9FLX8QagGz4nvl6MrqrjY/kYAQpomuGhzgOq+
XQ3OlEleDyrITzfTA2vv39hFqs8Wg7jUbzD7ii0y2X0i17Q1lMiADuWykQrPM5Xl
ey813aHexN8Rc9EOhZU5R2uDAXwu+1FpFzrpydVcRCguXrVB6/Ou8v6cfqsM3U1+
69ZZ+BnHlS8NBQ4zip+9BatOp2XOkOD7weBZ7COHyW0/Li1wlbX8lGob06m05Yz9
mNsePM5ED1benjoHqZutClNARdylleH00laLNn2tNQ+SJeTv0A/R2VpccMU8DIKY
fVnMEWa4r0t7gL0M2TgezNfIOaU8T2jbDFBA5AhqaAg59bX4d+R3itSuVsuQnCe2
u300NBwe+2YUuckjyfLPCGGFq8S5DPIi/xPtOKASchOiFDo3l1aiu5bF6yh/4HSo
747pELp7Xzy1ozx4j8QbkzlfxiWk5zXTezZVFqwFN8m451K9Yq+970Frgu6QvV53
uQ/H/GyAYu1w6qm6PQtHAihc3tE7CHZd4S04XzhYypxkXSgQz1MtqBNxmvgPyldb
AE5QHsvSs7Q0mpayPPaOCXviK9owpe/1KW4metX4k9Qh8Z6ONr0w9nPhjUlqosnO
dzoHBjry8nfIDEi2qkq9weLJUAb8HnVU5VqwkNUrE/5x6usqUBrfXIZyuOKQ/SpL
22OImFsxvU1KK2Mru4BN/F2rw3SV4wvjzQEv8R2csPHoxUrKf/mYRRCoM6moCifN
ojpLuodXtS/kI9EI0rFEp3TXIwf+Trz0MQLNmyHYW7fEVq7hE5blnxp9Ip5NiGjY
nxRal3rRtbkRgGOKTmERnnWlfDHAJDF3t9MYRvfLZI7buNdIN1ZoSuugj+pcFGGI
qnT+80QOXnKknGQanexxXpNv2f+XyLw48T0ef2K/Z5QwQwQB9Fe2GPJF5UvPxXRJ
j7rypdjBCRQd/p13RfkPcHm1iLSc/qpDztMpiBkfD3nIMjecaupY89CnB4YJhQ11
/jj7U/FAzAOu0NwSW81pBGY75wn7eZnMwChT3W4M5ye3hMD4f80by34LoGpoAcHf
jhG4/euhen2K2wG5KEkTBzlTL59Ea0v9oc7kaABHos1UNDupqyuZwg981kupF50z
1Q01VtqG1F/tcIT/vd3ulgOSx7873mp+AdF91ZOBe6IRJDJ7V1fFhvdf/7/Satcd
TeK59TO0lVsiUa3Upz1wxJTy/rxu4cDqnLC+d10Vp+dqWVU9Gbjelbz7EbL5vyle
/NO9KTtgZMxNyTsF2UFldiSQC3o/A7iT+IQewaDmNXU7SXXv18g3xSqZRk3N/ymV
vrHh9CYYrBM/qsxXqceWo9qZZ4ZT1cTqwZ5e8FVbgFm2JpB32PRe6CEq68IXDO3w
ilyjABU87CQAxZ9LP4+wId6Rk9QNbZI5110eJlJTXXo7nnJhEWrNs8ielzSB6rCx
EyhZWUa0meiypcPNZtzISSBc+qu+HD4AUNIx54pQL8+orH+sONJQVEVOD6kkOojm
a+7tPmM4IyIeIQIP1BBuAm7HHuW2Vas4VWfYSQipUwHzffVePBHHtr6HINb4jyB0
KKdf6+WKj/3hOuJFOrVBUl/V8U3nKB+f0nzFl3iOFOjSvcgkAUW8nk84nXl2fM38
9mG4St+L8Vzdt+1bZh+l2jkK729ZcMTMZWc17NWyPO70wQU02pR4roa8FAjoUwQi
nEKplB95cMrF2XMLzCOnQKUVxR4DSigIlAJ6jVYCNWA1HUJ9O3GkgSDNamcOgi7w
isvk3XK+MEr1ZbWjwhNTboFVKcW8uCTVxoNT74+u+vIkOzhO6Ogh0DsXoswCtTNf
EXmGEIocAmZVBdLPlwvgzuVgyRF9Im/3vMozTXtGm07z5+ixHc313YtLuTS0OcdH
Rcl7W9LKBm/vSilJVpFX0MasTgJVfkkOgU7oFYGCgJO80vsIvetZU7NeDZ6CTOlp
PWwTX3SmUbxjB1PgKx0vpUJb23/RvDhOVfKcL1GG6o/T0+j0xfT8okVlxWb+1jUw
n7T09XJdXjBNf0wGM3fj0pDq0/gYMUiDyUWrrs6bPcp3nwPtfhhZ1gB1f3VcwBf5
mlJpZJiJUjgKGjLb5FSUoTaSFTl+QXSkJV0eUYxdM35s2lzJ4i/C7HHYYj/rJ5BQ
mB4oyNVpNDnAJFzLEZaOO1SpXJ2sJgsgP5VkBHolYDb9PdAtI6nMfrYffY32o08e
d2UbtSgUc1pUg5sskpL8mRhvcvN2FvVS85FdOkqc09JT/LDFt6v2tuUPeIV4+x6q
OXzXvTDh1hgu3oMmO3guxPcb4y1pTwL5dYUW7gorElXskONegyrLxEklE98jKqYu
xLpUegQjX1jhKKt9ggrN6x14IdxIejolczDK4H3x4X4UTQ8Thx2wNn5ynbFZLMzl
pxVyAlFXSFmwsYBEr2AzeEnhk0G6MBl1Bbhtnne5wJgS8PU3iZIL0DV2skO/n7O+
ejZrj9f75oHWGkynp1zr21bLBaV5RtlUvoY9hsbZkRoRbPQ31NYSKHgfngJk4P6q
BQQfSRCfkaFF2EzVJ3sXLrvDEVhEHihfbvcEWIqHlaFY8b0LTwsnDAAqdZ3iQdou
tgDIEDxNrtt07rkg8Aaeqe1SyPj0rLFDvX3L5eB0tw1Zy/axqPG4aab2HganU/BM
6n1IHnDD5onQ9IY5cHGlu6ufSQetqxZwwhco6t5FMxtU3B5hmSFV1rWeOKONkIF4
zz/q34h8i/lFqERnl2jL55pZ1mHWEWGdENzTYkj4812XEAIydlpSRwl5ci2yAyOI
+VCNs99r3Sxnc4VsB3prDmg8a00PZcHJLapjkqY8cch+VgsyWB0SzdZQq8dRaNiH
mNgUHUe5v6afEGNyYetXmEg9Vlhfml46td5ZWMdirYjVCizPHU7o08RIJHZt4rga
IO9d/1pe5ODpCHAMLa+eNVz1/0MZqhfIhKl/phj66dQ/i7Tohyk+vQBgGu4r6L4N
nNpzEJXzkRsPtUPNpSJYgpYuTZORZ7zHk/ekYfW9ybkHdgdQGfySA0f+inIoxpK7
vWNr4H28WsxhZCqVCJUuiFSbuFZAm3OCYrPRl0QKhThZWtsraYpiN7Usdk0CqU9r
GiCifIgD10d1UC57norVSmpMIzUbpaAeZz9ChQbH11CFIYiGAMlI+YAgPY6F1jN5
ZFrLj65wZnAexkf03NNph2Xi3zfHOBgOAuTWqsM14Q94mcW98Y3Uw//3uGju+5g2
0vDPP7Wo30uoVvz7iQI3UZGw6nO0/tH/70oSoZTDvohvqDRA3Pjq3Ivcz6nnBQE4
OfdOGQlSRVXz+AUMHAN6hsVw3NLz2VI5zg4Soi799wipGzNijTjBXKbGGV7SelCm
Ps3236fxQouVmrtSKmAmsb4vi/qQS8KRa6WWEVZzZT3CMlgNdY/cXXyiv0gSCa4+
NdVQPGiFlUWrb4gVhQLj225qLlUpOwd71Am180RpkVNkOMNuUV+gyWVz+2aM+5Rf
PyoSwaYrvtxEdVpLIL1hl0pZ/I2xVeGvGxSH3HL3xaTQ7Z+TUdwDasrqw6RaZVLq
hkDVyheFtOBw5eHzX6pS2/xF0nn+/2IGJXM92DYesrDIYmqRVbWH+yxbnJNNszxC
DZUEZYqTnXG1JROny6qXadx9DyDh45ggCsmPsWICXlQt9zLIw4FW56uIDD2iIB5v
wHiNLeFVBb8FtaNPOxnFvoRGcDHoEwaH+Vfrq7FjCSr7TkxCTUi7T4kGjJPrEGGL
RTZagzKVmxDRh8Ha40cEGIvNHdKk6MYvU37YWbVhgnOzvRj3dNIbX7qem9tj03Rs
Q47hn5Rc2Q3QH89bjo9+gbGQos/4xrwQFnVjKCQ/1l1XHAtIjZ/OZo22mrLsOcJn
+yTqazYGsJTw/t5hfXd6JM91UoiA23sv294sz2t/DWLSehr7boD+33NAKMUcSOet
ecEvQuXGVo3zbMetDG/VebZ6kghEK/m4OKJGAbSzJukg5OHw0CHDXlXpYZdvFt2V
y8IgV7L78PJpWJoFSN3q2KKdMLcA/a66xG0xZffmgE1MtRbzPAS1FQbd1Qf1TuNu
4g7SOg6P64lAciC7SeRlroD4EdCUwxNBroLT7WRSj9H5lQCAnQB2CJWouQOPTEzV
Obro6OMp/DLUU14e2Ma1fGd01fkyX7Y52N0rGcRP0YNzU3mHyh2k14ylojmUGLU7
dxpIJmFX3N7n6VbUbTHh7GeC8ZmcsHGml0NsMx2vD0xP90seTS/Erd4jaNok/LRy
U2eIScUUXKbA3M5jEdH2TAKy/5ed07b/pPAd7HLxEixPUqXR6Uo4YpPs/uC3UI8s
QQLc3NV1rLu5L3zYDoiXPBQbHEW/6BBOgbTJHm47DyZfTjTyy+YrLJMWVa7qEWTA
KcGr7h7BR8O9RGCXVbWYfJ4CKBkZ5sLO2Q2XXvRehLSj9Rzg2AXOHo4bTnBKrlqK
o/EOYmu7+eCT2jjdkHESZBo/xxygN+ycFYoDWTxSpFcvnX1/uC2MBEZG5O0jViPi
`pragma protect end_protected

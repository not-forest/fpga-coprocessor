// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
ALXWPcdm8w5oyrgcOjiJtZLrPS0SLsAovJIBHN1OgCGaOZ8HW6am3r13SWav1P+HVnIThS6jh5wM
G9Ru1JN+jxURbUBfI7uF2GBfkVRc3qs6gRSJlQGNAmt7mdgtyv2MA7dY271lE3Au4Vd5DEW2Rfuw
MpHKrXRKMkyTfrLm2l+llREM8ipPqmQoDJHa8bcbsCgi3wZ55nvP7cQoRwssNILoTfO9dQNRQDIz
kTZwly/gDD8QOI12ScCHz8m/bOgvWjYovgc7lQ2w6SI7V7d2Rbp5R8tWVyUCdkPVAnINZ6u96Kyo
1EyT486L2LwYXKGDnkdciy9F8/cqrGnOoM1Pog==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8592)
PCnuHDgXjuWCoVOqi6kKsCuddS5QfcebcQF5vCFImzY4hgmOQE5iMPyRmIHRfXFn/WqnBMeYOlsR
YHWygLy7D3Zgil3XTDDWY7Fnjh2/mg8QhGACKDYNcINncSb7V+6k5dCtqhYNopSxCrun/Lwoejcs
DHn55nXI+uxMdiGJBX6zgN9RC7jCwyi+dvzjeshFWKMDChFkvFC0VXoMEAHN19miPlL3n1Azgr7W
VPLd5e0IRmPbWiivk6/gCqievCYt8NjZcZ0nt1PlwrSpIbFjbxuKJ7v/lyD51+pPYMln0lvwS1qG
AaFNJABJivzL9OxSjHOYDpqOi9/EiZOJPEdrs8+xT/HYdxjhe78bBpCtq/ZQwT2NEPEbN6uraldp
OiCuWGDm/k1kCzT67gG6UCdlToCUOMtemhd4R33BImgpsN7AR1D4XP7WqmgphvNHOiwGsVgr6399
wk5rg9B4H7P2KtQRgoClnDaz2yxWboD3S+1Osx18wJLDqRe8e6rX/xJeFu2RHsxldSw4Pffavq7g
Zdq9ifL09krQmYvcozav7QFrNfW2uDxC6bwY0BbC4k7DGO4m1CV5KpdK87PZWuIakyWiEY4AVXHK
aR3rXWmUFr5iigTE/4AQYIoAGKV3vv9IKITd0oc6k2ef6gfX3HxfK7uxFi4W/tX+VhIDwkVBQpxm
vQImsINmPq0iiRVJZNbC+gBkvz4yV9ZxpRnIM9+rRN4UzgYw8Im0H5+e1D3+tOkzd5oNlFkxalIA
OYUpRqBZfFkWViNMeJwaP0y5AUT3Ej8ZwroCUOKeeADfFieGgB3q5qjy2dnYFoBxfqIcB5lfypKh
SCVdjv8DAoIFpJhWcmhvOKHFoTlMvzwLKWaa/b5il12/oEGRVBog0c0AigTmbkWLib0JcXfuuj55
54zRWt0/IK1zf2CfurID0hnuEppRoQBii6ZIXNgsSXrgMFYHwBsTBLbDunuekPEMubQb/vIDAPGK
4riPvZR6Q981QjMuCwGgOF2wtXUyiFSjpOTN6VhiZQarVgiVMfmliAg74m6F494ax24SGmEP8B4E
oWSwM5314JEQt6QNotcCie/CGFPaNwGMPTXnrDa0fVHH5Q2O5ZFyshVT9JH86oRcc+51wyyx2MOV
h33qTxB8seZvJ1q6ByZA5k0ntGfFAkoKXsc0N6rPoGN+E0oWS26hcrw/4gKfBz6bFUAf0aTtRE9z
y/m5RdwAuK4Pphg78LCbU5ureYKgUGWG9+KModGRN44xTJZH99yzYksHIWZ+NRR3daCux1z1YNI7
F75GpeygocEknbO39+CbDl479oOYRrWZh1P42tqFx9Mh1DsBJYd69ds5Uce/b9ya9CkyJGIr7LIv
8An6H8GAwxtMjUJiZMbLZTO1pGOBptj+866dxUzguSjpTpgMRSyJMD49AGkego4aX2IUjqt29Mol
N6mlwRWMVlVgwNFavGPGVBNkt2c38b1a02VdDQVNK1BhuRPqQj95VgKrmLc4P5fuW5Qt1VdEAEF/
CvOcTYgMZhPIK3R6xQOpojwdgz51ZJybPKyOQRpn5qPzj2JJtC8jrEEERbiAm2x/+VuGgel6xomY
mrek8zJSEY6FccTy/NVNl70gnKvQOMtooQqJfhQ7H4zq2Wv3qQ4oPKXl9eOAdEjgAdbwkvDXFBVd
y8n1kipFfl4sXzLL4ttGJvoL7iPyEukLw1eBs7YmtrZtOgNEZnMXOa/JnFPaoRZ8vh88zNYK+6Va
Eo8yoLKqjENaVidTDWrwIcqFf8GmtILizPi6DFpqCzovd80dz6lfB6d9uGXie28en3ci4rgcVhXk
Jm8STNkbxjOOJCZrZrIeIixhiP7ffEBWIrD2VyZzP6ktz0Ge8G4ky50892Ax53McuESscHAzGFzC
MRBzT/fD648tGI9qikEbqnILWlYzs8pSMFFkAQVteJ6JZHCWA5nenD1GojMoNPOFtskkT2knh7ZM
vxc1QEeO/psmf6jblxfWxNenyKHFrfP27FxEzbXtLgYXf6oKfmPi3rpZT3MLzoT693gnNXc8QQSd
tBc3KcafsJAxsO7/klLQLh1+cABvyxARXUCdXpiauOY5q3Dc7+GszS926TFT1EG08c5hsubD908j
xbm4tvuS77JsgT5l+tjD7UZ4k3csxB83mvpovColLU64/gsDuERDvK99LKDiGxREi5lg5N4LGLEN
ZdfBdJYitqY35k3gZ9sBorQh3w7lIvciWp5DAFfX0M8z9jq4ItLFeSDo7Re1Y/azcOAYyqC4vZiS
MY5GO1Ph8+JUhwcp7/+RPxPBB2fFml18QUqrFBzylqLnt+Jj7meM0fc/5mIU+ctRgTFRqyT/jx1q
qXozuX8on4s3bdwtcxT6cK3XLPDK7Li0A3uIL5lFUaKCl8UoscPVH7kl4uX0Wz2F2ozt1Wqag2ht
0LJhuOdFAw78Bxn/8hhY0fgnF/dg+zkY3PJl+Il1ZMeOn2Y2tanbeCOWwsRcCmVUbM6ejnH2a9go
RhWAVHKWBldjKaaDFjjzq+H1NvbRBKPpTeyPCqXQEXHJAZFkYBlhHxx2z5LIop0hko1WmQwdfp09
Tf5M/WbtMTwbWK/4XKyKcCOdfO2ftYhwNe4ulIrsQ3UZwIPYXuOWtzWT2/7ljg8pDmcMJ31CU8Ac
xPhsRz2OBWLvT1Bap/haASbgvzs+kP443Metq2yvmevHGmYLSqq2j3sSBLru4iJ0kEueYxzbKks9
TbOJ8yYV2cdkFBEU5OjksUisHYGAuMpF8s5KSOlL5OlKgGgDpt63QqUjDB0fg+tallZdZ9LAFlLv
FVkgWeRigTjz7vMOXj4zqulhgI8rN6gSR8gX8A/DUS9MolmNzRpLBZJdRimKQGKZeqv5t22un06X
BjKI1lcMUMzouJdjUvZ8PYwCV6X5DRdLjuJeVOh5O9D88DT4Y5X7pEk8pvsXKji8j0dXEzn3gY90
QSUmESmlJ4sky+MKYpfvE8+bd+pkBEPhXq//wGNpyeEqelzcl2b0S2AyT1YIFUu0aDnshOvxN0+R
X80aB6EZJasHdmflPzlhPeF17e5bI5VhARWn5WzHzrp9nM4ze7LIeYA7JCTltxD20EyF4uSUMNJO
VnRgzvvd0hofbO32CsVHEs3u2oU9tFrIG609pH0ODokpU0lkdTopxLNL0OjQdYG1MvrJhibtoWeJ
gE+Lo1/m2jUq+OE0GDTZRw89eWR41FJNnYMG9abSKwsHiRdSS9xvjR9ox92oktBh/lrVoJ8c9n0O
ohvgf6sWXm0YXpqOjZFkHqnYIl3TzPpzk8YdaZOrsRjwLNTc7sRQk/1UjnXb/z1MSUAcHF5OBjBj
oTfV6MvZmPE5VTGKOqRIob4/rjLaQX9ff7RsKTo6ZAeRPAoqzxAM9NYxInsT83Hfx0Dr9kaWKVIN
BaB0hdrOiEhipKLNQUkR3jZ4Y4OAcTJM5F2qcuL4wUUsZWAr0NrHcqfpkorM8K+lTaz4ZJLYZYdg
hXsQhjSrKb3nWtaXIMbmMg9wjs1Vw9m/fLSgJ/r/ose0jMNnRZ8s6s3HUjX4/YFUkUl8znZpLyRK
a49Ebcu9L3f+C9cC/lQaD2SMHgYW8pTqfRmGaDZa8bCIJ9+WDNnEARunFWuBXsT5Rz93q+E7byf/
F0VpqVF/YyKGZE70OUKJ4TTN07iiR7hW3SeCFvrCUHU/Dotknn8OZq13ZKNHBwKLp7oNRBV/fPlH
SUy2cWUiwDOntD7yem5utIl9Y3V2PtfywmvwUfp8RVEQNwnjk+HydKZZVdRUN7HZIPdMVVKuq37T
579i0+LR0PNdPb0GVwpQsFHOJPXaFL7oVGgHZtSg4PG8ALa17+zEcrZ2ILc+f/OlNOSwVBgAtOQf
2ohXXQMmy7K95IHca83PZLudDVf0BVVeTMOEOOpgAf5lPH1GNAiT76AXNzt1eTTFYFApsF1jOssp
jxjkuW0bumndu+JQFgG+As40aFzEhyuh4ZYp7unZqIaCWB+9dRV5n/S/oE4WX6pWduYxF1hAkKBO
/xotr/Mtf/iUUBFWQOP9Pv4DgohDYAwDfdxpvUzBeHo2wh6jmBqr6WDxh0D3naX9LRi5UEYGendu
P/6jEeBJ6jVaL7PM3Mpr0SoKaSLuy08pK0TORXTz83uPMt2hHQn6GlSPxtJ2ht1OBLeGz4sPW0Ar
nsHKE5UlcuNeF+NeU5+BHAft4HbpPpJ5xUVwltLxD+/y/x9ZIsut/GZS6NzjFm7k07Kt/bwZh9nV
4GJfzP7zzKbEXGDkYv/K7aS34WbIouGo/qUhRvEw03V5m1yk0gT06UDt2TlXivOxJXau2dxFmzfK
7Lp1wDcaT97r4eOo9LtyIefCTuI2wc9shWg7MaLdt0104XUgdTUzJUO+UP7ZI8snR9EVZADBDWjs
7J66tKuFiRfAevIBQVa/5FAtp1Zw3L4rnk20uUVG4PngJJvc/2qgG/q3tXOc5mSFCFQ+S0QPm1E2
yaRNF5gEr3FF7Cu6enCr65wstnKOaGECzF0MgAOO0Ri8E53Fg1gYC9GvbzlZrNREP/jDrOAL8UJz
penuj6+6UzHWWQTgk2ckq8H2tejGHjyi6/0rYoMYidddhOebWB30KZXdkGtEaVz+G6PJBfKx2mtG
OJ/V19dHCkCT5CE9k2VmYH6LWiyHAIUmOBhYk1HWRzK9o0xIsymB4zDVAIeSF3gumxlxU55nzYfd
6INmE9lNlJmfvWWBCVTr1Ml2vhGhCNZzRz/ejrnsjp7hyKKsSqqYJjfMAk8LokYjIAN799+F626z
m5lUZA31DmCZSpmMCRqmL2YoI1XKG0Mrde6+iUBdlkuSz8oa98QyOOxzGSaTFC8KwQiEeVzYa998
sbY7RU3yf2PRIUKzsI4++SPs7CCmfTemkABSX7frJJ7SIRnREPdqc+co5dlzYvlBtqHodHs0eGBy
zwBgV25Jh8JtIEZhzKmDuadNeXJa8oPtF/CVpNLkB19zKNPaF9AiAGLbaTc3sS0ncQCyov1q/3V7
8SbEdT6nVle0T24c3Sg6z9QPX/RYiDCqgfXE2nlffwYJGC99UxW6atzZyIGQ4wSeSqrJ5rDj7cMu
2EYs0k4/b1h3ZqnaMt0KqTuaV1SR2a8g5dhmqhdFqwWHsQRVbr6pk40Op935bV5y8T4+VwrDfgji
uKPVuMJ8aU03eET4U5knUrPNTcPt5isRPcfJLxY720hxBR+Oss0f7lVbvWuAOnGjOJyUJTAzzMXx
iNaJ/SF4m7t5WTz26BYqH07hv0O2Y8ZE7BjHyakTGpHLzYpqPttSmVq6ANkO0ZbIuDWkl6MXCOZL
nIlyMVzaPd6CIYS0YDk6mG3AV9xSNNBECgyyX6XriudIpnmLDJPgTm81rTb4yWmfkYq9LJztEpam
hSj+tOATyD2jPT+99Q0ZUqPLGuiT9Z2nhKw7VQZJdWqOky106UPILHBJVEGWuDpxZjHFMg7dt/cC
ItBw3oej9WDo2elziOP7mAJgUveXQ38VOD0tj6l/lOBL/rqmmSY8q620wKmYzaiBMB6mVept7sw4
sS6WxeI1Aei5gMr0BiCRvIKtoim5BOMhD/41ApotsIgnZTquFv4bIb2JbPWQDS44pXdF7dIbIB8D
bzq595mXi7IV9v0QddVcapElgNXGU4kipn2dk3dvGT2K3BnEA+2kwZbQqvDRqAQwktSrlvIH/mpe
mK4+n9RlqthUayJog05I0x5kpVH1Ob0g48xlQXsnWo1/wX7/HjCut5rYqMGJxXDZ64IKgcIH5WGb
eYmsZAWJIogiWpCQpa3sxT3MhCuCNXJ361LaxZQhqBFAuyzV4fmOuXVd4yO6DHSc27o+zvAylNZN
Zj1Olvx4f4VHt3DpKEoXwvTYam0ZtYGddAlOdGZqMaVxkX7jsFfndvyp2VbcvYGxR4JCHDB2Gt+O
sJYmoYR+smH5P7PxyhIyie1htRnYlvcQTbvLzpRpJMDFRJYGrj4M9z304y/twDcBtzN2CK64O/kV
vvKQgLW1CSqTvIKKNPA4rR92E1Mj4qogdWTEXBH+yOm6RdFd6vEFvAgOYFfB8B09mUEs23rRtGvi
yDlMa4oMnk7/B6T5M0PQYt4B4KEI1gOUl4JtBA94hDKh/FFbbfqPwNIKjn5jucVa7R1FBFNYc2tN
T/ZmqRxGuRmA8TXD82nR/qSl0jCwAj3Pz0kUp87cOQOqVy1p1g8M/Yic5ioIWACqVb8NFXiQqmb7
0Crgjph+KememQCosovqh8RqE15Oh4dj5aLO4uQ/aegxk3RJeV3/pyJkCawqOQp+C70oZXSHPwZn
kkrnAjv6RLBV058SDOKdOqWFP0c/2OfoqFQzoGyUdQxtovfBR1YWx977IwSmRZScKPcrKwjTqHPO
txzMdSNIc3sJNp/1OnQ55lwQO/GxFPmNNn8DFw+Nuvs1NULhVFbUqJ39wAZBax7twosSe+/tGijm
DMaAfzrQ30geMmCWUFLdoZ4FE3z3NSLroA15Sa7v4ImvrcJvbgMMYbfIc0cf+BeIqBtEhwYsb3bm
Nd9TZmWDiv/3+BiZj9G27fLoCaEgHk/enXY/WKrpo3wVYFjYsDe4pQIc48l8Rysc7XemDE9fiKSZ
pxT7iapbaSknWVJBKdiUQUzBvoHIAd/o3KvIr07lS/0udrmFCIaspc6nDNzmqme3Htv8EH6LedwO
jQExqI6SkhGI62NOtG4ri10S+DCmTYywLT2mcPu3yk1EzFYFfb4giU5ghstmLGp3xvKTHjV+WUCt
VzZlZhT8naurSOZhOGJBgeSfS8EjfNmcMHv6LTwbpZTpjUYeLgEa6epPKICxr528eL+BaTuC2X5W
b2/NcD95sltEwN74qPeIBGl1/30pKtiXdHFSRWbvs/OxM3OUXUNiYLaCPI5oKEagnogMk6z5Cseg
x8WVmAfDrqswwgMP9S8SihSr42sdS2SKat0iAAz3IUCjq6HtZ6HFChRzGJImhsesHKQieFnezaJW
GOSdM5/l1kN4H6EdMr8KiAt2O7o287hSJq3Lfpcm74Yc7bsA1Iu7+/C1p/qMmZFfsKDKvObL4jEG
tKduPLuBPGI9DzXbGc6XDCo5VzaJ9kr/CK9aDHYqYU3SQqu0TT1wPI8icX0RBGW4I9NobtUBZfSJ
dmdhKznJE/UsvcK/GkX55P5gH1PPiEhZPbS3SCGygv8PujzsLiOxXs1Bgb0ZJDg2PyHeJ8kwsAtc
GTPZU3AstAxt2Xk/3xownzjqt4o4dDSPK4pFqVBQ/V35V4/MsXqzg0YybSWXGQjqjmpa+DB8pawq
/qIUW/ngfiTgeBPSe815Hh6mSRx5wOr19R0yEKAW4bS/4GC/u8gLTUgz1BO0SkH8wYifBnla7Iof
1FEdomOI/L1SOFl04WVGcX4A2FzqluXoWeyliyfvmDsm/IonIt8RtHrmwVgK006pp48T6sYe3rvA
TTzija7AFUQ89Vxn0sD8O8xiJi57yneGa3EZTHnQCYepyjSCl5tHXMICRcPUV/il/OdDqm52+NiP
7NC1/tO1Qkxbtsllw141wYDVjjo4DX8p/r3iA2gqnUcFUZ6hJW6RbUtwDU7nh53yvbC4K3HIosub
GjC906JSwo+jA527t169XFLzKWqemIbeJrMJbBMcsX4zyWMfPMiZJSeS9WNZi3PbGhUVTl8ox/e9
DXBxk/DhJqRoy2DTzyRcGiNXNlQMqVYj4hVcqLU24f05CQJWFiEtsqZ74myWZRFuwzKHanbOeQYK
X6nwSFqomYBuMMKQtHyrmtqZIHWdOEdZL2bEGy2uHicmX/wDFFfZjP72GR0w0II8DuKMFRCygFAU
g6+C8e2znota+yCoLppFHouklRLqNR7mRgyZyMPgRxvLb8m0ymMz85EF8ylYPvpRZPLLKQ4zP8Jz
qyEcz6hJGnr7VTl04ahERv+sdo5DYnTQZaZevOpBPeeXVDdubAHEPVh4YNvAeCWFYomybqRSzDNw
aWcBbPFBtdVwWFArQVaR19MenBkSiQ4jDqiALIqOjDpN1GXFyDQJMa0PcMpIElBp/Ui5auGd7rQh
qSL473YCIlyymzaz7UYeO53FolxGaThWbPikL1WMaBqOMdcvsEm5BidS4PzMUTE4G3Eek4QQtqDx
AGlPP+M17ElnZGoZnB3He6DqmZxqQHJlhi3ya8wZltFuwG8XBrOhMBmdFUy3VKnezyeDM6zWGz6E
SsDJmIspJ2zKD2sgd6gcyDwFEqWwnAHvNLBCqnRNkXL4yO9ysWpSnxk0uWZspoaN9tkaLOKeS0sn
2b2SL33KO73q8xe7cbf4jwqShim1AFVdIKdzfGIpnxf7qtmyyWqh7mFSOLNKUrzgP1Js7KdpxslN
JesrmY199VXZ2H+xfwTiSCXznlDQt2BZdi/RLpJutOqy+GklYZANxjyjw6rlAII/dZTdOeCsP8WC
NIPyPDyhBnIIIf8v1eUShPF1m9VDRpYPP0yTO8ynFDnMWjj1YrJF/1mcaWklZas+SAgO8p8cq5J7
olAojBwXXOZF/rAw8YmDpu/rQQbYDOl7/Rh/JXoddDI+hSpO0LVptVcf1Q87bvUWr5DK61r58ler
B932UQ8zlaJt6msZcMM6AFlfrAj4GqynYWfkSovHpf1F9/Ueexfi1ufO5BZwWgjmWeTQqWJSTWEn
j4PvFUW+p2bpqNIhNEVnQOUYD7j6YML+ZuCsEvKxICen8RFLq5EczpVIinwAS651ROCBUtQ2g5C8
6oNpIxJEI7n9zQDv0kRU7//DndIqhaBiKgfOujB1PRU6l/jKKLieysoAFaNDuqGfobrLHQdTLBQo
NdW1FpVRaUKjqhHLpSPcgkFt8zchR2MgyMtq/X7rzXewgASAQw69Ql5+oouLSXeBGqnJ/vQ2jCD1
7+57MsCytaNHbyiz1vZ9SQ4FdlJ4sUdkfYOjSKBeop7VIB1+tbprzjejpD/mjX+26sJDoi9zGDyH
y9QoxpzerOmzlqwHYn+DohW+cKrG0K+nen0Ek8xjSVtFFfGO5uJrhhxHTs75FZGEYMXHcsQs0wt7
9xQS673MaA0cDrMGP+gZEPJdh/5MW9J0SOAgrO47QSiWHQoTcc9bmlGw4mwEGgRldUbVe60eEc9i
/9/nx4+IeaJDG7ohuCbDv9JLP3YA9cxYKFN8AdLLs8DymZ5lES/Qn8leoKH5P5uXkJRDW2S8fCdn
vIlCypluSsPnpzKUYdomqBHMIfV+5d1uKRXhUbbk2Dr3l9MX7W7tNj3F6fUPfuKgkuc86/OopX6V
X4XdbWJUEWmxVEkl+Y23a+vLBi6yuyNzO68vSxZ0tPQUJS6puoG6M15hpX7qR0GFGO+/l8WWNp9o
muAsR3rGIQLuZKdyGggUmjUB5iBDp+BmAZRIzvlk0GjXKo9TCDHUHiV44arbTrc2xtaqPu11Vwy5
lD1T17RGMxNq8CyBeNwULwwE/A1p4ehCiw19g9zTC4rfNiQVoJHCmCfxHmy8XMiIWed7qQTZxVOx
k+FWplnGJakK+SBgX3PS+Fzh/vRzR0Xv8Mo2TP/xooWAYVJBpyJPiXyRoSN1NCEzolbnw9h3f84A
8gIZK0+z0AfmQ8668KJStm4+DIRZndLMA8s1s5MNUQhhCpE+YEhdEfRq2Gy6XKbxengltdCyy5wM
QkAXMWlBN5J8ewt2Bcuch1j+TMO3Y8VfLy6evcU80vAe668AVgkpd59ATukLJ4af617fVflxxEoH
Mk1Zaj5MefCULJcGR8zhg3I/GHLxj56ZU/vZqrbwIpEI0/WD4hmUXtuFQtvtICt1U1uWoh5Yms21
wVhHxkO3IMEt5/x1U1PtjggZUwqVsaM9sUtS1kc2TuCLAnMiHw3AMVdJ2j6yv7yNY/SSiDVUYqkq
LCh6kiqAkL3JmPc1SlqAz9eagu+jfEz6Zr9DIMl4JskxafbOljL8yJzlsdL6Y8jhqvJHxik+78Rf
n8XYEa1xoFIDu86u5lAaQFW9EGYUSivxwElmFMekF6Q5OGiTlJfum/MYMILNyxHFMfn4bkBe2n68
FhL8awQVxZNPaoMTCfmZCUnw9AaWTHLKeLJQaGzIjIfNE5pjXAMut4SQhxZPio9TV0Nr9qu2gm2O
80A1qn2Iog39vE1vG7IGJXhiRvziVRMKfeimk4uviPwhPn99+j46spoFiJdYpu9WEfSbg11c0IpL
f8E3J5mwQ0eJnct3sigXWdOw7lYFss9B9kdlvagxLWyPOeWBw3w4S+Ie1qGEUqxLPdMKCi84oexo
A2BdEhtfBCR1K+G0zjzllazSmgEAUA7e66vIoF9zLE9xctfhlF4RG94mZwQyoMZ5lKk2xMmVF7+C
JuEf79Yy6iEtAeGB6nuoGtXS06R8PZmhbd780qonVt/PeuqlO+PiHyMHTj3H48k5c3vf473YI2OY
JXjb0bwVJtd6wdWBJ5sWS11WYrvqhQeguClSTJLfKu1O7bI/s5xyUxCHgcUxrTepoMMd4Ip/kcIp
PPWDeVcr/awcXMlg+A66Lx7xPKXznSgXy6MwjYXgqXVssh5fQnEVYIfKKHestjuU3yTOdhImrSe1
1EiLCm5MCgd3gOjOByS+GNxQaFKB4s/t2LmNcKB5OOmTWgB8m10XutwSr/UJNqXtrPIZeLA3+jkm
p5ZpQreQQIlvzyJ2tHF2m0TLfnp6brzm25ptYscCNIKS2AlZFu/dEz8KYIRyw+NPqY4KxE4DxBcO
/9+V3wpbpefjkQs/qOiIVSHyxwBW2Bc/18k10nQx7VauSgLYHkQ2jiS4EFGGlSBrH+gAgBRdLIjF
+dYctSvUb9A7XqR2NDIm1acP+ZF/b1lfKjMLQQ1hBRGafEMIzx2iK59eaJPog+HDqwiA02nF+vXX
3c8ynsYJWt9FT5L+o6jWjSH6JbDjvhsZVi+f+Ry9XoRRJhqP+1q4mRLfxwevzH5AZKvct1SdWjY3
20DoZ/CaClgLzXt9Hol/8c8qRpqSK9qi8FRnppTfAqYNc3F8eqD89jkpdrDb11MlVJ17DdYi6+32
lxEzqX5GQLTNqNP3pwJPRWFMyVHCdKyQgIKmr4LA4KvGBAPAf0OZgmf31z+eAfF1yykTc9oDoqPh
NXGJ+s+/jaRzqWMLbs6bf1U3QR3uVIMA/R4qikbWlS2M+qqkjVrRlMRD1rC3TnZAc9udioeHNQAF
IUt4hTspw2GML6jrJT8Lp0WsUPvr7frJtQvpqgXdFvl2rDTcsxMWeOuRy52JKTnGkGLkwiwxuXgF
bP8M8M5zullJiKpOmJ6jP8Lok+j2Ds2GEc03Wlm4uA+CvUlgetajhIMALHipoL6K3cc64FChauOM
rrS/qPQbLq6MSutv1410AV2Z9vInJIccjRPNsrUPd2kyMHxmD1cwiZx3jeV041JROO/h6VoDPbEw
h8XbHcBYGRlWHYqcZ3cVScMvfRBdrogaVGsFJDsCMpqHH0K8kesQkBGC
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
c+kn4018Y3fsqC8c1BDvdGLSKq8loVyAFSacyvRV4h1D1+Efiv4M6FM7XWyTHQH+G+dmS02vwxM5
q3VOLT2VWqN871HBf5annVWUJlpYOPz9/VWhhcYQwS23zZDmfBkOb1xM6TEBoAn6ZZCG00mdzOQH
B2/y5EujaN7SJBbQpnKD/acMS3Xn7TalFMdJOZsYuMuGTGBqGGE45R1Gvu4z9A5XkS8zA8qfyJbg
GtYn+B0dlG/Jryw8H5qYarQmf5lRACKZExMmu08diBnETuMcR0MaozRjYBsvDA4YFS7NAsjx/eqB
cG1XsQN40yKgVLlxzxp4EnLaWaY+H50eMxRplA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 8736)
8gpeaADLNHvHC+djHuBUVqG2w6RmTOSlen2yXwt1wg9+HfcV2vVBFF/hpUN0bzb0LJe0LSDeTIkm
nxpQkXi91sXSjj5FTnvmcNpcbITNOx2JChnpLbG+hcPlZvhCz4H0qzig/TWbiaomrrSj7iKpvcsr
cbwW7ZrrXu0t0PzvNc8yHSmjQ6DNJgiKL+F40+o35v39h/yXtIbC12BI5GmQBduPVeXOp47Tm+nK
i9kk7MGsMJK+SvrcVW/BZKCFr71fcjTY90UaZDzr+vcQ7ENJRoHo23mINANq5+9fRYgOGLw60IYT
Rl9SFCOYlMnh6Ef2mMiq6whV7v2SG/A1teJrDKqTfEfK/B8YAsIidNr833KaoD0vmMk6LM4Ikj4v
YMKBJXMOJVFNC+d1TmSnKAkmiErwnqlpn2KdVLDPBvKLdUP+TS+k6ZGaM8HDODplfg6Xg/iONEaE
b9ErfjwvjNOeyQND0V6clBmzld/jsYS1u1fU6y+CtKf3h1nqL+P9C2UPap00fxBcp1sFTMhY8yWY
rKrIKa+5RGIEqk8jyI6Ufnz8ERFjn6QVZxq+XkJ7Shj3HcJn7FiFAzwrfIXNu46+WFMYDtScymKF
cHUjRAsaesQrShQuc6s2LYGvvUkf1EgJHkk1i69y8F2C8vemN5RHsIQ0OcJGK/PJS/sViQP0B1oH
kNPCNsZpJxPCOjdFktUY6sd+Oqn7w7wqlbZF8oqQRB16c9rcl1BXxchJ9RZTIXrK2ZvH1E4Hht9M
Z8NXsv3ssTunKOsYFF0dVGYDBS5WSd8NYBFg7TlWwab0+8YHsL4R5tNjqYSl7nBxDEl3+DA/DVly
rrKER0qpeyMmVhM2HFwNansXrAx1K0NxrIqbGvDVhFq7vMepaz3pX7q2w9un8VfXjg9B0fxw/aWc
ixmLBB0yk09jYHqtZnJU2BipwMgQqNcu2pCUkD3UWiKhI7amNqEFIroz+xSiM9Rv3r0QETVGAnma
CLdfK3zxnOmfemLjMu2nkr6dmHRZLBVquTM6E+Y7PIUl3Yl9m2+yX0BmJVUNB0ZXstadeNXyxkBn
yLCYpY5pxVeaT6FeFuungcfDAY6fubVkUVZCCsZkieyaduZ9ORpResVfRpwSUp9lQFM3GmaMUIyN
KNhSRdX8GQGMaUNJw2bdMxMmT7+fCiEu9xE+wUg20gy4fo08tDU9C2yKDNXAYrFDxIwr+AnaP/+3
HTYLGvmD/GYYe72fBopJD3bE1b1w9ZtwIN29XzIRrX74XQPRj0vzlBB1hSus/NY/1ywSbBlYNyN0
UNmgqn73AE9fya9ZwxAiHnVhHC/Irim4G/yEO+KcCgQkxB/pvbaRl55GcdwImnt7+PwCTtLzAoJy
6mtvmnKVpDrvxhwF9xmznHhYEoK+OOxVdgZSmFAMJDTNEBBzdme6C/9yhwqKhPlNxYj/+N1Vnnc/
wxZwSxCkKfCjVBB7xDaalsjsaSXsPTNGIdovYUKKjNf2PeyE8ik05bqAXXujgOFWxxdI3vHKlXCU
GDMeE+OUll/su2JtfBM2q1tlbMos4DtGVKFLZKQYw3GkHpbQkQJrUjfmkBL0qAjGVfA+eI5HfWI9
FP5qSRGwAkt9uW/iiFd/iHdD87D/li3vnGCl6xwDukG2CO/orkRNSAXLGZiSXNGTRuwwMZPRy05l
ifXCSYx0azz86zU5cgPTR6qMizw3Wt+jT9vqLxS+JhMG+rj51kBoIzD8PHvdJ8Bh5Z+69TP5zy5+
I+PZ/JwE51/6LmckECm9zp5wfxsYKymBsyBBi+/IJKyDmdu4DHLUcY2sHNWI+oo2h3P0pWVtODWf
5q1fRh39g5/GQTXonFeewr2C83nWydLgqYyIZj4Gf52o7cq+Hk1wTA+l8fbmpf67XorEVzQYz+mm
c5BahCZHVrYy3rVsMkDOl8kcTNRDfmzUpPFpHEcfj/+wbnInKJb6VDfF6I7hUjG/Hc1mcQQCViJC
bTDxrUlkzdEH4kmjoxLYpQ5G7KiP+XMWQf9Z4ji7gPIY05NBs28VoSjhr3/msLfOzR6W0f5nNW1s
b15KweVJHamfNJ8BbCG6DInUucl+Qqw03YhSgDi61I6e+FS5XUehuJoSFJovR77sM7yG2B0BWEUL
Ot9SgJ4o589QC76TrbfnjSmpWbj/tk4d3Am7LySsmpOa1Z4+hbhqzj7BIbfzrEazPyBtcNzq5pCR
CGPFa3KfbxNB9wl431i6WXXV98szRNkz07nqiEIibmV0urg+6ZQuW4ZnR+IPiReR+EGkcM88UV3r
WXQjhBAMKiEmr+MR9ORkJxAjtBgWGKBSiGktQrzdEv5kC7dMxhUR5r1D63AFdBtoNljtYvV8Twl4
wTjPJFVuFYICXuZYKnrLfgAVuqtBxVo3N+g+a+XWhOpDlElrdZwmXN37b2pdFLfCaWKHfaWNlUaR
BENBG3KbhHWqOgo+DDJZ3PjQQJxFnM1Z+SuDd+Jh3RiB9UtOiCnOx8mjjOPYHdpFfufv177s6Tin
A6LXu5fjZzO0orSoZ0E3kEy2GqEtR5c39Avue6PO3FaC792zU/orOkYGbw4hJO6rQgtK5kpuN9yo
TlQObiFpx3lWIVLWkHE3mQnfOGQD4i8GMI1mWMdiEdSVTDUPHHjZG8MpZtzpUSAUXTdx9UgtUdIY
hT3wfU4TQ5d5RvFX2l8nKj9b+azl1cGEr5wkBS/+jOg8TblqpA+pUILZBL58aWapwlUrxQxa20TC
Xy83bLtgrVn1z6zxmXC10Ug1TXO0litblIjZdkxaVV5NYp8an+12QlKyaSq8VxG1/1+DyFxq3Q+T
q6ukLiq4uE+HYwW0Uo0a1R9Ii5yVBsuFxQhDhCol04qqN+e90DGV9HT3KJr+96/IvrS6LjDcUsPI
kxxd7pL0qUwV/+xSqLSRbJQuHzkSJNBuAz5FNEVw+HfDDUctYYsZHrsxCEaRQqTMX1LdE0It38KR
NWOa8xkkL/hGyNB2I+d/nlx1yjk9jfipZd0k2eRMF0u33y/ugGd5Zumy1KJ62DSBmF+32njp7Iim
ghWCrD7SKM3DVPpuWQ1lLVzu29KG/2MbG2pZDesvkkFc/r+Vz4k2Jz4S8+D4vmqyJ+ZmlLJXPWbc
u4NKsZNxx9fHYgkg9e9J+djY0zLKRBZ8jfTNBlOoKO2o5TROiRI3GugPAUnBY/OjrAJzjoYvfeQw
aIWbqzJ74CSFyDyoJBXiVaSWe07GIb0ebqLgseU7IahUA90ATF8u5OqriIB/+aM7x5wb5eFEmM5Q
4dAmQoBVmcv6xAa3SJimVu+vd+iZhxDOX1gzmNUp6jjho32JZobD+lrG14CewKir9l7uTZIzPb2Z
8SPCkH784MErwiWDCCcHNLZbYEp1tfR+aqstm2uwMwlA+TbtVnXleHsFCRVQZ/pxeR2Eyl1us1ua
4i7fNqsJSMbPgAlkHiYk/ELvL6U5Yk20omuQ3UyXDvfpdtTYozThXuNne3alBE8e4BZWpwX/K2OZ
uszPUMjcVULR8MHvySZRmB10HjgDY/gJ/fmMMUu2gIhfGRjSVwW2lZA5vG49uhMiwi0708a1fuSf
OeHYprwEAW1nSbrvEHVyO6xcO/kRkgESjdMNsrDEa3fTvS5K8upPAbVukW7UwznWWqTm+r7A8Dip
VsMgds5pJJ0JGAfnW1wiGtr+XteGk03nF6wcT5eU5JM1+m54dLh1AtgyXEaYBadpb0M5en4XIUuT
37CvFCfu54rlzZqFoIEvSFl3RBPKBZFK8rqlvbyHUM5v+4+q2wjPNIyzPQEmz5Ig4GdGbN2Za/VD
2zBSuepqneH4SVN9FEMI4N6b7ZDM9EyZcd/eAot535Jf21baN8WoEb+yo4jHF09T95hE5NPLo9/b
605+mPs0YjI4Fg0p3XdxhsrT/qycniAO/jKL4K+sdKiFsrOhg383wG228xkPnaJOF1Lquo/tjN2K
/g3gSdnKLOvnxBPlYarXbQMFcCt29qn6uL2EJjSyp4pBAhe5JPDzDjF4YMSU3PAsD1lUeAcfVIs1
78e5ySfGmwhDI+Rm26P4JH0rT3LRjtxw7z1aKOXTJmAiqDIhtfOc5l2QB6RIMB+rQfkLZrRYqYqZ
HxS45U2kMOmFq9QNlt6Al2Phnc3P0AW2+Ijeu2G5AHkmuOPA8sjhPcz4bf8jCgMVqzmiRVpwbHtL
ATQal3Sa4FR+X9LjBMu75Onw5qAriXJz9pMN3X8UVlkxC72LGOoxupoBxD76IMlD170dencAAUCv
wxnsKYnTKcQV2sIYn1CWc/xjxWc0ld87F1lLeCSCIqM467Bg9kZ/PCUYA5ssterPC5CWAPQ+OX/V
w9bRP8etashJqeVB9Ubyv0iv8/xI7ouZOFx8NetYo6BHE5RkK1NIRcUJbYBvLEITnGig9sIItmYX
xrXDzj3y7xCGrfMWYGgCcH/YkHqa29rEcTQeEqyvvk8Rvt6ul+KV77tGWczK2k9xRuT95zw5Vh+G
O1oY0HmUczLD5mJ2cr6T0vYHn/kSa/3FPYgJcKnTf1v0/M07wG1rYt6FejGcQq+glkIfa7ToFf6i
pAeTPEMQkQBUEyqfFPo3r1bhVJfzmVTs8P5J/00TdIEox5cePfXszB76mno/iWFW2sz2x2XB13nS
2L81aTFsc9OG3/kYgyVeCTDhZi3hSm0syPoNzQrloc6MsaIPiq/BOerBIPutGQVyfwBRsDOi5POY
BUa3aKedWQqPcjfZcI13lttixvXFS6BPzSwyof73KXYxpmFsl4K+zm9oHaR1wT5VIKKKMpszFOGI
ICkJltE0D2neiNx2keoG66b62y+z6l1YRB6NNBxi+JHcipW5lK6gEIDF0Vx6MfRP5klczl9Ipinx
bPwg6eQMeHRPONQot8y+v7YXPaHBSJl4oygn17Az2knvfkLwHYV4UboJarKkJf3Q54XcdcQJxmYn
HDNBpEpf5W8TwD23qWzmoLJ6AmmPDDetrAyhAt7v8JfC5tPxWDwlCxNOJIfI1azYdpsGG5aFFTlC
ZG6km15qKnNNflxly/DRVLtR8xOAZecvEhJfIWJ1mLOKsdArsiiJqBhwehR2dCUztgsLy+fuBhth
54NKHlSFsgJyroSZAa/JTEOvUV/pd2V4eu3HF1JZehaDUR5ujT6liZweMFiOaKUwNmvTvDkZQkUf
vShg1XK6d6IspOsp2KXxSnstbh4E9k9yzauW/o6xWHBNlR6l7zV7D2kLbUDejtV6OtuuRm8+TC01
SHAgu8Utr/1sDsf4HSXIWs7DWP4dAMjQ41D2KoRZB4FQDYDv/SY0R460tWxNA8EelxvdcK8/CAp2
WrIjsj0Dg69uTJEBzNB/vE6JlyWim22foIRsYF8TEMVhwP795N0FAnjuBLpYMiJnwrwZu8HtD6sP
qlGtgTax62L29amwpXgKVfBoLksGcbckVOBdW32EldcArTcCB/4jZ1+BzzZS3s7I34P+BoD1HVq7
2CfBsOKq3T6V/wwCUQ3GFEpY1ovf7/lRLZ55PFcI9q97w6RwKPNfidElVD0iEuyccS7zKtuG1Xgt
ks8yT073vjB3AauS8LpYhsW3xR4p4bS8ClNcoJKQ5uWoxRikj/MYIhqFoDLokDxfs8ZkWZUK8WZt
SheKeNilxcxFFHFhbmdcPVojVGseP74HvrM1mgNlr5Jw3CE3vMrjBL0G8RF7TBtwg0rN9qlKYShT
tfgucUEEf4AzAsE668G5RK7pWdaO215zcrby6MnBhditE/qYab/IV8dckBkyQmP1iqOPHRVHYyuY
Tyrs1r2ebXLwHBmTfRWjKG4YAdP26wAhCheWW/5qfPupObhhdwHtWa/WG9Y4cfAO+OjE+pqOlJFu
+6Ze5LShBn8ki9HFkX+pgqB7U3WduVlNFhiXrranrAft9xVnCm9kUjQVpqHRJqzkTzAjdTYFJGkA
T8Uxb4WoAkBPyvG5TvjtYQBs30BGOUqFqmOTC129C2hEaRUhHKTsV1mb9f13O/XqRoO9k9Mk0HsD
C+q1MGYOLyrEE4bDPRwbZpbIgNmHcXgz5S21nRsRorrUCM9WVem88VEMVm8mxOnqepXEgtfc/cZI
RhOrpPD4SWeStSWoo7VGfz4kl0VHzkFii5Y8/QarKjajwksB1Qif8ym6x9JLdVfxhJhnhncK4ji8
J3plE4dZBXYwt/DLGgojGa9e6VSzn2R5apAwUZEwVemWbsVReSJKolrCbkoS+fRkSaP3KdK3iS3i
wq07/5OQX3+E57JdbJFCAauWfEwoMmfSrjki1MlVAl+b+acqieesBDh0Zd9Oovfho36Ox9oBsD8i
/MWF1hHbqSZX/B2G0NWAoXGuJF0GYv1KnITB0LqL3wwtWVzG7xcnaUYcSnrrmBaBttvARPyx6Yrq
t74p6PLLu+YcN9JcyCKl5aLtz3aJF8+W18rxe3zw4Gu+rFi2iGfYFpAmPgHuoYBxti5qwC6cMNdf
MjTavqQ7cNjjWCCfHr+MMg26cWUleX4YuImOxGWunkMzP+mLSDTi4qiphxfAUomF2BnZ8/95dt73
6P+tKK2uPRjSVXG0pSlTyQyUtfkGDsc1XumcSlYk3Kfb0cPbQFt1dCH+qX5Z5TblpT2w6l7P+B3+
TKD6+No/a8/aOEdBMpUjJEvkfrFSNBm3aExnPf147GuI0v+gfsPad8gTvfTE0M83e7uh6R7EE2XN
GXmPKsd2WDtKZx6MGIAO+yeYJBWeVmoL9LGEzcdSaRXTpRb/4kXY9SBCBOtRtAl1qRTHF6u4W8Ey
TNcXxWNFznSAHxX/5Gmy48ODgchVA6jxUI4gnlbaFhqAzT+QAY/ivd5tEcndXvpRBKfUi6iBoBhd
zMCCzaFgnPvXZhihjyXnRaNA1Mf/I3oWG59NFWb/TuVR9DgbQ5PqDTHEFtemxWUjxFxXwPB3JH0L
pwv9vDeCwFk/Wrp4OHhrqZVyG3vncneSvRm4tanVlbneJm+35mZzjF3PgVvfKzZeiG+U3PSMZRIh
69DxbQn8cNFxqT9rG6i1yIWuuQ/QoUk/vbG8EoAzys7HI87rBqCrvl/sgFVkvctcImJyacjZmJd6
hVU/RVjHeQCsjOmlC1XixH2pu4758CTSc0YasoE9D21cX71Evyd6Fs4bdPTLaoEb7cGMFJRcsiAD
yYlnMpJo6QAYXDahDa3cIS2+JS5LGDnOmbpbJ5NHuI4ASygAKcuYcRkI29ESz3KUsrENwDTOSP1a
aQQ0OsunItAlEfeTmP8SBZtUmvopO9RukhJ/QtTKra6LOh3EMth880i9uBsIkucZevxvurM7Ey7l
/d+55VYmWnw9r+wyOaGlZ/pub5arFuWTu89PlcXsXEuDVOJlEkvp53r+v3uqZfrHmUzyqdJKxJ34
aqEzz5lbrbqLHIwZyD1f/PiVyJVtkNl2zer4BGhI/vflffHniEkXn4esfvdzj1T62SadvSnIXwJD
F0BgUngw4C4O7egpwxPqjq6zb0KzzyhaPLvpGDrkfyZy5byZNF1eZW7NfihKLt1+MkCCMPTZuDau
HFAtLdxoJ25Z5SeIKkBxcleq9A/HK1vS63JAZ4bnYm2Y+eeGx4oHEdKTTzgrPvpKEFNgXFMsKBew
plVT9DXZnrvFchIy+NOfsTjw6xKohJrTf0JfVpnKOCW+zuycB8M6+8A9JeGIQkUpnrr5t/PkCdHC
aEZNmwuqP0oQMrLTnHTc5t4OSR2pptKQ4I67xvT/d084Q4EtbUYRu0b8MXycdvXVqa3crPumvj5S
yQGp4+aBM7TuiINRlzjtVmrUNbXAtDD6lBNnscFEIyXE+sQ8JFAth6TfkD0f9zp5E89OrPHrXmuj
g9BJLjSmx38w1KHCi9BWhl+k5nJaGbkKYPJoFgfykPw1wDVQtcd+QN+wL8MHfc2Nhbgb0RenxCw8
uMTcFR4lK9R+OI9QATvN2jJhwhXX7H9Sk1zJXcdsoNQmz5VsuYTzPWNAh7VCOcXJ2WYcTKdXyfJ5
FTwIOj/hyD9Z+KQ56u1a8/yS+Ovc66yz6Q1lCD/nzFNSKjgUQiYszeN1xM4//fGaHL0esBAQ/6c/
hbYCRw+uhhWWzHZ+oxyTCFx3l3SZSfaKwrnf8dmqj7QzFtJDGknv/0cnN/jY9icg7D9tjKMN3YoD
lguPSDYVmkd1miXmbBhteyJsjfTEQwPtkvUBo5kLhT+9IhWf1Zs5UwMYqySI/F5VSSD9suk2cUD8
JMUvn2GlQwlIYU9AJRdG8nvWQ5Gt3SIEYEuNSFkMYM9toENIzT1k6TvZBabVpWsyZi94fuzSw+3T
2/Sen72OhV1cJ5uUiqvlJHY1s0mouruA1rBlsQJlcE03nhAmSuJVJIt/1MutwZuVwvl7arBjr9SM
vhp6ygcgk4iX/Lf1hFhx/kS3rvhq7Wz0eAH8SPc0idStMOfUY6V74jUv1YtG21i1L9nEIv518T3a
yqnoyKAfbcLmr5maNaSU4e0B84Ib4pcQ5vyYXGVfYdlRmMpqOmcTbNKvB3h2QY/kvQ5HoA+gw1uo
yI5Jg1VQilcz5fTXcswJfNjwnpVSXmvjcMreU6KxYWoclvzjtEUyRXNm1tjapxKk8c7GjXKYKa1g
vAjFlxSfr7tRmrOSq1nbOIEm7TeJsf2EZ+Pb/Uv13X6BhN0CSwpmFuXVEUKZsA3SjaDdQ/gag17m
P3q7p2TO4HAEomd/Gdlg6v7cf6iKZbaO0FEt/3YvuSP/zj/iXbNhs/JxjVM2YWCJX19NXWI/ijZd
y1MQ3Wd7lBuVP00uH17yxLzuptm30hkdMfAZce3nIE1rfx3YkE07mfkI9a9Y0+chLXilI+qW9RCZ
s7dUujC5h5k6BDfnDUKCzwN3BFJXPP8yyqh4HYviq5b5bN2j9QQPHQNapPtsTISaPsd2E5BY2utR
aDeM8dQsUX7Ny5u5J1kja0q10vKYd/uGJPTfJzTY4+e7AvwvtV/qPdxA3soLIMqEE7glSvp6Yjbk
XZDVqXYipJMrXRy1uJJV+OQnMivYBo/B8osfd9cG7W+4oBGVpzObiyme0883c5B9j5PY56Vn9Sfn
TB9xC6SpOeZ2/+klb3sXQDvxPwZrv+c1VKDlG4RA9YWM2u3JNAYJjNLmNxPJQd9tuaFEJyq0hU+U
q5pQ0IvVJTojzn0PK+f89FLwejutfn1HCsiQr0Ho22Y/Zx3/5gMWBLAeA8ZoXZhhojFT4bPRrVcJ
HWPw6S6KHK0z4S6f0uGjqzCLGWeVDUUCpFfa8ibKYnucD4YmV05Iy7h+uSuxfVITt2QVmCRqupSN
XM/4mAni4yPLVAmhTc3AuQLdzfZqloEvDIUABb0mn4SkAadDgqDsro3hviqFNY12MrAZGYES1oxy
p/IYNrf1QF8XmviNTlI5DUpsG4CE9wPpKkYx/mWJTauY6lL+DHV5rs9n0PSjCdkXXhVommPIUou3
Xs5pCMMrR/QvuCVrzu2EOe17Yhrxlt7FUxdcnbsb0tkuL0niKAedfrDgmvByUMXVNE/nMUTC2N/e
0zO7Ytd427g3gUZisrI5uQEo8dJ+3L6ArCwDq1aFvr6cr6f0FIQpvsnni6ZlbCf/LYZ+ywE4fRue
/9qf1poBZEPvRf9Fx5DKPC1qBm1JcKPsAoBWC88Ptqf4Xbxl6EEYOUP9IMIwwTlCN/4wMEdF3tlh
ZuEQZz6n2yI1U1rDr++h2sFaD/gvwIXRWq4c7nY/He4aGKwNqHaCtR2NseaEv/17VdQsrAqVJ0Yx
AFenEFhusX5nW9jRP7JeDjglSXIzfn9UfwjR1mZGz1ZfFRETF7Hfb9siZX9Ft4W8v/WPAm38e9st
y0IwVcrMA4EVtQwyzYzJbeMAjax+7aiH4fyKlcIuNerm0i2itXZC/mWlq2SsQJRNeY6Xp7IgLUmU
PyCHeVKECOuKquWAKD7t7xPN8lyqL2iGzbcDDfTmkaEZdc96p4y+Tn845TIvctOrHSwGagb+IWAm
aOg6wPIsSFeit5ztdFMy6MHSmtlHL0kZCtFinGqvNWFsIXKe2fda0CCn26jBt7/2mNnT2m1w+oXD
xAVS3+pZ3UixypBEQiQIaIk3H5s8z9ErI5/x7zlIA2it5DaJakP7kmCpxZPimEcGYcIO88sTgaoP
LGuAJrwz/UO2SLVIC/ip7RrqNrYW7z2RMouUPO11GuRjuzffDgEDJxKQvoVMk9kS7OsL9KlyOMFN
69Ft2H+7Zdy/cquUM2vmxlAIkpMEPEro/kjPZdlrS4kwcIxKscqzodar5Jz9+mmZILuR22xjsxQl
PzgQ6gane9G7b8xnN7x0w/7wmwArUV5yltJ8BJbx9/Xj6LNsb7ZPZfm3la4wkvrlkUJhUBJS/dK0
IFRWeetnDL7+K2cX/BDX5VeYUaT28U98ubF0rAxbVonTQTuhNHL19dvo4ph2cwxIPyCM3VaEKWqu
mZa4Wy/N08yC7e4Ta8zlNt3wnDQlGY0FscS6gSOGxQx0x3t1VgIxjOJHij7MDQ4HQoOq2fIBhNGB
H8absIxQjd56bL+QEq9Kmot7BbPptfBr22QmgYTHcvvB4mjIrXu4YftOOvt42Vlx5fUR96GarSIL
YPpvC08haCdKZJ2C9ixDoWhHwv/tLQVrK3cPtiXcBwldoU5onWV+RnUVopGtOGXj9Z/vf3O2J9aE
pBh6RZJk8w0b+Q3CLpNbVGThU32rh76FJc4Axb6fidrt9+TRwYSkqvMWvH13NC/aEc9iWf5WXMjK
aN13rYGPt40citeBcXTvbP5kx8pR8QNe5dayu/JkXjXPk9g7QypyXvbdWNVuQlvsAlrdf4B22uvv
2HjNtzZlQA9PGxdGCu8JXseYADtKosWRclU4mBsu2DPzFrfCtDCAXPbBT65HOivFKwseUInwY7m5
9Hq/2NnYi3Dyvuu6QvLuYH6Hp+6VRTkRmDTpEwx/2yo9zv9CwfWx2Sh9WxEuowcRoSMPkTJGJPjQ
p3/mmjfUM02HpEW/MWTz399uIKXqoApFRHNTAa4rWlze5MAqL1Np8+3V2v9mDcrCMOESSWnImUzQ
KpMO+C9AC5WnD1O26gDtUccV2UVZ9g/7Fx2oOTaer+WtWQ85pjGvY/aSXakfq+zRy/SzjN/03BAU
Q6eud+TswG7x15NLGiBBPe25V5QjPw/xur0gdsO5ChwfoeOp0yXMhmSvE6kb3YReBKUpn0rmq2gV
tV8EFfFTfzYZSPmGk9Yaal7h2G399luM5WzsKDYzy9pnztJjyYwrTzLOBoACxkFOhMFopiSHoQxP
DcJC+ffnLzSOeF8vh5UyOHMLi4o1pgTz3XUA06FZjmfsc5Wx5SMvzlCO/C2Eim2ian5vKiXucmFc
goD0FFwig1T50HmEA9wdZ53llmLASvGBJVBJDlV8DRoKVB8TJeWWqZpfgpbcpPK+8kFojMw70r2E
kVi4VBbY4cYPhe4O6sQq+4mLmklTR6e16A4amGUCk6sk+0883MOwgyjw0huHVY6AxXmFNlQK7/++
vWMulP8OD/KYHn004/G7Wf/k4l9y/vubWTyQVQEAiCEAi26J8Xt/MEg8RaGGHaq2JrMDpccRkgvd
IuuRCH182oGR0hYFWkm6G/AI0pkiu43JD9DT4b0jlC20BX3jn/z/Dbz1WEXAcbLSAUjt4hWL23au
Ud7jMMj4MqobN6I0ZrSD
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
4VV4wIUIVEGpw3ecCT3EdL5DHKEk6QPz+nVjYT07VXkXax9ljlJGj9Q4TMGPwygd
YVjK3KDyP0OiUTmVUUBiyv/4VZCzyyJRx2QxIh+lygQk9wVbLZaKXLVYWg4FBXnN
dsRsNo2C8/uXdTX5z4uGbsZ5wlAKe+Nt/5SiynSkniI=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 4528 )
`pragma protect data_block
aT8oPg3oqPR+OklsfNsS/lwqgmDznrvAW76QpBkcUq69rQqNk9vQ57+r0Jyu+43T
oc+/pkeox5PuFaFtvor8KwUGuT3W7tc7UvOXEhXNwfK6B4iyEYxSJPeI91c5IZCC
+DzrIswEDpDNATUuSTw/Sl8rhdzVtVKXtEqBkvLHKewYrhEKxaH6l0gbnt0Rt1EV
uF7+vv3rYsxssbqD2omHyA1snushMfa2+wUPj5aQhl3h+dpfnkhaNV7uLW0jjq4U
gbo1yPXSA+Yt1BLu5XPy6RqQgNknXr5RPR/JAh7lyWQsGbrKghEzlxK64TJeFwDm
2Cinw4YEgnkfdeMWhb2FMwK+zrFa5BaanIjNCyfl3bAstW06D2OdFr49vxLjgToW
AqV9bZKyxG52DEJi8LAGJHpwiFZ7ZV31eW4Wo+xqbzzDtTZcVe7/1ej2o0z4uXq8
MU9YOZYT7Xf1+zJjZz+F/Q9xmAnnafrXnO59mDdTenGMp3MFpeclweWMmjUG8cvC
JNZ2BXPgBl+4C7KmIJgHvDqpaeXE8GwwZA/ives98KcAVPfPqJobom2tn0gGpwbQ
/FLvU0sZTJxOvzzgqFsthkvcKJDeuOGCeRxjKYyAjWQiHxrfVyoAJVnyl5USgl6k
ciVfIUQ2M52JkoS9Qfq7Jmbe316tO+8itk/dVz34Tsnq+9IPIw87rZVNnWo/T1Gr
P5L+gMquych3ct6aZSRCp2pOLXhcawYn4w1udjXXSiq7+fuocbQ4V5S8OZ0Xr9z7
yDWeYX8nd44yV4FLw9nLQy30AOd+ROgdCL+MS8MaJYHwVyl/snBmdO5ec6Qokmtc
NgMRcu+sRplF+0MM2pGtb2g8u4QpjztZtpojSrfhbGn3Wo62cdJzUx6lyPqNoVSf
sf+P6E0kKt4/A4SLgyvNGAPzp4tmgd2NDLLyukso/JT76+voJ08Pj/s6AAXBjq/f
IvJ7VQUXIYa1oPAaYktNUn0x6MQ+w0+iBW09kJKy3pLIPu19xRatXeVsFqBA9tY/
sjnvy6UsBerwWVDTmGfUWSl7o5dJoAd/9eNeNa82lzvxP/yYE34NGZ/0cZzkRc0X
qhftyleU5a695Y2CO+2F4sOhgyyfq1qBss8+E2qT4shMa49jLIt+w2yMVZYguTAy
fu5zxDdDyE/lqDfKenp+sea4HnW9ne1ZgNzTmcKEtUKjqPc4umu/73Raaytr2yig
U77F0JJCvQK3Z27XuZmd4BPaXRMJm3sqgptb78lQgsW5nvTRrTWHLythHNnNAzIt
dJA9zDqQUFT9TSGF4yoabPllM0Q1cmXvoIR0H3daaOI4btfH25HOQ3h1Dczr4TWj
ml1CUk+DlmohknbIomL8tqfTgaxUBPpbcZ3D8uyuO9RnO3rL6SSSEBPtXecY9PX0
tXi4SuoZ+5XFwhDFny6UJO8iJbkG51JBiM0sBAV20Z99QKi3bHk/iu2EY/7Ge7t2
oGA7qjHpWrgPmiomjVdwgeXZ7EjIbwE6bFxUyqOG5s/3rzcXTJQ46bksC5FWEDu+
s75s3zUvXmC7dJnlQteCUjctqqDm2CMtnyfh0WnY8oT1fBLLU9o/o+69IR1q4BZo
k72B64zW9HLAnA17FkjZ/jHYmd54M3yrFRWm2CoCpwTmrMIDmXfqJjzE8Y+8kuqP
W8JWdEN3FFHnulqbNRP35KuF9kJztIUfwLZzcactp5dM8DRgRyc3KFBZ7NuNf0SK
WFWDOF1LnWxOvNw97g6bt2PkAFIALXd25KHq1Z7cLfaQIQ4TXAXfgfV0emOkbWE5
7rKEPgIvItzZqis+2oZt9ezpnek+TPddj2GEwtzyvjnDAR57iFG/TWOSv5IYDNE0
AzQoWzuwoEAfA9i8FsKfZwSO0HyAk186YSzHpLIszIGTqsg2+gabIhxoZIPsTa5R
PjOthiI4b+3OXrryvgBSD1e3wfJMaVE5k8clb4v2+/KzWayNxnn02WsA6sE+tkg3
ddmiziSQ4DPauDKwYUbAd4ZkhAbwHiortrQnIAyyMbvsuB1EbM4EBRV5w7/acLrN
hn5lViLpzUhECmE99gWPtsFmsk06tW4g0b8xiHGwqAa9kfg25tHUWfUXSXVdodKu
fRr1mzgGNKIh5LUMBIeQ3InlvPoZy6FR6rGnw4oMfK/2YPvGyXhW0UQm+yHaVB+C
mXkHg161uWn5Ldqm+hgzi0RP4N0XNla+48Y4AXDMKkptSg9a0OajF0+0yVHym5TS
OO1Rbtu+aOsE8I70NSKw52SXPrD5sEjoYOAyJ8XOkwyJaMWd3SgM4kycOSInka58
aGRgEilVIGORSUz4BT77ZKdy6P+inLZ9aGDmWi8LJM3RcSBpcY8YCWsl8BbffHIZ
NHV9U3Afy2n8MAVu6nt2eDn6ecgrv7/5EsPFIfu7rK9BwqlbFMPp0wlGt5M7Thng
qnS0EBtqqzHXl0Ue3LJEisyeDFCF/FgmCDNepUKnj4NMv7nGk5W1wVudw7UevNjQ
N6ShC3emcuG/W83/ZpWgsy3tHAl2CQI1J0lAXjXZXJ/wcb2fNAFkjfT1DZ/Ui47X
j6S1CedgXxmVZz6enNX3eajhsRV1b1a5QyJ5aM/KbFWQqdKc5tN6CTHPte9Ag1GN
aBc+KTaypP/92R3cAForSvDBDaWCTXR3WPIl3MuFIslKk8z8Ax2DpXfad+e0t4Il
xCN6alM12Rz80wIeUFBccf76IXtnVRhtqg4qUQ5933r4wj6YpoziT8OpwpK+AcGl
BjioU/Ul01h2nmjgMpuv2yJR6OD6sWNnziItRb4zGIRGRbB/kdZtZz1nQIJRf1td
CcqQUSVkR3y+YlS6RB/XRGYTfyZvRJsGWhf4/aFHvgVqTP4wjt/kLyTAsRcZV79S
tIZGs37o0hPU7PXA5CoFwrePXKGtykxQ01LiwSw7J5oUaJi5oNv8Z8XUMb8lKMD9
yRVLeSmxVGj0r5xz9j5upmnbuf7djqKdwiXqqGazxKqGHk052dTxGZxtY99/smwF
D+4l+iQaKxRiFR6FZ27wQEMZfJ8qogNkWDBcz/fFW86hkUtQBe/dnAoMUzbEPofy
cckaP4OLJ99NfMBF58uLyBe91Z5q+vFlWioh0cpE9SeISOpB8f0R8cnF8/++zTl1
hUPjgf8HhtOv/tYrWsMff2rBrvUexWrf/hsDO7TOP1wpoC63gM7aLof7el4kN895
lBUJ9ZybCIf4CHxiiCSJcKPgo9eh3W7SACbtgdf6ORDfMtIPeS1BSHq2p+RUOZfH
hZuUCCao2o5aLVHnm37oeVi9aMZPzJcCscE6QmYtqxzW7M50Njsy1tXyOYgYgM7t
bDWQWMkTmjkWwxgIuKYdTdOBlwilf0oJoY/Udhnui1AoBxsQWh8VmSNInbNThRHX
3XtiQQVS0xP0Au+AG5mb2o2tElmgb9FCBiyEOgiJ1NhHpnYCPTtnon1ZWaib90dN
Hol/1o1xWKudv8VyDu48Rdep7UY6qH0R0RVGuSka720grOiiLphId+q+ms0Gzi2l
VF+eLTXcRvgwfNu1B8qZVuoqZStUpVPB2AIybwIX6aIPgtneesInIVWGu+7rMz8u
YUBhYbPoxJLvOKVSJSY3J+ckCwMDHUeScZitaSzKegAy4K7Xa6jWsEO3xZ9+fVip
EUiQFdY8StnbDk/AqxWuCVRlbTozbbem0ocZes8F2YaWByIPk8enD0V7nEd6h/90
2YlJiPWOOShTrEphzKF+grKWKRIeyeaZbfNcf5K8XDAFd1naBN334tE4egajAIFU
15jhYkowyVU6mjfNBwrTBy+ys00YOQHI7KMkAXecX/Wj3UJd68t6idOBDHELwXbW
KneHO1Jr4R2KlyVGAhi8lFvPQ1UgZZcmWFnucYxlMubK+ndprxBumtftTDsLnusn
DZ9dSqisbN/VU7kbSzp221+vKBcak4W3w1/iaK0V6cUykswzfESKAyKV6J+ZysbH
LTwfoTad90MMcDw2lEIMuIWm1CzxA6vTWXiGTVs3Mx/jr21cGMPWRInMUU/7miib
lrsfG1dU0DNTIPSMSlxX87jTnWmPGJAVxNU9+W1Uh2ZNaSQ3u0U+joqIu0kGkquQ
Z3y6gKUpIAEGr5+zxo3ZoySdgIOmksiUswt48QwWvvNri2zI4sc0waIa1ggSnThE
YchLggEvhqHpY1c8tflPXvgwhrhqza8p88oA+8u+A0pHZ4QZerfiDKDjeN9038uo
/b6qx0IQ3jJsDLxK0fViLNdwO9rGWcF1IePtMyRstaKvx3fzWtoS+A6VLLB181oL
UsicdElh6b7bXMgHzNy+q7sCbBP5ViYt5J2ZGtd60K0l15yN2NVItbRvNdjGgfww
8H2DAyO5jbs10XF7saQjyFDiWDDSM8tJhWD2/Nl9JJ0mEY4nt2o4tAyZqM/Ox+Dh
snD3xIQB4DHelgYO/JGo1srnjR2ksnSq4Kq7yHFda+xTgCDUSYwQXnpuSWT9zJTE
DiEWsHEgTfLyszsXQ3KO3x+K8/LgCCQMlvlb1yVcDvB/XvXwQ1hrJCjfVBtVwruz
OS1iUb9W8dYVXA3YF1fr5SjQ37SiTiGlrUZ0r9cROeCDn2Q6iXWxTeBj2cJ0p7Zq
og9hLVaE7UZmpCGupB+KaaqQlmrCxw6KsdEeS7D0LrLgyxtjYdqu+cb9gUy/V42W
ZkJbmrP/S3J8nMnI3I4DB/VIWSbS6607RpFAmJaiHKs3piEH9C63/EOlBGs0x2qK
qPoMauLDWrU/DBQLpYhy+bmz5f9ly06ZHy6QTu5pibcnPjR/B3MrSVEFoRJHB08d
0tpHmrcnJBCb/NumnJKH8BK3+6jFscR+MzeV2JRZGoXhx+f1xe/omC/s0JG44US2
POCBGazupKtxB9zLiVkjOX1ETbXXtZmv1pCdBa+5jN9YY6QZRUz+m1mPXUA+ZMex
WdOVB98GJUj2jVTSGb/4yjI6fqrbojHR6976sX8tFGCj0Ph+6IHfp7tZOdcZfbot
8kG3ceOyKsANjNc7CB9Yi/KFawZbMJob6GICl9msRZYcwlSxRNfDDhSUG3H4HWfW
fj2RkGGaL/c1ls7WALHhgX87oFqjNJ0oj3/EXDKIhVfIzxnMpagPaWIl2/xPZ72h
K8iGexRrJXnKPO99/jXBCHpGPdxzT72xiz0Pr2FaZ9PSpjy8cfWC5aw8uP73JeFD
HEpwvTZZlE1moYHssMoc5ZjYfYu3M6e8ThKj9jqHhU9veW6WE+pK9nhB9UTV0hA5
S8MPmuTAeoSYT4b6HPfL028iUrjCl+p3N1T5Ji2zB/iQYpt9+4itI5vtDP/MTGKU
JZ10p6V1csBe7emipo5ALCc5MrviMiVsLca6d18RnNlgZMIs/yU7zhJWShnCZR0L
DMLotrZn9oiqqZE7kUrJEN1ujgDR+rG8Up2O1/UVyE7C2qlkcZG/9mquQjj/7FUt
sUcxBaV97NT2Cv+5vp7hLUA8aI4lQ/Lp075YNx9NhFZfZdQVW92xOoTHkPjSnITk
3TRau7ALDVkWuhgTN53xp+F+FFNcrx7b3YWhzDkr52Xp70uK6cg93dERE9iTsl5W
LCudB7A3SCoow/Us3VqE7LzYUAlwUxo+IhvqHV5U75CTcs5qiB4HZPL0Va8gHfFk
v6tzKjTkKMnA64DLkOJNreWWRrk9DfXy2CziIAVVfEXIXqgGB0aaDViIO5A2vTMp
MYXKYgcPp0TVD8Ifb/WnarPAlHgWMWp9jfyLwPo1wKU3ONhG9sJjbcXIj10MtjAg
h7jbmEPG4Q8xCehIbmgZA3WopY3xBYiN7EQMj1RvtLy8LXLQfSzRujZNsfN864Ys
WNGwCYiDYXBIh0A091T0Coj8T67jySHAiA29F8x56OQpRy3OCtvTIMIz/e8ZCoA5
thdYrIh9VRs+t3gDH10eCw6sCuR81tsCSuRZQk3hS+hj3QMKsKzmbi/zLAZ52iQ7
n+JmZXPi60bUumeJ2pV+xg/HZYS8vPka6EsCbLnd6zghrqqgvbOVYjty5NcnkQmB
AReu0ZBNEWDW01/5AuzwgA==

`pragma protect end_protected

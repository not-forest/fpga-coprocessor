// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
O9fn9BVDhtVBcmTTeUSvn8fwj0M7JbcxF39DMCmrn8oEchxGCglITFuI4/ceauZC05DH1SNLJTBJ
vviOJ+6ZbPQf+PDwz/x5/c8z4QNhZPxFhLIov7lcwebxH1ouuL3mUTEWv95Q7tmqT8FsiV/5XFBy
ziDnNkfgyhjxWYQak3jW3ZAyFO2jCZyMkKFOmamvESERbSzZ1ewv+HWY3k3A3dmvhPTwv7t/f9IN
cmq3oREHxwpF++NGpAOJExrYRJPTzdHwsRsH50g/hCkRf8AXJCqg6YqMcMvYUHLlOhi5il4KHUKe
aXtI5yXUEB+LjbU2uopt2QC2txH4DCq2/I1zUQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 9216)
4sxRJY9CIOhqlhPm/cNIUOGeye47v6cDFJNCfrqbIa63DGROX2xvoKVl8VVTZrhHhMf3oeNiOC+S
dzcysYA6rvwfJpCAZUzh5e7gthf6/h2IWmBzJt7LrKFohkTDDTO/voGR0oCIAc70pBljLU+QJ2g5
9B+pNxl/KFe4qKeRBEzaykdmr3w1x1Pnt1kBcrFhapp3DHUXdUagmV0rHSHqKhIBr7/ana+M9JEk
T7Qie3zNP1CWVgdEvYzh+U4xSgqhRwYm1f26ATGky5w5et+ZsI/5DG/7HUxxDE3nxNh67E5OFY3S
SowocBk2MwDAWVb+KJs/5gEjZk9fjnXMl9NIS0siyfNlmZmL81XH94GoclQOqSM6lsj4TdF4qxsX
omnFqee53jWOhdLetC0RnDqJqpx3CHfAC2T1A82h1BJVZRhWoH699l74fOZ70ebiYbJNAHEKj4Q9
FBxJVbeJMxP/nhQgOnpHLzCqE/HKELYwXGGESx3+s8O6FJLAUcBS+EBApW2BKXLsMpgIu7n85FLU
sZtX17af8az+0NeLWpGMU1Pi1oxREInhg4n1E6gy/W1CNSXJtlczvvmfofX9KAkIarg59U2GKJ2T
dlxccrYx46earw2MpAK3sY/h6Q9htlajkaPvj2x+4wXgDisEVXMDS/grW3yQ4siM5BjZ08j6xNXF
EQEhH9nk0HeM5vb/d0DgMf+hA2eUbK16WBoC4WxrYNvU011j+8JjdyGZl9vNNUXmCfFA7Q3xI9Xx
DYtjcwE9PbGXxxMJ8OFxKxhpgSNgyjNS64DpLHwIfSe86bdq3L0lT2k9x6SP6lbrjVFJ8CfVncTt
tfnzPxYyNoqK0fpaMugF5fko6fxNjpbPzzJbYKZ+HPhXAn2bVrjT+6mxaz8x3jGaBKJGf9unUeDm
0MhXm9INv1bLV4S/Tao8OIZ2RFGSm+6NqXHzDE/TY/Brwag0vCV4pBADbkNHwRLdVUlN9IWS8sCZ
aUtV3Upfp5l8i7hpfvRA1WLCx5oedBxCFLTyKVmfkIO7V3OXUG3n8iL7MW1i+grmVaAzj9trFcck
Sgi5QilyaHRg08bzGpIeKoTAciti6v0sCp2iBUMVsQhvGWdQrMOxGoxXef9E528mZiO4La405bpA
pwiBQRB1ayS8cJnxEYoCVUU5Wa1NW1349/odRcwsQ6u62SCFmCr4krqUJEFp7wox6wydVNrTt9QK
KlHzFdwiVQqi75emwH9or7vO4vwKGvAb0QdJyYT1AUvKPNP/fv3I9YdvzOnuCGxRizQM5ziyKGy2
uHKXMHb/O+ixKEyx63jlv7B5f5yPehKeGcx4X2asnXVhU8MS9df34RXILq8YmXjrWpwfcunedvGA
c+A1x09nMTwTYZMUG32T5pnAbnSx5LMlx4XHniczMkINf1gBvued9jr3i3GkBCRn8ts+oEPieMqe
HkxeofiX8kzDx+LYP3IMN2zlqw+I+ufPV5rfu62KkX42RDRSIev0Y6RUo9tA83CX5ynf0BCrtPmb
OlJN1N5moEvBGSqodkvkVnc/H/OujLPFScEYhg0L2Ykn5gXvcXGRbUtWvTd5OaMtW2h7yhS9HudY
DypZ80PUCox3We7DRN2OptPmMVZD/xsxk0noU/E3UW3g2KTt5Rb5k/dX/cHr93KvM3dKnh5Pwyig
9gV2Yx+zlHpLfYXjno6ztfOu1U4V4CWJJAcR58iuhnjpgne1ay+i71l/mHBScCJwbonCgk8UNUZQ
Mo4j6fQ/58bzMH+skcmh+uHamBInH0P1FvgamRe6ysv8E3qK+8nnlhnxuMYDyxHriBrtdVpzGRP0
DKByTkAIyiTpyUeVwAqgAMqIlmbfZc9TUNq/0bsQkkyjw1PS5VZVk9Xjd/CP3DMvE/AanJ3oqsdJ
WVz0Z8i3eQ/hSyKKqHKXGWLBbRHSpjiXlaokEqle6ypmWM6QPHCCQFhP+sTCwopZMyH3hgd+BLOT
Xa/i+ilDAOUAKqcnCnnXuStgRAkndjzsEqx4ylk9IwXHv6VqclWCdWFwfQfqjsJDGVRjfqyiOR1q
fQV2ItnBNFwC6KrmbtKyxRSxVVoont5jcYZTNEYCpwyH6MSvgnFaya8HA26NHWFQnF97wb4Gy9r/
M9czfmaL3JnB5JRes07z3fiE/ywkmuLiJbwzsb2xKrv9gwgkQYRK6dtSEON0cxj8bMgHL/8xDz3M
VgS7n/YMxNNqmsnoULa+M4IQtKOt2o+nUJ19qIZgrjmurOrbFLQ8R79rTgVdjwHTAJcuJQodSK6t
We1cMY1EZZumknqdf+hZcIiH+/4okoVqMFZPtbsGkWK3kCT/hKKIeeKTzCfXKLxpkUCK0tvlN6mc
plI0lOwndumzy79h9VkOWpCh7Hgm1lx31/kAHD+m0sTK26XMgrcfB/54JgykDAe5bHv6lHSJZ3yX
uvrGGnLMLgxkj+7dmV+jK34kUOSAo1HJdcPBKBS6gYXZ5kL0ptYDFyTWcAjCFX3O9ZvHN6zEEhc7
9JOI8vQAgKCut5XYJLd0UDjVLCODO1s81SQ6EvIRWnOfTiZJQDh1VatLBiF2TDLcaK/HN/Q+ZEBG
ALYbuGgIVtW+sYd17ed+68g1jvIyLDmUQ+HVQCq8foeCwa4hjXtNOGY1S2hu9zgSlPVVZJk/NXLi
J6/iQaewS/uLjpeMgEZJc9XKIWO8xT0TeX27ODIw24RJha33wuhdZeJVVElQoG83VzyKUr6Itr25
9JeRszJCN+IzpCpRbj50IONuEIdoF4qb8agSlCSxbD9wtwC3h2bymbxegqs3RWxpQQ4kRyzJ6fmC
+kuZUd+2izn/3wjSBdkfsIf9nsDXoiyJojjVYk/c42yGIYkN9jXNA5drgUpshMPH24hBC0l1XNGJ
7qXxldDGC4FEkK9RJbJCXTkhIA3WsRqUQ/orjU3dgotwyfHynPIPFwAZrYO7yZf0EGpvHx6a2bZR
VA7AEJS3T7vRRWsbqu6/pwOch/onXzXQYnTsdigOxXmMWgle6si1Fi7vpbRTCXigVfEufswNeFkX
oYEFfnm8ehjiwBheTtebmllMY1Ko6FUl4VHj3ExrYsWSSNCZSU5aXdBkbfshDXo3yAtQLy84UfaX
3Q5ss24dP6mq2+2jijnNZYGEQjC8MWIDOjj9JPI4vq6eAm4I7vz4qMuJi5Boyab3qeJzFqHKIFDN
AAccuCe7N3B541s41fZQST19vggx0+fqpt3R/UctWIjedyaf6nvJBSvGYcHQH5dARIJkY7rXCPNR
yv9DaTujgjbWV4Z7SJlMDv4SoFzWGroWPY0caOWJp5vpMQmtUpcnLPGJTgmAHy2sUx4PI+V2nJhE
ySbURw9ekyNpAnB7Ie+qIw1CnFE5sn3yhXDSfeQi/RTI5ZtuVzOROG0md0MXvDS8sVGDphTJfFXV
mGnMXM5NYeboQXOviMNM7ZOAf+p8twOWK9ZfsnL+XCG35yQXkZYY8y9EeA9EbPhAv2TxN74Yvrih
LCcMc5cMR912wVyfDkRj9ei6Nctuwgo0Xh66s8rDp/RD0TIoJ+BMJ49IdLUjsBDGfnWb1Wz60ron
m4wg+cugywkdACcfjZOpv9Ba2oTkraG6VpwfpvhQH6hWmUzTxaDf1v7eOAbKYLQo/nCWCev5SpeS
g3p4yz7AXNxo7clxHmm+LzVfUyQD2eCmhjRZ+tB8KY1zofzb/sceOKqLUwmJDEQmKbRwCNjk6aRc
hOT2zvutgiH0nCfwCqduJ+E6Zxg5296nChRjkXxbsBdtxqHy2MVkZy3yQYp1f3/L3SmxDhflDmHZ
pZyeiZP4eLQ+ua6R4ApwwuiwC++aH8etT1/+tvbHSKj1zXVwFGVPBJcRUEptGvxxfKI+jR99wjQT
ABui7YjaRE7k5d1H5OgNkH0Pr1Z44YY2i5J+nW1rCslRPOOF60/buXsrUaEDBEsrGBmX63yEEZJC
+EjW6Mi3uqC+ji2XsLgTXmTyruAtbJSlcBTQJMDGYGq5rH22sAuNzHf/05uVzk60aB0OvXl8RRKs
JeD6j6kFYVO9Ny5R0T81cQ3N69gt8MQpaywbeiaFCYCtH9qz19kkkWcwfQkpGKdLw85pR5xhMXKP
aZEdm2hHgLCNSmg7tIDlxBgRRy0YDeT6Za99ccQ7IApXMV/k+POjk9w4oU6wWZih/zVDSvdajk72
nKHmAsn+CwYKgKCvHMicHmVfJAsLY9ltc4GVhUO4NKKWOeNCFk+iKoFY3g2R1u0wavwj72k7aLpC
2zwZh+K8GhkDuMmofLB0ziySKJ0KGjmjx9sLM7d+0DuYJFRvlpBLBDddG94E3EjMjuFw0OEg9wVS
C35bNTOardZNkwA4PkzqXgYaUwiCrmS9mrs3e0awCxkl56+dJ297EiVQnXSo9x3aESdb9P+LGsRR
mUcm5HXCvBGXGCdRdLEcuUpiPUks2lhyFq5Yc9hQgS8kCksLiorLaxKTRYGZPjosB0P0cW13HGIq
tnGIKK+qJ7q6Xg9MgGwFO7kj1rgkZ74Tn8p3JewSSTyRDWEViGMKUReltcI7jmrHeZ2fWw42Z9Tn
86r8m+vG6kuqAnV5/hSeuWhkoegbLdIwx+Kskl/KCmKue+0yXJLJ8fVDOoQ0umjdvWGbukEQ+39H
5xpeRsbafVOQAhfeAxHrprolFIcM/JbkfQA0O2EDqcoPQIJbBNyH5gokJmvqi9kFCV9PAzo1JcQO
6KSeP41bFwstPOFKv1PuoGmgeTQJ7Jwu6cITqldGIPQY4XZr7vwxRsUfbxzVKI0T5bNdAaZAa1Hm
teIdPZ+YGrp6G4fWseSt1Fy4TyeR7nA5hiU/eZyV4RjXJCO/UVk+IfPS025mz42m++SQBfakEpac
Ggn0mUabyDwtG4tAhRGIituN5stQbEOw2l3qCBLfQQsH21GqAQ4INFm9HHu3FC7kQRtkOwCmstas
E9s0LM7bhElc4Xf7HmRPs1F9Oa2/3HGh/PLQuJUlMHK997tr3zFHDf1gyU8/05rQzLcS1ZqiOTVB
WO9s9VQuhxoSJ0oJFxn4iyO8wKE/jR6p/bYS3lKIMqebkLg3LEQFpIVNXYnMOTB3D2uJqBAgD8TA
AfB5goLovFw6+4BhEcNybAhnIgU1ZZzZxoO8NqEdKXer7CXOITXZOpE3KkBziY34KEKgq3B4ADAd
HNkECxuLodNg0nrSq58/beYkNNlnGOGZgUri2hTqeoB+xXUmBN2V42cAlWBx+nrmujGkW9bvVNfO
wmB/01HfxTBzWrIyaFYk28WVXmIHYJIkg/Y6A+kNLXnqp8eeCfEmYxDVHgIqxVy8mzKbqVUhtZww
63yqZB2n+yBCSWjro4vJrPikvbHCXii6pUuaLsO6nPs1fP2wBFXaWUzhWmfHNl3W8no8CMrDxLvQ
+8ZZi6CaP4ORgXk/PLngyTX2/vemttRYFb9TRr3TLro2MwSSTHB4Lk31YGEVNjNLXxQ0f348j6MP
SrkdyvLj5D18hfVQS+CtarRd3OWtVaM1VjYLwG/QqDiDF+wBJ6cJO5ZiclcDkTKQ0NCF1Up1kdhs
/eStqmW3XDhvgWcn2qjCOVjzZfghS91gXwgZqsIFUx8kvgEJXNnux91AzNRs+AtV9YgDwqmZLKtM
oUBZ+4wTkZOKXznMLjPZBRZOYWM+VQR8oKmzMNjCFgk4r4OgzAd/8r23KkNnMeNSLaYnitLF9Mj/
hv/u1lVsFOv1yzba0FLcXunGXtTAHy5b+I6K0NTYujuwaBeicSDtgeh677TrPayDwR6BNyNbkFYD
rRhumVBP6o8Ki+HBfOIcv5De4mAXywA388P2YfQr/nAujkP9dBPoGsLtcBRDNBiKDTV3ArEvil3u
W/4GkVS7e08z5xzGxbyG0azsKB0X6+pcX+2BlWBKsR1KUFtO2UpxzIX/3JLXHBtNxg98XRQvHtGh
cOK9CcZWT2VOY9HjQUIDSsU/5FlTZrVEBNsLISUgFIwDUS9Sg9keD6KvtxiWz5kkxE+FVOmAKDSi
7uc8vasGM5VGxJDkWbXczCdW9giEgUm9DuLF+WhkdF1bjONmOaz2lFwWykUrUBH1lXbQ1+oI3SN0
dgZmqK97vOrFKsVp5DPDmP+viRlWdmDB7a6AS/HGjCurHw03KKyNslM0P/NzlSM0yIpQ5hORopMQ
ZirucsuWu0HsU56FTw5w5FVtfxXhQC9J+DC8kKq3KslTjTQ6tgPC2wsElx/JYgGOyp8gCkaMLga9
rkbckd9qXDt20lQmpKdzYuMZ8kOn2WPjuVFstoWGn2oISrqnTQbqf4rXCk3FtZS9Lpcz88O2s6vm
Dbr9R80l6U1X6EChHSjGKXoqVABq03H6oIhArnF5tOJdZHJIgC8lWLJbzVaz5kWbbBowrlDG19mu
TJSZFZ/BQT9D2wHpg3B5KtddZmbCEInNrFCJpeW0FUkY0rZ+Hk3YPD6Lf+K4XT/YL+N+qu2SqTgH
6xnlBTpRqUtBRJAJwNeHDPOLTPmnjayaFFLemuFaD6tz3wexyv1Nc/EmLVyu0uIBQTcnlld1fwKS
UOD2Og3sc0Ey37PmXkLqczmfdT9mlJeweoEFUJoWv4R44aSVbmm38y8WXKqpjTHzBlOIWhKYOEXC
BgDkLTyrdPcjz1CuH17FAh6MyYVpbZx4Hq+d52qUcSPXmG0HRnx4eJQds6dxcmxi1cTtnz6mM9hV
aRgduw+ewqgqT2ixehcU6fZn6PwTIZSmb55KcA4V9SiuQYgXnjuug11MEblSQbjOYOeA8naVakbM
icEE5HSl+RLtDwx8GnEqlalCkg2wUSVFPSlJUe08v4mMHDdUj4llPfTPaiN9+mi5vh0ZaHPwDzH5
dw1WQ9U7h0sNiDHY1ymGuGafUz276Y01kyU4PcKRs41PiHYW+w8PwCF/qSrFCZ6TB98BPp8KGGOj
UI8Bts2mBenIrTJRoinMhoObF4Pq8OcccrzdkugECxESI59r3hXhW3T2rjqTO1PvFG8/nNhhgMuM
yc5Wy85c0XdJKg8LMjhi6GxuHyhPrRDdigBIOPPvLAC5IqEr4CUnz6BM/rpYJoidoupGXJ0bskU1
ygP29MlGi7CsIp4AChdlIm0YN5WaIzh+vNV9JOIrbjgj6muqmbyt8ID7UdbFcKDhvfgRdQBDHhH0
r9YWg1dQuP7Yb7uuINeA4Og/qeFNrrOZFS4N9mfEygAxsVoJj5hZCds80AscEQ2Tw4apFrYR++dW
Jhxao1HLBAQ57OWWCKcbmyjGlA+b3/C49XcMjtUyX74erzXK+sHkoSm6/iDCg1Q8GMWUNKm7NAsI
rHeDk8hiY+SFgsZ5Fyb9L4ZtJYaIWuDALSWp8kbltS9zX4GxwEOtK4uEhz+pmPMdwQwPwPw+fENX
hzuheG4YWavdMUaE91FXjNp9NXIDE1im1VAd+v+z3xtOMDivoxKDze5toZjljcw/BqGZjYf+oatO
uX3xJmmaephTaj58FLZD6DDJOD4uHTl4R6stj2vjpseNrTdqnaIa2/exD0CkNvZhmReyvJFVilzA
RSY6f4AXygkPsMCvcQFV25TtxMW1Q1iM95r4eSdAM2ujJVvDfeTjhgvp8KAIeXLORTUHISItOKr+
LCPbyvGiRAxZDjPSQPN+A6A8ZBAmGE0OJ8Qpkac5UBSh1pQ3+MunkGAGowzQXof0d6WjuD47Cp4E
aN56ary9dW0piXR5BDmEbzsyv/dwubUNcP67P9nFAI0l/xBLYd4jx11pYOXI/m9l4gFVqW/GLy9y
N1+XIYCYYIRoEQKY6h4V5KQCCODjfAwki7yfGvz5w5ZHSI79ygmghBfGXWwOGjVh/Oz6LODf90TN
WxFF48zLZoY9pls19lLVwcgrNKfkf00VUhgZck3P7Ev95m8Ij9DW6RYoT3sTgol/avnZYppCNchl
9WcJ26KX4Kaeuti1Vh9BoYIRvf+rRrpCcWbvpE3ELZUdzAzYu0YIQ3XEggJshzSOmQH8LMqW+Evi
HWg3HxxBIu6WsJix33uXOnZJ6qC1ayi6ln94sh4LKn0+Xk4GnJckjMeaXgaSkLQZnB4WU645k7jl
ao5r/lGAF+jjZDNTCO0f+QGyZD6ODTCRxkMBwKjt2jQ8l8/Hcw+Zjd9sDT60v1eXhPtky0AcBwIR
5gbtxK+virxDa1Gukj/tOp+YRdvmV3XcZEnGh2iLkxqZAdowp0hRmqP7fTE59EXKAG7DWI0p+RDU
kF4WO5Cp/HDEIs5aSHh70VugmMQtV1QAXO7EPfltlGRKYvg+pjkJk8GN8223ljfcCEd1XlltvFUS
OPIFl0APM6vIpKUJPRSKrv0EXvv6AJXS1x+KHjpfWfKzjQ22b2jgdLP7Kqa6myRp7T8G2eKpvhLW
+xJcjdnqWYKpS+ef3iFEq9qsdJL7T7wqF5rGJkZWpdBmxbbx4hRoHi7T3GQ5WcID93fslwTT78Gi
N6x9PhMoVDBzuopP2dl33hBZIE3KvLSrNLhM4WW54mnegdNHWDZVoWpavjFVFQd8tbS5CwAcCj0Z
9BGc4GGGk393XD1d3kn2mPp7Lkm7vVChntuy+pbIlbzc4OMeB5EVVi6RJvUCrYKtaGetcbgPqs7G
Asxya9kAJdLFevc6YlazXWVpCBV2gvMNCg/EiTKWm/Au25MQRZYW5IX6NKaZM6a+obM3bNgA1nwI
90j1787cPj+QK05mt1HhNmwUMNHUaMl5u4vNz5QKJsxn/E5RqogRiBQB+fEPSxGWRQ2mprxVpZ1C
A7LXWwz74yjckSB7GUCrXhLOq5siydPflJUwO4wJ2nqm1W3AqW/9hQI8pAgITagWYceenEcHuJ7O
2YTpdbGcS1PivahlC/rgp4/HtLaDcK7UXEx3QnjH1NZZVGxhjv0mDgB77bv9+EEEVg8vv36uBpdR
leKUU4X6QMSpzeg/fFRLVHXAes2vEuoxChYt1QSjknGe+iEMwclb1DPWAWwziu+r+6DRdGRfLlbK
RJgxCAFpcidJlpZwPjIq898df+wu+dDL89nnJcnwyJsBDrrqW3JFGEuKoy/xhoU4/N+S/kUahhs6
ADH3oclpINPH6WDOQDCrLax7G3QlwqCn42xdYZF6loHFkx+MZymBM6UmBlzeXUGQkHNzhM4GWEG/
JS4rENl0Gxr3A6ZhlDFdzbwfGQXjDvCxb8dbyH2ScneTF0FUb0F27oxKUdxonJmJuKbK49B4LesO
5Go4tedG6C82EQbIA/9GyAhhbkvdu62fQX/1iRK6pOsKR7lLIGFqm/43CvFo7T8oCpIH+UB9gnln
C9ME1x1bgeGi518EtGYguNetmkxcfd1qAyCE6X7pFSmJHVZMKFrpvrPq/8xlYd5G/IbzgEbf0QiU
p+v0n2iXj6b+Tu7gIUV9RMUcL78mhq8mlcOHnny1ODzFg2yuWxTzqFLoYBUBtvQdnk/oTteY7eMY
yQqFSpNRwGz88XQnG29fknovZI9zQ128Jux7ngrtcUNAW7p8IUsG6iXFIiD1rG8tovgK4+UAFKeQ
uyRnd5oZ2nnxCBjfNJu4H/MpiXqueUAFNovnDwBCoNVLP1ZIk47lq8WC2eWCWbF3c4qqnuPaiYHz
zQ/rHyez41z/P1ntX/40BgisbemG2L4kMgzSJFx7yHFTe7MPABbnFEaTDHkztN2e6svuTpB6yoc8
0Kwccc2B1gmJudPKsNX8RyET5VSdmsYbSY0QO77hNIP9ALbnjccffI0cwbMVQFn26N+2HHLNbbXs
yjZpWUhNqLEj1nKZXG7C2dk6mG/NPqvLAjv6ixBlXIxieVWebZkOZ7eiiWNoAX2JK21jSY0LkzF/
l/6xfHrotjPNPZPsjxUu+KcsUeHXPWcA4THcreNSnFRrmZ488QTPZf+aYr4yXL1YRiPR3CfJ03xm
BYQ6MoSOxfLaE5Z6jcMb2AzIEy92Gqwaqa0wqwvBTY1ljrkj/WQX0NeQOZqjny3nnTZzeurBJHOH
wNfk7oGzPwieQDtvN1aj+XEYcarBi8BjA/xQSxlmFzjBY0iy7PGjibuZTFq4iGDlBT92lnG/hdEh
pr8jDoJzkpn98L++8qbwBSF1OJ7kKpzESvZtrnpfvjVMDBw6OPlEK6uwcFWXt1yk0h9WIlGpAaFl
h/+Hu08ATYR0hy0upCGvO0p0/iAQYk2yX03NdcJ/YE1QZmMZ2R9+7+HYzt+6sP8C0GgAzgjgdIc5
rkL4C0V8MmELc81O6UKfEm2/yt9qdrKlj3kJkKj86RcHsWCj8NcId3eoFyOB7/CG+U8yZtkT7vVM
/diIa9DwaPj6+gqpv/QDLu1owPtybqw2i8ZAnT64fJOR9/04lmcogBV1itmp8MR4uaOBkVu9rINo
LwsISmlc2RozfQppS6h771/qDBxLG+zGrq1s8u7DgTmpx2HjmlelvdaZn+Vn+ME2RyOb299yxDaV
r0r/8zStP2d0yOL1WkFtcUFSuBcN46azU5YckWVgq3CY3OTDGn7jvUOu4uUTnCq83PirNSZ+/0G/
mPVBOpmJ7hFklJFMhKsD3LYXi9h5xM7TstK4KrrjNSvVe+5EZVZxAJocn6AVgJeVD3teitLhctHR
8VbyEHdi6mMwPaOnRByIv33h04va7ILBAkF7wSL56KRo6yCMlz/y8BB1uGi8QzoclS4OuwgoCtQZ
hGsBb5yWkUtlCD40xdQsGSeYUctISrXyGOT9Mb8c+qIY61vKXpGHP6VRAFXlm97TEZYgj9RMpIen
PvRWGhZFiXs9Ae/BzlWbVbUSVws5M7wLE0TvrfD7um9otz62HlwJcXpLQf/MtYrchZAzaSwf9uAg
8b9VUYL+MX0Pw4sO2QGIJwgzVU6tBQGUpPV9uR0lnj304x+rVwUoFjBn8C0Ga2K3DWJIlTeCf0O3
woS1h7wtSiHULLXbeLE1BtguxC2CEr+Pe2HAd8wv7FG3hRbXLSIpPeadGxo+Hge1oMH6CsnKlwRS
XaZqlN9XPvZq+fmhoXxU5AasJl6j9PRpz/x+K1zLuoRE8/lPhxqtz5ycZ75AqN2BNItKasQMF6wg
OSqS1PbTk4NA9qy2twOscKbfAFf9dmiL+RA8eOxZrWozFlbUGTkUKhK/oEuUoBw9wbS1Q4wuYzjY
A9QtnOYJ3bUSJWjvq2zX7ezx9WHS8j7oL2izzl7sBMvEsQugXmr8vX5uV+0wuYDNwQ+Cl+kU8zPR
cCtkIMTE+c+xhd/gDNvRVYOOrfzqJb7BsiV+ZSdLDull88mJVxdPD3UkRQC+luzLscgpjF/Blm4G
VoX10mxGky95WSrlv8x9tzjNQMLRXj9LGRH28KH7UHRg5MgCPQzgWF6Glqa9MdxQ0RblC2NqyNG2
mNy4scTcBvMSr5Q1E7ewpqCKiCJmz751mzKuzsvRMuT/A6EBtig+Yjm3G7A0+lKFbSHIVNdaH17C
msLO7824Dh/QZAcKRibzCTXBpS88ABOROwaaf6CdXX/KIJTRX+9T0YDxZ9ebeQn/+U1c6Rf5vJgU
YDLrqXf+SrJTP8ewQa0qypjHbjMcX3CpW6Cus63zusNqQ7GzJDVdG4cpKnHXnTiGhpnQJ87wQnzg
PMkEVXpAWrBZHQoqciWAmd06mJIkh7+MZxN6rCbMLSBq1qTH/CpLVP+UlGEAUuh4/ATJYv7vB713
StUQ+JTGUQGosvIcWIvaJRhHq6kezDvquSnU5Pny1QMQ7xzaopLmQ8unOnu6pGwJCNO3Frn6v1fT
OlrwJIf2dZ9hR/U46QWGLyLjbrc63fq0LrzqGNTBGw+K0EwaI+K6zljiDvkFbIWgkq/2S4mk/i1G
HeQm7vTfuEwN4yNYrHnvalvTY23fMJqGuTubRWNN84l1G0aiZtT4B6cwSoGTKXnD9JwD5/8k36AH
AIoaHXBLEdSLRuXY2tVxSxWjicJweonySJaWL86gknyE9ZxZIe23zZheWYEZTyf5LmNO5ZeqhYDG
dDPLDv4p4wf3Tl7hQiEzNAUgAw7lbOzTGO7l3BO6s6jRLwAfN3cdm6lKx7Ka65+Ko3kQUvZVVwYD
BImE9x8t0ySWDVNApTFXSCU5zSS3fc3mX+hXqemkyBkFQAoBfpgDK6+JwzDC0RDL2Nps3nM5GdRH
tWQy3jlu6d/TT2fDh2CpD5r2PBmMkIzLeK8B8Hf7stlD5mY5zlffm841NeGRiDW3xBATo4m23wxB
8rQ/fbgzV2GAAnU6/Jo28EkZHvCVS4zGOluI6Y448JrxU3ZgivSp/iWmU46mZkeTE9QBalZX7EAh
KodRSuFpttofXFe2vX0X285E1KjneMvLAazBUGodPhdIv8+vGuYb
`pragma protect end_protected

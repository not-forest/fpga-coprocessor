`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MxwmZlGb6RXpjHifmdHBjNdJq4ICZu0CyfybqD5ZUZHZBn987TCiw6QooP9TfWHh
EaUS3d+Ta9MRVRuWf1hh41xYd6Dg72FeCDbwyRyHQ4rVWXY/4ANuo+rtPLi7iaeV
qJbV5GleP6tGAJTdqIvVRkkPSfxq+xfGX1tVJ+G4lLs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6272)
JzDTPqbklBVE9hzNImX4avZn0QkwkuA0AfHMhSBYjz4ddanKq9MD+7tn2vG6Z5t1
Y2KFuE9wHZsdMiv4hIt7FHN9Q9Q0S9zRZCUsQ9I0aDixL6XZTA4AzhRSjuUzqtgK
JzrkPrzfz5C0gGRaZRuJLwl7UGNklUiVyO23NJDwUirqryL5xWFeTnZ3wC9jZXcg
X3PRa3zyfeWLp7pCCwQOS2Li+P+mgueeHP/WT7ZVpjtVjyaDP/M8Jzii5aKiVIGL
rKvsdJwV9sgDvjf/i3SdktZzF23Qn/PffEVBHS6nrra/xxlvx0lijAiUIB74MR/Q
BNIKByxj8G6hKfFoNYILPiazZ89QZpDeCQhGjGw3U/3xWt4eWm6j4zkJpuJKFaYM
uHfQb4a2aD6nOiwbkHAeVcBCsYP1UCGlQBU+O7/CTBLzP0aKyba97rlT3Y0K68Yg
swp9GwjThA6XwAImjb4UH0/gRCDVX7KpV2Ps/Q7e6OWt2tD/UJzKkHpH1UUqz/CE
bVxC40biluYAc7K1DhjkJ4CWiJWupl6qa7E2Pq+FLDtyQ9kY+1QgdOutDXOOWIMM
EI6lqK1aQnsumEeQlFs7aTogt23g9YHbJy1aCX61P3jfU94A/HN+Jwrul0VyX4Zl
J2brTK/aXjgAvkIoH5yDjBZ11O/MvKGgvsSkQ89xva5cKkWqQa8/N/QZu13ZEeX/
5wmLbc0wTGjD90T5IkNIykKkCfbf9+bTfrHxWvGodK9JDHetVZXsNpQh0W29YAtS
koSo4QIc/vQE+rE1YmSWp6p5rRqMX53eSxBFx5EiqvEPyVMiDHGmb8eJcSZ5OT0a
Qlnvx81dX7BGWg9R4h/tX2zFhAeabuGR6JcvjLlnVIB57PugC21TLtYITiI6w0bI
9uc51UuzzboWoQCFWgHmfWNZPOdwOp/xirSnFUSEWmOcFD2vFghGD1VP0D7XZmQ6
4d5nZKwvv7v47xVgsrf78vEOUrAVpbiLr00wOc9DN48H0E6gUZRjPMyusZfh7qty
C0+ivWQkgaWo2Uq9WbN/XXmA+w/iKM7w9VndEjJJ/PGJcmoRfKtMg+rffUBvzOB1
WZKzv8RttO9MlyrNW6wAzSL+gYb19RXofq7Hz5kEE3XJAMM0Ss9XsfjqohYrzPjS
y+oKRiFKKnfXrh2HMSCwUJfh5Q35BSjjqvRcesL17MSZgs98taaZRY4MjMkF9lM2
3vp+6Imz6kU8XKj5rUqvsCSzZRZudCjMIa/bozSTfvouuwT7Mzb6WDLKpybde0Ta
3YxMAQcp8cVGvSNjWy3bS7r2CAEnAOyHetNOEKvURWsuN+/rrRi/Qyx9Lx3fLkyk
O1/+EY1/GCLuEEqc2Jp/A3XgSctZ1wCd2DpJkRbSSKwA193b6rt8EaCNqIHoKadH
QHTVPTcMtpb1yN/Gp+n9IOaU6hbo8DAhE/Qy690TbvLIdm5SiBevdrmnw7046Dra
TZ7qzeI5TYdhLc1tGLeidjmpX7pMqitVPvwhesPH7WOP7Ys1UhPTaXpmfdzwVZbE
1DR7fG1TsOdmrZmGZy7ThDjvlIisNuw0IdfjCLLngwkhD4ieulGj9IqT3iJrr4LQ
gfHjaKueIP39GvwiuOzc1mKH2XZry8NKnJsWWSUghfc0miImkjdxomfuqx8zUYxm
dfSLKlV/KCOYspHYFxBQ7FDz8GdIWQz2XcoeU+hXbf2bZ6iyZt6CquUGpP1D4l5f
8t2r9zOY9+VSvL/FyfiGBn8k4R1uEFqJ6eXDMktFlTdagBUuqplJ1rhXgEUccHhw
55DM2UtIwwbLdiEYK5zCtI2ixx40nx3AfgIGmR6e2G95uj397NEeb7p7AYdwcg76
qM8n+wbYMLhuorYXsupNJ2QHVlQMEy7nB767nqK9yUYn5ChXFgKN/5vGXENQvoZU
isjYa/WjXdzrn2r/7lzejS2heUhkqjXA2VcYQyFAaTD1wkfkdLHHJ0F5LSAIffV0
jzUTaF2q/3FqwExaerQq6XvujI1FFrALVgjblYAW6dbVr0RHzmAdnTcbSpHSKRQC
FoiPnekWCXstvFsuUF1QbYlnlBhUnEI0WS1Ym2DaaQFlU8sbBOFbaMjDaVFVwcxb
PaQbbjg9u21Oy5ZyfehN4sljSpwoj8xfMWHkU6TOlwB3g4v6z4l+Rd21LXKbW6aH
0Zl3CyC1f8wyfb3RtRyHYHyuKd6HIMGuaCZ4od9I86VBLGqmTx8YSuKQs2UqnEey
sj1OG5ukiIW70lOVXYqqAl3AQtXvdyr9zsqL0eBDlhIL5Qieg+2cgcGIMXRHiyrN
B2K79tZt3RiH4NHPvwhe7q4TzBB3kTtHnXtwkLGFnAOA9f1LUPGeXmTiabuA6II7
JT0nLACk+VfgjQzpo3Feoa9sFdyaelWdaZvhsPaVkwqo3bmRSDPiSLMVpaoxM5n3
d6XOk7AQK7wkA6iIFNwIRilqTGRtWsa4MC/Uz6AnHmDHwyScoJmzVqbzQIIYFN4g
+hwTxjU/J//OdMJ/XK2ZiLWG8dn4lxnyz1hBYRKVO7RCVIFlAuGFnSTHf1kbsD+E
5193Qr7LXV/5h0gCcYH2df2PPVM1sQUUSrblBDIt41UneR3nY6gafs0dkfCBRe9G
grdlcOsybOL8AIt3948auRrwBITUsFDNmDDnA9e6lYH5SfpUXBqKITR4UWATodqH
jpmWwID0VOqiCCaG4OQHXFBZ8CfBaiwWveu2p/vRkGn8mEnn9lLptcVZbjRMJOMY
dXhOXB2p2mPsa/ICq0D+ypBKWha7rGQ/mnbtUkVeqDQ4TtIkUipkbbym20p74e54
DMFE29I5A9D/o8FZmPe1a0v2hpuIbXkxWG21VjpSRI1UCxl6kDovCbjZaxBqsCyR
gTXiBimEuHpZ1fqsdkzlOd1Eay381oYSBj3ZT2+BWNqhgYdut+b6PsGz5qTq+tBg
iExHLaSYQkPPgD0wqa4CXiY1T4q9F+7ON/nNOYAk7Y0s21gdorneFt6fFAC+coxG
LujMpxrEirfRXRCoyTa7bmI8XawL55pxz1ly0MuFXSJGXjbt3sh3htnUklFXcaEn
qh+RxCpWHxHIr96M6wCa/FYvqGUc0JUVSew21V+58Bf5K8CISLWzxHFOZ1soilWX
nEDf9dO9a2Oi+oPVDx2UCVqBSCj1NEVvXPu1MekyVVmFmARVKTR4ZzHKCJzfX1u3
x5T6MEhutA3BVR2pGLzff7tO6B2zKWtoZ+ywzCo0OA37jTW0p/gY4aHti91DZxnx
jGyHpRsI2/9PC2tpV+C7f18k5S8FxT7pAPrcC8sTSg7FJyRmnsAnTwEqeb5jckZ0
0rb/V7raS2ufoH5oWBA8hs1uywOVYJG6Jjl3/qWf2UTjBeGEbXMfyc70reKnCkE4
ejBfK4TwyzgVz5hDetwT7up8GAqF2P0aMQgcP6nBxbnAt+2j8sbkCmLw944xZDqq
9C7YHTVIDcCf78ByyiQLlU+1EIAhplvpNMKc1GEFRXqYvepeOgzMBXISx+UCEa5C
lRPQCgzhzq38ryfUaZpjYZ0C0PkiZSbiu2xEJHbz4KKXp0v/sT5v5tsY01cburWZ
ccSHqQzuDUhmKwuAbypDu3VG2MHvgQQYOue1Bd4AEKbwJJ5/87uGlkC8fbyYIP9M
dH5GoAYIkkGsWTUQ2m3UQlS9ons7bFsOiQqCRBRSH3H7d8TGRnR0j+A+RvpqWb39
D2Zoer5ssNweoy4T5xi4SZgiTMB8RLK1VepSM3gxUQAkBpREPjP9629ICEEFSrV2
4c5SFj9NCthgVnZAWlJmvh2pQeY5o/NzxpgK4meqJEi8Dw+Nd3o/ZBCKp+mJXkkj
CiFipHJoYCg0r+X1mTnaCUvlJpu4wKHcwt0yPhYB7npPSUh03xIJDYPvuQjf8PAN
svM+f5TDO8ma4T++1zv14wurLoas2PCE3SwQD5ZKYHN1T+6XB7yEwOWqtkINoRLS
NMoXVVnwphkXH/VNml94AC2saJY/QCBfQCB/X4Hjp3DF5H1Urc2KhoruDW1jTdHh
Lf57tnsWWrjBNrGBAxItFUKWPh81DtLuxgnWU0XA8qKNCslwnbGoqNwxeqqjW8I4
vJvpQ5aVkrvOJF/o/fLul4V5wSu3fOldB9B46P570tnOACOSQ3lX4oOgJY3MIdxo
xHZKZVvU0R0TY4RauRHF7X//T9BIJM8ZjIb6w9bHFGKyFuiG8j/w5F7ljU5WdcHe
ZnxxeIuLXRrsHlgSlVyoAxdmFjVNP1SUvFhNQ7qXlOxHqlEaWsXfJG3DWdxjZRhG
Z8fNSlIRlu6nrFVExpUEmAHQ/Fxo//kiqIKB1apKtWxCrZWBRsJY4ivch/claDfu
xEmSqos/oxrnZCl9HSjEgiF336EAK/RNYyjZzc2ae9viEjnrCFqrTNBBHy7tiUfy
bzSuSBKbrxDddPxcYRq0U8kiIDovQH+4Gbt/KqnS84moGQwbxbF6qPXry09KjIcw
ZbqlUWFzuIv+/kKcOOIxXJItop+4aydBRP+8eAphMxA4F/+NoDIgBNILMTj8PKTk
pXffUens+l6S+vql/swe9BvTp39fxfjq0/lR0g86D9ueD5qYz++AWc6QTH+fVvRb
2HLZOEEhi6g/dNkcaNkacr4aVOnSmbzwpZYGLI1BTD+LRbcQff0kDTxJPw1JYB8l
lMN18Sog37N+a1AQVPyo94XN5rIWT9387AKGw/VGIiip8qua0eylIxWiZwwOIVEe
VnztbGH1Vm02D/XTJuw9yN3vOYJI2ZNFXJEdVaaUDW/55xmK04KruR4Tnty42m8I
0AxZW2yH3/eSxoK/kwNxpTZUY4CMHrlXS0xsQwDKQT2OZMLCqw8W5K5DCqxTHC6z
nMO445DuwyoW9g2iJgR21r2UPl/V+wHeefylnRhgMQZLOOp5Fb48ILG/M9YDjVVc
9qB2m2HYT4RW7xivC8NTSyizQbwkOQcGt4tu/zLgyaTpqeIUP5V40PrEwdp4JpHz
8+tjxXU2pvXP7zayBfMgLMFpABUxkkcv4RHVP84kyYmm5GLH39ne+bakxFHCZmtM
VquSuySgR/yTbxrvSuZDez7p1Ww6ysqUSCdJRLobRoWc7Osa6csL/xjcIIYvA7vM
NS48BJiWUF0ikrCAElDvSI43ivlSJdifHtx98Gz5xI+DIm0VSznybIngLO3e66EO
NAw/SdWO5Ep3QKLAtfyt0LjgqK76zQI6/S45PcBx4IMTzTsU71qRwjhVmsvPQzjs
1u1i3I/pU/S3QXEua5TK1iqPdhYBzMwr2w0+Zocou0jZaKutUyRL2SO6suAok7Os
qUmvEAawqqWKLVIkt8enLQsaroEf4ZDy96GOjKtSxDcl3B3U5ck2l1cRl6bUgcDf
LaGWNWNrCunsGlFUuCDCqJexjWOKLSwnu+Zb5C/W+tywtCza8P6IOPTbtriAM5qS
Lgr60pEOCb4EiepY8IOPo8gEFqm3tLbgZCu5rCdCbevrfCm7/WJZsMakojHRaNdU
Jgu6bvftPGj4dZrsHjjjwBPuOCo/OpH5YKp6uQoSS4oCTuCUErLck34v/Gsvu7zo
GMAw7eMgsp+AX5gTBlsLc8thyRPpTj2Y1ZbL4V7R0sFAaNP8h5d+fK6O+qs5sRvW
P6UMmxt2sedOJZf+HlGBglT4Acqfw+7q/os0DfWGS+V/Omt2oGzmeZBIi2fCZ9AS
5DDZ6kOgL3XTX5nkODG/+Z6DsDDRqYcnrzPh5KalgM74OJeJFCZBEwfNxC8IHnpR
zICtyjh3kR5iLgqF0x0qmFZ6E2/GqbneTsymYRuzmaTIkVhbJ6N8mYgWyQPXAFRB
1/Db3jLHlzn9P1EgPrQGJ4vCGLkU8nGA4Oi7JCuAtphhAUF/jvS8ksxeTjrkYtHb
pfoYA51rIbQGuLXIoxSBiGEF4+s8aJtfG/nnAJcQ4RUvldQpLMXuQi+mcA6U871L
dgdyInaBxv70gDZ4sUXSMrK1Ue0o3LOhnRNZ+YjmLhBbkilkFqZjWJMAAtfnaOaP
zSQfi8KUsWD4/LNG9mhoKiPku5Q6KEkCYKtk619/pnlFwzBZkxHgwQaQ4y8uSjk1
dmmSyJibKQdLmRTvsl6GGGOp9dX6TsrBSgoxgttybdt5RORHg1g1afLrloQ7oqRe
MU6LsI6TU/40R82oOf8up5CltTlfqY7iYaRIaQq3RzpANx1cTtiq4HlYYTgguHbG
vw5udmgVF0tiRe4OrkORUoG18Ced8gizzapiHsTIeo6hAf8WGKay/yOokPWVnA/o
Qg7W4shBXa1yQgPnmyD9Hl8XqtXfO/TZqlUyPflpKTFoWH6WirQp77Ua5pls44i6
gkLk4P7fb/8vK7eZSHEPwSxKXpWbeVhNAfj7hS/bCS5eXg1XUKvtBBpynNK8zyAx
rliEo6fmxGW70yI2Kfvrf95GYJY+OETtgdF4iwnDYphIYGhYGyhCxT9h2DqAF4aX
NFIcmvBCsSQEGtSm8XMwpKYNyFu3tA6jYYReAwkNdfVFjJERM0NwzAWKSqD0tFdi
h2f6zNjZZfEzZpagBWvfinl5NbOUjoGiHPVdxV1+gCVyZ15AsNYcGFmMp4Zf9WC5
X97fsEy32yZBJYInuL63vSdpq0nq+t/gRwJve85/HN30qHNQof+l2AviAvF/z5JF
5LibJt+bPKYRvGTKAx1MLTkvuspMAcQe9e8JQ3NCFDW6+Y8hAglRRFryTgx5Bx8h
neFRP7U1ARV6Zr4NFaDbl1sJKWwxjH6mSL5Pb4l3Hrd5At1lunvUiRjKjTlQYTne
n9suUZ9ovCa76NvVR9GuKRLwub3w1xZqfM/2W90nwj01MH+5EEx7dbkcCK9qCvbr
Gldd8qpCWo4lnofywUzsnMWv6gAZJpkIoCWqFo53/vW9pVYubaGdmV1MktWSgCXr
6qHJDt3ibl9Evs7P16AMvMmWnApvRI0Ne2Zv+Sz9jX3hwSirtRNeF2j/MXA3lsF7
pcO0U14ZIxbfnKdgw31nrfuyy5/ZZV6BOWANYLWjK+izk5dYqd1G8pApnqo5amRi
nSkORdJhpKroXi8lSV3gRA9RJGEqSh4l/SzAl4oFTjDiGGfJjykZEa3MY45QWY3g
KyOml+rCQVJDJ+mSe+pgcPYhPq0Soi3W+R/IEfPT9zQ9ey27cDV44xRWuYYSUZmj
XKq0omaOYusLKrR/o06mExTnBn2ZfVkC/CsMXUakDHMvA/oq5i8K38YRj4PTneKp
9LbdreqCt4Z3WUuYoiTvkg2+Qu6WVYeOZXINJ6xBr8yMXmKChoFr0CWgbcRTEfSm
1vVV9QU2XPl7hn7Xhv7/XYELTy2q0JNmy7xW7tEc66K3OACsccsmp18qfyX3MzDC
M8kUyYgI8z/XmFNQ78fQ3E8NAh15F185bk3Ctkyt+0JVMQmuHPw4Ti1EpexMIrsD
83ABMbh01fblLq2O2ncLTEGhg5Q8Xp5U5bhjasAZZT7+dEQXjPIkrQ9xtZBwD4J0
g1k6VYokoISWasfcxiOeP0rsk1Ro5P2nfGjH9F2QgzTuAkMklWmay+M8PDuzZ6EI
KnF+ceWd7ECCLCazM+I4FC9LGRIdQs/NAWybMTFY/kbYKvsAoHC9gDY07f2Q2NcV
6t2E0mHcnfknIxmg0u9yM1pyalEVSjJViZYstlDDujCmevpjoZGH5hlG61wEilp3
JugDjF2LNCzph6aQqvLOMs1dbuGc3OjEPigQtgt3WYkuqTYAXp5kGQQF7HKOt0xF
ZWlZTGnFwDLvmxtqkOA9p4qmAbwKGfqiLkoXtnPLTRNk7VfH1vfamMSdUOHAj6px
NZxg5lLOZYz6+pxaLjd+hE5ykE1aZeJqwTz/4vvcDJq72Imvxe9kCinhxkNl/HYE
N30eeOYmii81hXhyFbQVXMhZWU22AGWoFajkpvI0s0o5ttZBwMbCEQUc0gfGPMRp
12KQI9Yu/MkRxWhkS5hP+XhBdz0EDIluMtle1A00AVQVfHP0mT1pmUB9/Ca01Lkh
L2cdb8c4VWZoE1qOSobo8NRAAm4f5RYoKLCDqwP2RKkM5aUO79oDrrhYXDNGgdyw
3a5Gz9JdIcVMFLIig+pSL1BYdAbpqEvwWd/7Qyj+Q7S6xrZ++t9hQjnrf1FhBHdC
gM60Wlxt9MIXrAZePNP1Pp/BQQy7rsikjsj0N+iwSNBHTS/b9C4buMeb19hI3Szv
nBqqDzexER6m7XhE7PlhmRce1D0X/krJZS9sI/eDln5evTyZLc15FQjffSKeumnt
kGrMWryvdshkLE1f5GUfqSkkq/Wf2bwExK9NeaZeCYSTlCl1jCfS9QGRw9D8nehY
07lub1AM0/dgYZelbG4rnVIqHGaK2Yjp4zpK3NwrOAA=
`pragma protect end_protected

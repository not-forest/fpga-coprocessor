// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
fOGiTHQFflz2jzys/GLT5mHoH5FMVeSwhSD7fID4DO63KuLphqBKqWW1EumQIOMQ
YqgigbUeS3q2vBKnNw9OVGWdeNaxrkbBG1zpza1x0yp3oQYSd3jo/0ao+tjy03Yh
3fEivIjDHTut5BWeiYUXv1NFaTJ7h8h7zCuRlIpgd1cG5V2QSCRMXpDCF9DBzgt5
CEyHlhYqf7vxJOHh7QFoJq/D9Ia2upaBl2nd2Hny7uReF7gREknybuNv57AWQ3Kf
yxFQcjILQ/z08SVKZf5uBZoBjapqiWGvZ5DQRXHv8aHNcffkVUryo1tLk3wQCshs
PnprnoWqD1tjBE7kM3ungA==
//pragma protect end_key_block
//pragma protect digest_block
af7tCoTlqqo+eVopi9rWV8OIaj4=
//pragma protect end_digest_block
//pragma protect data_block
vKkajE/IfMQrjCmHJMoFwMphkkKDEHb85QKSSjReuuHiG+ce48d9E4aNe6orTO/D
f4ZaCSxkefR2kEo/TVZgFC+cM9Aq+4qb27KaMHL5qw5hug54qpRdlYnWM8zrGbu8
q9hHFO+V34ibMP2Swl12HJPXYR3MVWy9Rnntp2SkPRKkbkP0kBFcjjQVl+or1xVW
8njO55bVB7QPk/lrJfCIhSZW/UOkNrUczpPcoYdDdmFZ90OiKns3H1tMZbGc2SNt
ITsnZ9IvgLynr1pQT5P20AKtoB8i1w9TpLz8md4miVgd3a4oj1tjcbiZDdcrNXu4
RLq48iKtMQaay48BL4C3BevDKl5D8qyhi2fua3SgnS2lsZoUpHkxXy9FDY/2+O3x
D9Sy1Flh29o2DJ4N+F/cbuDvHU/siOh4SNKCH8KadeOF8guiZMpN4GBs0l1+LwYu
P3AJdE6NICfBSIHhh2Ithtu7svlY0ZPsyMA/bRhQsLwBc6q4fGUHa/bMwImDW9hR
TITqavINI7taneyaV6oJef47f25DGdB7ErFP0xpSD0BdLWzGSLm4gBoMNJTa7vhZ
tW1JdhSPAGbb/Nf3vCbkecjdhs0X2tZ9zVEQhSYv1hNu/jDxmfh51Y4n+vgvhT/y
AXZWXIsxxOb01lAtn39FXdaNENonIFuUUjlCOGExRi4okdX4sEAgeGu5wquyXAPb
VY6yPzR+aYnbu82tlVbgt2rbWt5lLUngX2XrVjTHVtnJE38uguX3GODizKKmJrWZ
cL0aro/dZEnmTn2W383oD4qFIC7i8YqPC4AL3v/Fs00xf6uUxkO0afis3V/TpTUc
aqbkjWvw0D9Jd3ws07OXJ5OvBeS5yEBiGBJf+0a9yYrJNceJB9d9fiXgaOGuDICO
sprjx+FjJGddtqw428UDIi+KdFV11IbY1s+vwhVcYDVFBxnAz0EMrW7xs7PuP6dF
1+/oxx4r6+GajOGvAKv/MTEAN1CnvhyOCUa0Jcx56MNMIWSnCr35jXAky8iaZg1e
oBDM028o0V1fn91aNesitxje2IuG4AcSAPA/hTyGR72nBx1p4su8Efn/6ALCFVP1
XHjteB0q3FQqHUkLSxGsZV0TctLp3Lao580nQM/YyD/KzXksWCNyQ0LbiClX+Fut
4RkLgMAe7YaPCJzA5aQ6u50CYNdzfavFMJu0h5ERi9Xd19wAGdCZQzJLboNz3GZh
WTKlweQL+F3eLqXATDpROWc7wjpWdziz+LRdFwD/ISk7JdbHHaMGjEaW7mlDdLpc
0FXHGRbS19FMWMJpCsSPx5aNo2JFu17WZ4MCSLxFkOThi/em88nONAeyOUMq5u4v
hosQoAZf5k2grP8mjnVfcYDMFbNp7JRtUfJtgh150A0aM3bgtdxfHo3Efc+HlQiJ
hnNYbvW9W+e3aWMJboIF8qPZ7rWi3s6J0CJIKhRWUeffqvzP1Eh+pP50tWqd0Of4
rJDAeimtZVtqRrRJjnVVLQExtWmTYSs+DAl6jKV7UKOVF6pR5uyXuJh18l6iEG1g
cf9V7/8ZDPKOooT2KM0uzMuhYrNEJ0HtlkaiVS1ixt5vwkvltkac8s05asyyicW4
4h6eiRBCnQHVuAi5a9d0jwSjKKMvr7g2VwtokUaUZhla3JWg0SLqu7qv3i4zAhJd
kert1Lw61bCdd1qK+jTBxbdb2SIVFE/eP40CAXHve3LY4ywHCPjEIznz6bAuQLHi
gt8GikPrSunpsL8w+tGJqm6BXOzHYu7us8RrXC6D5/N/yOAOrH43D0KTRH33dHox
DRnTeM/wRQP6otzidYBMTpLzzzDhmK7o926NZqANvCd4jG6xKpIra1X14YguexDl
UyKn1rk8jkvvXQcbqruf3nwGeJNOjoOIMob2Ey6mu1G4tLAqoibuTBSDEPxY3JQn
GNnPG+JQdFeBrmm9eKRvfyyQr/dAIQ+g/zJQcJ1+xGAx6VKLsIBDR6ITnryyUrTz
iT5mIDd7m4G0do7hKO7JIzA33aIIqw7zAKU85UNHqE6GbWg8lrj6Pj1i6MEWu1Nj
tpfCdlFRJwFp93B2sTv/RhZIbk8Ubeg5CmBdRdNThqyYgc/HjkC3oWWVQSkSWyil
bvAp+OBO4JIrz8WEk8OMxt3dDAPhitFKLk0bmri5XVHu9hYXrtq15xXhmK8gdAi3
w1qxC7W2Bz5TKVKYhkf/sAROZg5GOk18yHxsMmAw9p6Dt7JUKh8OPBVl60cF/4QF
pcDtiFZDEWFBnaTa7XieVjkcQd1UVFm55hqlds9rXvcrrE+nNDOVfAkQqUv8pDVb
vma56kevWv2Kw3gnv9mlUgseo7E5RAB/x1femB+00fyjVS4Pt4HlccU4lzjQoRk4
PRx5K/4OS6XtRa27aXgJFTYwcUGYHHVRy2HgXP8306eyYklVVTSpa/oqRelB7enM
VY/LzowNWD4Fqfp011xwy+PKA1Lvl0+joGx7DaYDdfRp5K8PzBYRMi5WbazF9iow
/ZvRcs4cFLCqbQW9D3FY7cmwO0Wuj/6moca/Tnsz7+88PZF4Y86YC0h+Yq+7gbvr
gUrVURW0hpsn1xkdo+/gb72+7lGynmBqRyCaTO9kemJPCBhBiqI2gNJ/+Y2IKTI1
AYoZe9tQp40hxhK9xfc3DBZvIwdrRnc/3eAULsFrXkDiVNR5I0Zsp+r6oLJL+pFi
H67ZWj7ADIXRQKjp7ePS3PI6UUPvROqxbTAfpN8DUd/XjsAWjGXotD4ere9oyA4O
J/oqOFu0h/uyAN2sxi7MoDnRaByvOKx/4Nv5oDoUiQ1OyT+zFLYCiXukoEELXIYP
M2nnMkS+Fs+CaEu7EQv1yqRkuhQRmijimYA2TXCiJasT26vq7j6o6YJwdRoc6aTv
g3R32tuuQJ8BVn455jRB8T9eBUdMLuThndU80j6eJLUav82ZfW1SjVoSpvfw1YkD
DiFYMnrbtDYQup962FGe7v7qzp4Yj1FoPo+jDNFLU3+XAnzaQkb5Kw2uMidim8Lr
AtmT6qE9mEgtG+IPfjmhpHb6G12KkdATPNb2en2QsvDut27iqmgJkeJU1fnZQ2NL
2G/88AZ1K06PzhJPP645UzAxpy8S1OrMh40XV8JmzKKoR6ehknwTm1pz+otgDD8M
K5XC2KPXthP6ietOtw7h4LY7irWKcoJa2N4JUvrKkXS9W/tBLRG88kRTnvEwn9t6
WiTK2RQBr8fbg7zF8G4W2WnoKkQRpNs61nt+pcr4zCx5etNIjp0BKY9hvlaYBxDd
XACtbFRiWXxrLtibVRUxU7IZ7ufUxjkgGjlCa7nMpibEjk1R7cN2Z0WbeqhNqRbk
bNfztziI+ls0R6owGP6+WnLFHddJjGyfbOtRLEFViex1KBYY9HcvJI2unb/U+ORr
ZpueGeAeDFj9bBazBi2ppNytTEurf0/tjV3hXYq5fjN6bKpZ/AbkCjv75MSoBbWh
Zafuxa2VVY0Ibh4OqYGvkxO1J5pugB6o3FaBh18sajjrV+kIBuS2B780z5bxMdK3
KC9QfBxITTvmFPRU5mFA+FWJZNUPXB98jIPWnrrjw64qFE3N+OI5ocPtRvSGtUNq
57UTZhu9dszpXno0HYPsh38gMQxIihTw5ZlPJ54AIkzqj4YWWPeE8VpBCb5EZhjB
bI7gv4/O5gmOBOB0sclH6dRwev1PpZMPQfbOoswG91goqlyECH912heP7jqkqyiw
BNZDtmfZ0Sl+z5j2amw9QFanCGcRECk059WpMwsh1JWTDMolLhCzuXH4N+k+qYw7
lQzwtVMTA6+dNlNNE1AHpcK9FBNAS5Al5NkG8lku9bDDuGWWuOaBGXOhvKZzISXI
snmMcUcXrlw8Q+w4zqX8ZVdCUkmhwigaZfSpwAelqSmW+blk1MJZ5cBUVXeGL6DA
+7Z8dLF3piXNmn6Lt4KxHWv5ev1aGVHIiQJF3u9h6zoZ4Ddh61wRnilrTIUkeSNv
Nc3r2s9hvNBWgEQUBl8g8JgyIwxOm/78RKzBAIlpbvuGpIO20m2t5ukHe2t+szN8
Ogn8T7CpX3i4CJyLBRj/waJj8llRQI92M7r7A2LdmZZmdbwf+0y14WNnfA0O5u6y
FbWlt2AXDEvHLO45hmMRo0w/n9gdJ/IYn9l6fCSkOPDgsifC7VIXQ7qtu3u9v6vl
Cde0eeW/87zSU+/Oiapq0s1n3bkj9iALE6v2DdfOcV7juDmmPmMhckNKVccJKXYp
H+2x2ZBLv+2AOgQg2DLWfJZ0eqGXHcW7uXLrhcEzfibiA6XWWW2oZ/upoh74IBZY
PLeF64Mbg5sVvJJ4IQOKyJiAWDjMH6pmx/IeRQfnYKzI54uxa7nMDXEFbvYXRCGY
wWOHntwvx2naRmQuuQ+kohbmmDwp5fcHsIYdUGOXhdP9KoPLyoKbKnlIZOcjVvmc
txNFLRomMiImd/98xdWbjstnNmfmPffPa5cRHLIquDGzHTMYeA3vsuZJ377GYWzm
MKfuxkiUnHY7BqDk5qHc/p8Vwutg0XN+IKis5uVs7zXMo1F9c8VOQrQivY7M69h9
NP9tOKDYJV9fQ5Y++6ttSxX1cgwGTDX1hJ7yIk+6uIpeLAa8usKdozMgEYvdEMg7
eJInsHnK5ergpFXCNLtKMnD5MxJApKkIXJnwhMYP16BH23ebz0i/ouIHL64MtqVk
lrCEDrXCXZoF6soP/dLmHCy8uc2GfqFMV9zLa3tC75UpzdhhDszS9RA2M4oI5+8y
ZNnzbQXMuT83qwYIcYcbxRYWHNUORfc1Xb9V9DSRQQFfTX+qrKAjeZSZNXh9pUob
musnNbbBo7rMhUmL1KxAShIrscAiyd4wU9x/4IJrukGRmNItg69h5vugSDY09lZ3
MeS8UJtHmcHg+0kNKmOG01skAsLCieNlDdmLktWbQd6rLSpybftbr09U4H9LqPEg
pQjFUA7CmO/q7gS5OKRCFqqqyMVKR4ystaU/S6WxXRptTKblvMRhAYuQBU7SHD6F
ezGObirsASd+V0iH9QXLq2FbcsDA0GTDt4IY+VxaLVoLB5CPNsxdvsIetAB5Smsc
5Za1EAkMbNOV7dwBDTlv6JyrrTMVTbJEDeoTFT9KHUDSiZNd+9WixQwkSiBt9Z8z
zIapvsPYcEthXu7TzAkQBnzopLY4vLFxXMagaHTP9LA9veOSTn49+L7yRQWvtDHD
rkSIakx95KmdB7W2ivfqFt2Y4TvzSD1CDYmpVL0x7+QOfMZawAKGaT5G/3MV/ESX
M/fzfsYmB8/0DeQsKWuVghS1+AYp+VVwbM0jLoJUqreECs2tRMRg9oM8gWY0G6I9
sW1TkzCF3vFkM/TnA+RQOJ7GHI1akzix2vmGZ9VG7CX05AQnr1zbMNmzk3AhVTGb
6wyjOrlzv2DHh7GWYl+SWu8i0vEGycAKBkXcYpC0nJza8Q4bCWjRRniL3aiApafZ
KMT9bLaY99h7xrSn5+b7bNtaAU0jwHIkzsswpnEjlEiQL34FNn9XUXSG/Aizg9Hd
ifQNq9reeXTgZdkJdH2GcpiWXiMsyeLLi12N2+ylePcRKT46iIW2sfrGogHwpCa7
jWDTdERFHMaa++1NXmvqBJ2HqVzG4xWw4xe0T5CKCptaru7+QPCzlLy7NM95do0/
zz+r7x6n6+QxJHN5hWKwbtAYprEm7MC6+keeFQgqumUOR15ungNkf7bP2hJEo/sg
Q78nRSAsKIyrT88zydl1iD37m8XaUxdq3Vpa2zhAKkAnPO5qqS1gSmwUOLIm4ZTW
C5ZuCDEoe9DVC676om6mJR4URxQIud/UJicfMxfIshqUqQ45EZTCzmKRaW6S3Q49
YeI5fIcGNex/wJTXBmejXtaR6lEimdFnED40kcyta1nDpcUe0MDFnDJAll9131Kk
HmpPHvQyasGJkm6rJ3SLY5teQtM8e+lVLTeUZKy6XYxvWUe003rxL3HY1pTkiTNo
zGo4hFkL4Ru/pw3pxf7aG25JidkY65CKIHrRNs9InNWpSiO8S19FDc5OwsISwrlT
FHep7r7JgxVCUWk/2qvJ8W6RV4lrXNbtaQrUnIxbb3SUHrKl98cHgoAQBrJXWpo+
9fHjTSgvavLxOCvb1kZEvDX6/BkeqeZPQ/2hwe9Wz8qMQl31RB2+tzEBaUYg/XFY
qGPrrLt54M9H7CiITVAeYAGAy8BezK7qzFalxO4S3uh78gttZer773K18yOlhS4z
kOhrrw2Xq2n/hRS9NsJVclJw3YbxP6F6tnoWVPNJRXW2MpXqpBHGdu1+/D0Fq3C5
tXKnhxmyjogf2MZNjhOdqZ2KdzOYkTYh3pT1BdhFvjx73l+/m2RtUIfvjnOMwCoZ
M9so192kOJKQGhOxXKNAbgslrvQ8965nxlzdIKJ8I1IZ1hAHrwfgjanP7WSUgXiU
2S79EDa8NTVE1/sIFhBExP5EjQMtODzFCw2gJ0WJJifv2U99XHdSuaH0j1MBksuP
5/kw234d07HuWkhiNrr/PqCgnsCt0MWilDnbmNrrSMWeDYzRPbA+DMp5Q6u2oi+5
/XVdoc48U4UJJfX3gc6xAGbxmTDTudu57gX/D0EIWZ1CpH7plgy/fw3GcdvvuMUE
dorF+6FYwmO8yezVJCBZ2Bd01N9POVq007PJ1qPecfiFTG2ZcmgD7xjeIpk+3huy
K1rHnhGpUXUHs2RutlbTCRemB07Tp0lBX+kylr0BY7jI7tF6DJ2ZAhF+jLWJyLpa
ibxMV6hRpdrrQbl/3g+IL0Eomsj+AX+QxFMh5CcJ/mHF08DbYohPrXQ5r9G1v+/+
r+NvR/2OOB88IJv3EKsmBs4tCOmsD2V7UmDT47S5Z3jrDOywCkE6s4+kJefIS5u8
PZ66Z3NI5EKczjGnaRD8wHgBK2UhiYLUddYwGyaUNyASW1ddlk34YJOurK53EmLp
Q4gz7leWM/z/HuqyeBrbV7i8/xiiCxGETjgu1EoHelJmQpbSw12SAqFOHMNTHO1M
26EqeeGJfDXXe9Up/eNJ5jMqikpH0JcAOMxybtV3/B+VQAfEwjN1RBzxMXAyysF3
/IrzlGb3YD0JFhWzr7ihzK2VXCA7wCQc0sFcgVeGd2AtjNTfFyySIRk03vEYM58R
kfvA1WedB5ryvDNqt6TZKM9stunVHaMRn3+eEBIlEVjq7u+SNsoNEl32+Hbh1mU5
KwRdZs52N26du/HQ9p3nBCDl5/etgI+EnrhuSyTnFS8SQmZUw/6NbM9OcvQ+hgLP
gcnq5TePPzJXN9Qlok4BIz4g6OYRL4IXFGaXzesxPTSl3hK6zSoE/Uwa94pXNAvi
m+aCs382u9M4eHBkRvwS4psqxs1u6XLQeP6yQ90UFXucEwb89XOVQQP03p0g5/MB
yRmShklmwesi3LloMfUCCokYMvaahUqOTACKriGDmdxAVZ/OoMhr4gio2Il23fqZ
eEfHgApY4OeNhNGXG4lA4l8lIpE5WYVUNIgY8n5LRVhSTi6zK53p7IA23YltNg9v
xRrlGP5BgAl1TtAjnN2LU9B6nY+DBrpxynbWcFLiGmxaItwTn9P4m+QQt5b7g+Mf
V0m6v5HtKZnqpsipzjDPSwaxDxYCb3ibskJIpcfnS0m2aINgzRo8oOyTRbb6zmXC
acRla/5JQYJeRfiG8dlx1/dJHfeNtfxwLrjL5DVcjMr4YC5hQVFSUCsqqaVoayu5
0WLHZhXQPatmTX3MOFjt1JpPJMd6ZSOAx6nEn0EOBtGRO/L+CVAPie+lfgbipjSV
+LGYduQPGwt4XnpHwz08ig8PpgXdWNtrF8vSAUXdoxqMvOGhkMnG8eJCh6YwOaRr
7Ihkw/muyFmpcF87bTgGw2J9RwY0HTtzrZWL1VyIJo5c86DQA8F5FM4BsCdmc46Y
dQ7z+1vgKRwLcOTwO/4ZPZN0Fs/S3+AO7p3NcExYcxrtJ/CVzTl50+55EC/AB83z
Brl6ZuRy4gRFe25ACgv27xLOj5XknvJaYJb1RFMXhL3OiGeblr5SQ753fjUmwhzP
grlRhV3eXfs+wc1upidbfsh1YiIHiF/zmZ5ie97RbtOCJvZWwFyl16UTK8HPVmrb
PrWbnYW0+hoLkZiJ6V+YhH+fHYZ7GiwXFhP2Ek8PpnQq/RS5vdzGVXvibHNN9B/p
ND4OlMWjoXFJs5RghiN0zdO83UbLyxBQkZE2Keohe/dm48mz0upLMiIb3ox2AkMl
op+X8MvqLUXOgUbpoZlobcBGxc7st3jdX3iOMMkk9FCoKFwJskspLifUrkXEHayj
5r7PNWfdultVkCKRL97O9PoLVW7mdIBjpZ9w0eBCzwsXz55ziBLyaj8x4mzLGqmD
mnz15PPU2g0mE/Tls8A5PeZLTQgXrAeVk9YpAaepQ2dDbNouXyzw9VML44QrSpWW
N5qFKWUpp3itxok8vQPlUq8HwBjn4obSFdOnFgZYsmp1NfjXjzbhMkm6K5JUs9mz
O+fXtw4TwkNSteBYRgs/cbivBwd1O1RcSlKE8TzDDZKx84UU7F7oY1JEGtwWV6Gh
F+XJaEF+8yLfIHJktrM1tZIME8ZCBowt5qUCphACdZHW+id0X2c1d56UPD1Sv30g
Dv0PX4oG8iAYKaip4VAN7hXjWpzN1qo6S9hmglSTV8++5f2+4M3CFWpUvSBL10gp
ezVBXa8E+tVF+gIZosUMILY6xAwmYdOsHNVp+JyY0VBrJLUidFS9Em3S+3HUhpIA
8BHc3iGYTp6rm3B4wDq/iej7KTjkiJcfuK+52UwfDk7v9D5DJ6o7iC5YFPCjeCF8
PJOJM0StRzE++q0Afty98nCl0oA4bNshqZfwF52jZ4Gz/6QBdaIa4fqHWM6MzQQO
eUjDIvG/PcJvsbYZf219aRuI4Fe9eB5/6hwAMTcBWUg/u9ZKS0YRIR9B+JZp/Vw+
z95mUVXIEl3u4MO1+2da1FZZDVKJM/Js7kl8YcWpzKH6luFKdxgJQgzRWF9tzrBH
JHFSRXXv8NWSirwAVYlXg/zjxG6+9L5/QixSj7kv8WSjZP/hlAfyGssfEnZwSv5x
jt8UvTegysT3gmUbeWVEcHbUtkR7NSsreXDuPmdg3EAvrUF3yMx+y9TK3Cj6fZBz
GWb+M6z/oK962vbA77nZeYY6hpqt9M+Cu/+r/3f7L+rsbl/VQyySbQlw6Z4VVx00
+nkB70mtBZ3yRGoKCzTexlUbJcS4EqztpTzO93bgxfjb+C4xIMct12L+QP1N1PG1
6d9nFkC4dbqBtn4QuEVzfsSNGpZOFwXojLDCJ1x3QV7qN+7SiP8PNA1MYfBGo6UX
1ldyM+J3USNYiMfm/m0vbmXGllMDArB3sW4/RN+2eCZMpLLaq6lDFpFeePGdAqy0
mTVI3FL212Na6HPPvtvMcKVX9qKpQd2rKBiMlMGYaDs51LpQTh7goMxFEhOKCmPP
RtuZtvLLilQSkaX73JKHsJaasvaH97LphdK/NRp9ZijD0c3az/T7fCZW7JwrXo1z
KIBvW2k+9q5M56MR9Zk9tdZJ11TjUwGa291FyRKEzj9JlvtpWl5RCB6eMsHVFX9Y
Jc0I2/E5NLDApU4EUE9GEF28uDyibGGtiGYPklKKlhsk8jIOeM3zm0yH7hvppLaG
H5+4JoKtRyba7dki/4Md9SYJbjoHwpV/9Y2yiDynPe93MZavoTJLiGIPqblOT5Hb
bIic7wopQdrVwz/DINeDvjimWARhGsWgwo+TCjP8qtMx9L07NOimlyM+ChxFA+9j
bJjfOVCkTrKo75m3VBcp9dCAnFXvd5d3pvIqpX0B8YNI8Fgz1xy7rK54gpjkbPq3
Vtd6KuXfIiBH7+EoXh9bPVAMsCWI4O+juGIYJIkecGQnmHwiwZmz7Xh+xQ/jSVOk
dNd75S0vSnDBZkOXNvJbrThhhSx8wv2gYIxnQENmysY/5u6pgS5AlJQdw3I4GLMi
cj2n8jw9rlhsuG+UKo2Sm0EX1QC0UczOp70TWcG+CMqSqrHn28F9+WjYgqyq+B5d
OJbnsAezHKIyYfd7FiH3UzxvFTQ6N792M9+YXx4scnrgz1YCjgXWw/parDC4aUdf
tSoWJ5ed3qhgPkK1+72YcQi7BQEvacv+nBEwULM1QOJdD2Z58QVo5APhobaix47a
yv9fVQGLvnVRrzrlkLTn2JHLYFjMR224SFETINsSKdk90zEic2aNYkmE5FkJXlkI
3oPst8MFLXD3evYe530y5J5k0LTot4gMKve1zAbEgdUhxSpV9rFwjjB1iIZmRfFl
M90kF8o7rSbNrWSOEtr/QOlyS4fClyZefmYfTy6wvAoFA+OHKj+pzC08Ez0jehp6
c/ulRMJ52/DAH+CmW4BZL54ibqM154qC4ON9m5FOy/eBfton7TsRzJ7Fa1IkBLCr
qNcG7HXgDVunEBISHDklvJqVBXWQ6dnmufs0ONwvPWnA8bcYdJXS19nEWkM+GeEg
zFHNC2UdjMI3LMey0w3pkkF6rDbNgRyrOr7CBD1e4DvrUPSbXooSBJAJ8CA7R8G+
FnBjg2aQK2LzAq7t+01czWCRn5qB0EpTc5YaI5Ja4KFLnqb22SCLlEyZWyrvo8Eg
CQE1cxFOfcs+Bt8c9a4hub+YB89u/+sZeL36KVxuMW6E69Sccxml3mjSyKGWBJ0B
vtJbF73vVLRrUq+wlUZlIZLcBEOa6UYMyBbvcjgmQm3FU4jS/4dVakurszu69Pfd
VEjydv+vOwA5WB2SWhvfBB0PbtqnBB5zMC5as8ZTUDyM5KfWRQGlAo1x2xZEM6Ww
TAgbMB5WqxXcRszgISTS7AuC0PoWkYopocIQUIfsEQ+mDthdu2DqYO1IeoIS7LtU
iif+YApY1YGrtfaCwPNJJ6OSq7Nx8+Tk6eJIbMW+GjeVLaItcsdITnxXwqc8IMYW
kiEbjadlpnP7b8By2AURDyLGsFqX8q8Bjeih/oyC6QXphAxyjQ/9NDuk5ElVJAw3
1hNYqtP5u3ej+Y/FeVqFUYfpZ4t7Inbu5eWk0Eq0IUGIT3T0rJymEBuTR1+vfGQm
mYIEuV6S3i9sDW/4GfZuuE+hxX/5qJYDAhDoDvbGyiV6UtXIZA1/CVwFlwhHFNQc
eNuJ/kVAAIT/lhCg8A59mndWlFaNy55QEk6PpOMXx+5NCGEULVu2Wu4vZtT31fGf
/oUosfZ7muFIyBMzp2hfPUlgcrOkve8pxIlQheEBswOCFZ/GBAbMtxpG0kMLxGbO
O3+G8a4AbABxzHE5ekwqg+D60/7RELgD9Vmc5uKGAZYLamWl/vi/BWGrFqilNP+x
z8QO8/mdF3bwczmz/nIcPnLWFLMHaJ4Wb/GtN/GXt4kQYlKpstx3wT4WL7f10Thm
cLIPDUMe93LRS0oH5zu614SRcOuUv+GDCtM7SdzMJFEaPkXXlVt5GvTWro4twiLy
pFV3yIAINc9xKD5VpsSlqDCEGjJ3npXlGk+zTVTBl5Tu/EqmnZDLc2ldJWGO4gg5
eisU8gIRXH0sd3MSyTmzco2QizObAXNNRVj/Ptp8kA2m4lxlVXUwItUEhtdGpQ7k
U1xIYddgYFLQZgSNDUDM0Cggn5S6RaSqlQzE8OwqAeO42conVwhjU40yQVvkhqAo
mUDRoWa2OrRjZC+yr9wK9ucuwRMFLw2Kn2WQH5TalAcOGMyJP2WcuD7ULBsL5imh
fBjy0AGC1LG2A3Z933iHvP9nEyU1n+cN1fe6DE1mU+k36DxzaqrVcYA9r2AbGEac
MutyNP7tOoyfgx9wKULNhGeBi0hXmi+DsgN00hZKFZufoEQgSQKWMb6gP4F0ZsPk
XQmQvPCvkgT4wVLW0bN5a0unb2TY94u5PQ/bjUSM/dyo79k0osp8aUyPQVp+T0Ds
tGVcGwDMZ6UXekaHduqo87QysBgM02T9uUcMC4QiHG62rl/c/zUDTVw2e21kDKMt
/Ggfyj4D2IBt2HNcN9Cx45bHSQGVLTAOEcxRSNCB5gLTMzUFrLvfl9HNMamJBzr+
9eugODOcYkcrFKoENe9HlCaUMMH1SsmN5LLH7vB7gZQMKNxYPdoYeJ58Hzc5dYJf
rHnc21oxz8g2MQhjMA8lv6Y1dd1f/QbU9rU68jMWq48kfHT19j7WZ4dLHLOcBJyf
sUv8yNlKn0mooJBjtv2VTSHnGiHQXlpoc7DAuiqeqCFgvZ2BuXf6ZQqAHo2chyQ2
tIzm7EMYegPNN3QFV1g/gPFaZd7JzerqpS/ihxEgTPX3pPeJwhjnyVTNDtz2O4sR
CwuTDglp6tt2l3GD5cLQTqdPgXTcEY39VbvFucOIQBOGIEvc1jJSYIpXyW6nXpCM
fOK6qqDH1fmsn3km9BBGQRchTv9PlNR6T7uieIP380IsXmzeOMt64haC6eVOd+Lv
6hvlm7IfBCSl1lkBcXZQ5s7famS37rRql/O32mDIzpButuAHiGf9uIcjXAS1EciJ
Y6IXwhSkNSL34ppSjUjIesaZJ++d8CFRRma0/X2GF9F46uH18KQYPLO/IJ054MQJ
05EdcyU2lwI3344Tex9vy7QFfo8lAM7vxAFLaHgWDQGOjkHHpZSjCWXVKV/UAtkK
lrpyVO+zNKOzAotF2g2dNFwmgK/GtrcVBzhk68OhNO/7sOkvgXmqueC7PbltQV6y
xkXmn3ZYku8kVH3Bv0P5P3IGQB0hrVygzFqQ3/LRuW61p0E/eOSqZnxqxkuMZi1b
3Y+mptvMtzeEmPk47js/Y/SU4+16qoCCpCWH2Gml8chsklRmzYtPcf9s1Oev6x9f
YViwIB/ixZGIiSgQ0uvT1SxuoD+tRYDuwnOnaMxhZf67IoJYhaB1Zec6vVJY0pMI
zYeoRsvkcaQfyRVtNLxFJ8Yrr+5wgZAX2KX15X0CqX7v3Mtt41qcH+fuOClODaCO
WZwBxqanXC59xnCSCBGRWbmmoDuxaI9m6gC7ezZAg1LpUSUfVwDoGJ2+VJ6/VXrB
Af8UEp0KPp2n3W+a0Ufo6KIZMQv26VlNKIQXxDr5Xj+Tcpcp1+rPKFK32wMTp95I
cvMzvMVDhJ9Ca77p/HPn1kgsV5VvG2UJHLuXB2Vd/eVtVXnU94sTdeyJiJE+j4FU
jaRrQjm0rvjI6h5kISlRVjBgWOzsQslTTnq4hKPCKU3WZJaJbMNh+vT6mIHkcJow
Sw55lpkKogZiM4Aqw+qrWhvtzi+rSXQE4KFWq4zZEN2FqE5W2sFwQ7IkNIGEb2PV
sXX3xO61NIO5kShOKRrF2x6GEkUyH/PpDQQ/b4Ijpv5Jo5CIX3t69LAvX8qv8BvS
0uNqeFBEU3OEVjUwhoomY8jOY+k22kA8vjbf4ZqP8Mg1PcmcSgP66rVFlI8B+Jk6
PvqlqRLXD6cihzVTzzsytE/rCJ+13cR/z0sn8uH1CSJ5RW835xG3u0Q0IRoEZGPG
6BVuxBU7NgO3H2DJRA1bKUmw0grkxEXo9lkOjsC1qRmzQW3OPvTptB0CngQORuJb
q23C0TE7h10Olq6nzXoytNdOGmxqA1b89O22nm58CCDRhwauNXK+Mj0wO8OAYEnR
AwYa3ADWiEiZ8EQ0aCZuHTClwEXdgYJeh2MkCGj44Cw7o/keMqI//D4L68yocFkD
inKH9cxyhCGFvaF7ZlG9lM65JI1i+Cg2OVidKNiByIxjogBwOwWbHs0Hfy3fTxEU
QGEHf29SsQBeTo9DMlxCmfZuqM0NVnIzyhbdyjgSb+JY4pIlDB9C6iEc27EX3iPD
IPRq0zR4Y5QrXFOWZOeoR6WGMg/vWtpTXtFyWy0yJItJEklkvXHtsk8Rwe0M40XX
zMW5CRfDjagU1aNxaklt6lZFtDgaWF0i5OK5QbPDA3hBNsfdFbGd0oXiJYt0G3Yt
kAecd8268qFkEoj6botBIoU84jrvaVU576UdJYDOyyrMJ/za3zu3bZA2FpgR+PTa
+gZyejojN+49GXcl537kU/5VyBQeBgiMzFwLIqpna8xYWt3AjuJ0BQm/U2kbxoXy
81F5BajzvAS7G2LoqaGw60dI3k7w6d17pfL2UBD4mGfZ47zBC9s7uU7d57gz9hVU
CgPAGNp0Z136ZVtm3V+iDDPhSyAutLQsWqmGx8RK0Kw5sRCzAd7Y7R+6VmRpJ97f
cAN9VY7gP9HQEkJxNTkhFc57wqP7POY101Cv/UfIbSnDTcTfjY61/9nTJowmSrfH
3y0flz6iRVJBruUW1FlgbqG7oI51vzDHJK5IJDbXjXAFf6q3+VJx2TXfFCuVcjdG
xXGD1bv9uU2ocM2qOUjQbwPMXY9fXrOTW8y1xegTx3H6ziWz6mcqkDUjZW4DzyEg
CwmqxXsj5URfRo8NvBvjtcCxoL4U9PPeNkG0eZNwKYNFwRbTtLv5blCqHrv6ouvE
Pf5tgnhBnYJN+Ij5kWC1Km6wnupZCzX+t9I3x1rDx3fuW7gfY2b6KHryR+JEeptp
JtusuT30L9iPathyHWDVBSgoi8jIvGtzxh96z6KpycjTd5Wfi1qjkJmVLsgF94G1
am5tSgKeT7Nh2vXu91baSz4Y08iEGmvIg/oABg2cW8gZdHC14lsz8Zfce5viIOb9
PlbHQrhWYbc+sNW7DToVIjvBn/LxTy4zb4JYJxJxqfoTR5slMsVscRnKfp4uGaj5
E5ZPjeuUfEZc+KoYa9/FBg8bpXN1i2MdZMvCp8qMiC4ULoi/z80LCf1CclmgeubV
MFWv0357qHA6fXjvrxlXmlC641aXvi0pnXVbix8b0pf4TuiJmAsQSkiBWo+GS81a
3/OW/cqaukc669MlQNVZgampG4ogltuaCf26D32tyYG8sXLjrUHmHdDPifa1+CVx
SbV5Mkf5snCdOquEz3CJqSPzhfbEkOLAiufi/Ojmj7GyuZNyeSWtgq/WBJt6tdO3
a3sZ5AKdzW0FJ2nGGxR0kH48qRecYvZa2ih7sv9ZWOPS5karI+L/ZuZpY32D6wDN
v8Iml23IhM7Om+b23gTjlv4SN60XvQf2nILsx1BwphLZFzggTczJX3FXlBb0/wDy
dB6g0iYgcu17QX0m5GNQZaqPyFsNZKbZZnnFQSGk5IcEkhgPburV2NcqSu+YZDXw
DiCVfbQVaj7LBX7XenfshFPPeyk9t3DJcPCPijUmsc31meN2Cq2MzaBS2XLsNle2
9SBA+t+jUTATpBkKQqfutEexVRX7eHfnrrjfqbWPsZxG0A8ZNngHRd3bkTRyOGkk
+eT9NoriF6jiOAmrlWt+TslA5ZX3SH2Pt9UpL8HZ9Xuks3IxvcqhuItIbyxxGmDr
SegQITPjVdK558DeqgA84nBQmrNVWVKDeEq55Sw4POLHXhFZtxKTXTE4ZNiCHdq1
n3WjZNa9xQlTObiVc36eO/fA+HSHCEW32jCxIJc/HkV923hQUdOFKZQGef+4jH4D
iqy0i+qJU9iOO9DZyKKRpknxNIVgLWxIp2aay4zf+oDpo0rhp2sow32cPjIkIqmS
UFwDZCkHWzuDAwHCmhQN3zn+roQHOl9hV3GoQ6wpSHZygKwhnRJtJJI2MLbWfWP8
BMTz6NguRit3O2qRlTt6qazhi/OFsW7DqmS2xERK/UbUq4JWOZgPuxKh2jRWaaWO
Q0hwO2LTk13R2etdKy/WtEYrlq7w+oMVdwODVyHgtQwTCRDl6jf5FQe2GKf0+gqd
XVZVDbnYhWHVvWi1Sm/HTOoNTkl49009mGMdhfXsx52DMddmRgxxnt6ElfhNunkk
5hCn9QvuL18rm2B96Yh8g301q7jOX1EGpOmBRMmQp7R7r+tYqCRR2J9pNaNaJFBI
a1rPyVSU9Tm84A+6sbk7tVu/RAh2gvpw87VcNECktFFJMAchpGo5CXenicDOMkz7
+bDGvG0b4WKageqkvdfDLA3kFKzIGmsUl9fn23uZYUhFnXstkv9mrSQSZBNlz+zl
5pUIVU74qghLI76BkfGeZCBFI6Da51eN3O8w2/yJ8PIw93coOtYmeTu/ibfyq1Bv
roMAmRGnOd7q6/Pb+5vDW+AUp+SZdM61B4k24/0QrfPyqO3vBGHS9sNVB07YdOem
Gfh2k1lzdbaUVp2oAoIpXbco/Lo35gjeXR0kMbdd4oUrcNnL/ipCHrR033ceWFud
IXVH92KM76sdaCTjRh4EjbZf4a5uf7IEJ5D/y7I9XjNl+MEuhEj+9CpzzIL8SmD9
qJOkFB74JlCoB3gATNzyXSc2LJHY/9nqyi6/YDjzZ+yS6Fk5t8Ogx2AHilpyaKVV
TARKpb2F16YYMecHmFmCZ+lImObI8kCtEx1Ie6L5d+Im9BVyaEVrdKHij3jYhBYn
/e2txOffv5nACPljnmfkLdEzjax8rlPT05bWNH0CAcyke9xwxjU5J1R/4uQIDh9F
9cJZ3HHKz7BrHXrYpfNkSF4RGyT2AFN+QYDS5D0H9S6oWULFs8ol8AqJ2wb4y2Se
cmLV9zDYqmdZf02+k4wWU96CgBQkd3Kuv1KMguGeSXWwGG4oLm7dOetWXW8xjjnL
HXV5YgqJTgxGeGnB1h9W1LIrXKKkNKnCMntajcEtYQoiltPLRKCVNuWh4E340qf5
gBbncUOSny4FDaci19e3s5o4LIGiOjREnVWfQXSeCIvrRBSPT9UkicHC8hU0Nup1
KvPkrGIvDCmxU5gtUvRFIWbx+dkt3sqMzsFzjqNNG7l1iNj2OotglFiN+uNTrw3Q
LkTMCTF5JuJ5YOJaRnGuPn2UK4rfxL0wsvNwL03ricZrTqLnRrEPStVkzPFOgpir
fHk6EELVJ2q8jtAMTYcSLbu8SfeMmPdiwa3WKlUn867bOLeyl8eaCwW+ml0Y9YZY
wYRhpd7InTETd2Dce2s1eTAuBhkzK3k4/r4BEuqL20B5xVABs5xgEYsBF9H6m3D0
63sV+CqscNEZd3q2L2I8uIEWZ89LFR6pfKdmuB+UR7sa/cJwi+PFFPSnHjAXhpCZ
ryYjK9aFNdyGQX0TCs1VPutVN3MEi5AHsu4gWH6Z2NXDVQ5QTH2xTFWgH7D9IFt3
P9gFadnoNWTImuVdeqCAnMQPrNsMdPIFGDwY6CQIXbyYQ8C5PUVXRjlsomVc37VB
ZLo9qw83tJqHsKHcN7GInPftNOKd/AJNClhy1X7MxcuTQPA8DqdPhVZAgUdXlfyo
dq8VfAcpe+2NB3vqcl8O7rPlEFuF6HNi6bS3W1aE3GFMK+fH5vzzY9/sPe7hdF7w
QVfTZHbNsp3IhV0WyaXKXwb/vJOEKhlL+TCG/znMGvcbmSnpkafeYkDIjTO0Jb1k
C79GQceR+sCpziDPM7seTINrKUkUouNxxTsw0koVr5IUML26upDTsnNyqcmdKhw8
p7ALrtV9sko1pUbZSNKqa8RruqlyH/tD/jfdPVevLIstwnajKMcBPtgyQ0WIjxok
RF42YBkrtGotBs2v20SJjEDe7RfOChbWCS39cMSDw6xnEzEUeq5ulnDtQ341KRPz
2ImhS9Ik6cWAK9FCiaOpCG+4EQhguRQnF1vZOXVwgOFfHkpLVMk/nUkbxQIJC97N
SAGnsSZ4quhXlPlJzxbFX0+8ZwAYaq9Lxahc/dGJ7KLJ3A+UPTJSO2neANdPX5rh
bjqZf7mpY+5GWwnbTJU321f4OhOHLY+CuXTH2WYDKBY48gPsp5GT3ttu/tGaaDSE
pj9mFp4mruIvMeoQg4r6bqAyBYIU5rYfaeMwrInWJsjoc3vcQfUnAc6dezlwdoxb
oEvKk4OLxYJ0fsJgc3qPFINjY3FCoyy2B+14fzdL/INVUwwhaIfsrBiuhbCZ3qpp
UYt6w3HVgdyR7i10zH2eehw4QTtDf8PcovTjyEs6eRvRp99m5+DxC+yGBWEJX7ZF
hWeUKt1G3+O4bT/W/Pg3FuHMSbBsnUgzQw9qYgvcSeMR5JF4E4HKq4XSryzseYj6
Nu90YFjBt95HtSA1M+rFL+VRB6roby7O3ifi8M5b9w9M+nCdySwiEyaSymsuO/mo
3bEvtMtP5uA2reP0Ijimz6Tnqtxo/JT6czxmKgg1HNywN8R++uSsXfsQCJuadD56
TrEBqPh2np61MMEQ8CB0TlsoS1jhWZX74FAT0f3ZFsxqdCtPlKFnFxtJEcNCPwee
uMDm4vITnC6h8mUDZvBC+VzD4qAuJjGTDyEkAjJj1it4zUlxZ8o14IXpjbOBWePL
EX6kSgTnr3W0XBIBHcghmY5/7Ft6y0Cjrv3aBCO1rLnOFd1jhr8MvDB1kIWd2eaq
w0+lOHLMm6nZLfC+nDWOhypxYCIQvJr1Lw5VfVfOCI2UIHqJvPSJMRgfoXxvnejG
4XF+W2wq1YrQdz0eZZDXg//tSkUwWxmzVb3h/fNl4gOCiyQbYx6+aLw284bQTJq5
Vrbk388cJRgMsuVVSMh8P0JdyEwEpmuQgTYwUGt/IipIczhYbdQXHx3TskrwpdTz
WuySmLkF27bHCw32ouSkB/S76/zvshvewGTLvF25Ar9+YDnnhPbN7bgGIcMKacVH
0eg23LWkisQ3bFdKGcrTXGAbp8zunWqAvPxuoFOthmk1brOqPTzhctxActRZfacm
BxEZ3hxDAJmwN7xbw4Lh8AseYUwirMOuP9xrMlpUasbRsq28DFbjTMmKYuP7Mqrs
L8u3m+PIx5mlKWs0HBj8Jy0N5+i2gZbNYkbXy/NToiCY6qMQlMslL3MNeE5mP37e
CxOAZuAo1dvRCOhqgNdeJEcZUD/Tpafk0G7ft8w+sotEb90UgC3RJr4zuLY/eE5v
m5O0FX2A/EkF6ANjtj4MIKxOrP4EzWCDdcrFQ72PilmjRioHZkKx/w//tUkk78RP
AkWd1+5F6tDbZkj7FiXgjVd0a9Jd6XiIiGW8p2FFbM1dTORDkoByIvCDTL0thP26
zC2TBEeh9m0Ddnnv3ruF1zZ6wDiwbfcmgEkkShoIqydQ1NC81ZFDHXtxfbRxyGh5
rM8D6NiGG+FRbOH9/FESwfLwpOvkumRCkSpciN1pFRA7OhWe7ckgU7UCgYfrlKwB
Sws6BP4Y5Qjujerj9E2qSTD3dAqLO9J9gOxhk81lYsUpq1xTq51Fq+WoQAePFoOG
wZJdJeAsvQ0/liDtkOcjwe5xdvQsY3wrDSDC2SQ6H55JoS2WRHX0cO9lSxhpBc1L
If+59bJrum2R+PjvjbAyx8IR+BpfS/0OJRfYZsnBwhEN2PjYHi+GqRMA3uTFoRyt
rlGyN/FQQQVpN+YbOSKdiWAouI078N671+M6mGHCQNdHYRNEnrZUrtyDWVnEox/t
dpKAPBSu//CpJl4wwPfl63GTA7meSzo6rHPSnuIcK1QFvFSp4fyoM6oNi69NleLs
qWT5P4rygknt+E7xRsj8LXcMamTiodGgFBryocUR+jjke7rQ/MjwrzbYcAlTdnTX
IPZcJ8k5bM6Rvvi0lWkDrX4CfpfyVw6fcw64AYsOrT6aoEzmPGzWpCrJNc98FdbQ
AcEuAv87hdTygqt8wqpggQq9cZyuoSOWgNg89ntNCMVJ1A5q7WKoSNdPDOsereHC
TiqCgaECoO3nDISQrxHxTvkxNQgUnzq01edE6Jo4Q1MnctVSN0d2ZIiwRK6J6ty2
xcPWNKGnTBQQ41SuwgfbiEs1MAez9vrGM4uzLv7sgXfNUcvsT0l7qUayua1ft9wL
WtQWBEV4tUGZyo0f57rbwx5Jmbu/XUf65vKWmnN0WgaEO+QmjzmnF2VQVsYQElPv
Yf+x3Gnb7kJNm1XNqnureE5r7kj7jKOnPP5fUh3KEh7kFgvqL3coDV/pSoVxuarQ
win+LqKjOgHxmDKWoNnEpqBgGbPpGaEzi0yq9p7TgYoQof5mF87uBlyZmMGC4u9N
mjohijbaZC/MM/Uu2b5T/dt1R8/4toM0566BYUrEMdqH1vn3wht9DU6eC0HiMA4I
C2Jb4LQExa7FHRZIhqwKIAH9pStRnejuOukL/KZFfXZGW6g1sHk4+RrWhBijUnaF
r142H4M4i74DBxuB05jp8/MHXv07vBAOIHsUrMjKwGVKH465S6ASw5uNnZy5Q99i
MOn0C0K83lncHOo8Bhh00Ajm5tguryunCtTNOPm/AKctPW7Yw8PcqbAyv9kyM4HO
eTP/pSv8y9njkvu4MdX4ronaqqJuI9B4E6kA5kNa8u6aRjLfdMHQOLhwvnX5fXGn
76GlzMIh9W47xMb5VYnhjaZA76v0KeI38VP1zrrrrp5DjP7uywLxUV3Xx4BIEuFL
uWOvlJ7hQzNLZb+WbAxN+Q8U42ip9UK571Sonjgyme2lOfrF5QADnTVBWwaWFGPz
7H31B8XFYelr1VCJJKwitB3d0PsZZBczeTpF49GglrCmrxYGJVQ1Q7vQVc0l1Qco
ugQ0+yW0/KI2ARnHYsWPDyaI8gzMHxhtSi8S9wNjg0fJELkgND8nBeFpLa9B3iou
z1fQni45ah0HIubeov8wo6uwJZ47jVBuHBHbliNrC3WxXvyRhU3Bil9xOx1sF+M2
ZyCdCOxBcunFEqaRRCrh4i5CCqeECui8lrAQS1y6UxboFAZFoBmLrgJRUNp0GD83
SZd4wEo9u0aRQh0Ytsa9mBXLy7tB9xIX7meUQn9194u0z6Dr+fDTeubSOP37PAK3
NdPNl88rERSzX32g0m6kBOuRTZU5wkVkuari6pnRcApwFoE8n39YkPfkq91FhnnC
MDP5Egez6uHItiUPVynnaCS9V0rAN7+p3Wne25r+2PstiJBoexE2Hk0aObHDp9ro
Ad+l+208UJM/3ZBkPclIhM6N9xKlbcxa7GDeaPBnFLaZGN6UtSA02lpU2N2/MCNi
iS867JgHowMdZitQq6oeZP3OeeO9iOKUDR4+JM5A5t1OcDnHCRtzxAWweR8g1+9S
/SMNS7Bla+uvAR+V2r7l+P8hnhnub7QcReA+TUCaQlvUdHZPTFZ5r1nFLInam5AD
FEwyHPZLIoHn6djyyDV9V1ZsRw859MKDMRi6/OoBU7pY1qMIM34IIgPPtaspxpZY
//pragma protect end_data_block
//pragma protect digest_block
yLQqZzbz02QNAulDDAsQrlup4oA=
//pragma protect end_digest_block
//pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
EluQikk5tXzsCVEAubyQHlDpw5ka8DXrNnmVTOMdk2bF7y4eeLwI7DtwpuCW3CHA0ca/1yRUpF6f
6U9RE6C3XTRaHHGZXwOS9q7Ie4DGJse0Wxoh8nizeSwSspYATQhqAIMgRV7dhG21VChfe1Gz85cp
vXAtcJ0AE2h2tw+6UHJVS7IPrD+GdH/pkcpFYj3eaqBhxdjXeKqiiD2aQhDfMl6BN8hOxkknBX+4
rdKrRPU92rXNWP53+6e60yC2sN+JQ/jcYoUvbztARVJM4ayAG/lzPwH4DoFVo9/wJlx6jVb3EYGp
KLkbXBMMmot0Xml4F61RwBHHz2zUYvKZH4sDRw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 22096)
78gwlQJBPa1C3jON/Y91x+fVueEDvk9lJY3y7su/pRHYTwfwjZbL9RZWl1FJCf5iDGKx8OrDFRN6
UvSNvVAroJ5Oy/CKCVElITylJL54O/TSkwNL4K3MLrps9Knazrojq9JLS+qWpedEOAd0+s0ypjzx
o+InYEdUFJfdeTS8e6lJ2ENoV2257n76ytWwnTUBOUi0Xlp2s/cZEGnn9MdRDUT032X6zCgLhEoB
XAoSRdZEwLyD/A8ouzg9thsO/pA1TyAhrKVHyYsyAWMq2sjO2nh3SzNVSMrGZ9FUEt6olu+U4Urw
eIdQ4poncOfzYxDzlPn6YlSEx3obwunPACuJ8wnzikcqhDpP+cqX5Qos5DRhZTDA30by0y2xWNDP
U6FQtCMBaWzYmFbO50XhX7dsMF8xblnuuD+ey7hatmV0Og6TZSqo3Zr1IP0/Ff3J5ZX1BVL1jHaT
gGouKlRe8TnrzUKsyTYWzpdOOgTf1n2hjtuib7quleYcHgaY872hkbCoKjwFISPhLnVGViRIjb9q
O1ncxgd006Dex7UDHyen/opKRdpd4hATFE2uoEDr2Oq17Qf5iOvn3xVVe708G8C9+Ic3S+HnX3gy
iCOpzCSOg5pKV0KIWjfSdPpm2SCzieeG1Nqjp6iZYG+X8cuG0cxZH8Q2a3z+crFVCcTDJyuAeBuT
7p7oBKyWqxlq0kDiYXGDZbRbLhPOZJI1UvbUfKg5LXeA9TZWtQMB9lCCmFOeT+9auTH/82wvk2Is
UxKhqAtyHL05VB4nvZiIjsFniLpLVLTrK6LrM8zlF2wZ3l7eRgiSJKjX0u5InArSqPodkx9n8xDk
+qHXvYQBQHbEG8MaW0etlhQv8z7VGo59CMfiBKrWoun3BDiJX5tTuROGTDRBESCMHX2llCgdTzhh
hSrD4gh0nQxLAhfR+b5CfzZC6DE89fbhCb8KWajx7tAp7dm94UuiOJVuoPrsbFEan8pz+VvDfvvR
0P2wnbgKabijp416DdxVt6ka5lZGHdX7/WcR6QA6j05SXyFEj9DwYcptTLQUxQl/7pA8bZHFhPg3
CDviWfFnfY0fqtya1sqgnIe2VeqMFX3fa1X0eEuqPnjXq3Vb+MuHk4iHbgi9qZQBqIIHl/HpOoY8
cFgGMurchNGIxqy5lJZXfh4pFSw8iPW9kGtxvEfWPi8mVQ8K8dGSaWpUH+kdnJi0orFquI3Go/wG
mdOGNVTocZIV9B50TugS57sIpW1RnpJVs5Ls2umQB6Kk9ADFFgV5IcmKPrqQvbgrhV6CPjo4A3vd
muWNt1MinlWrCLZ7iasAx+DosHq9AK+/MhF/t3i/pMabMJk/Gluw2h0WBl8Cjn5O/7rB777ULWMr
jkG8v9VUc4SOWYTeKBFV9oF66cUlQcvszSzCpd6giujNuZvzciErgWGgdgyM/vLXR7pKBfIldbqM
IBOpHEAQtpZAS4meM5fWSZ4vvt2mF6QIYd1fCbpcM+YrNj+zFY12Z94wm//4EV0NHHhho8PHC3UK
eLysG+/blZ6isWAzfwJRBZoRO31iAzP99m1UwtEhe8DdWJ8Oa9l+6dkKYnHgefUJ4zJkAH0T4JTl
JQtZ+6Fk3TCo5D8KTyTvZLphgkS5Wdc1KwzdpNbTPd/4OHUFs775lGMvIhm56P+UBYwRadrl3O0R
lBJ7lLXtHs+F8mxbuf2M6Zw5meYZB9gQ9l70D88B8b81/scRQS4w+KzQ8RfzMyiYoF5kNlk7nz90
m6yYGTTYKnI03Nn7u30Qyhg+LIBQVVEmEqEwXmrwTXod87ZfO+EDcx9DKv9D4phoKRBZj5MbaqE5
rQsa7osuScwQpB2RoBOzw5RB3TyQrn9ASmMT0Nsu8IYO1eVuXPxGZUjwSa918oG+s4ZPXPfBAcwJ
6OMB9kjKnzmByQHT+0F2ZE8aUt2oNwx1/sKJWpfOPnHBRzLVNwRZ6pbpHFiT4iOVHoUC+sMRaYnt
0IOprtJAyguflXqlBpFqwSJ78Jt0kz4D83g00A5LZra0Uh2KCWVcAlRZhpewzU6rzwHBLLcmL9m/
QGfqehRFYtXKbCvjcumNVpaXknrHHZdPDALITNyHP57vGOGUETS8EHoHhGiYTP32o+3Lnd4owfG6
GTFEM7ru8+IABLUKDv/4/wYmOAhSJHrsdbBlyMFwkJVcZeqE2uSfOFwjl42aX/DKlARjx+RpiIa/
MK3sLg6yD9/t6qX9v1j46uUarER+u5xc3EU+rvYy/HbIx91nlMAk+SU1T0J573XPYHkUEjITaXP2
TpYhp6HgHVWv30A8NDKd8CoqLliC0SjH8O8bAYKVy5IDEE3zmnPrvQWy7ZzPAyUZYoC9lXQyRfzP
MVE0P1SbAaKGoZchMHJEp0cAC9EczIr9UpcqgV+eAcZNDAI11SXwukt2Bnr8YB1/y8E9MiUNg2HT
q94X344a4D/XH925G+0ZhWFn1qOpF+yDqcC04/WwWI3S5+Vfb1AXtp3g9w6bV+mjDF9I2FJzw76X
6XOMJFZQ0Y0hoh0FNM4GsWitR+LTep+WA/C9qBCntAtVFdsWS2C5xpQB5R6ev+vP/ZBGhyugB3CW
mB/LAEOs0OFlD2btgNerKmCG3rB/2M+oFSTSGuN4AdYY7Ay1TCfVqROHYcuXSublm46PmGF5CY/u
pl+2wGRBtmPND5ahK1Cw/KNJA4bd3A2+bVASYfjhf+UvpfAqbqe/fufFFg19j1IPSi7aj3XIWDaq
lRypcCXKEMdlUuzeAqe03eT7Jmbk/TfnndqIKFOPo60l7wjhg4+AKAY/FOdak9G8XJPf7HU7Wo7i
uH9/yJop12gLpU/Jo1cljnUwas1m6p/d19EvbU9ElAVFyzMkhQuPVQS++anx8alV+JFqpfWCQPpj
KwF2kGzHhMNXVEtQzeQLToD4C1TZBBOFHVrmsnqWqDqA4ZxPyFwPiMa60kd+hHzXSIkz4Co8Ll1m
6e8yDrbkpJ03b40pc/E50fU5dSzTbo2aMJAABfJBVtcgsR3BlCAMTUsC6eQjlMnejQtpIBY07SSx
QTRuMgUHxhMN5LtzYthN4lauYeNCfxLmAodzAvsVCpBx3PjholnlLR7XoD0+iSCKh+buE1uq+yd8
8UQ0wnBGdPxWl0iZpCRmywxo5Xgq+HvHHlCNpV6uea8bLAcly1G5kynZ9LYf+89PmdoEKZZiMsl+
8VkX0Qf032Nd6ZOlPwWZ9+nzSx23uYlm/YkKN6cKoM0SscS0GjDJtYMIk7fxING9wELdJhoMEJOC
gqyhL4pgzFSvzSzEoKOZdT8rE0rgNPSqlR+W8soeWXp8yUO/nyd8eDE6E8r1vhGPs3kwXeaJi4Qc
jw7QtYdnLBhL6Y/GBOQbV4tXJCCXvipt2uQKXjQKpsJK9sbHC5CKf57WCBEQm0W4+56qtu207lu+
ADswbsPsejxEoX30qnaT58nJXrGtDS1HVCTp8naq7XzYySGPtixEh3vXnE7/HFQar+5T8eZdySQm
uMCSJ4bwEYWvtdps5Iy20S/oO7T/smOhqrsP3RcVGtNNs9qvIbNnMKczHwRnWOlFZck+bJTJI3mW
BOx+uLpFcNF63a/cxvnrnJT8HTo5D50rP8PrqHzYutwHuWGezTQef1S9iUNuJHOs6pxcugbMbuNV
P1sladHGeu3oB0jFFOzHmmStxbr1VJMMlhgHCQVnhExULKTXA1o8hAjKW8pgfALXI5bxrq14dU0j
L+RE2xUkOj0VkC2rDidW9LttwaQVV6VRCGZsVII7Auth4CqTyRRr0rFcHGDbohd0xscoC0kZ4wBy
HXw3pdGl32JPEa+8wxofYdI3lYep+NV9ae4RnVZutZM5ICuzl06Qga7y3474VeBjoN9dStiTnAbK
bVBmgoHp97P0ppM4otFxb5usyxCTkrEE4+JWjRRPTpquihuDspjcLAaXqW5Kkfqc000+5Sw4UJ8l
XkaWTliC0CdxnzFjq88oyCOvpHbpyDy8brgZ1zI00AqG6KoQUUnm0LATa3k8WwaaVJgnVHSosobo
yrKyLLa0LD4XXJynCMNZHdONRVme+cpB+1IPVgrcu7W7L3CSSMPorviOnVrDBP0+lluJ+tTRdM1x
tfGZxhqJ2+wfzJHeWjjnWJcQQGHGQi3iBEnrcMKsN7Dtdk2EkbR7hEFOc2ZwyFGMj/9HTyei0cSZ
5w6RyrxOv6LC5toXpquuNofXwThI50ECIbha6tNU7+Vok4HD+7G0ViG3/2QnhfTqTKbnLwh7xW8e
dsGsUHShdA3lh6dOBkFBwHLaDNd+bhp4FlKsADoTCGzR/sDilDi/Tg8lPYo1wGeec/P69zXZyNDP
3jdDh9zsGguPaMpncYSBmNj5HLiV5zM+2xrG2z44p8AlRgPGQvdJX2idFtVBrpK7gxbX1sNoiZ+t
/AIB1nanWoT1nVV8SIjHaW3gnAAQduuH6voCy639ewKIGSCVeOUnFw3i+dgcFoTKkmKP8pUk4vjv
70UPAdFh+1o7AeQIO3ludqsMyaGWUf9AfZH9MCgShBDuzs6qm7WiKGLMTPLjI2j3MWUweQPG91MK
TZi2jsif/vTXnE0FFxSIhkwovUXgAW1X2Tve/eVgIAC0R2B6yhLwkaSA98BLc2t4ff/v8zCX1IxZ
poakhVLIY7T+VG8O+UIeY8wr57Kb8yao/VA7IhEv1m/9yKt/a5htgg23dEgoaoSqHDtAZVRwQ065
mDYDCUjH8z5X6WGI7CTaZlXZ8277UA/I8d9MTJP7JklEP6pH8GSP31s3WQPT5c0mpgI59DC0Drh9
LIUjgTYuhOR4MxHDpByShG6Nx6dwhofyx1kxf0n9IW2aplX5g19G/BJtz18FRi36XBOAUVHR5N/Y
uvdooUosgMB180roAknUEfWB07zXwAKvs9OBf7oSMOJzfOFedeHBkjAUpHtOlceZ10j1Zmx594tV
H7qno/Qo3LFKgWTxTtOb4CqX2tOY1JTprcbY95Kitkpz7rvmUNNuOLli+x1DvcqywnTZr6t5LRr4
KJfRtAqQx73JqRRuCkXBB+BiOfBHKzhi8+wqd9ZyM8a593kCZllTpni7vIZXwM54K0p6N0UR1eT+
evgXLWnePOPR2xUBc6ZLNStMZWo9gm8c6sCZNG8lblrSSc1HviCkvhLht3Rz4Xs8wQZ+gVrW07Qk
O83RweXGFDcpYQr77gqbxvMujHdlgYoizaP505MgFuwiblMeO9IOtQeBT6IM7Urho0JTywjZiOoF
s20KYUQlSPkTLsxhdISeBpTnNlLN9Ov4N17ZWPHVbRyeWdW98GPrEsenvjuIIdY7p5SqK2GyyEm2
YObqLv0Q+iTfJo5Sefh8xFsk8JVMxS6c89WrlJvz2GKnxZfhfjRrJluUVNUwvALVfEClF2FJ6uAO
ikLYFWuhXWb/3GxmPpvRv+hlesr+Uar2ABKBT3u9GwQ1AAzvz5gkU56j1KuYPpZGXbGt8+H3v9vx
o2leLq84/J7I3JKxt/bueB07pZ68Yt2F7bVgg5RlJkV/Ob7B2d5OMt+sLs6iLHE94rKwR62VMifg
iotRyoOa7KbMC0/VuIy7GilB5v8bYGYpbJcKOJK62ITuFspe0E3AxiET1+EW841iPhU2gkWCtI3T
Myt6glrkFo7Kiiut/otFWM0BC9YJ3I1aj0e5SmeBDDnpmRTL40H4V7Aog88H4kQGcCvnupPx1NOj
opuq1Gdktyc/J40IkJ0J49UhKQ3dp36B/TBCl0hQ96PF+vKySZ95iWOOmScnaaAMorY0LBbtOEX8
ylIwyD1rthGxakpbCTZSqhO1i4d+wzewv9752XhCW255JpLbFe9LSmBopxCrStjKA5iFjpwzmJP+
kflDfu6+A5ZciefoyhSsFORAo8J4tBtPTsbLYzARgsnutSYU11RvmmaPd9tJb23QSXwa4gMp3AlK
8R7nPMDo2E7mYK4FGGXDMnKWTFh/ThVclbVrdv6IhP11NsO77yuiBNwLWW5YWUdL7Gs/9HwbFXJw
yd5gCIWOZp2yEFX7OvzCc248Dh6TcWYfmsQXlJ8crTHmkCDyr2yUP+LY9y3jnGTbgwfCwAF3MtXH
1nfwHY1D9LP2Xrvv+Gd6XE76XhUQUcO62HzXrPOHrNKL9ChH+xM+O1+zsYNdLDxYl9FSZuiU4kMv
+d3tM/60fTHOaBNG8G/c/6IDEXeOvDMWIh3R7vgPoq+eunAsiBUUqCucJ79Xvq7lL2hPJro4sAHi
xLi57yD7s+pG6L5h/9IBVAbaYsExnVAPGUFtoEkWmgKFLTKBORPKmRc6jlsjUWpfMG8D8y8lbWuX
MWfshx18QRmqV+iznnqzn0T/xQlGfP9GmMMxBrAEyUpfvWPIrilLRBzw3Bq+fWQoKPF4KqmdTJqC
VuF+8xSzIESEzzcpmTag9MGJCxJDaFvBHjznls/2/3Akl9vq0LYiO5V5VpaDIW9BcihBT93FJGIG
EqD5LH/5rWNcTXB+SlmqYRiRz4IiQS94JT8FAVxPIdlCCH8XDN6n0DrmrkAWJ6B4dvI6Cyqmejwa
0l8ALfrkiG9FGbsJr9r36V6h3kSSxiJmPCqGwNrY0sailli76/UELmqZHiKsk67yDujfgdoIuYxZ
KH99AiEwLIFlvDVZSup1T3lOIpfWOABeGSdjR/1WlC5VOnhUOPFzkJIF18bCCgaIGrAD1ZJz07bQ
QgbgsSGtdQlGFQeLoRiqSa9zx5LVKbV45cZp2fdgLp7HjLcutioo22G2PZMg76OtAXUfynnc+nrs
AxNZnbg8WylxF61fkWNM1w1q887Lgid/M9Pm/FY+f9FM+gZfvTIWqfyiXYXm/LLCWVsNKxp0dF23
BFDQxCQ6KTISEtoj9z7aO982ybkNNytBvU73c7gqnUAbOHuqi7uXpCZxeevZxysJ/YLAjek/ftTz
RIIGW/H7AIuMkSiV7bhTIwGZ+GcP22HY9JGI66fT28CEXCYrPJQd3I26c9Xi6zf6aNYf7686AXkC
y+2zeUhwyc9p1snqlN7z3KEJsgjzj+mubvaja5ptor57fC8WnPCOHjUqAguCZUyfJlWEH3QjC6MI
Si8uTdiE9qZivRZ8Pg2BSNksICFYHAFxHQb2vpyd4Z2ucY7vkp1c4AseGp8pU/glF+oex6ewqujI
GtRNt0PijhKrI+bBw+nZEm/eB++gycG5IqI+308wNv9yjlKaOex1IkbhT4a2zw6UkOtl2FV1BN0f
7vl5u7A4cLdv71stkQIENI5+X1v0DvzX2mjspHEoDIZ7aAZCIlUPlI3z7R47+wTGGkKtvNwUuMkP
jPOn7aCaPPVF7v5VObJsZVjkzKk+uY2rZAr6wp7P9qiNF69TOSGq2blWG8nnRoX+ID8U+0g5GArp
w5oeDZBRuXnTkkaTGwPbABJGtbX+ZY6CD1R4UQBO2cGYdpGu3N7B4QS1jlMtINvAaeHVbO/j2cXW
MMPs4Grfg2NkjpVixCYGj7nCFzOV82MCj9w/tmwqRvfGZPGIl4bAeBvNA5OYiFDw37wSlnxc66RV
1l6JKnuqmLY9YsMDrfsYlH709Xo+kYWA/Bgu1SzKZ8XsJssQwiT4y1wKOgKKn7pcPbhIe3R7igW5
EZFSe7Z2N8nuTYN1ExtdR7ra8DVryAeF7dbgL9lqOpHxuX6rKpNJNx+9J2WEslXsOuSDzzgwZC3w
bQWDEjq+DkIkLGGhRaKUcYhasFcaOIDXhQeLNt/G+Owx7LdE1S5Cb6g/FqkLF9zEFLpdHfzZKiCw
9LNKBrSceMOTFqkyR+T2lwGeO4cYoHRjibXY3fdRPeejUy+LdQzQnpP5v88hHi1a63B+Z5Nt8zDX
xBIxFGlUlYIRs7YslHAZcPmuu7byHsles3EixYweVfsoh4STgRe9ehp9g3wyl19Am385wDcWBCnP
a5QavjMFqhMuNqU+kqPsWTsxyJTAChT6+lj48kxcMqjZEnG1v07ihsr5P2lcQAJgzgYv0zbyb/Ar
SSAGySA1fiZGXQfYLCfMdzVf+3S1OTuxtt9PBiWP/8kZ9Z/tUYcRPd1Z8IN9YEa4lgKEeruCJV6a
sYtkeJSzPtHo3sE5wGRnwee/FUMQDINsTYVz63nAClTbxZdu2ad726a8eWDJnFn8PT6dPBkxGMEZ
44TpniI3PK6mjmNmJnyFYuoatkX3ciD7t0v1NEKSr13cabn/Toy6cQRhuyOuCe3F7i4Mi1awrU1L
3nx4NCZRoT/kl8M8AL7hRDk6C5cLgSRRPsRe/E8rQBbSnTH5LOKesQsxQ9Fzulsei1+1WopuxuwB
+3OeT9owcxe94cb5E0g6oDppM+gduZGZttRsKVgXFuiozX/uC50ETb7CKuhCTPF8AZ9l9rxg/7v4
+/NwBPmlaS+a8K6p7lWsebNy1P1gW3hE6cPitFddipC2uwseKrW9rqcLuTf9FBEgz0J1j8o6MpPT
b/tGBY9mo6UiW6h9h4XADrIc0y7uyvi9wDCbnGv1BG/3+/3fvVF5jtWArwSTwiC2JWZNoPMJSc4l
R+QORJmwceT30WCslt+unEaIuF9d8XxKzsFuBMZ41B2c6sKZ1oWJNsVsuGc4yuLYw51iPee9edqb
L460plbabJXmW05vcAtkqFOEaZ0/ryjE/9QcUxU39SYdiJjZkOyhtFRCkUY8xM31rzZHPqiV5DU7
9oO/aQCG7lrjC3BTojyLWFEEd+1lcePEcV6hnKo8+wG6M7IRpthDpc1nM9rlxk8sGQLl3mmZoKek
uTy/t9GtjrD6s2WlGLFJb+AagOz6/R6bfnoxAOGOueEbmttTz74EbZXnSAHTO29Tc3XgAhTNRe58
gfC7lhXF5l0n1PjKN+TzXwLUs1sqlD3ku8Vqi8WpK6OcXryJ6761PlC+hxTw6BwDhJC+w2jejbpl
SDsQORZSe/l/QZ73w9Db/8dXrK8+koV/gsBWO2RsU6ZBIBJUITaOxcA1HD8/CiErAvsy2+EKlli6
ggFHF7WFeZw6BUPi1G6Dew2KsUZui9FvlMJxchD6BBeX6gZb9BTkuhk+PQFIiuxMBA1t9iVEstPi
mEYmvJmsSu71cxIS2YfZDlxOpROCobjczlYHE9OwbHaKBNkJcVbIGbCF0WkHl7PLSlzP/iKeopm6
3jab9hp5DSpf14Nqy7oRsB6v1zY8GVKXHLOAdMHSqe2DtLbNueL+Y9qLU94xCsSBNu3tgXKtdcZa
EuPO+I8yoaAtsiF5JC/6q++F+leObSpl3Mf5ePwFTd/58X7f12B2YAuPG3HFRNhZH691rtscYNpN
lfGnrP0jxQ1yaccFOI6XpFWBa5D7rxEHGPgBcjRqsk65o7Nk5q1E1dcyiYOIVFt9sZ3ytITVPgqB
S2CLN0/Uzjta4PQvIetSsGN9TftFhtcGflAqT+AgFTjsMR/xBHkFelSPBYQMyfDxVSGyOmsPA+Wu
xj984jop0KlbCtsrtuvlBQ8rzr4L05luRHytnmjdvSem0Nrc+TdV/VH9gjUdQZnEATKonUPLScsK
nKK26uzITqAubLIIgZx/rWaMxpXKYaFbjHipOqk0i6Yr0EIOQbJ6yLyON1r3K4sHdu7jQ0GzFdo+
FB7idnjowa5nMCZwwU6HhgPHGQgplAFZlJGp/3xyOTp1b/1j2G5iV0AuBRPLA4LPzy+ZQLYu/n+J
3AFU5LK6vzRobQH4s1gof/paGdMNvCdeXeqvbS8yIQKizB/0LE383wGVz6maN0WJebiiZuwSEOlc
IQXQ+UYgrMano1njtLRaLGBmOdyljOgE2lk5YVf0Puz7I+KvTasrqK1TJnmZayKHqf+R9zT3Pea5
xXyu19MgmH6YX/WWAPH0gdHx8BnDKA3ZOXAWmj69m5/lmVivS93G5bXKQnke3GltHVhobb0L1+dF
KDVPLgmNAxpi+EGBRrHLVoQEIYwphgTdleLwl+PPaY+T1vn1aLlGWBMfRkZekwVpEa9Y8opTC6nO
P8xF6IURbOY+Wt1qhMb01R5MedJxEk9+whtVd6UjJRkWHMXIfBjbQ6cWVS6KM3EpjkqCksFc01Wg
IYj080Gz+xLpB0ctKsuq7XISbaw1A7JOGrtM0nyXiixBnzidL+Wuk3HpyYUviyLWNo+9gDRqN/FO
Xl99qtA8ApZ11Mep4KJFEpzYxNXXqjCTJkoiNCconW32xEdh1shzLN/KbZz4KaoAsiejrm2fzUyR
5fmrTe/EkibjoMbW8v1ot9+0V+wQAQKzHzHtCZ/qTlRsUy3CF6qpeCOq/9qvPPHmw7RychNxK4T8
ZAuFP7JlJn2DgGuP7vKQekmEggUUcUWIMERqBk6G3PGIMelJS2vaxnhoCt7hWtwfIHHKVNxOFsP4
7c6sVeZ9Bpc6zLu/kFnh836/t/EuubG6Vub1Jf8gTYh7FDKUx393BhSv9lgeTwv0r4hYV6XJ1ZiB
f44JzEHQHA9EEF6ujaYwt0lLiwqOEMraNRgN05yxfjeFIiuDaY5Zka67PYZ+4PIRj5VF/nam1Gzo
W1ee8Pyg7oPqpN0eNKKe0wGZQfDXs4cRt3AZt+Ol/HAHlh/kjcCnOSZDepgdSnSSo1voyxMwUeqC
zA4d7qkRWX/YAUtGyHvvCkae/25Je8eGy1tS8W587UMlclvpXixwKZbzDCi7MVdKeajID++G2sUG
heiWil/Da0XwYJv9CiXVO1p6ssv3lkZ1mk/8/cHd7VvMJqRy5CBsi3nUXNJC/r/Fhlw/tD2Jr0QA
1z30yIq7RaLTYSdK+an37EC5wQkqLUrHgZfGeLSfzZAVGeeG4ppFWe6N5KVrza+TOuApWgEPbZyq
YioLKPXUP+lu7kTJBz+q/BED/N2GrqarcuTAipIY2d5fIL35e4CqiEajjS/RNFVrDtPcA76LSvLV
FnHX+sClAdJNgx//z6wwCO/ln7yjNFzQk2LZVMfPPtdqatJgHtUVXbYnwIQRc9bRxiMd/LjBAEDx
y6JGVQio5jSctbAY+DuCLMi8HM64IphO3jiC1ogiB90ISD2xI31peOeu/9tPT2EzEBexh9RBCLoU
43Tl3KxuinPhTWVZnU2tscsbamXOAL7HS18lOoZKFeifcoFuJN0bKIVLAosLtadQqksrvl3eHvP4
fee8Xu3F+EjbflWCXb64kStmivwRy+CT4OgUpX1n8c+ZsffZA/lP2mpGgNYsKq8dsciq4qMFL0Wk
pcNuHhesU8+CXl0HvhbmuMlguyq7G6L1Z33ihYyV+EmLLPIBU0K4v8vhXWlJ2mP9HecvYPcr547O
ltJybbj/dWRco+DR8/alqCehwhTP0Gv3mQRWBr2kqp278hhX4dNCCkowxJNNMjZKhQqLFE6CqQEJ
TGLYymM6Bn9oTrez8GH1kOpe+w+DlDzNbumCaW4he9BaX0PGmauk48J9oGFFnRCyGn4I9fMo9v1Y
n+Edl7CaMHL93yWjgk6ZHeWm5IhXchHKA176lwudrZr3p50Zki5wVe6szQc7s/CIpKvu6LeypNGe
E9JwPL1aXYEzR7VXkbuyBITLZQppzbAw3UMP/QRH2sem7rpZGUAdTRAcbbA+akGr6CWD12VqcmW/
vubJcIOQL5wIwppYosu8H/n2TpKGstXWuAFZidd0DRd6uMZlBL6s/p98JcxB9BYJfvCrH68KI0jf
oRKfD9b8SzpSRS8digDY+bH9ON2lUJFxVvthfwlH4eXt3h45inbw5B7QRTbJvQzyMtzvyIgeqbaT
ePEokbPqRNoYnXybZQBwGGQb7d+N1cknmKn07lGkoQqW691BjeyhuWsA5Na+YwUHRHPx6Uhjmpgl
MoxOpSdUWP508HUoBYdvrDEPbPgj7CCdhz7E/O2xzj7pfshU9oicmaRQHI9KyKd0ffjd6DwcQu3v
GnTV4PRAodFLlYEDX72rvF73f4HHyOZEaThzcvvx9ds6i9VcjmWs4hBBmhe2ajHlw3par0ZfQv2V
gQHpdxENvHgp//I8xcTjD88hzGVfPHgWGicU9Zfu6OtExCSSU23Uhh7tIq0ixvhKc6+g63vBxS7p
ME/fYNZ9aoMHH9bgXR4pUoF0BEH7tmLDoy35n+GT2jdXzoB6jXPBqo7Mn1Skd/i1LqwHft7BOAMn
LQSMOmuBlbSDd9BpcKTL/Gh6yr+C5GMV99cLTw7y9K3mYSag9uMgbwxe7i27QN8cfqwf3ONmNr/j
KYQb2ge1Sc+STl0nZD9zpaOYDjeY7IkP/NC/fRWFb3hu9yW9cy5uTSyLScQLjT2PwCBDlURgXHeS
CyvWfvYjAw4uWhxjxL0qxgotH0XrNe4T9x/hpQb/n9DPe9GRxXPyJxs14WozEVIZaIoAjwgKjjBP
WqGtcIOEuCepbiYpLWhFul16qoZuj3k+a/nZZXxQIzrRqsXYpOgT8S0cUdOiKlKwuAGa99+VLW0k
Z3EMXEcw0RpEH5xGHntXMNY5qfxtkdzh9qGHFejyK5MgeyPUZxiBSKEhphG7I/6U9Pf0sUdZPRb8
XmiWzmC+iyfXaZZa5VBsMQF/E/kdi2vDKJB09wc3E9Mt2Vbltfy8gvdMItDmjqI8os5ZY5NYEzkI
zl7nZ/SoDQgFIxWCPyB0IX8RXbxkngR6jRGvF8FeS55XjznEge9wSJqKLKOmcP9zf3SF5X8aAGLn
XhbIE9hlWir3/bFj1USnNTU1uQpkyEuMPQfZvKCFSlUNPBSsf5T5JX5dopg63fqIcJEmNYfryXIN
gW1uIUGjTULvdVffsFMJge+T56j2TSRubbcRS5iJnGPxdOQ1emV9Wki55SODEU/ZAdG0bgFtXMUz
+TXUyupANwgymcHohDojjv5tXfD5BkxJVGocgAybo6/rU7/ZhZ9ngM2rDc+REXGKppGI6wxBCvMr
fSTI8rlX3JwKWhCuxyeEUwHh30wX6aRjuJBMkj69j1elo/liXzLqtaa2HK9Ce23cJwCeHEhMjvKn
hf+ICY2oTMsdNwu3B/9PCvHy5CfM8PtmfybwvIEh1HY4Szbd+bz2JNR9TL4IdgciZ2U3yyVXFNe8
E998c9P1MZu0SRXnl7vU70WAJwrnlGTOOdY0PAH053ut40tg40CeobHrl+IQg2wca7JVrxos9T38
UpZIbfHMorJfNLaWmWslagKwov+whjGwBPt6Edm1MBUxrl/rZgf5euseEu0nvsRyaJ91RgbN9i7B
3IiaTi0iIG5slgBCsCIDd+9fwv0r8onBi7b1G32sK8/ZkWYU43hHJlpuZJedTmlkQNo4NkAwxL8j
xvc14cVEFGa5txs0Oq+YPARVASYZMHTPyU4xNzWy0W1G9h8EQNSqXgQU8ZZTUnBy6KJFpkOYEeJT
sh8ADwv52ZEgHf67BF0phFtNRxOgv67/MowrW1aY0S/kOxFyuGJMd3aFmXjHI62zNiUk+6JkZjOy
4lII09BjfNcOswhjwQl6OJNDK/1N1KI0xMM9vBP2pjt3Apce7AfNu+vmFkM5xGOqUewiDynqhxki
8vXIti47LST4aoe1qaq1vHE1xpEU3sQ58bYX1vaJWZac4zeK/c5Y5JqhyuwZjHAP//uVDsz+KXuQ
sjEHwqmLuqUSdK3u7xuw/gUdG58Q9vH3x+nwIX08m6oRMwHfDyglhp829CQZFjBxDRI7roH/oA3J
0mzPCsdzNBHgcgeuIuzDFdUmoM/PnbIAA/UYvIkbc9SejHXfZ0xHv1sKiSePsIy0bIRSoAm2RmW8
gVf2u6Sq2Ygb3u5vDDO68rss2w11Ax1KCKj2wVQ8Z9DqQ3u+JYQ2mYHfeyyjzYI7xyHbq1iVwoKr
0jl5hVmFFDl273NOL2psU/orTlIopCw+dgkV0ElEARYiW0SA1LMqAuVTZqK8RmVUIS6L56Ahh7eF
vT7OO5KoBpO2KPDd9LXKi79g3skxxOlSdclo6jQTCra4OC76cYGSXJ82thBhaoogIb6SPmMwnzS3
fGdShCywMo0tumYsYWwqagrl5CYcUHYo4ge3O5FnbbNlfaN/Z9lKVgo/k0Lyd1wwNiHOi02ceXH/
nqfZAZnU1LUVy5G0rTN4OKUVU/Bw/pXeO9uCvIMv1bpJMK6UIErDYvzP+5QzdK+blItiSV3FRVOI
NRezujv9VAashKAM36JVriIFy+6mJQU0gKCejEQU6ABdT75igfgGY6UxmYq4IRBZ5fLoDCZ5ZA83
HCVxgJKGulQ9MPi8BV9+RNVWzN8tVUS2in/ZZxTpXMq+aQfzz4VvWFsPjQTg8/ZmLpYZcUZSYqQ9
VHNyjgqQZ+xYR4nt7Maa9/7Xcoc56rzp8l46JNA9eE7Yg1Qcmz+ji/clofqmC9JvsYbsCqQ7zczD
5juFD7D9TMRtfPW91c01kx/U1oHs+sWTkAR7bXpesvaCu73y4NVc3pM57pw7Hlz58SU8wcRlkF/l
vdrBBkLknkd4y06rEWKw4f3IEuKK+0NskW9BWYW+3FuOfzxQw1BStuZzkHM9unaFo0G97chu0gmF
JxasJEzFKAR0/bQVt9GBAekvpU9ghKRPv2v3d1Mh0VNw0knkJeN96AwED+J55xUVs49Ynq8PCTax
EV0UU50gG8It4/qFfHQCgEeaMLh0RJRfX7+Mv8VZ4vtRjtMkEEFBoJYrDL9s7+gzxZZxScghFyI9
HGvBjghDTOlMIFS5iylij+Lj1pyTvSI+vCoT+dcXjYNzh4yO+JZNJxUzaUKiD+lwjo8MpEPFm73O
UPvJ9wQ9QipMgFotaukqJy2XNeTaK+ilZG2BzmJW9RAk5a1e6iPGoyJtAfHHMUwOBh0IAqx7EucH
WTeLaKCFI6bL/ivuFVnplkmMem3Jxgp9xLyDzk4eYMKEXrb7oz4LAqX3L7T+UVwki/PkugBBP+nD
XjojAw0KeGDzG4IVygNfvg5JbcqgCWYrQw5KmqKK3qiV9Imxzm4e3fU92eyeiYY0jqL4pOlSVDCK
BaZjd+tT0RWPqE5NK+NkeWUYEvI6ymTkIcVf2lJ3nwCtXHn7KpbBhxSlLdSDYWCiSxT984fcSO7M
c8YjTPU4rQLNKHkijcLrBI09HmKippPV095fUxvtTzqSdluJsi45CqvpDRcEeEpXSIWxEZANyLng
rr/5R25Yz2dNFN/8I28QyF9gXNsfgjbXri1yqbOdNfOalKQLgum7MTwuj4y7uKmd/QzLHTuGqg7V
xJpoo6c67IbdqIp0JDRIG2gHpygRPanacDa1ppT9ONpzWUnZPa3xHqmRHBdUF2a2qTV1PnsaYkO7
m2Dt+SlIOum9+1jLCMMmtMZgtKW2GzvbPQuOGui+W8eZw3yB/EgagYDeBt9U0UlGvlvA0WP3pQEY
GCNyiamGEQfs+MNp99Bfq87M7QSp0cSPCmc1qpihEDbo2rxewg9AjEpIcLo4CiMbhONsabxxeaj4
cv7D+SKxHnU3UOckCFTcL228YZfQ9rAJrnYbLu8CZEddxIzbe2c56Om2M3tZ+t6HSFyvIy6rPEpq
VQYPDfvQc6FL7HURUL+4GF7J+zJJvfBFtvYabclUdWrhyzjAtHnDluqd0nJTOQyoH2rpcp8rtfRl
oqiwFm1Yuvt1kA6bg2/5MdFV6Rv+Ey4EWhpf9sVUUTQAkukOjRunkobuK7SdXS5u/KWTmmP8QcqM
QStG45bhbZ8eCivCtEXDRpfxUn3KhOPNkwMHsA3zhT9TWYm66lPzxwEDsl+T1ZljWOUmqlKtd3bp
C30l5IzP2PbAE+EcUBlLhYp8giIMNit94k4YkIWuB8uiLZsD+/RCdSQ8W7AUIZtdJkcx6KTf+Rc0
/06WpCqM6n1iVWsd8Z8tieBMTKgKXX+OI7te/c/LJX/VTBe8V50VyHZwSTyOfmvQrKmrCMq/tCsZ
DdBvi/UyEMd31psSs08K0LlCeZ6TBs9Y1dUBuiIrGaojWPRnKAVw3SaOB0/CdLmXVixOnUaCyFvN
f0J6oN8mv3BCawP5HNhHDRLuJuwNLAPhv0pDyRqo3OVhbSLCknHFluMV23ot+hXtcrMP8JFxOWgL
d7li3Pvsta0VGvPkvIgY4Aw/cIEhvSp07cIHQPJfdmSuLfYskbNtI0wNLNN+0xAKBUyQGg1JO3CS
XWZRhxUEDN9ZWOywgaZYN6w01RBdMgb6vvdDhkXA36oJRVfu5GetMViFYQDHnfg2lyI4EMIe6HHI
j7sH+jOT6Jb3qouIft9rGuczKmS+QQgAUmqBa0kLF9Bbfp6SJ1r5CEXorHfRPUAFDi3zQQaNgehJ
olxCqB05cPyMb++/EK9a7KiKl+EixuGmWGvbR7K4c3wRPRhNQYJ8i6a1ZsKDVCfxtZncHCdeA5BT
MHEVMAjAGCJ9VYihinioGH2rwPCCT2RriY4oNvwfQoKPIk4kiSgUPNqKKA25i/jqba3C+yAG895m
iFqMXylOIgIVlNLL0kFptvdcAdhNcfJJ/ct/Nubz4GtiVbtUwO4Rnux9r8wm/9EEMrIyRGaiSacp
OGkXW0mS/Zk5hMZp+OnHseBcvRg40pPT8dVKJEG1lqolm8Do55J658RyFxihAx4rn4kCYpiX6paW
9gC1IwWzwb3w+7tr+uVD/e0RJPTyrmbJbhW5VxmUDUI5VywgXJ0JQNjB4hzuxGeLL2oQ4bsdLPZ6
IBLNRgwNf225jqJffoC2ySq8e0367M2kgcLXh8eRvAClAHqSJs55X50W5PnTdwzaeVSFFeLYyskl
ywKgDpb/mTC4QOErTQMJwibfoK9U8a6WRpjvwF5CxcvTxeEf6I7wB/QoqLMflvxkI2Y8bw7KFG5G
LF9uDmd9nGU5XoE0SQK/xJOIJlzdscJ3he8K5FdARUWliBeG/fm+UsRHeTBC3hzcDxuNaz4ZKBxP
MnXHmdYeFFPP/xWSkHuK3jVdAQMui85z90ugRSP1ZlmGNPUzXcfoEoOz6mJzGXU/alzrFdR2GWIl
3/B8X7GU3/o1XbNLybjxJ794qWU1d+JD5qN20ne0dBzbjOTMvVKleKsRJeuIiFVvFK9QUgZExQha
9KEb58oMAxigf61VRGq4Ha25haLhhqw27aJSGzB4RofwDak5PS9R6VqaIGyah1rrJJ2Xaojy0E1p
jCXfVecfARrysGyAgjlvPYFM/iWp2SJGHqiVTk2Ip0IViOHlKhiDz1u7JYOijtrx9RQEkDf7yD2l
1HjfLx0IH1x7n8Q+1ILuDitaFLcOrVw64vV2iMmuLwxima3L5Xh8DDkUSHQIq0FJ84U9w7Bo8VnY
HrrXuf1APH3KEse6hYOyYJZYHYpnnfJYlSj2C0SPTDY3UqV3AZpqUGpslsJ7GEZtbhSVf4q71IuD
a9DKTfzPW0C7jHXYBxzM4wj1l9sn2/GxoiR1B9HIqxUvmCkdabVyKJQUMwQ7faGAgQSnRcwmiEYf
mw6t+ysiH9jEpk7h1iyWd6SvM+6B2JJSk9hPJECDInEnvUIKlOJBpIhkHH9c+OJLl8KB/JTwF0QD
Mu/jSWpNEDUItWTkh4KLyzThDHQMgeR9vDOyohMVy8kHIlZpjGlYz7p5oPSNULX08oG4Xdq3nMud
3dSppPAtaVEtK8UOh730IaGKgZej5eWhWr0Fzdk6f3/KmJRizdqPaMcHdHwmzjWmudfKXsK5IH6V
ttc3bFdrRjh0rKj5l2M7rUT+1w60PHj+IGK9jjE+AsBNaGBjUL1ZmmDIV1kUUhPRaQccVEicJqOI
e2qKWgsTwHxC2KvF4G1iIC3QL0s6K/HaKjUfOSkgv+GMonxsUrdLa35RJWfsNyL4YFJvrDR37pWd
OZpaDzETjSvjMEU1++g6QL//2eka/RSTD9YzOwomcG+cc5/IvYZ+s3F7dhXx0ODUrMs0rHWjXM7v
LchdDfkA//lAS/TNYMXir3gsUNR6PFP5aB3cUEfuf+iWsJuLrGvdxQOxdmk31Goo7YDWz9io80el
P7GN78td2GwT9v9pqhpI8LGi0MZ7rEDmrIDN8oeQHum54VARzFbK5ZicCRsfOXqVcYiliLxv7LuL
OoMAsEereB/rku/0HCja9F8uykxvZGmx3ew18aD3/GqLq1YmV5XOB+JGU3E7prwYKYP9PN4hOxkD
8j0mjyjpRJ/LV6FTP4kjnBFEE0uE6uYJ4gRPW2XDHl/gqxpxjFykklYkK+ry5HZyZWLKEBGqRqRR
PIIB+on56CKxKWIaTeOcJEaEPAy0tFFdDzCTbS8vYKV5NIkSZzTB+jing6NX1GjFvDm48ZEeqXmE
1uy4KaNfC+ZqOZLjBl9S6BHdz/JjoyLlcnY+e4JN8cAMupblKfKlN/fgNkGTL/QTWMLgaGHTspzI
EpyKiyeuaieDzNwIKU5Qb6KoOTvWw5JcfWoJI3EaVRA5yui9pZsgzDmjM5gvqv49SH8GHKPN3wq4
dVI22peh790IEhYlD08J4a9CLiDxyR4DJfSgs67tNVTLM1JrWVjpeCO/y2LKyjWTtjL1rwUFi3rX
t5+DGxKZPjfS/kfcFg+46fB2ZjsOsCYOrOwf03BF80skgCgNJFDZOANCmV7C9ogCV1p/k00mS862
f6zpYcxOxHDPZPJfjn6hanDaXrgl+10/NjMYPrEEgxO4rhOlMP1DtOr4qltAupIP+ppjErzSjl7S
NJQnnYq8WOMdDDypYNgBU5OxXUN0UDMOKmKGfXIHYUGLaKyEmz/2OQJte0O3WAlxPvsY1gegpQJa
BqAFQOefzCIzz2MrfJL1JQ4rZpO1HzXSUv4nnwlT39QSEsacPBaPk9EmuQQmVGvlJbhTRLPdmeWM
nmE6r9fVvizw1vlkm3EQZZkf5w6B8HyVjXeUW9rrTOgjAjxnUxzX1/0EoPu1R9QUebKA5brwxTRl
CkTumIEMVoZnTPd0ITW681DAgh0jROwQEvrZqjuymCroYzoY3ZrkO/jkY3gXQy568rvxaYxABshh
skg+4Mjy+xXyP12mgVBRdvSLhcPYt27MWzDnoilgiX/YtAWwHT2s05XzpVAYprdKaxJ5sRyi/ZUh
4pXbLzuqbS4+TTkKup6MO4jmx09QOt6h5ZgrgVSOE2iOE2ztBsaDGxEOX19YjQ2WTUBCbCkl+gtD
BcuEFeX13t+Pg8YuODaIMrJ7JmErdHD4CcWJHGXJmCo8Xpp5wO4gnHSxVESxDSc2T5rrdFH3/j+d
+IEXnzdw47negRCXzNFqBU2O66cTNl8q9eBzLADTiJkChU4n5+zR4kL6IppFXZvVQNIntI9AkHlL
5lA/CCOMnfC7YlV9GUP9lEmQV3f6gqx8WW9oHWGGy/S+FJQC3MaIgKXkuO1qcpz/u20TI5iVtM1w
FOleObcSiIt16X5tS9iwbfE17kok3cyuam80gfJi0Ks9zsBuftrP6Hkxn0AJa5sdj5GbIGMjmt6G
2PJxjse8hWJn4L8KscSOW9Vesy2f7Br3gGHwIaonh0LEL0frqLvTWF0zK14xg+HdU+xDXQ9qAdnP
BPgi9L+we/9kca+b42vemtzRFVLUirvcBUDSghFn5lxZdwpMXpZoC+A44nG0s8uqdbb96dcFhYdz
Yw7s5Q3MKlTt8MoSF2gh8P7RblCyalbSgby1wXFviIdZ0MgFsWl1UcSlchZCeU+j1EHst4vlaxc3
0vVGhl/P7+Ojc7IYpWh/JZErrpp0NbRsbJZAO4Ut1PSIsOIhG9QyZUMCWR1pbNonBL5KmDOfKiic
tH8hoQchSY+OB1ahXocdak0abOOIZCotldaYM07UK/WuoEiGzpKjZysFOwtsYBRaYt204HLWuVD3
GZgQXpkIogUQlLw7Qo5xhsHV+OyLthmcxnlNuUpKvwcx7of2BWxT33Yv+WRdkQSaN6813BWo0AKv
2PND/RrxHKpXBPNH0KrkoThR60JOsoYLA4vqeA+Sz7CX7tTDz9ivKXy+6zKaNUR10dxilk6kGXqp
iONF9bsMJHKRampBi4mSEyTK2+7qvpN6j/TChPhNUg7g7Jaxe4hSNBqDNmEqZzGoX7vtyXMo4yCE
jc+uYjZFti9qg1OLCe+CgbVxthKE16XZS/QGaVrFrI/cmwEvXmk7IByfG7JzJB87Zl0y5CjHXrxF
cjT5QiInUIugkJPZlcqcowXbruwpl26Z4q9kCLu8NiDquJYFJlr92T3uR8sdlz4Q/ypj5lVYW69W
0AX8wHXelzplNpS0a4a9VTkHEH7/u6K+7R7hEsjh5MooK/JfMtnE4lHwTdSknpjCDEejOGy2SQEJ
H0dISp0LbW03pwIgOjF0yJkQU3JqX/CThJlfISjXQJb3BfxBFlFZcPDTNVSPa9WGn9DBluW38txd
Klxig2lJhBfladPejN6j/9nPa0M0lJgEsWJy02Z7EmLseFmUNX2Dqa5VVHjsyxT+zGzFMFkLWoLr
D0gZ+H049GXzFsIY+XX1GHFib5/TFjPuCJn/H+XjqtqdH1Sf40WIdYomuHhwLGi30XKb5qlb6BwN
1DORXIeOX9oN4qbG8M+jk6K/y8J3eAtAjBUHCbsXpRoNOgF/3jIKxbV0b8QSLXX/ys+9K6V9/oZf
GNxA8BMT3VOYLi0DG503uZSapzFyHA58DSy7E/WTiQsmm0RsP3O842Pw/bMdZ/mOMO+pwoedqgVh
jUvAtRvsRsYDB14sbe3NiGLc81zjUccqHIeocXYbx4Gd4NCkMMosCF9pGDcX3PgdEqsVs/PdOxOg
mXZqFE4pPcRewYsFeNSASwxC0GGvh7CYL8aLP4V+C+142s1qy+yAD1/d3OMKFg9w9OwbnAR5wAah
bBTXxNy/vcLpvzK7+pQnt97lA8sbbvcrLej+BphNz/ZePG5WQu6dFBmr6kic1udlvhTP6uGWSjbL
B2FpvCXAOBIQz7EXJIJg4PkSnUt614hlPXZ7f/iZXVypXS6LR/NI1F7Dk+Y+nBtTfJOb9rHJ4HEu
ZmNhaub+V0iH0g5+izxRfXJcACtmQ0prElB7woy0vZrSF7jOECZfAc7AZSaWLRBhCJGJMGUat817
LYtWAhnWFzD3fwiB2LzRP6OBLeI3CHF4xwD8rsMc8A8XpKz1F+J9Ohg8/16FwgQt3IBiioEnoG39
+2i4wcioF+tVM/Es2TqyEsbnBkfVQoBKirTJyNcTYnd/+WD+T34DRN88ZlD4TRIooqWSx+aCRq3w
YcbUMSsULZSwL6Ulnf4WdsMOjVkJcICF+Vo0wphMsNYFd2SMhtbcppQYAu26A4qHdXcAPUDN4nHT
NZZrfw0jqvmaHRQ9kOkBQUvM+ZbB+j4KZP5k2VjOhUr0+kQq70cxk+2tJgmceJPrh+8QQNJPIaVR
jR+w2FCuhfvNO1SmeSPRc2oWaMZFo8xpWkzeDpJxQoG1rY/kzEawr7t8BsdbGxRycp7uegqzXNYa
R7pixFb+2L5XDiixiEvJCZOGS0a7gpHyNgjVDlg4W/I+++YgN9Y/Y1GkdUGt7tKtGiuMG6sIQkk7
rTdUZx4RRncDTbwTxMRdS2Le4dedfWxHwjGQXJ4SBHP6sRQEd15n8Ks3uzLU8w9chS/wuP8gpder
Lw756DhHSOWznEyu+CGxBSxBM5DWoFUJu6Tdo1PIHEKl1Fv82DWCPnM9nrhobt86IGEco0kxdc0S
a+FR0/+0Q9//TnKcMwtIywslwpX4fYKCDwPiZFJPJgQmz6Z7Y6PBLqnJlAp8IfaIJ4pQLtK3n47H
VzGrXFpHm5yVT6tkFCtrjh2GLdsth5AxsXZf8WfVyh+1ZxZuAl8q1793ES94vHrz6t1GnI5VPlYe
gqclzftSRGyGVYh2fyZ0OJDUsHnZLXtBUa5VL3H9aoPPw4YqX2YYo18MBSjIoir4Pt6eslIm1Uxb
LQjHBcq6qPmF2RXlgkpFytxbNuPxpsrhp1wfUjDIkOHKcxes6ybSxSlKbDcS8vxh47slefTcwylZ
uLuw8oUBScagL4HR7CqWOw1eL1V5a1Q5kz5NkBOnhmCeBFqluRPXlpXVkv+T4FhekdK8xQJOFk19
apWvn2NH1pUgvKDgWGmn9Ko8ysrR+hIL4XCtp8O9fe0G3diGu/0JGV5jhOLTtlbjCzWyS0T0WbMy
rF1h+e6pFzCaksdebzkOARzr7I2vIiMSpPTLnsAxCbHJagCdxnxifI3IaR+fVw//ah+RuKkpyv7l
/9Jd5QI6W1zoNUflsPQlBo71RCDMnIILrsb5xM3D1c0UF8qXAead7FLswozCarZMe6MqeCPs5sAV
fHpuViuDbOqfH43mMHK03Slgnia5Mfj6FgxkP7FAf9dvU4PJAO23z8EFcJEEdz7DQjS6Yxw0HaYP
UFN2B3Frc1f2gstGIep6rQZcDRorho+Ck1mwG1D40D/IqSrJRx9OjEZjx2uFrKRdQv/1pXcLHLwG
XDOdgE4kVmv1alWIdNAf0U5HF+8ns6aMlgTIrHsJqFSmJ3cT1wX4qOn6jb1FS6s9cWVtZmJlUmNR
PgdK/Kk0Ibm4/FbZg7ENyPtN6JRJuUVtzn6W3smkhPV4nglq4fESQmDi1esUNFUHZtcLKxfseoGD
ghHGp5RHWkUYVoWqnPnAjZlHecJngpnJkVYjGkNStoxNxSkvV0KizUqDMbMZk9aHKdNAPVVQtAuk
HMh9Ly1a+GZkL6IW2aVpY5+LSx5HxRqW6hEyF98LKHNcot4iqjV7YQ/2PYn43CSyAz1W9I6mHiJR
WCl9L7UxlAwjLjfx2NHLu7NZqsymGQ7gCdr6a0u3zkPXSyyPCpYNIwaPXFrzJ53f1lFLuTKdxUSm
kIfJIlsNDd/Ve4C1X6n+Hl9/JT9GvtEhjm6Y9IkiQ+OGV+op01Q3gCYHeIUCKk3UL3ETk8KZGAFf
VosWz8VQpDlZANeGcLQJajhGhsdRVPpf70I1Ho3QF9UJLiViQOjnSkFKgK392ZRhzlhO1E/hC2G9
WmSsLkPmszBNtQEfVFMcj3ENozxJ7ymwCZ6UQKOgCmJOpmpg9CtnttPFu8ux3f2O0SE27Nee077i
WGeLORD8H91dDluwO/ekPyw4WHNDwL1ZMGHtP2lei/kNQqJMW1aXVmKgzG+hNgyk//DBwhdkF/FA
mz1Sw6rdT3e9F/XtUkFJ2Wg5pisZd0dB+XgwwiDpfW3Qy/co5Vt4nnFT9Yq/2SnutmvSl3gsRfRS
OacGqgx4j/5+X7h4DTgqcDIoomruxD8d3ZaqSAXgBbvOS+yI6fnc1dJngGyNU7Bn6iqCsWaV3Qza
vzGwpIvXC18EYF3Fsc8p/rg2LmhiJS8EsqUkdeqSwvRzLx6gbVEQ+4oaTGq2uUT9scrMOuJV8n4T
MlO6PiSVxoJkMdy4zsJUitOMB8PKTaZE/XwKoBWKJapqaM7eMKqsrAifYXLVdXbBHxYI9LvLABUU
JicGxmm1F/EzIuHr7kXlCDfQPAJPGpzfoJM2hhBxPOFSRR43qe8QN4LwNE/1q9/kxnsCyuPw9OWY
7+XMWsXSSUje+I8wuriamaf+rxs+hZwyRazK3EkSeRAwLIjteCmfFgoJX5+FOSs8F1ewpX1mgTsq
eaBB6Dhv/GPbFQbPfXxYVnf4E8hm5gJiY57DUVd6hUYiV6NqUtZE0ZCwUFe52qozW5qFXV3oEIxY
E0Ir9/BD9Iu1XqQExtoJo0TztjMb7rsAQHLkdkyW8g/8+RxKyCXWeLd8pYXZnYnvj9KzcjFm9Puv
JnRAvPPG84kl6ruH3y/qt9cr0de720clM9c3W7RmUuWg6gWSoan871Vpun5DjPSQFoI7J8o/1Tbj
1+w12hVLLgNj2y9as3JQ5ZcnVCRxCxmiigtZUKk72NIQuRQvFQXvvUG/8y5B1BUoPS8ONo2u+4TG
WOfOeINTSXeMUMvEZP0Ns/JsLC0o82WZsQvFwW2Qgy+xaFnY/2Xthss4kTNkKwYluFKadT2UdvPp
UkzCAcgXh9QmMAbM/zlw6jbLFizCjRW8AgvRfpRowZdXydolGXhhpiv/MC34nSFk+GD0RazfIJzs
coQCVmmyzja5JD0Hvdv6Q7ye/0Tdt0V+Pev9vxTVpw+MW3Opygnm+P4JCkp4qpNuNp34RpSiz/P0
KUR0acyd0YBpDnj/rq6+WzJvm0RaG0edjLe9EXSRXdsbmk8kaBSrvZYgKGQeMZ8dFMcHk40vWkLq
1M809vqwPtySmjZwN0d0q9E1bXKgf683ejuxl/8hKIRhH8gBPrWGZTTo9VaTr3TTHJcrkzVqJee9
Bc2yFVQWURLUy6tZRtEnzgmak7jWHbWYxggTzkOfGAP7T3XUQ+TDZspUZfpsIugJCEizMFpsVQl5
U/HF4aE1r7t6cRe6AJWFt+I1i0A19BjBYb96bd/IW3VeY2AhFg9CMbcD34Udr0PWpmYrsrR/e6Uc
mYcIFuO1ykO26ERLxq8CeKAITeMuDQ5ZQC7jAOVWGXZ/bwP36YAqTlh5da0L9kR7NDCxSKIwQ1oa
8ZPougDTp/KYkFfTZLEYJnY+3uNIqpivTolEVAcuwibQ74akiv8LXKP6xdcztHEvSQxVyK8pFXNR
eeUkAouR8zNRnpbmSjEgbsijkTZ/RvLV16NXpyK8PMnUyOiMYjdZ6pjaKEJGASa1yKs9sK1nZxMa
l4wzWvL/fN4Cq8d05j8F1eXavMt6RPtVqFUjjP9dg8nQY9aszdRWYk6RX3UzYOj2MgrygBM0itqU
ITusBblLeNpZBgRPAQ5Bx3dLj0zw7ODEj88mDc+uSak7NTM4/9qC27uljvmnsoF/qGiY8ZkCkOTO
wHCwoc+odURbMqW5QhpneV1ZXwt+moINXjXv1pecuOige4TgHY4IyHaRzUS45bRzyoUEzkb3NblO
dslCvCtP42b2yKLb6+xWGOzqBw/sbUIhDzxjN6KgTcVWMH+dvAObk7XKJO6AT1v2jGMuB+OYaDPl
I6f0idYLjXeHQkWDnRst3Yk/VCY10xHDbjV6zxSctlAhqMc80v60i/tgPr6Z4bFWhUAb5/xKfkDF
kcL7NkXTbpj6itT2qRWvWncyQsB1l+Lj+oLy7hAQjjlThkHa1+9kMXCL9R57C2Om9k0zb4/ZQoxh
1DlRhqMvorgfQrIN2HcnKZCod1zw54UnJ//Rn91AZSEUTwo0gvdIyUtLG4JUbeWPyEEGi9ZL1IC1
5+6OzaavAVY1BtPE0ADIU6O2KVwYY+f5LL9l8pg/yMeSEgWVJBIFWldl4ZP6K6P9XTu7rp03/pbS
7ySVtpkzWDMmzRY9BJ9DT5iv2f5ZgsWa/pr1sV5J+wOM6oZd4lmli9dMLE3O4Ah0cJ9zKjkKXIWX
psM7CTLtkMl7+WGoWFXhp6tPldUSVvzOIBw10Ocj+d45p+JlNrgQEC28aWVeKwnSpZKRMEOh0OZk
aRGGLEkMI36LvQCbqoH/FryTkH/+zKIejAirWox2YUJLj7kxhA3ElXfN9QyWle3i5SupNC7Knv0O
xpE7VnyI/fdAYuNH8VZECtkplWttg3vdyKfi3+bg6qfCM9K4XufrbbO9nrWGequvrffy9ntZ+ESd
fu8E/Pm6RWrAl5FW/NTEtH+tDnHje0yKD77T6XDTlpc7wTi/9QKByD712fk8b0ySk9bq3+WsRzfK
8qk70n7BhmeBh40dABdWVMCjHbn64Ur3e1qFIffJrbNvwR1szY7tOKSS4TiraQLL9/LVqtJypNko
SR8t3Z0LoaQZLcGUKfIkwPaHVFoPZS6E1aYSkVR7HnaFr7sCPfYXdgD1tFqpiJGdxFKQ8Ga85/g/
JxsRFqbBl5sC6xL8mlqLGKEQwXsMPRhk94aQEvQy6kAHIePhxRgTRqdVlka8mck8NGBR7+FDiAkO
9fFYN6kKbBv39gwZVZC7FiOHfse4p5HwPSEI13aVo6uQgIgqC7W/dxC8whCqRhXxWyDvMR1Hp68t
h2bJkdhtz2hV445EnIRwpYW1Qfer9jqj4jUJhBbR7SkQ6avswrEzElM+svXNvAOhXxWIRgmhaJSX
EfCSLi7iA4GOxph3NvNukR5ncYbX/4idhuWfee5+PEbPy327tqWnVGBXFD2DTehGKXRL5FvnvrsP
t8qoMdGAVW8wtTnkTzvzngW6gdc+7ZQzMiZmvRJufs3T+bFTIAVfWz4zFoAxw5wSqvtYjtBlhxDW
YHe6OLyJUcpi6qWN6JfXEV7K3ieGCclPzRv0k/6cxfpltMjCX2dPmAjJDkFVb2HxofhcjFeIWdam
oGUF5HzK76vdAA4BkRI5EmU8a0eYxOAPiA9Sj/i7rioiewfivnVJZFOoHFGxjBvmS8SdG72MBpn+
CxPN2GXlT1OPRCgD578MYn8J2ZzBTZGGM/vev/kXyOfwOEROte/qbdoe3Jk2GJaB2knzBTGilsYo
lcWRL1SWNzZTEIbLPagmkmEQ5Yg7FdK3KhaH06wAIQPIlQxzfEPUKO5vDlvFshrsEJ7Uvlbxye7k
InXMDhDOMkQa7eEmk0hffWZ0vvYEHR6ftMktjKhOQhCXtXtTqbKffAzXrZOb19aXHRpo03bzwbCO
x7ulGUd3rb4khRBPpKhMlorjwIw+hvieeCtxq6I/SOK5sjR5t88tSjOI2E2f/Cwx8aocKN/nItr/
Kzun9fXPqgxVNpHViD23Q59jagkmwt/jdnhB9BEsLbwTrDUkU3cIdi/hA8qygYHxz9qpLQaDhgOV
nzhGEfVjvmD7IECgkrgjCYXDpfBatfH2MSZ4LleTjPtYDYyqQ6PLDHz1W7nu66cD4qiOOwMzM4Q+
W4Lb2OEHdc85IFMHvuDMkxdDDzXhKFyz0KW2z3+8iQYdXdlREnfqoSA47g39lsjY2kgH1eyIcSLf
zscIBZ8jkT24P8650H5Sarmdg3ClS3ZezubJm7fIioPoKT0QANdM3qCDF7OG7oBPN9UZyxbQIp6J
6bdDDRrYDRSSPUC5KkwjzU01sXNoiuhU8ypJEt9gvNUir1fIfG0m2zVqbq5UxnqLecjmVprkXy2q
1R7q6b7fEVOhPHAHJ0thNL/Kli3oCvc43iNlA3GkpirW+N0JcEp+r9xwuDMSf4RI8qUQucVknwvv
YoU2fxfm4jdybNHBqdPkpnkJojm+EH6ja0UH/l5J2BUQLK03tR71pxH8d26P65tjYWzTprfWoNfU
KE7UYtUSKro8TR8c5nE5I/0xmpugeF2WTz0FdDXkaO0lo+47bDCm3qXzIb+y1R9XzJVRaqsmblbk
kRJOapF+2JeSbJPki15xF2q8hXqmEYOl4vbHviT/P8t0c6oVvzojXZGMtQ3O2V9YQwTWELzd8wkK
4nm6gv6KY35wQPOl4Ib42j7NOZLJhUXQ1DJoFwMQmHksTn/s584YIRzQc2cwhCtcpkINIs5ivONt
cG5CEiJBf+yWg5IjSMMQwz1e5H6QR2l9D+k1LeTb3jJM649aude0e2iH4OUiYetcuOTDkd5VtfzP
MoRacPIXW9YIssojNC6dHSVk+p2E7XW1EGrrHyWb9aXH3ku16d5DqiuA8G67A8UefAQRMw2U1zmd
I822+dn2OcPy3l2TaXI3Hv68uqXVRZIeCVhN0rWob+NVU7HLNhdTl8K/eiFY3EkaUx0K0q21DLtZ
eQRPvnQ8XNkmjiLD8UPkfXZfJrgp9h27dSBOTm1GBrVNhE0n5JqblZ87DZBa94DoChDKjKxvgYca
3SnhE0JM41r5VTpkxMqeAvHNIOtiaYjTRXU4vLvQQTnUJ8CUoOvz4jwqHJ7QvAlPs2Q43QqDfsSL
5s/ViLzJLzw0v6GJbbI5sPXh9PpoKlGr/0y5kLJ0HLFKBQq43qI0pxSHSaaa7Q9RXO3fjjpbM9dD
W7C5tlRVMlu/TpXGewfUZiMhdWE/f/uXQFxiEO9C7Lzk/7sAJ4bdc73NJPjEs1opC0LNseGpPUGv
zZK/hf1CDdZiJiYlPPY8mDd69Kl1Q0UaeqvkRwHmGo4Jv2WprQaTnGUWgbztGAlBSDO3cPtmaSlN
ysIOtWHF4lEIXBG2zdtkzTJOt6Y1PHbwVvP9p5MFo4p+3Fi6+OLvMQteeCvDJdww9QSHc9Cs+B5Z
ld6ha3ZLN803VPtzOKN2A9xUuDlNE11cY4U10jEerSeMBG0ceelGrqeHKL7igaKeyykw0MxAP68G
URF6GMxdcRjaL1H3jBo8hWf5Cp1/t00B0BOHa7FSldKSeZQVTWeRmf9HEx+jasdLrHmTb1SRi+rq
vEzyuP0sESTnRXi0Wg4c1wxF6+o62Ouhs1+j98nS3flmooqNe9Jgjc8YXv3PXUBjd1yhCBHyiHJ2
7nmmnXykGMijsobUIcfkuiUM4fX1gIEYCiE7e7tH6pl45SCbfNDosxzjRZAscECrNCzssF9qcoiz
8TD2j3baeGhy2dSCnx4VNdIkRATGrA1noJIJyWAzeKHBp3QoF8T274Ys6Xx1qTVrw62sFISFh26X
PWWwf32XTfXhcgVMuUmdYKFkjFk0dwI7ccvqIRQx9qTJDLyaxiUen/M3dyHdb6PEMpG117poLpuf
16hI7/ppx/4wxnCycEXzwrafN0FxjxdUtabOix7U0jKFHFawaJlDnOHCRZATuRrVVI6tTPIimUlX
VZXRQK6jz6DNpB7At+pQBS1ajvwgOL8B6IV7pS27fz2Eumv7g6/JNRGwrpk4TWEaDYxFg8nKwTNp
lc4AH/hqSC9jQMpEwwsxc2y1lqWTTw2S2iathFJFBwWcEn/Fjki1l7NFg3SPrxvLREw86nHBxt14
fRD2+w+gFsMZGtYHnG9VyIWDICksXljDSZfcDFi3omFYFjQKKjuIXUKGwS2OavFQh1MtAzvLZFdS
ixfz4ESkT8GX7huh2T2PYiD3LSRONlERx00CXK0xDPrqCRG3/TutXpgwhqxedq43/NhNfhtAekjf
9qlhZMiHHuz0X4xxgFi93uQq5LeCc46vZlhDRlg+RdwZDwNpyi3ODntSCIzxRrfYA8ct+2G+YHG6
5G64NWpgFVyXSJiv0TX8uiTsRpzCiupw/qkW6FPVliLaIBWvb0Vaanwy2i7S97RkAzQLaZ/wWsVi
ZRAjrYK7/k71cjAAAqUozqV/zfmwt2Ag0wwIpHG2fPWXnoPyScHUB0v1DQxR7W/Kx2DK8FU/3n60
GUjQBiTz1kBB6tV3qQ/opt5FD0RnQWBhuwzRtKC/piJ9SWuNCdAddpO6S2tLJBboMfNoZRXoQEFb
uGmpwDRFhJedfB+Nt2fJh4HnvBbuYxEdn6+JXKFNvaxhaFBv9SE4c2KjvFk4PyGNhqQEGSWgg0vY
mRUz8sMvjjRlXio8vARMfOVLcwEMOBKUSA/sYSicQ4ku4lEXZHXpaOy2ZidhsNV4Ph9SNeAvk3b+
65SPBaEbRp/TNrzvffgdGJ1vBG5TYmhLnMNp5sgCFS3bJncv6cgZ1f0epjunkI8gBi437uLD+XON
sX9tHTqiHpN5QFNUYb6Ovayt8JIQw3+muk9Cugg91XIqpbKFtrMwUkv7FlVs9UT6xKwAAbpX2lkH
FkqWA8iydJUM/on9EWDrs7BGkA8kgX5v7iGhwFanNPpSU0jCv058fY3qVVIwHEihuj561R8Gn9m9
f36ihGfCHV7Ih7099XiValzhhJsCmYZUXc/I5IYf/rZfGlHg7g==
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
QgdIxnNVUf5qhC0x+U9uLAs3cgs+qKGu5GA0q/T3IIijNveLHj5e/L12JJKoy97W
VEVUQIBnXz0v0opTcCSlesMquD9CFcOI4hWQDzVbHtE9QtQ7s1+VifiaQyDxi0B2
6ozovz294fscGD56aTsmdY6xg2v7RpsF2Pn9Smf+MO6ndTIaosBzoMU7UiswOo6M
XrYhqYbA1ZY4zIbCdmg4AesfxjjHjajSWA2qthqVsQmHfY5USkAXUjtGzhjBeoys
dLGzI+C3PqI+QW27riOInweZyZ6ENMhcPqKVFIRKWEqIh+iEVJJ35+wc2aF0cfX3
TNk4LRswP8BPMrGWkHRwRg==
//pragma protect end_key_block
//pragma protect digest_block
jaZJGMG6dc2fBraglsDwHRHXk2g=
//pragma protect end_digest_block
//pragma protect data_block
vP/HvGx7mgtRs7SH2gyqor5t9RMMQT3Qyw/4RJYcmW3a5wMiCNs59w3GshWtaDxq
WOXK+dCOMQo24aD5y5mUIYM3i3yu5aLzjfBiNMGScjA+SAgr3bliD8ZFjgpVswJ5
xKkkSVhhOE/nRR1tgEvcc75qF0nokjsyuKIQVzE8XOQ4qJcCC+d4KQwaok8BR/pI
3BrRD+XNfExwNKTZt8s4f9IKfo5xrUzQV6j6f5uM4vWle+yCuVxHnOAVEndxVHA3
iiqKR+6saD1jfv84KdNtqWDD38VrSxllMum9M5krVwHikT/BQjHL0DZ94sxgA8tU
BgcVRb5hFdWWolHDm91bBJLwp7foUdmvkkoxcXN6lLW/mRuOTCrpIYNAmZPFNeVw
qPlglA++3D2UAioS5cJ7orRQwn/d3BnUH8u/nK/ogou09X2dGP3quTZ/aSy2lgRb
oEukC7Jk/izy+rFAOy036Pdf0JZqetS3H1aWGxzwk7PT3eNzmg434hwoPT2Gjd+E
Gbw8qR5hfoxfp6aGLlyU9BRn7dV36/uekkjwykwx0HB4SxJMNU/OYYjQ8j/eudqe
O2QgH4lQVmwZrkWkq3TWU0AuJJbp0PxOa+fkeCSmIDfSgNqGrUkVCZq5n97pzeui
vnaFr6GzdiTZ675ooxS3YYvcXEP1OFeoRHeD9TYAJlRuh1vgSzGasX1DZ7JsbCId
zGBBCqLTOc4uFAiwsMbW1bBYq7ykGDLwcWMw/8jp7wSN72ZDTcX2DaTv/p0Fj/H0
ES+LDSzfxvBvyVCo8jP/+FfjK7ZJUFb6SH3MbmIyEUb7syeiRZkFizqUIbEBBfum
lqCabShFG4l0Kh6SzG+hucLnVKtfVxWpYSxAFsOjn73bwy0tMR1ILRr1nYA2mpNR
Sl8thBNGRZlfI26lg3U8hXL5Tp5ivUulJHVl157TdCk0X4TOBGkE+Uk0+feRH6mm
8aQaOKsdgPNaTK43NpwWPKihL9XzD1KgjlZFPGhasLTG0h5qVYA1UOwUTgvZ4rua
maNgOHDmsSItpZ8Use3cS9UT1CNi35XhTLYWMg7JQpZLGsnzT4x8YZ7p7q11nET8
I/Z+lPFko+SSJ49co3Dl/ynECp+pQInT0oxFhp8EigVsRYJ7nYV4pbn5dBEFlTym
4zAtSKZDTidn3N8JkfvlFhbkuoaciF9jx093dfsnEv35P0HzINsGlYVWi7FLFMFF
VYjCwVpLUgTj+RkTwiwj0AHTVJfahIpHptfCKMtYa0SJjyvzl9XA1SzU+LZSP9lZ
jaleXw1woA4OTmURWFv368C7p3T7QmShlSZOuEgQfThx0xPKxCF3QTGVQTKgEEtM
pB9JZJ6AvmMDHX8h0SkDFJQ6gCys+eqvyLLrSydp7mx1IdzTrlbfNEM4K68Uf8p0
wVUxXNe2Kwir0l4CAwnWImwapUBcOWHLDbz9uQ4zPSGF/xbp7pBGgmGs3SPY7mLu
+B4WEfN7lTIUCKjdSPKncqhWy9Lcm2dLuZ2PLxfDqpR790oMtFPctLZA02uyBsDA
kbGuL6P8/mcsJDmaRuSUyBk2trw0ZzRYS5PsSb5gDnobj0poRwO5qo12GvcW6K74
DKWjFyI3uYJzU4aP5QoFdb0RjI/Q+PeMXnMnraTm0QrTUpbmXREmKpSPE3BbmyLo
4/Fore0XIo/jf454krI1GOg7gxJk+QLofwBAGpRcHvpdJtZJ8Y63oeuNoeZFPpy+
kaJV25wsSS4gp5w7rI6+KjgwAaaOiDYSHhbPGbwzXKBdRwlzYIoB4+QlEWC1Y98I
FzTye8pd81BpTKnTXlDlt2V2x0I2iXZmVVJ/aK+VN3lJNXX6pxvCUoE2Vrfc20se
mVnAy8dxIhf5YiCt7yERylK5AxM0/wR8+D3N3D0URNYlfq5miBhBhPbwcB1Iah6+
vDtKAEO4RDvrc8gecnAvssYJ5OvxPzGS0IPXm1fCLNfPSRcIZ6SskRVlC+cWT52q
tZ+zcRfFEAe81a/viwKGMYKAg3MXAc/ZgftuuvMRkb9r5VogDCum8CDtBxIasFTt
0Yvpmu078ydWlqnFdeaYl5fhcj2l/wIzAHqp1JhPFKhpvrXfFPKz9YVWflN59LJb
gSm9T/9EdNbjZ+C2HZc3ntw8YKhtAS2+aFreCJ1LhxL1GC924NjUO5MC7Bqh3lSg
sH+0F3r5DbKSQxSd7U7WmGR4kes6wb/odxcQbs2c+pfbF5dAF2AIOP7Z4NBM5v1x
6Pk3DVqOWVA1utl8wg5V8N9/ONBhV3vS1A8UncVTpRrA4f9QlgFZJ376DqJ+CpHh
LHjRzsVsMrlzBb/xRLMrAkYjPeroObrboiFnlm+OMSaYZ3vv0OCHF3OkDeMWBMZB
ckOW066Lr3Ejnm7KRwXNiWr4wjFcKCaj6d2pGf0BwkQQeTk7WYVIBdqqhbM3JI5r
Cd3Li359CN/x92Jb8fN5ab2BtHLI8s5Ye+fgUiaUr5hKgl3XmAElIEndEmT31iBK
NaYgCt7uA+7QwFddyx+kubij47AHKCJ1R+Xja9D2L8hLovN5sTlOj1FdZIp0aQ43
KZPOdq2+EXntuwv56crhepgWQZV1xgtA21mUYJtsKKCxzW320uXqT7urt3d0YX1j
wZqp18CSmjy5GuowRoYPZTD+9qziTzN4svgYN/dLmM+IRO7V3UlX5sjhQ3NZk/8a
PlIMkufa6JezIGP3rykDX3TZVqUkyy9XGZEeYyhAozEUAZl9rKu23IV5kPMCdnWj
YtFpxi2fpy1eArPe2cCazKUGK75cH9g3igGHgirhHWEDEfZcz9B9IDqcpoJh0M9H
wvLP/c7JkceBxVyaPA7TfbguNhISjaG4ibLCdbCrPlKes0fFNmbgQi4W7b8v4TEu
KSr45Hxi4fZArVlbxd0LsDmpik//rs24JpRBUFSinZzqYYPPMZ6dhNAgSSW39H6x
1yH0bTWsEeaMIlbikot9+ScNYozQNjA7Fb8KE8LV4k6a+K5VzRmCDea43fmFVAtf
0dcaovIac2fUp7Gl3NAhFlLLmQSuarBBwLpqaybSP5RVL3EqwAaBEUORLpJEws7v
XRY39oFHiRp9ibpEHenB3ZqUBUFrqWTKaWZrCg8nTeCiMD8lT3aCJNe/gnuB84DW
anT96l2+8e320DmKCgfZlbh/znBwucW1SJTvfuFID98s01n2u4KmOKyjkaFThqkB
iP18MUGK/Ee+D+oCMi9domRNo7Xq0FEhGsUOW5QEFW9EeJvRbAPQKVvZQXoVoEKy
g4MgIBCiU8SGByh6/2sW9U/ssHv8DnlWCafr4ES6hnDVUZ/b7oVaxl6q3BKrtMZ2
8ELT7ayl2nq7SVqBcRTKz5IPGmwVM/2gdYeSl09bNZJCvU3fvbkMC4olPq8HTin3
ZkxibhsOQENTNTtY0QMvzVZPDYq1HFKW6UOWugxUmNq7iuZSkUw0vmtWPvT0i85u
zsKBiohfLmH/A3/Fn20K9Ntg5NWCYJ01Ny+wf7CQrzzne6flQ7C6ymLyiYxOkaRo
QeTydkNz1eqSFMEaSXX8U53hSjXm7JtniBHgHnk4p7URhbdIVfW0SwbR1OPgiqNp
WE++V/Fa6BuWPxetm++fndLw05MUmNPelqfZ4iMQb0H2poadwVHyBABRT1kE7S4M
6j4IFtJIj1a0ohBEMiKXtkOb0taODGf7iyptvzsixy/s5EvlhRZTgWEp/DcjNwFd
N9aDZBo37ASqpP6A7CjZZeabTGx1NobrJyrKbysMclBAg8iQMAXOJ/h5jhDAS5cY
eK7kMvB+XNyUclwdsBYpfJCdqF+HudOxCXcT78BPiaw39HsWukxRXe+PdB8QyAtD
YAmLj6y2PyZWmZiw4utWzDpsrUJ4dvTcnG5nC3D5JTCB8VOlfpMzQJ6+c3HrLF5Q
hTafXtFoOc7prwb8uBqPc/JUt+xebX8PTfpcZvu0c4uISxhRHP+UK2O3daIpMEnn
xOwBVl/49n8kUdb0p6lzEKQt2lbVoX9NY4Np6s8kKAu1X4gDq8dQeMSFYqIKe8r7
dMZXtOnbgnCHlpVso/wp7u77V6RsxU5FswuVgshxGrAlbcEpmZ6PEJa0wNNiqt0T
OnF9+M0EpWQhk4JEj0OUjlk6x3jf65gS9P+zR1MuA4sTGg76o2FrClwh84hD7SnD
DNGs7Ibj97Wmki4NKxY6WbD4rgBp6xT8zgW+zYH5gg7KcN09ahHCgTzdM4m+T+zU
K9ENkaGnp0j/z+yFVaP2BviHFsAnwwcUSDYnR1/nKsN+YOCbYaxzadKskv8+QcXF
GrbOkU0XeIfEUk0FKhVwGN5ly/amek1qMisx5SVw313pr4JANYbJEM6F1+SDi91C
Fc18iS0tOCCEqAUnzKBY7JYmDY3mgQyhVEc2f8HOmaQkvvSlgAuTazqBXx/erR5I
ciIvvWq1WHRCRApe1L6qjWhdP1z43/OBJksuBVQ0zdBrE98ID1FpH2sd8RxxZ/ZY
rJfrqqPeSPto2JaIzeMFQBs96xuRy91BudUn3ZJYTKhgLu+vEtoalHYW5P9JYkUJ
ChFowEqm5F0jug2Dp56sW4keWMcYYRNRcHjxZPeDsLTs5WBbm8viAYlrmUG4sxhl
0KbHAPBnCO50vyvWWNQb/abq5VspaWvOlvim10+hAu31kmLiXq7Dyz4+zUQ2LyeD
jbJHXGnrS5CCHwgQ6ipxhAOtUTmIoeQdG/0WdiOYwqDM/3e+Q64rb6O7lh6YzrfH
7BPhLhBfLUFn6Br3SP2fBG7dDiNZ+l8AQS9JL4S3X8pRorEiDz03TY7uoh59EzMy
4AgYmvoplxFm593wDsqoyT9i3bVD/3rxG0p5rpmJ+9UrAHBqQKOsOAyIIJKhpSNG
57DzKhDgDgTlHBVxUWpSON+Gw2EfTJewvOsf61b+tCyzSZkR7UkGaavdl7vS6ce7
rO0Q4URNjKEmhCn4392HVpPGUfKMR7pI0MUm3VLwBrKntkxbFoOAvz/+uzixgBSj
tIyhyHztQ0EKnl7frcClw0ONgXgr9Ns7E9BnxCKu5uU/boQZkF0YzHU1dwD0Eu23
vvPlAoj5187MMQVqm/4HbD1h4UlmeHamJZ2AHAtwZAnC0ESyCyXuoehegMHYphA3
TXcslV6ZowWXrKIGlpP7/qtofeKyZzBijtqO6nJt+Wk=
//pragma protect end_data_block
//pragma protect digest_block
yJYRNoMfce8EuTzElc8vNMmVmQs=
//pragma protect end_digest_block
//pragma protect end_protected

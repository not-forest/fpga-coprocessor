`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
VC1KLP9hjrD80jVKGStO7HrnxLYuDdrGf3ufJZMgsfKwev3CzXZ9JLoi15S4uZyG
JPpfUmu6gQ0gMBVrzn8gVRv4HPg3Sqam5jQNuFv+guCzK7fg+XLcel+jgtWUNT4n
mwCMEOYKOBi4wPQ8D61x4VrRXlu87GNp6ElIn7EJDeA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4608)
0MNOtOgUPuxMGFyeYrQIEaP1Vu9Bypl7lU1ojLcwIT/E3IX2Ji7eUWyOMMSQnx7q
XLeyn8AJYe9TBoTQUrYjEvsVcIz6tgxXV1KzBR9SkSn8HyH1ZJ8VC1C372YpBBtf
ftdyd+TyqB3vlq28+p7KGHOSpJIWBRLEQ73UaPQIx6aAfiDgXcySnUYyBcpqGKbN
GunOplGHQKMD23FpdeHbZJzGIp1ftrEJ+ycKmo4aDx3DrlqF9aEuppMWSU7M/wcA
XnCuxz2j4vWlmYZ+KYLViq3KwsSKndpSA7XmNS3tUj0O3UezxQkizEbcrZ64vLjD
Y+MzBWUAT97vgzaw6YIRDNDs4EZ/geSZVVKJEe25OCqbsCbWETvJt3xC5PAbCEn7
V25fsisVA310a80WYiG/xBDr0/GRIpnf6Pn9DiIj/c3GADrVb4T/c6V1ZTu6NtX6
aubQl+QW1ZCoQg3UAB737PtFILdu5rfT+XH6RE9HSlCu1jSsiivSq+lwIf4aBbmz
vPp/pK3svPEd1/J/s6Vr2dvSj9CG1iyORLa6dQP07qcvfZ4fpaBfW02Ift/URX5k
kMFtDhGPuG6Xxtn2tEzwdfLdgOpwkQ13X9mh2HlJbL0VFUq+raaC2NM9IeHA16E8
OCL2PZQQzWYDzRZWz3ibLgTxyF2u8LRUrBtNtled2lz7V8YC6yxNpLLjtL4v/CtY
2M6lxHVjCqWoNrPwP+eygZQhTx4VJJP81dfvGgATKebIC/FawOMUdpZ/HmDBqVEv
SbXoyHZ3RE0ncuSjOwxF519Nz54mZqBC77dEvOgnfhYjwCRgYTqhT+CjNGuHa6tT
DCMc2TZ1mkz+aWdojKPAd6pIg6LnAAFMoSY0zavP6UfSSX4hHvD/VAsA7cUgqFDT
HQ2ZhWGQ+iNZpTtYGP74ZFXdFtuI1PkvmnZmFyoVQyDHgfjr3H58TT0VhwFxYI7d
pW0LW1ZpvWRbYQmMedPWYAOryz7x6xhWikPzkpc+UmmVTu8ZFVpoUkfQImTYSfJN
ca3FF7/8RUpi0AU2xwKhfexVxyqsRhPNXelDs9pK0d30vN05R9GEuiBkdHoiD5zS
kAW1AbXJoHh9qiqRH/WUVk+cO/qL2rPd6xrs+AjNuEB/2FuV8yxDqHvgIhv6MS2X
jeQXH33IrvVEtA2K43EWOglK5MQ59pnDmNX2XdVQDMO9i9EOy8yHf6PO302bil31
Q6Ux/NfMGJNgqL/3KpbhwXjuRyNqH93u/Snh1Hm8hmcsyoajoaK6U0Qet04H2bdV
0ghlYqhwGUKCkP4Yiu4NNxpa4cwgXofYK3DYfk9hVmQUhpLweY7Q2y4421gYSGcq
fFS+Ol3ouFRw5jkrKl6uO8/qrsz3WygEogIVWMgu/Z1Yj3jGosZNupWw5LH6aAJC
Tnu2WuF2UyPyI1OSETp4cmDyt0HyukMUzZb/wu2YALS/Nj3vIh2DZVX0aHGxvvhQ
VIoogx2BvRncMAMirkvQ31RpGvO+aRsYhBLvYn6OzwgmZbIF4+jcrTrZJ5lCnhGm
Q6bRjAan1t7KXz2aVMvs065CuBNfSFQTVNbuieor4e9loYtyMELtjbYqYdkzINFk
eG95C+qA52ZgC1Q4862WWYHXqbqCpgaej2WsI3JeRBvtNEOD5jrNVGGqQGPLeZ2E
C3fjJOhtsPWKJXTmM4uQPdXqlLoPjiqIiyf61rcjSWCY3gMd1QZh3xNm7uRXnska
yjX+RdeGGuDY/vGjuNJSNXNJWnCkWYyvs4RzNu7ZeRoAApE5Q7mOxhAQfdOmnmFa
/0/03G6kUIEHD+hLlfekH2bfsfBEqqj702FSGWmyybBNyvCQUDK2NHvVIz7usy0p
tuCF3oopXMYmnYy5+2Vfpt3UNUlBss/8kI70RWzwGsfdnYIkgM484Pk1/2W7lI8t
8Us9fnAbGDG6rIUVjrGnm2j3ubZyzqq0jXbmrYKRGRfha/T3oCYVru6O06UVIZq9
x+aMtKc2oonNVP5bxYnZ4xbfA3zkYFHYX9hLNHz2NgztyRu9uQf8mP0sOGPp6Qtj
/uUQXY6ndnkmXNFPytgFuhYwKuxUe9W4mgWgZyh8yNoYb+1YGUNmb2iWVxyVJWBJ
GwYgM24OOzw55P1ZB/c/qccOgTnlbfSaFClusdGSNscyTfqLOA+ciTQ7iQ7P4IKT
G5phwOKXucLcsrC7bHwwdHvimakq5N0z6/FreWfnabS5pw5slKXDRv8x9eQ7v0vQ
R1n+XVerY9WQQY18qHJX0r+55aX2616KSG2OcFEbYQYtihE1VyiBF/8zkJ6Dka96
GtlbwLGZOmhFF8BSE6/CBRRZ++nDHgt/TSLxeGz8tSAnoBtmgoaufg7ZDhE94kRo
c5lHUcsHlfmufD1IVaqSPUAicFKizWysS2vZ5jYXy49vztSrtQzsbh9T1DoY4QF9
8VWGLKxfSVW/4l0JEYEd5boLLMJHUSAawLpFIH1dblHWe1LtU81wWmseXutPjfdu
yjht9P7AQp5i2+dB15t/6CA8NTR6vcUVCH40090ma95/F0cgG/Tb0Mw1AlAcVhHN
HubBGKsaIxBTsdr88aj0UxxKuauLK+wwQ1tNDJgzyqbjQl5CsXWzIdhfu47bH64l
W9xe7rKnF1qk0Pl+h6LPDO0EFwLRF4tS7rQIa+bFXea3zIFhEe+9mHwSY0sumi45
HWuxJOuHKHsFE1ceesOE2ravU6JKEoXkRfUPv2X/EE2oHRe3Df5zVMbVQIPudm+Q
eRlDfbgawsTHFd5AcQsfAtgDhxY1/e4B4IGrhaP9mv/SYWQVl7yjqQvRg7F3VtBL
b9INbOiFqC9CgVDf9RZOYB2KGtOqlrX4klVK4wfhvZjASxcU48N4vXlCjvaN3Fuq
rf090SUKOQxAqBr+fFCvOsd9H7CJp/EQJzuuLqDrp5MYaB5fellE0hSk4blTn90P
/Xi32pbUykVOx6Ut+ZuDQMveLtptkK5uywLTEomk843LhP+2quWuHvhykgWy/rys
r0QTV1STc14ONPxC4tqIaVkLLBHDdDkprhpG/4zwt2IVBQvG/3m5XLxHmZ7pp/Kf
Nv4Ohh2qqNaMCnpgEhbuf4NF6ZRvsmrhxelRUlEcddSmXQJYnKX+GLQwNwOIbrhF
2QFWKwCkopcAw1GJsCqqVeXTfRk/r2JQTI4JL+7+riv7UPHKqsfbuctJ9E/YHkRP
cjQyIr9L4mvNVPGLDASVuoacloYMCQijyI0YGZJmlTpFlt9I5JChjpUtk+OoHcy7
i9QR/gaBqH2uidgrq3OG2KVDw9ENMNzYZ35i1N5Z3e+m5TyC3zysahOv46Mfd3Ve
HGeQjYgMokzVURncK7FKsxpk8Frm4r83sy6JqsAWj8tC203Lhu0/+3S+wNz+VPhZ
YAPudgwG1LNsyFHeQkiw3gBfT6ikSDvcNgFwYSY/H6UlTv8n1bz/PdC3YtL8aCG3
tUkFAbxhIsL4ARgLR6pjw3n3LHw6t/oTxsGlGqo0uPPdBVOlsy0QzXdaR4PaZE+s
wufTJsMFfz8ZhWFP+UbyoItpi3nbycgEtF14eqHfd+gnVDC8N5vIgjxJa6ZWs+bs
NKN88+EUPTTN0SdeNk3S0+Di8RNU9WU7GECZnquGRmgNxhMT36E8mHLX/wRVP9ZR
p/FT98dLKwXQqgST2YJOrx0UBtBwrjpCQpWTBhAMiSppg4zFKVm1vwzCO39ae8H3
qOTKhqjjQZcRtER+vILxTgY2wWJW+zqhZYbjYb81P+QBESBcj19BBBQGjWoDm5AU
N0X4I+rZS3no0jsI5dH2FLGfw9h4ZsaRXCCdK5wkdXgx4gmdrMtPb8i2Xb1oZxjH
IXt4TQ9qQeLio2m/+ARbVQIutWTDqgprI9hvCwuqVz6KlZv5lNafQ3cUDmJG6wMy
un8r21jbJbQ40CtNWdYHuRnZ7Fm5/Ip8bNGl0Dk5r10LewIdFKNiZPf4f9KXg1WG
C1E7cN+pNIgBcywezNxNnyjTydQwyMXjDgJ1EFM9uK3NZaWbenCqt5BG9DqDlEe1
w1ILaBdBjI46N4B2vkD+1GmXBFqIduCq7hKNfaYJgUkEf0xkcyKK3nliHnrG/yrF
0RW5Haj4LMLu3WHD7fkp2Mnwm/n01PIfBoqikz7PBu7hR/WtFh8NBc42U3b8gq4s
GFHOaGQjT+gGGCw7yArVw6V59k+WibAK+4WZMtYdfSkehpVGRDZobTQKZ/MmQUhl
hR4glFHGEYezdm4ZeRcRnu5zp9BC98dj0uKPiQczAawlYu784QMHPuYfmukyYSPG
u+aZw2g0iVQo/Y1jLgLnpkPqAih8KM6Ut1IqEBOF+7UQvKEV21SWoPPiYvmkw/+i
b4UfUl1lHlKFPdb31QN5X4muruZjULxX0k4t7xMn91S4yCXrxRK+jrd9tbOlAhI0
cNijEMVvcKYbdDiZBka4c7g6/CAGeB1CKd6hMLEVpGZiSYOfiedvV/4/e+AT7+Cd
JrQ/QfX++hPomD3TaU1ggECexsekmW9t50v9OGmoQhZVxcD3IYSiD9Sqwh027LF1
W344q2PGZhSTuvwdbjJaB91Fmw+D9fFlt4hjizAiL5lSOJpzXcPxmvmPUlSi8U+1
crs4R/hurTqfNaxUlJFg+fnQMhQoek4r3rha0cemtM+x94j6Jq5L1R/CsF54q8oI
heRtsyq5xR1G/Iy/QzhOF8BtbPJLbW1JPw0ksf4W1VU2TkbIYnXVf3WHiXbn+qgB
HsTaBwmYSep8lzruZAY9iw0HD6GJJIjoCjCTnsDyY8dcAHxcP+RyQ0NpisHFTxtk
OypODnHwUh5R+uo1xvEzQn9N7mqHYldrqW8xVJmF5e+NUXspBjbNdEpQFlHjL3jV
xj1P2+cVxm3E+lAyK0MqfjinoMC1/O6PhTECMUczeQ2DKkVWsAEoVatRK8ifpy+e
ubMuR8y71dt+irVweGSbQlAjmfTQclofP2VcjARzhdx/nAQrNkaMb78es48qYB33
Par08SUsC7fKKEf44Wx1ZBtLkaT2aWEKC2s7e+oeCfBQnR7hPx+e79HyavEh/b5u
cAFnn0JcF2WrmGO/BdRw4kakg06s9iinLoAjYfPTUkfxvRwH166B9Ro9kMmra0ht
NyiZwDzNzjBlenf6ZGzn69ywu5Wce3GufkIc2oATxQ9G4aZ6z+oDSg2AzGcyR4ip
ToViw//TPxW4OTwB6OHDXJXwmpy7YJXUPNFEMsTAUeIidU2Zqeix9jCgPw5V4AHX
ioYW8vfqCUfu2BBOx/adW/zH1cO1n6lVDO5rfLUhrRg3GYqgMyv0amFFrs1UJKzT
xtz8FoIz8aNmo9rDri56kA3NXdSJ9rt/p+Iv7OmG0vDl4rBgx8yXwslcNERlQCac
2RI9gJrUpFhEhqUkvTBhN6MB6mTSHJET5ljyMYPhj1oFlw1rPTatjDQQmmh67blK
IRdokUb6z/YjaX9vsIkmCu9TEbteYnhuJEwvVR0bT8qrx5/THICnKe8j3mdMFDra
fIF341ETE0C/uAiaIgK4w3u2BM8LSW5uYp4EuAtu/BNSA/m4/GTNX1APfSJRyJyy
uunrSBB5ajfGJaFm3lD/k8CDQiv3RK+gATgPF2Rt+jcHqsXOG1ASp/w+g+uz50SG
sF/YvzAbxZLxJuMEDYeNTJIdK1ofzjT8vIImnoRZV4DdAsWogcc54Fp2D3rcjPKw
1fgCfKosIW09K7Z7ofiRBpUNoLAYxn+G3JXuCwB3jphnzO7FVyJC/DCKz3VOmHBD
BT/+cQ8TBOGabh8A8hr1nYD/Zj1BKpMj9ZvYNTrSx2DJQU+RtacojAm5PJFVbHVs
k3pm/LfoPi+JtxsSIynpf9aAFwTUx2ZxDv0Kp6C3dsqLcTTG3Zi++A3E8FapBMBb
9VvhsOwi+xi/0AF3qv82K0x3h/qLB8Tgb2HfljNv7JGExTgkoXz9BZdBg8m7H8Zp
HfrOR/O/lDxYps95RG4ERr+sfOTgihHmjPnzy0lnRvKu5HTE2hBjYfwSTS/KZPnb
HwnLgzvplmZTzCDD/j7uh7BS+6eKUcmnWMoeRh3zlQTRbY5p6NihYG8UebLXDdK/
Cbj1mgGEhQgg229MzcyJXeGyksTlEb1RFbz4BxnJH2aVwdmnOYWdYx/p+3JmzdN8
`pragma protect end_protected

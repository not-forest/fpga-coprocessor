// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
gQKWKArxHM77aSbqtPI4aVRmuJZ3mKalbemqUCDPqZGjsmo+KyMN4winBC14SRjS+g0Ik6Ilic8i
qPEX4SNjDe/qKucUVWrSCatN1ZziRR6RW3lXvyI/NcdFknbnTJHw+F46QvnITnQblkjRxIi1F+It
Iwpb2ocvw5WAAMTb5sFoc0owA2/kX/rBLLoD9yPbQQ5cUT53YHuNMmZdjK13UkkxUKUa7ZHa8sGl
sL8Yk8h7l0Vg+AIAGu4wxgDZmkA/CAoe6JJpmFs1vJc3/8trX5zel+CBBD8HCLp5zlXmntYrLjNG
god54f61Jx++TVf/DBTiYfB+wT3kZlwPgrSGjQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5440)
npOty8URfSJzp+qYKWDRlYJWlABehzk/H0DfYbmufbzdqZQycQet9TlVkf2PecOM6UZV7p6GNk5o
r91xTtbkVJUVYHMAfOqiiU+DEw9q6u8WIcbKAy1rBBzV/4HkKAkG92JONXyXbu/MfCw8RpKZANpP
Xi9BYktWZ2s2tCnU1C+ourvzzDkzbsWpLN3vmWTnK/LBL1AyK9rDfPNUzy2575HAAHcImtBHq9es
Aff/v3RpM1ToMDYWKV0RwzZq7ZD9JLEwtyZCLth/bKiRMbGDyQjlRf9i5Hv9y0SV9ocr/DmePOpT
rdO+MZBqDEhJunvIumKXXNBjLz8i/idMxFpj45FDnJjdHPo4xst61uAr+eYWK3F6MW5HfOFb+T3G
YyMSybKjEmsVwli3ir8LsaF2CirsEml8iEtw57A/LkjIagzmzyfixWmLaW3WileimfMPe7smDhEb
Sw5QqG14rp56APGz5Wz98e3q9PHxXcxoKb7n7e9PZ82D/DM/O45DHIwpewpvDScD9ZQfM7lwMzTj
Yphs/RV8BnCoS1TexopTWdvVM+CWTRnkntvdIUvBBHsxqKI6dztvxDgr1STf/gf45oko9XkF1M2u
tKc/3DNALJzt21Tui6RrMjIdW2WZ6FI6461jIU+IM2j4KMWLdS7fn5xtHYdKeKgnqpYSXZo9sAzS
vH/Hj563Rl9GjCqmPxrgt4yQ5+273HsJ9CMebpDkMws5kuqGfPspbmTltQ5hpfYgjFQpqS1UPafK
DJjsS4y7VXtLRRGGCp3uFu0V3He1NlGEsYGfeGDj1W8CZ8lcxH0emXE7H4yJWSzAPx3DYymmGaua
zlMses9tFRvkZBywUHRK1f7X6nm1al+hP7NYIYAn/dhJ/kVwiIqqK59U7VsQbdL8GdHHzLYfQ3Fh
GifcbOGX7ySId1dhTq7Emj4JjJLVVYiNYUpq2e6eNWwl4tde4KFMF8ygnpOYkmFMmJRi2i7+0tAt
E6P82BfR4o1sth/V6NwOhTOlI/J0oO4v6CHPInlbl83q70FczbivmJ5jFhCq3Pes0rDMG5NvIcrG
u4D/yrLeNd4JocKAaORwSRNjzqAjeYVQwj7hJjmreuJ3wTExBg1AUKxuv56V/ovSZ47ezNuw13/1
EK9X9NXwBrMA9kMGfDnJd4k3ZAPEgs9Sn3R28ZrO1d9LZBpGNqi+IBDtKjH25XOj2IlJWKQF7ui7
q/7Wh5rbbPyeW5wCX2XBpLcLv7vz3ik1MqLX1cW/B8nlTL4oXcfjaPDLAEeKmMFr1oVzgvz/lKPl
gItu3sBh7W6Q3xfAhH9Umfn+R20+HPhryQLotu1oA1mfy1Z5d+Rm+K8QN1fRpWjprq1ZUBX8aImJ
eur2hMMFdcs4dLJcFX8VXkpP5UjO8g0eh2GB6X6/oKu7bR0Jy3SGB4cwbXYSzNqYDozZyAraSc2t
VaqMuq3S5+I5+2tf8O/CMOT3CJo13CJbIwvVE+3EgYJ0hCNmg4VT4w7VinFsxOOPLh1KVQPgPmfb
CKXZ5fYrjyL5FnlsZXY4z0QqPxWJsvpxhou4xhCbfa+Cu/u6rSRLijie7MazA7m1mzG51OJJ0T9y
LL9BuDnveolWsNGPghXX0F/z4wffIOc0sl9zhN1PixI40j43U8C82tAq6Q+dZDLIfvkVO0t6GrNS
ABHuZ94pP8ly1Lfwddw9bO6hju1CUuTPC66cAb9lPT6zWvWdmb2pTlxgBQ0KyJ75DndhRoM8XicD
7ibC+FsQVg6T/9TIugYbQ5o4hDwGPpQd+RPSJAMt53ev7OhT7KeUPHPL9/sk6o7eH1O+F2HPeGfX
qi4701iSII0GfJt/K4Y31LaGL9EgKgtxk4JrIkDA49Jw10XcQVCiXsGK2XJCO3GIUtJGz9UYnx2+
i36WSuEeV0U+WLHSXHWNxnwQkySiegB2TK7UYqsoqF7r/xOcTrtUlHP53SHZGHgVeG3KynAX2bVH
TsAD0kaf4Lc4UMYHNLr7xT9kgvHzvVKtxRuRX4evGnnlZRMedIP1PVvQG0WbfeJk6xTGAf95S+7A
hTOJWZOb5VOXEMsPhLqS89vqpN7TZ5HtnsSi8j9czWNsr4Fc+eQDJzSobfh+keDEsR8m5THjL9x8
d72iP+FST0KKeF5wxz56SK6kd0dsXlchrteyub5i8QS9B+1BLjHKsGVvfLXFRFAhmH8XP9JjfzVg
mu+LSWwOuI5oZKvxFdRJ5S05hJSma05wdNKRjoP4o+EaUImRF1sBtmUYiBtI7/XjtWBhrNKQrHYT
jvsSEF76BzdDUbfX+o8mWdpANPSch+JIJrBcKfzQlTrE5Ui6Lh6xJme7IbZbc8LfDRC3EPs0bh7z
Xsu+SAXEek9xv9kHPuVYp8tHAKkJUjpQPPRMA+bcLWse+ugLzX2prUxKwpsTxtbIyUBt6KegbUML
IGEmHvhiAZBvpnCBAmXCKgbN75A1Qh15NqPEtpfchDRJLMK+OGBbuMnbXERcJL/llNjUGONBYzTY
JpTYlYjbTmF6LacV+Rgv4YJPwK41GTzSkV7wOJ7JKbuuy4bn1rCXQEAGWXz6f2+vFqDkpJ8VwJC8
EL4W2bslZVX8f0JRjvB5NGw8nR+lABMuOYs8ODsgCqQZadsbcosQBaUWPWpp1rxF+ENI14P3wul5
WYuCN4zNXOpgCgnnORCYl3KcbVBVAHadEV7CgEtj/CJILm31xD4QYX37wlsH0LuzpF7XQzIK/rcY
DsB0PQIkNPMGkGm4d/vLKEJrHJXCaTOE+fb8tbLYyeEYFNBPkLf2TsxjLCyMXlP3X6a3eSPwWxia
7It70M7Fojy8tnAlw5y/585oa6QMGpScBoK5o567Cw54ULAuBAMhe9Mp8ASkuzdpALIf+rfNV+ES
iRjlkPFe/6quqTiqa32KjKwzaZAbrJhmNmPbd32d60//t8ChaG2932geLYEcSdnnvbWw+Bj/U9+1
qQZR10IKYyKKUaVt+2AXtlS8pXr+HRJClQqeZhfmzxhLcTH/5w8CpOtNBmcVAtQkLPE6eQznKfXg
lyvhd02TMo9WijwE/ajpNoZ+GBJscefFViTONfVTdiwpsd3CJYxtzX5cvv9JhuUhibsvtUa8sOUX
ha4H6uMVJvb/D5/Evu4+rOJTxi0wU0Wt6N5H+d18T9arE4cHNrqibICNEeqmY4THnZRqJPdIm8/L
sDMr9MWV8MFYnYvw/wPYHgLZtVhzP/DzncesNU49YsgsjvIf/fOnh97CANVo/xZeNp7qekdlNUgU
Q08nRywntJ1Y2FDS2C/05ARhTvvmwREwrRxbViDPb0iFwS3Kjos2Of0e+R5mKZ6Th3J4bvSgEo4K
xM8QlDVOeqF+pxhrq4VekmAMblmJw4jqq8mMpx8Snyi2JvQolBb3OE4ErUsvRWzM2nVmNSThNUR7
dYzJ0iOQ1px8TRARZafeYRKH8DkLrkNTWRpGo3ZBP2ti1lv2sqtyWf6EJ1Fge4TFvKE1+/LAhwNc
Svup4cB77iLk/IZ97UN/UaCLUhcOt1IpRGUaGbrnoHw3+sc8ROgZpN6AL2Le6lGKGnGwsja8Xryr
FRWvrl0mDfg/M+ifpsPL5XQkKqtJVnX5Xs8ySN9ZObj91RSpnCPoy1aVaSzlJxxMu6w0OHM8OXF7
xSOqurRkkGhHMmxaEf7DsrlcYznzR9poAQBwbCQaMiRYjBZm1fmOY/xXb1rYdnTpL44AJbjupVu7
ABwbIgvBlxH5gLaBom3LO3BitXIhJMNs9M0JZHQq0GR5dBvCYkt5SV2P/kqJgn15SFEToruVV/gn
369ewISII/fPClCqFgmzaC2XJfnDd63NKtnQFQahIxTUVCwEwDsUx7HHMDiGQs/7445yUFkiqaQ7
gPVSRbR4IOin6W/+yNdX5fhgCOh3SkJEqYB45Ibtf0O/39uY9n6uytkOkkdNWAGifLShsVWQ5CCM
ic3lGYK/DzFkvAK218jzknWY6u2gFNIJSP2yxoiF4ay0sNgsxOnGIVN9HzGM61v6ypC8W81lPhlH
3vA6bm1D9u8DZ5AO/XBEQcSu604svrzmVHt0YGztG7KHNvcDyOGyi5QPo4tKwk65JUCWWBXk4r6o
GRzDntIQgyCp9qJaBbMNcsVth7TGh/WElN0xXBV+qsKebee3P0G9vju0qtqvge8DxSAAG3Q9l6fV
a2jsrbTHF8r6b8S4HZaSJDEzyPIP1o+IYcG/+takXbfkumQTpkgKWneD7dQBr7ND8Bm1x1lqfdgy
PFKqo7QvsYsHKRzzfMhstqC5Sm5/a7zSnhTgLgtrW+v5hjsjO7Y/iRcsfxOSAumoUMyYI3QcmIHk
7IIt9mjHDitXrDWOlqLDEr8tFVCLra2oNZs197inqWGXJb4vc+CJZr2dIiwQpARmkszqrDbSvzfk
/VLZFBSQpkpQSClBkE8JiQtnDYrbuoJfSUeeY+PtsutsFuocjyY9DSlCv+3bycsQiGXNr7SU9N9Z
/sYTEaxdvUsAoXZ/qeIX+8L3GmAVP9aoOvtpOYTnj1RrcAQBKzcYoHwbcjVApKxj6WdPgGKmpLUb
EqJE0U8rHv/sZizymKG52+ufVvLWJUHfBZrVUCYtOsgBcRHPkrHbq80S+vLX3Rlr4iEHtpS8uoRs
g/0QlGePq5V2AeLbX2qvoi6I15nsNQ3kj7UXb+8aoCiurXiAb7KHgRGNv3GuvPjPTiiLsXxymwZT
Vzum7JFmwkUcbhYdEPTWoytv3eWvlCscFOBEqNWT6MjaHAD1UgaUMjN3kPphUQrff0EawmhLesVl
LoVugo4oEG+Q1rjPOFcpkg6LjReDqVCU62IiOXmeI01uDQRDWiETLtTKr1H8MZklQxYUQ+NvSoRb
OPjhlSg8U450xuRzpHZUPY3sCoT4IO5fEECP2fqR0dUO44FslbYLNTXNcoeaHEIMc8kyA/ZYzmQl
ZRQAvjvjg15GVR5kN/3yIqP5la6gjr5/e8FlR9l0st9F85CY8jJlC9HankBi3ZJRyGBvNVa5DBp3
MMwfrsnD32dr4jg2/GAHl596fcMbm2y6Q+gqS5B1gyzLfWZaKX7jyKHKOOLeCD9yDTvgc7aQIjAo
IMZde1GY0ZVpmzmWLiEP8Bj8mRTsCQOCGq5nrs49cWv0fF/VKFcre3UbfDiqeYXDGrO7DMpZApkJ
TBvNx4p5MoONVjWpuQL8YMqT1T2Tbj+ImsrqHMM2AkAWKoJyu/ZMsmzZ69Ee/jFCFx+TcEYdcBtP
4qKKYS3G8hCWK4HaGCWjNJRzA1qXgxPUlgMRkmgSJvcJ2yZ+D0TLCvtYoM+9ITbWBKkfGiKBSwNp
wqYNXkpP6y1nyWhUQfNkE3C5kD9iyksHYqqTCz7BcYN/tCHle1NmTrqhCzmveEM/MlAem0e5qOqx
2aQwuyYsaB/CE97DdWnRtrfC+U8wgm9YZThns1oNcFgxQoFs9eq9fjVUBDwT9IQUQO8y+FOUhASr
s9W5A7qJGIu5GfXAbFdZ8I35MEOZ6FPGsWsWWbDYtBxPbH/LZrXHZp0HZbgF/JTlp4XCpuPm4F73
F5XX7ZMQpgMkD/1spVTfs761hF8WtAuV2ej36pX3lcWFkxKJmVR1MIj5GW2iOMoOL2RbgiAuNCIE
JoidYzKm35iDFUh1g3XnLwNhgk66fLKcS7AOvJ0/MPtwDR8KmZ/cit8ffXswALiMm68TVJppelC7
GXOkSL1e61zy7vTmtK8NgXi+BoKm78/AYg+upNMndl+ueaRhUO2VtHI4ZwVvkemwtNLoFUAb6kXI
zqvVzh8/IV0mc+zvPUL81ixEte9z0yAcpEfduwQ/GZljG9neu2Z9Dj5XkKjAkJHy483MmuZ4NyVO
pRRPjeSpteZ8Y328T14dGriRt3zo82y3nId+zAnwVFCCpTZzMKD4EENIHqe+JheGQMZi0qFGFvyB
gDUTkPi4P11Ru6R4lHU2AgYLl5dUk29IVukOCCpSme7sI7hmh7x+bSE2IfdEkaq4Xecucc0/cATT
Uum/NJCALyjVCM/HjS1GaQHjv0KW0irlM9MyuZznqLv6oYo2vmcOy1krJPTfPGVVlBQHjR9ai8Pt
pN00Gddn985wk4aAeiUHhWd0ytQSK4a8fPNpl8cQFWCjpOdRPMXAXYhojH3GdlOw6XPZXG/fMIoA
YRD1HxyCYXkedSCrQZpPWt1S0hh7iTpja65+uVWFSLe9gACH7VT4SZBK8Wo5gcbU9+o3nlMTYxmQ
GdcU18B9ynSL9lpZclsdlmMDaUt175ULZWfcMmbigkLgDcv9Uv1YtE26HS7FvITEdB0U+5bqaPD9
nrrZH5Lvyqawb3JixCk3erD4+Q5Ndekvh0D8GqG3TZiwf7R9aNoGUd+ZlNqh986Dzk7WDPER6ohV
V2tLXK/kW35GIcl1/KoJIK4tqVrVI3eoVqRHxMcdwliQxChBaJkwXzHUr3VsUJUz2SnOy+BHufNR
+930BmbNZH9ZYhKSMqYJGvllbCoihwfQkToLy4t9cK1+lYhHr7QkhGKKDgJ40cg/LhShNPwXL3q1
iqS5fq+yKDcGt0ntXOwY0Omm1LOSrVK3aDC5ft/Ow3QxMZnAMlwtJFyPXkod2JtCk5WECT5i0c4Z
Y3D+QUaOcnBEq2KSu423ee2+vT94Mu2BvpiLzEZBYeUqoKyIUB0Yo/FPsaw10YDshcwQrrurcQ7Z
vvD4uE6lk/UiWLS+P2LEtVHCVnfIryQ/07wIBh0X2hUIX0w/ireNi8/9s/VSB557YIz8SOaKkjPm
hYSvLJcI4OnPCdZEWp0JtvaYazqMYBfkxdfRBI+IofklHabSF613iXHmRs71qr6o7NZRcgExmlhS
G7E2wPda2+uB3oAn5F1vqIYJPx4Dl9uXd3HO6xaRyMcBsh/XB/9TxBc/w8Ue1Mkh+ARcCSfvMwg2
srYJvmcZ1Il0WNM6uZEiKcTpqfhGiUiDA1uI0k30S+Lmq195I58rDhK2BvCr7t0EL4nJCSod7qD5
nlbDvqIkDge2W4WmhneBllrfOUrJ39EY68x2sZBvFZIGAGLolb5hXrum5hut6j2nDiq6lzTPiSj2
0pS+Sqyh8tkqD1XQ9WX0DZBuBQ5QlaqFkgBRzehEtw5IVwkC4sA0SJOW4f6X8oF9bbrhaEkFGeEd
Rrs13JRJOC/pkOyGWyVcHrKuYfTQQ+QjZMJ+3pcnGFX2l5YYW8uFNtP+sqc2E4IgiEjg9W4OmfXS
8IfbQNhLNRpSIeY1j8eD0HX8I8S7r1+IOA==
`pragma protect end_protected

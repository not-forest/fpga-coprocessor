`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RgFFX6KsFsrBrIwaYS6de2rg69iEEqAb3IFX58wTkNfivNEAcBLIk00IQHIouHui
LHuVcYfy4wxL4LnbSveM+Jqq+Y54F3eljiNyK6ZTYRjG4LL7Nc/Ouhue+bH/YMbt
9f1oiqx3UU7sldxJGoHrHlh7hzCyAKHf+6QBGciJlRs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6496)
VtT93CqDQDnkZt7rhxC7SriaLE2wygY4YRwbrYNkIvBdw8NHV0JH5XMRAfxAT5gg
NRmFU5TaIzf+DA2YnpQugvZJxVqxfpIuo53aMowYMqt4XNeKdZDuEwSsrkNlRA6d
Rh3CQthXjzDmo0HefaCqyU8OWjdYUjm0FAd/Arw6PgpBkQUsvKeWMpUQQ+S/ZXKa
RwvDlE5hoyxYzfk4x0dPhT33qDGDbzYOxT+yMy2trvHJzmpypPrbDJk/VFOYdMQU
fPjYfMwemFbaDAJYNKE8WTyION5VtZcbU/ylIpx0NQQ9+jkg9o8Oz+KOdtQczrWW
k68Soy3Ixp7bUXTpUjWNm20ALkRiBqgbLX8DFsoWx6gRFtwtbju2t1MDyDKTFgiC
Fq3viWDWgT/hk6AaoAXElh37MPDST+nkPJV8TltD0TTKMNLwRnbDWWmGzj5/QlKu
9PLoZD1X2wBycgZjRzQ0EjUFF02wCNYpR3h1vEXWr0oikmO4IrZW0irjRFPWyuIH
sPk6mWhuzeion+GL37HzeX0uOIyzQaxEPRZSctNtvlbG1d0oi5UgNjESMGQpMFcx
w75uFStTXkeUniFF+WaYeIStqogjYE9qVpZ/G2lPq7HDhxvbjpoG5ITlw5AbP9AV
WQaOyz48NKLf6QkmazmdufrCeTNXu574ZJVSIGMOPnKrGhzi12b+eemdXXfZXjK/
e5dV3EEj75y06Ckj3ldNpRmoZcg4PTHn6cpO+U+snsR7iuSX8koczZVHqcNhCA8q
2gBtnW+QFtC0OxxbPETma06VTgvh7Pwou4PCNSXZn+U7MLPxEKYqw6b+9tpVs7qj
towNR/tZC4cKSShBCkDvZoucVKD7rshAAX5Yl81VmbnaxJunWgfesuUN+TlUf7Ro
6G+XAtqv3GD+5BnocHwBGeSOPy+DOHwW2GqQ0laYpA2fPlKEZFEZ6wmlwGDt76AF
4a+fR+BzVFbEEA+5Q/RCRc86UwA5myBe/iHo094LXGM79tAxey7QSvC4z3pq2d39
zks2IrDVwTBf9d0t7rla/5xOKmhImFXRZSKVv77E0YeyFbghG1qgrlXKRtO2S2JK
3p372dYP56U4jA9AOIbWIoKB67Zwhew6rtolEoHdAlSZ06xjISjAiLa5JtCXA4Ib
o+XGTBOuHs6+VfJ8nCuUKzxqOedk2tJn5oBwMCJVE1WSr9MFA8/02D+UIIKPvBAV
BuyYaq6Ixp9aL5UcVDSpESRcakHkycCVNaf2TVQi8/rHCy+ESDHtuspC4PtOFVkT
mAGqn+PGdzhlfqf6zdH79/AvaKo8EQf2k4rVrf+FbTH3CNLKyoHTPrK+6M7h6gFT
4eXKMQdXDcfMWMsfG8HyErgCcDJfWmfNTTqCiBchwrw6RF8LKFCqjd8wuKTwEBGR
+lGAcpv3yg+BxMSxelTpYABzTsvWx29JsYP8B54nK9551JEPJjGCfgYjYBVWSM6W
GVzEidsn0x7rBsNxiOJDguL5wY1HwQjjJlofFTYzCSTVJBkf/ocU/8I1E+Mp+aBe
56it2XEkYoWEMOAb63KIrLUxyMHncIP16ZCwvv9gVRO+G0VpyHxoWE2OgBwx+cjc
hdnjHyRNutn1gZi6JlPb3CztvuVW/7rzYfLRQTWKXSFsN1RNLT0A1eEISq68BJKt
UTkCWgCaZ7zyDwY0B+e0ghNK/MuFLCCHuQ+EIV8ktzH3GQMBsZ67EIfEBUPaHvhl
FGcmv6vDtB0UV8gkHkr+Cq35KFfN+SU9t+jy6KEKExwmkqqWXTB1Gc6DOocMQpoi
IKO0KuYK1/vchi44s5Preq9ICb6Valrt6aqY/0C3KY1iVXcmaGMuJlOQJmRgJ1jw
i046xzcfV8FZfDMyh/gx4qq55jz2VHWAwjAf9P9fp+OyAztgpYDNHDfI6ZKZYmEA
zP9vXS7J2QZOgOAb3GotXCYxs8LN45pYfwmtNHDsbnsQGNjiVipHgx+7iJ7pjy4u
pU7nklNVEXpas04sUxm7K2t7F2xCEbLqXzEKg3S3OBn4+t0Bsuh+/IpiN6+t6w1M
u5AAc/d8jQKHmdkRcCLQvMUibx5o9I5/jtxFT+sQhmRBrR7kNXQyaKgwdh1f+txQ
bpJBkTfjx5xwDxu74lojUIxEKyWY44kiZ8ZqdGFHdibHEfSeRX79dYHMZH96Pa2C
Yc4brBlAeOshnrF4GPKt1MdTDuBuB1jC2hFOFlVFVc+Z6yEHcEn7ZIoM20QEvoPI
SQkUXHDkyD/lrigZd7pcJF70HjXieplscTHyV2bbsvCqDowWLmjVaMJ2DiWC0oOC
5JV4beVug8rO0vHHoFeJqMSBCH7VPTefpuZNzYf1BSl1cUvh0Rl5QsbDs/C+SG8N
XztwqTqWGlKL7HjWEHX5c9UikYkXOhzdr2F176L6PoxzrRH2AePC+JfHVUS5Kkvv
Pzx/HeEGAWaBZiYNMlWgAIGk4Z1Tg9OSp1XRYjgjNrnsMIVEcRavfBYc1nJAdaL7
yxpCCZCIP4suJ2qIFZHWugIrhaTb1FBreaYmM2Q26YMcffX96hiGeLq3yAgJx1fs
zAz7RLydG6HdfDWy0MkKLH1CG/Ohhn8Mk2UrhrsSLjK44P2H2tW3Rqxb97BlA7i/
j2yiaJtTZVx60ovq8jxySOJfZYQI2fYSiVGr3ByOvy8ov0zRccRy1IuKhhyk7S1B
nbDZ9p9raf84s++BCPnNaNbYQRQsXjvtGMUaTKKoXvBSNa4vX5XSy996fwvOmTC6
4LutGTKmxkAP1XrOxnInWBRdwxHRE6iYwmlIbY00iLRCpWbDeZNPk9ILc6Rzzq6M
TjuuJVVW/FALVgNxTl3rFufW+LDg9edf+xBGHzcSU1ewQ2u44UY/OdneUeeKsyRq
loOM2uAP2hQf6my4keGd4aJ8fkwPQVpEqSeRzYrxuxEFvP1bKknXKu4XlIxbTEN/
RzEDzUNAsrLMvWkzkRC1O4dpTRnVXoGeGXSUN9KKVLfm0W85snYnAWXPQfl0ej/6
9V2Eu3DwCNWMOmdTKY4m9/DZon4WK6ksT+crRD7vi+bpnY+2SPIfPlataE7wRoB/
mQtBs1yxLM2zrRRqq2vFkOOUmaZVrHbnrfD9KrBwA7uYj8pOUxl+Wcrbt/kYfUUX
ZO0W28rZaT1IoDZdywsMORkiKC3izpJsoVpzpNmJzGyWQvykpTZ+OQXuO0AGMmHE
krayMHozcYp8HyFy6CoM086WpINi5h35hCcg/4m+bHRUsEsWohDIP9gt5AGReMeM
lVh033NG+jZ+Os/vcMx2sPKBJFJSex1lcQTo788vyvWdD3c+OdrbBBxy3QebLfHN
ZuxgmPCoBAwvH6oGGoqLGf2G0DSAhREiJClsaQewvBFJ1gE+o9JZRVB7I1e7jGPA
o5GlrnNHPBUE8UKz3M5ymb9iZoa5uHWptjxEAHsNzarRusjnuKmEGMf7RSBDM5nN
s2HRE3ZMFDVZ34MCJnVHMctHmQ7PCR6nol6Qgv6eZBXz2ds4wRDMXhb5evR73B++
f0GLpCgCgq3q0vB2Y6H9z5sakNgkgcs9lVPEHkIJRoTo2TiOfAy/80paAfzvPumO
X2kcdvVZSq7EVh61np/qBy863YJSdy+wLCR80rs5sKjO67S71rH5LT2FJKl6lfn4
DzZJ7lLqbVhPL5pr9NTRI1it9ToGbw7d6K7wc7oDbm5xgeemXAT0w4HyCumJLyZP
HLLXPfWjJNvEU8oLReiVPSQ5Iy7jZIAkaiBpOFGdVYGqFnFOhj080SlKH8AxFofE
j+UzaGu5yHjlLQUD2RgPCyEb4leTa1YWlenmCCK+uudQi/2PaIzv+x/41kNF3LSS
+JJ9lWpqjUj2qHOVLigA6biSyJWlHyj8E2M+pAeyKRQDcdST0Kw5unV72qjRg/dp
piNtiXbWVHsyAq9m2s9e0qGSXSuoCt0aB8vuQ33QzthlmtHBjJ/Ye5Doo0WHdwXI
8vZhMy4CaSfKbIm7PLUI4291VzbLj7dkRvnDuw/S7CAqsXAbjB9CbFo1UtKU+0+Z
qUS8nNG/dyxE3NhfRjT7SgPpt0DcX/8+tk5qoqN46WGAhhUG6isrpSx0ANCevKm/
iKE2oKwfWVjDwbWQwc++W3WUhgq755m+A9fdlMVXHucvYfjsXortumINwyEYFo56
Y2CBxRa+AWHKMbYCASzDeXEzQh0Za5NfwS646Nh07lOFnH91Y4/+TJs9YHcHRn9X
RPHdiHzR2FD1PXTPu3IHv/cBwTKCFlRixae9eZUIR5u+NzZjC2xg7KGO3PvCTe/I
35R0KbligL003wcwzSSnOPPdZFsIemNlvV0iWwc9mc3uQWjr6aeTHlIVR6pnNoIk
cIcAByLzAXUDYmzv4j5DtGk/7cTiY+fTQF+88BJNjktQbxd20zNyDPk6ZwspApJw
shsj4FwMTPQx7m+y1bkCqmLpzpGXvUFmKUau4mKZ0/XjTmQr/rmJ5N1lBXZN0eKB
O+lsm7owzFAEY8eaekAkJANmKhM+nGiKr5L/HbO3VPkvr3/xCHoyQCAcVVyNd9tg
51FjEm25zNOKmZUm06J/Q8xgsHTA/wzE0WtThGc8g+TLGZxmwAlPY5rGPdofhyLn
BuyBPITBGj8P5k9UluK7shTVkRQMcpV+SMEhI4Ja3rlK6WFiSBg3lvWsOeyNQalg
s+JTAS60Ci+2VsN5caJMghfGk3kw3kU4ksry9t06r/KLubbqeHZu+/jvOCMpKQqW
KGavjjyMvejW5OU7YmUJ9VclKdfK4xp+a8SqupDZvRaQABcSdADJ4zTZM1bCy6Rw
Vo6VZaWqme//Xr6poYFZ6Pyx0CN/JMaIaQQP3ZYgsuHr/cQfoBNuJOGT0yGAXX9q
vNHpxQByh9Z7CTUV6O6oyB9tezEzinlbUKCWM/VsY36HKqDSc7T/C6q/026wWUHk
8v+HIk6Z0oAW206ZNmRPHh1dAkGO1os/fivv/9p/42oBLrgtziOcMUIQsoeRzJSC
vDMxO8/JzyzxIWploNZCXkf/ikIEo/aMvdtPBRodokUbBHEQfxrtdZqRoGIAELk8
jtv94YJJMWAqufTNxvGyeDMM9WfXrDUwMPtTWJXjxcc6PO8qmaZvNKv2bjHAXPC2
huiCComd9d96PacrVTgKckUIuJlYsoAQLMmXceSVWsHxMrpc9Lo/43FnLcMeMY17
wA88Qoojv+N+AeEWbHQfUilDTuVW4VUnLqMhJ37p9XmBedFIBtmQqfrO1YUvBFZg
uxEVnKi6T40/DF5DZye9g1Utgs6QGYDyickXhL1Cj5W+Oj037pIJVSOl812UoP1X
42pcSqGyVgdtG0p/v7oZ1vxkpJ3bt1VTtBEsTSQd2VMfVIEjm+ExZNEUAI+aVgPk
2fRns/ntakjZnnElxPCZ+VPiXGFSvlnserUxFzoYFdZatsFlcuzRlfhnzvDJIcbo
fw/vDmLOJAyqOeqr0OlHD7qWtlkZcdzSESjaXSZs72xgbmGzHD39lAsqDgAQffYX
RKmGkCsSUyz7DW/wbDzB2Yg85MimhPZyJbthWzs/aaolYJcf6Li9MtKCvyMV713N
7t2rTe4VmmOOXsak4UbiWt1B/NTpYUB/gkC6js6oSQ6Vhoqv1PJ8ubPygzHqOz5w
X91iELIymJ5ERJmD1NGcya62vQ7plyiVZ2XkTmcqyujqqq9J/HW8wgnIXTLwM9Ot
O9rDXbcge6MVfB64MYfEnvXdpC9zhr/fL6iiX2TU9+/5jSNhMUrEN7L4k7Ybi4X/
7S3nqrBACNG4iff/5Bz1UTKgrLBvELe4m4IhQHCXKJY+/ndygbFlxqgpEp0jT7PU
bu2Ud/ynEN787J+Q+Syqee2IdIo8Q9ixBu6zyVOefNyecFM2gbayuyHWwRQkcFLg
kLg6PTikk5bAAufa/eh1LrNwPeBdMC8kOrjmcSzLCUrNcFQdTw7YNmzxgU+jTP6p
cagJZS86mnC2KN+YrreKskBC7Qd5roRKvlhPopSPzqz7NUcpxAR5wXFNTzc1/Zvi
R3kObdmsobbRkvjxgk5WlF7I31WGaaxu5UJ3+QHMWDLWW5Q9ZlgQ5YSAkSJ1tEoq
vWbaYK1BX4Xusoq5FiZwJbMsFAmRq6WhQbEzTVWnGoJb4lx1ua+2wmZD5+UrwzSy
GCEUHh2m8olFdT/U3CjCej4kWktibAa781RMA9y7ZnKMewg6ac+nznqX0U2LIdFA
IhCAakNZs0UG+sg/BkXLvNQX0A5sKjWl4THP0X/0wDeJ9+VoDGcE+AuP0ISaP5W7
FHL9n+/fFQh0nHlfjOg+7pwJ4oqeKyLQ2iGthKYV1BsCo5n6Q/HEBM/fcu334zQJ
S0aisgoPfu186Z5m1P+E435GDdGUMTgxYIiqwjWqRVod9d8s+qgorCmEeQnyzZc6
HxEqJpC9rCG6d3Z40dKHQZ1F7jHSni7w03ehB4DZiTBVJjK1xtlcI+6GeASknmmF
9xo6q8DOmzINOPtp2EJk6DSqvgwYFrnzpXRF7MuonEExhVNF/WZa1YQPP9pwYa+i
CkLMasmNKdk0XQxnhS59u8eCt5ChF17oTF9IECPcHML7Ee2JdVgvcKPdeeqH8zd4
VxFpy435XTeAMAUiILaIw+ng6XGqgeUlxrFIx0/CWM/B486iO0dpJS3gfJ1NBU2X
WiaiHVIcvBUoYcTkhFQs+Y8bT6voh/QShXN02Hy5s/o6UzIzXIDU7ozKlnCKGADz
SXBqjYwC2By9Gdv8AJtAz0uflF2MBT7puFQmf38EDyPmTJi17rsSmnHcf7XkMncu
DSSrbEkELFuf0XWq9UaBlCb+irDBA1VBuKGO6YMZAyzjpg6V8ab/aJWMq8MyPXKP
QJntd1cZJ8m95tturbJWuh3lnEmX7TY8wjKJuNwlcNxEELiItF4Aql/IceQgXH/r
fQoCQt/s5xwZcw6VfmJhUftYONJYwEPnAtAsT2fpuJwF5c5hi8MzgvsnRN417Tza
C8PSK1DR3CtZNHvwGZIyplinVkmJIFH7gC5/2UshGwSDiDdS4vEzFYqCtdBeh0u7
43ahsWf+nael1vghzMK7iwCDcptLUoIOd3Z8fDkNHpcZBJ/q0sf6sVemq86nm3aA
3CHkIOwzne2Th8uZEDZ2iQ1WAsIg+ybWBgOvc4BCC7Z6BDKWiMwzIF7eBP8wVE7V
TxeqV6kWzg3q1Rs3VotTeW6Ej5RIscYxEvgZ831xY550YvInCBHpWu3Pk+RaF+1k
Q0bvShvrd8R8eEIs/IS83VHa7bQOCimQI0rmntTXgEHl1FgoCHDDRaJ2E6dd6LDL
VuNi6oVZahUhDv3ybpeZGE/782KJhcttczQF2zWtvsaiwy2i2qbvQgp8Dd+QPM7b
27raDcfwDl4cDPiT2lyhvL9yxsu+P5Tcgzj0v3hWAFwYUc35MyPB8BBVo9/qYo9N
KBrbIYti36nJI//lklxOvy6yoC/UR431j+BA+woETQm4/RjQ9L+h/LgYXGHV2lQg
FcPqhAFEuCbTytPh1gjqbqDmHLFNWttEvVpSEiSBou0mmr6t2O2cZpuQoUzt7a0q
Ixst9AHIYjn2x3cB3EFvuINIGzLDDIvtTx3zTUyaSOkkvhIbVeGtJYJ64f7RyjRg
Rpr6+yFf+16cXHGDh6YefCegLbaSSLOERzvc1EGgcgfoxVm5xj2JSEV1+QkAMC5n
GI/IPv8yQko/bmAxiA/aXo6uCbP5P3YPLZR/a48dCwqE0IntwSdXj2CNw5KI+ZLf
IjFPNtyly78T/7WJdVgDwchTYb8cTWwkl/cJYOWHZw4hsHl4cVsBuTPlWEWifObt
gSQdtAuxsR2OImXSSm2GC+TDzLm1RU6HERZ+Y/F+USmAbL1Stfljf7DYs9yPRATv
x8kwOEc0LRZ4OpwryFt06QQiUg8mnZx+Ng0Q+HAXqdxd7T2zkm5qM0J2Fep+8DHo
ORMaAu4brUBYp7bwVWmvQigQ6K8314LfA21NjkQ78NsZty/cMDwn8zw/uCKuW9Fx
p/l8Aibkiuusi9fkHerXAkDuCprj2gpFDbrf6j5fsPCPEahpl4DhFJl0Zqiu7RKp
IpmYv0Dd1I9Gp5Hcc6OcuIr7kX2b9qXjCYRjkziy7gDXqENTxZfWcR4Qd+4wvSnT
WTXrsPFlUKgcI0GA008b5fDdTPliEt6gLKOYZBrXU8eg42JJ7ng47LMmTfd5gykK
UpsSksBwnjygq7We9oTs/n4vEszEvn/O3cl57y1ymQ5EIdBPomeUJq7aFq4XQBXi
eBisRFcGnjS9S6fQCtIspC4f/m4sVxP174SU3mqtjCNxmDlNwWVLkrzLesZ6EM4E
RGNXRAezOvuDJHAO0x3+tyl2vtxfqZzMYAJyjli9tcPDJlaDpI4GKbG3m4kjq4fs
Wdyus3xSKVEWlW+wq76KV3tkxBhA+Dj8c/bWen77lY2z+oX+1/z9Qmbhq1MXjFq/
akEHyQfxf6V4pQOReDlVU1YtzJgwjxksYr++/jX4rwILV5M5Yx/Ot0BhRjfsTk7z
QZ/comTkFLTpNuLRhvN+oWZFspBPWlwqxEq010DhU1dAXITUpR2CtVKbGxXhVsam
p1ubb6FP4fa9WWL9trpy2deKtdus4fLKKk6TK0qbHhHm7uSbm1FW4nq/aItxrbtl
VghF8B2AwqohxSRa2LS8xQ==
`pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
FhYUGhJyHsZF/12njejtBlfEZlEnXEa40QvUiCoAllFrvwdI/ibg5uwKA1j4C4Xn
9D01wM+ckJSyPOYw1F9YzEEc5l56XRsOUSiNhUCe2Pkv5tovKVm3o1FtC+1o27RE
T4Q2sBKbiRSUwg6BvkhtdrMMct3693bhtP5cn6kCXbY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12128)
j9RqAWzFqw7NBb0wumbZSLfdopTCKoXINHPQG6FaCP9Qq4TsR/XtX7bSL9js+55P
zfSVZnwYCrJIy+MbsFcA3Syr352colhsBg7lLhpfYl0jtevRtRJyhKANQsIyYlrV
JjutFNi6pmRWjTkdLkjBZdMpHIHwRQV8SbxgRzp2iGVoN3Gp+vJSdtWIrxtZQn/1
K4gLGiyxwoNi0OuJeb0R6SzcOZ/6bmKfsOIQ+CcRBoEz4xpvrR7LNounV18F1DSA
xD+0fF1IBYtCeswV8LoDhIka9mb9P24uwwF8kMGKjKA80TGlHlQHN3jC3zsYASkw
PBbm/A/oJu6E5pM+Ga1tbq7t8eL8aLxwUuqsk5P0nzNDNLAVFz/v4JHgDO8HZvXm
jYIRoWFcRdAHnpNANY76BwP57cm7e2T6yyI6jpevuXxRvDOn/zc0bJimv84GAciF
10nc0/iZU3ycWLgvILUhnoQinqaAU3xiclLbAQGDGFxvZDN7jvIPjaP2S88b4wOr
3T8XLOATsqKTCZVjuu50DdTIVY2RZrzhKHcSCTUucadaFbPl3RBfE5CQcRY8TfzQ
Bh5M8xCIcU+v22HNzFXmnHTWVmVMzA2FNGR1qIkW03uPW6cXzVz9oDAmgA0WWo9/
njSeeEdu2oNF1/9XU2eDhXzp/020HFnQ9iiMXaCrVQwR2hHlxL50T6leSPNnNKiG
f6tJQlOKi8t+jlNvepaadTQdrq+Vxs+59vPw8dAHU8K+dY9tIW8Cc6TZuXd6Y08a
IRmzUW9qWisOzzcR3MtD6eaTmge9fRkHX9QumVlNvzvXl20q06Zm3j1q5cnrIatg
YDx9hOHfye3PhSbDd7j0oMJUohr8/XyO793QpJZ3juOj/RQOJHCp+R9O8NNIUK/4
eoCs4djW0fFng9x1uBhTUxyah2AUJYg88SKnKa5bh7icGXyoWmb+LvtL1nfsuPXe
X/sIEJPirDG8bh/kALQLiSJhQUL8LKOu/QLk4L3c0AgC9uzMxR1DXKsXXlxo8ObR
obh0I+ZdgalJ2rvHwSh1G0BauS1dEFvMSTlOvt40pH5O1ueqxI2+wPElVnyL36v+
XBVp2Fb08V/MzWOVh9c5wTyT4AUFLQh9O6CB4GCNMy2tOmFbyN0X7/GbQn1RiiQA
GfK03MIicDWW6D0VMNXopArOeuiodSHMwTeWJsmbeS7cJakiyMuu6+EbYpyyB3RR
YuDdOGV+/UIxOrO0hcCUltbecn+0HlbZls3nQN2DVZ5dSubLcpfUkXjnChzA+MtY
OfzUeWyY50DPFyEVYj5M/899ONL3GVTm9SfSORmM4ufcu5fsYbkdecPhoS6e60Vz
hWhWXlvbBItlTkNfq858hbWVe+5yanSWTT8lEJPPyY4Uap2v4tlGeJMkCp7sR/LS
nwXpgW8FSUmLRYB4BuGvZId9tWbQjzp8BCieyEGlTUT065jC4Nh7jchklHeqwvur
oZHDAhdLtUQJjMPk+FMYlgE10wO0eOtUzy1yYckLBskgQj681vd8jopdsR3fOiIG
mYVm0oZMJuolQ1xJVt3PnVhWLKxCw+YcghtAvAPLrlNFm9BS1qzfat7y3pDE1dHK
Ba3gy/589HdBbIUqWUd2lPBp//D7+3slIPU7n6tefso33UWrI4/gBShlRNblLabU
PPLh20VukZVnwtBmWa+bN1i5Y4aei537xlfnKAnP514kn5dMPlry3Qvnu5gGJw7a
EHQaRXkcc60Mhd+3In2YY1YKJUBJ8NsvCKi1vPzdQi+jY0OQhcv2fiEshmKpiMML
STViH1iNc+1IeBh+JKCQkNzCFfjtQQfpN2zqTIq30nwbgTMH78iBQwsMht3/CGTB
smWMpMHd9FgLv3Bx+UQuVnm/zH/oWiMXrOld4XaPIe1mi/j0BKiZU9BdYnmTZIwv
eZmp3TgBapyNkVS70PGAJ9tTkLVtkCrB4rSf2djwrpzQpcYVlG4ffjX2HaSZj7HO
fqdcUVKtlRzCjYI+pupX2MkvcUdv5RhXaK0CqjrttVGcVCeVPNJwnJvYHLopqum6
WiLiNjM7vVWb7qCFNcxfTQcpEkSfjg25Rz/FaWWjltnvc4re3CNUMtGsQC42w3Wc
wkb8nj3HJ069tJ4olg9UhJVCsg37DVzKJSWH9zGo+FO6smquWCQbPRE8/gv1eM8n
pf7U7cUct9xBjWUFi3U6YLFOkLQapDezRlQcY2hV/ZkGk1gfjXYgViLG2m1/qLEI
WSfNz8usQujiSTQM7ufQpXmHh5ZFgYlhFIXaEMfrLrmoyuNiDUXfk8fCPh+mvVon
mH4p9J2NN8JDdMQ9y5Cd/6lLm7X2sUpArAs1Pl/Bk9hV7kcsPCl+v4lPu5EQcd7R
4g05/7ddEsAfQ6vHwExFpk1uqgB+5uBEABHbPgF7vrRVhHAfpHpN4dgJqqYHbVLA
iWeDtwOepl2R5OX6o33Xfgc41EJVnl/nyhgaaFLLgNVN5XWWrdGojiJ37/JRL2Qd
ddHWVGAo8sgJMyEUCPsIyA8FPvXgvwsGeGkcZIyMukobP10E3hV3F3dmXey4P933
lCOkTujiwvHWjxNM/L5UZcPELcLs4ap8zWrpAHunKmdgC6ZQ4g0vt/wrK5+yUSfJ
0QC+Q3qLABZ1OWBItcDPJV/3hYEPOkTu86U+mp5SDt0i4QC8hQ87WxeL4iOfvR8a
37RstMm9EGCPT+l7TPDR0dkGbsnu3YhVkGv0bmopIa849MWxXNZaIQaEqkeKKrmZ
qKi5CmaS+LKlCWULgzl5E7qYqt1JhpABwAdmWJoif6bjkXEYsorSFmLD9GqNrLDI
BOOoNM6J8cw8sX7Bi7VEHzh8b24uVPcIFIZA8GYzBAk0o9muVrUdzupMeiZaS9E6
4hIixlred0SiDA9lJ07/oGyYNYRwfP7WF+6xyH8t1ZsW1yrP0vwzhczjYTkRh7La
kn7lZw3t3oFc5tAYRrrdjuvhbhMs91Sk5pVcHLJ1v3hk10P1rFMGr2V4AaMSJ+py
gBIO20xP9FKqRHXm+EeUPYSpSJazrSeKpUY84aXIzyfQcTOQCgLDtQ/xk2Mj+Zsq
jCx16G0HFuQ+xRgTyxx05il8ZzcWpBnjKxXRZZ4B61qK2TbrJlGQ9os5X7OLPX5Y
EjafYsoM/7mAObkTw6s0bBp2tfRqIe21TBT5MviekhI3oSqYvpu0MJDSl9EvNjcN
pcbEdD5U6dhI5uhcmNsx7xrywqRIG7PsrykFU6GoZNOBuumNXMjPH3oUnrnoV/rt
eCSU+TVHuOaT2OhmJ8pCrzJxhTpoNnAzmdKwVCcbTNZpQ1hxiTvtSt4JD5xUuwg3
b3QocDw5otmdt7qRM19FlkNTo3DrzeDkrVN0l2hH13q4hnwzVh4N5rsLrXQ0s8GU
ECWC47fPvBaPnuDL5HuRccQtgFFPuNSA2A4D7dEwyY0TTYSCGIYo+8/W+bfgzQg9
UD0UswHznAtCyh+C+58ULOvKEIaOO8KwELLQGKeQK6qsJalw4vseLRKgjD3t4YbL
4CFAu3wvfgEzxfzRyYKK9B4sJVZae+zbiEPe0obna4z/V6KG5KIYLaubqj5H8J9D
tMfXVFLz38WdKFD58Cy2E5JtI/jSefpp7gfvZWVBQrlQABwGNFIMyLDNwVBtfqwQ
qUUldm9GKaWzHhAiti/SU0TsZgIjZlemeZyTV2gyizw4ZfVxHOrBaZ244I6zzsVd
ly65KeZjaRVEeRvIZlms/MiKDzot8AW6NvFFkBrqeEYdNrjWEJY6uY7vOVLenE6w
ZFGuVh7ZP11hJlZsIXxP9ywH8Ujo62yaC5G+guC2cStctzCLklYIN2l8iBREO21D
mhr7WsfeUYdAk7s+XmYO2Yh77X1PMtfJXvL8hrGFfyoxfukgojKl0S63dH8shAVG
V0cI7AF5cpf2dxypYogcJEHIY11pYUYrpcXgbf6CRzBhXw8UXvTcyTFgAgZAj49E
T3x6zPB11RubxSErTMtnYeVG9+h9DW5dRJIhwyD/d5rjY/A9u1J2/HNu+64f71gQ
MSgqczJRu2XKUSCR56WQV7uwZ7yid65Ls3KeBz2WiP3fVba8QpvneB5wiXvuZjs0
1mj4l2fJanGWm7tLwMTOpoP4E8CsqXXRu9XT4uBvVyuHvTlKBXviYY7BgqdDnYnf
NvOg4c3ivXHBpo/brCiqw9fZ0lNSv484oFmNZMlVJWn1hK7k6kxFX4Um75jN1Kya
M5V7+xNAZqiYWNXYqAuiQjvF0IqHbfp3rGe4P+iLg7U6NRaQIWZjgnaNkbCFm/tv
E/fEDLmi7vg+LIKPqOzk9uiYbXTlWqSYoyeyqBN6L9v3N6KixhRO0G3Y29S2dz68
dkhbZwVbFsmU6e0QwsPv3aP9Ob33RMYqDU+bGTkkn8y+4kW3hsubHwc+bBy/W1Mh
aV0thpveoA4p2P/aEZawxO7tO8VwYMWnek0+MS2EQFAmZ529DLk8WxsqEYV4lNkh
Xya7nqjp6ztdczf9hQUeGhXpE3CNC7x0eG0sjaYE7XBW7NxqrvH4sKNyxQC1TFg0
FT7+LRu96wOeeY6tIB7kf3GCmdOTazAeyatvUPzXQ1e/OK4BsEnHETy5cyKVecJO
JAGUkPCZqySPi1/oGAQGLdOqJdUflRixY8/Nb8onGg/MhzOwAYLX2pf6W4fLAQVC
6u4jfzAPrVLzWsu6UbAwvfft9ILu7F4JMcYO6JbOpI//zjC5ULiuXc7CCvel8EHs
kRP++lwG9b3djeWmQwBnrhzvyY3w9Qz6bVtq1NG2vdQYRAN85TrozbDKAwqzNVxV
6HEntvI4EI2UdVml4Qde0qmdcreo1hm5z0EvvtsxB12IXP5GCUSfE5v9y3FAHFsD
k7xSSqS9DOClWIx9E9+5eLs3KUtTQZ7rYKVSMTeCZl+J32LEJT2GIHNEqthQHscI
ZjMjZtqwLA4L2sPITekX4MP7cNrqvSCt78yxLTrW9YgEUmEW7yikMD4ZR1+FaTtn
/Jm2D5kGQfGWJuj7NHHShsgrX6lA6SsnduRKjlzwhoBoDzha33vw9eobHStPZHku
0o6Q0bdarvJBbyRUQWrJAeaugakcb+ZKrW9rqEpHCVoT49ZZF5V7I2HlTEJj3IKX
A6o68vE23Zvjd7QFHOLTxGQhnOx4SQnk7LzyRXonWNKtbNB38nLJifSvjoZ/qnrO
UwQdun604GDQdDfH/vPYel/p0CLO23cLBcjmvE+h1UgO0e2sihvN3qjF7eGFkbUu
DDp2R6/xs3zrjTjd2oTnlA8p7VqtmkoA3JuYyZLenW3v8RRSOtCqkheHKOMkwOmD
JxlmT922rFFgm5RbzyR40wc5VL3cpiGdVbyTKA+D2UP6uzxOi3JVzlQ3sfXX6iJz
UaGDFHA6Ui+nDvID0ontITARvyRnro+PyAdwXcyxtuQHJvoZK1vNeoJLG0jFZxZe
XHza0WH4qX0i97v2ax7V8xBi6G8V5X9UudoFTdiaJSPB1hkl9tH8INheO0qUen1U
Khu+ItNghx99yHrZWQKbbM5CcOi/Xo3QMxRBJrEivR0fSOC1a+vJq7saStZX3Kj8
ZhLZCfbx8rGmlJF5TxjlL/TrUj2bw7a7FhCckRzukIG11kUQzE18VTab/L0tZVzV
7FkulNusq+Uij1gzd+wCrrAIUxE0uM/KLlEaZ2aT+OgHykVRaAS2enxAxLqBYGnm
Xrln3VY8wh6wqypfVuk5R2Qy9KkdzoBhnU+sGitQSSCJUvsbNBUzvzSTjGyKzxVo
KT4y/IE+qXEp+fbWUJZHbMevp/JLIufFcAfKqSlHGf8OPc/oMeakEC0OI2QIDJxb
Bc//kjQXSRlidQo/tskrsIrhU1a8t536oTlrO72WNbVP5o88CsGA/dDG4R/w8S5X
UdX7VJYqsjv4okeKGEB/I9jfyRE7rovZLS2Dnh0eu31kxhtjDElXz1/HO6qAfMsF
ywAshp8flh3BIxGpc16mI1XaWiNocBt+S6UGtN1GcwuMGdZrUHL7COgUi3BrM4n1
Myl0Q+uaLHiXmD52dO0fnIknkwnsQ+zHefxNUiN1zK/UMWrprrIKcFz2OjP+gQuV
C0LXjUkD7p4MBmhZfjckP9yfdajGJPZbSFnAliuhK+L0yB6+N6M0qz/d1TNQyg1J
vg9scvHJMuwzIZuuuLOtKTiXQJsnFCmLudUsCVzSm7679KoFzVGSVGBbqwSULn6l
rtSgMMgfgjT3f7brzuTmLEP93d7Z5VSbTpUKqFJr5uShHaRVN8sDpoLrMTFksuY9
1l7FrLQX471fH/QzhKLUNUKY3CbNYHYgkzDxiN04r8RfChue5TDTA//JD2HNWJdo
dQNkiOylHY08iGJjJnVUsC5wjf2aeQZA0YnbDCdV7zUB9Pvx3BUQTA1p8Gqi2Wup
YRRf3wuxXWrVd1ISvWemtUvZ8oqGjdM1cAsjI/YcgZu2fhVjI9ygq9BF07jOQpQ2
3/BKdWKESafE/c/CQNe2KmQ7DQSNMiYFChWJN/hu1siBp4kdDRZc+vkB908JCaeD
hJnnAVO7q7JzzE7tVAuV62VeZyT/1tpuaulpBsYA7IXphgzkgChVSbyq/xxpBIFk
hQsxDDQrYR/KTMGKlCPdZhQDth0sCTYm0qyZKZ7b0bFXeVj0iVgHwY2vrd4cYj01
D7tuYy+7dgKYfnKqJWWiTBO4QutssjvkkOzgMA9n3on86Y2F5P4h0KHS368RiyZ4
M+fhomVnYgGwLLWfZuYjxhovP9ZLwMEpgtKn8BQOR2LY7HyhXfZaIAB83jnRUnGY
40UKY4tRac5LI2WgZavnjzhe5SO15M9qcLfSy4gBRiNTdKJm3/f0nt1oVN17u/ew
Ry6BNhjR32ykNbhi/tOJZ9LRo5xx+ILZfcT5wYrbj3xVNb8LG+I/tsyUjLrFqLDq
C1wlNzA3ngWQJwEqZe5gSpYKJtwTWnKt6/oaCUzbM1OiF6DpudnNsJea/n/ANmmG
K2lvGdMdLfqYmgtIaQqoXGcfiJ+crNGvv7VEZh49MAtN6781U47+dGLWiBayPgMz
fTZptutjRnTWjSYHe/3FALecHpo+43ONNhJobdvR8CVuEsGU2+V8kTkzZEhh4xmv
WZFNeiMeESnHt2mtE6ehb2rw1ZslmAr7EgD6hUwdmcWRS4XG/CUTLhy++kpXIeym
Q0wW6zFiIysYxa+onveK8BlvjzRyXC4IiIr5aXk/M2gY0f/5Hsrlx1QZ6lvKFBHd
SBbiqsUFkvwzIcvabnrtzlV9o5MArD2CUMg1wr9vgdNKycfzGl9djS9RyRvJo3Ha
lMr9FWS/PtvLwt+EAuvX4773VajyfFP5m5rNVDDfKKLy8lZbKOPWFa+0W2nf+zR1
n/seCQJzI+Jz2NzHHxoBqpUPCUQgxNsCDePwZ7ZV/poq3zGIUS25MSB6vL9MQTk3
h1UKEeOny2VTI2aiRUIbdLge8jMWC6VFZV65U+NJbgYiq6rEXmCBk+DNiluId6K6
btYZjcqaLqknpoUplxWGRcXOMh3hJYNBbvhSois5yxjwXtmF7rmIeUv5Ap9dftMK
X4677iKZXrwi1MSo9hZFYpsaRxNuSO3pXiA/r9WlUeO6dybhOhNC26wR4sF75WWE
S23TIti0JiemCOujH2hPcK6dqrYlJ0lVuh9eTIEzqs5MKvstpL7/zQDWn0UbnbZ8
YTk/Iv+AD3Km7UCWYTo5S16QtE7Qbv1qIHbaooZ8CNtR6OJnwScPXYTXAfwmR+Ls
2QP+xsR2c4GDrzfZr6U+CKBmTlRLiYJYyyvJE/ndhiRxBhHmV/DJzknMMqMB3duR
Ux5ZwCPx6S8d2NJK6y/CTHo4g6i1+6dJs395UAFNnYo6lg+vj4dwYUhBaZRFBAL1
gbYR8JPpNKVGiprQMY4zZ1R5+9E4mQ2oQIdFijTrVo1KvklGothv5omnLvIT1Ka4
qUif6pgfCqJivn+02wzNA1cxrDetRkxxMEMuCS+b5MUrQrRt7BRENEN7qPGwdXhB
LggBpXjYWXV3Sisv1LYcBD+bkxI2+JixoEhLlKIt44Ir6qF399Vpsm0mMZTu7frm
3+mC0aMi5+WvCsBJyqJuZ/4uZ1kXpfyaVhLfaM6wKFeG/7uAvJWY91C7WrbeA55S
ijDUa5Rh5o3zN6FwJpm8EkMcbCFUnoJ5xtDyxEffDWwa3QxPqpRLnq9TMYZM92Kc
/SVElyZjxNJjRGvqkfsqER4MbCgQxaGkV7RZYCB1g1tcFHzOPRpI+okyCsTH9AfV
buRSUNN8mmDyAZXdw8UPiyhJulblrbHjjj4KHAm3k5w7Gmj4VB5O9806iLb+Uutp
mOH/Iy1KXW+YuatVhaQdFlm754GKLyEyrWDUUd8txSvWrJIyC2LFTu1Aj/Hb0+wE
IG8sdRIkDwcExxPRSkMAlf1TZHyFCc5FFqz0kd+KnVrBHfDbTIfbMQszpEmZxd4t
iCCjIC7paZrmY8q4nnVnbxaZdALYhxZBdkUep0k1ucob/CQW5aut6ySW1b58SJKL
Sp8+pCGRTlbFowOAI8UYBp05JjCR/uVMPw7SY5bYS9/1zkSoC4DEOohBZMJu087m
QkTgjNLvyBgbV90nRatrDvHu98MAJM6iljwhDMCCZ+UFfK+hvMp1O0/BPW/5HJL7
OxgI50tObSbxRPZZ8euB4lp1bUGQyAlLoJZRgvOujNhNzqk3MbFLsv11fHDR0Qzw
eqJIdWlXdceCbQVAXu98h1qymKhnn3gtDm0EwmL22aN8likaO0cCb0rwQl/mvUm4
Pkrd4zpKnc6Uy/gk3/J9KWJ6FNJ89bpQtv4V9mmuqqB71r/Tm/8zPvP48spViLtA
q795/ZWsiR3wvHCu//wdbHH9ZDsi+ncAw2ao6+rozwJBHQz1c53sCgNQKVdTex3j
J5jxLK+DjamWrlMbffUuok5h6T2yR6tmGUElhA86p5oHxB14cSohWW/F4qN/5fS4
xuhuZ+7hejnr9En7uhJLo0hmqahUkAFffx9bd9I0degvTiJetFHkBuhxDOBINAV0
027tYByQ0kzf4butzW3hubD4EZT+P9EpT9NsMiKgkQtBfEuUMhNczqw4DL2AeWnl
BMoGr/iwIkX9cBVHmJY1RTQ4UbCGkKoYJWPVAofteZUY8rsIi0mtySujTvHgIiiy
PlXS83R2KQro32VJH+by1g3RHQaN0MEkrBF6/qmuR4broRQ0eamo4Q5xU7uJ5zPa
O6j+OOgloJYH5J9rzrtng4p+atuid8i3i7zmAn+UEEkAChYqnR7wGIPFJXYToflT
iDXikg7TRZwONM9aiexzYlT8FYm0eNj1jSGI2DiPlpB3hIA7XNIx5mOfPhfG4la4
cE+JiMD71K10faQeY+fqMpXF9wrwhy+YSHMlmi+bVhwqWjgi7NtYTyE1WqAB1FAu
O40BCXhfo1FqopEstWBI0WzM/ifegv7SFa6SWGU2gxkc8BCBTwtpiOw932KWH3OK
Y257CDwDrycadxeo6TaewK3ZfZtHKWCiJg/9wRwB/Ygzon6em8Yh50Bq6sIxb2b/
qcKdk7Pg9C+QrZm2Yy8ealGb6xOzcg2CVgTwHPraqb7Fidmj7FWXhLHqf3e884GZ
3cAPBrAstnRSZXUewr88N0igjnBhNzHwG5TOS+/mBcJlmeUotCMuZMHz60OtcqtN
+xhs7DBiNtMlE85mkxwjakZuUV4bqSA8MQubdxE5/dsjOj0n/TbyE3z+dn4Vhwap
h70VDWS67HBT1FxNP2ZOph8KIm2xfAcEJRejH2gUTP8NDd2/86uh3yEaM4/8Gi+T
7L9xiaW6qvxpYkLJKCaznhiGEHtTO1jy5BsCGk0+gMhqaTBEToZAEV0596eylACl
1cHJkf8GRN0HcuwqIgLDfmygf+0xBQB+SPmMPA8JG1TODVpBHG8KUy58qMZ3g3aD
3KeTT5+krBt2QrN1I+Mb2mfXdsoQJk6RKHy7OYTe4sGZQr0xJ6lcC5TubzBPRar6
6wDCzcmDUyNewSq+dkZw5OHgCp9F9iPOXTENzXeBzTUfLF0iy8BhqY0FOLlUGTcy
a0aD/GvuimeaBDYnbq2inIj+Nr/wk3tX0VRWoEi+bpt9TBLW/IQ0xCv/Up0rtc4I
pDn0mcsn1GYOCwoErOOhxEvxHGJricKN/YchM0xuAXaa+6SM4waRCczU1vb6Sh+x
7UWwxxk0p9cArutONL2T0I1JVeyhMUP/zYgtVoGlynUvqmxO2T1GVTpHirxPyGMi
AuUM0lrAzMg3Wukpx3D0wySIJjbnduF6OV7AgvydT8crtjJH7zabh6YQnIhrIL+v
kQ7Xl/yBugfTDCCzgeYtbWB4CMS0HbRfX0WsyQUPvHYkXAmXSC1cWklN3sXWvMek
mENOn/bsdlF0xROV5pUQKSOuACsjPB39ief8f4eTsX1TBPYuzbETm1EMdLovzPRE
zLXyPxWH+EfV83ZCwtVhH+jvYMC/3Z7zGbh/chNJPm5S81kHqSqWEJ85ByMC6yHQ
eTFpguTynhqNuOFc4pI6ul/c9ux3XI7UTe7gD72/bp5+iH5pyioQallSxoiBEMud
DbovYD1mGAVdx9HND/KQclgKD0UJXUiv+KkQawWb++PmplsB8kVSLCK9UbuaIZfP
17aWhAgv1oQEm+1VW0T1Exj39WSTgasNWHNco2nV2hKRW0i8zDqATDbx6Lo2CA9F
7g9dTLlgevEQ6XpsJPj4UlYNAGTTk6FPCMGX9rpEnp2PCP4eYueLFrL4fER0Rdx0
Vs5sLDGsM1YRYCJ6jpxhooVtN34HqL2EM6QIP69uxwRx/PFRKTm1k781ZBjkkAZn
fRewnguQGIGtguECf84gV280HaNm1qmRG98KqI5OxYTQbgDrme3U0XcwQNRGkgxh
vQVx3z6U3cUT/QW1d+pSMkW2L45RZKcWo/3GSTToIiQQRRSN2MjCkn5rNILjattD
9tTHl+fVpWFFPypURs4hhXwAmpnpXC1hn5M1UfFneQwJhu6ju0T+pNpJFf0oIjdu
bf1w0ggqgUmCURCCv07SxKgGbadjfGgUBuuGgzz3NlkxmCZq5Q5i3evGfO28+qdg
/ZabMSMME4NCfdoQZKs92zm59itmlc6hg3z7XDPcLgjqTwgWU14mDrMORqy/pvFN
5J5Bp+wyReRpuMuCWYOEVT9EaAlP+AGn13bHCjsMoA5k+WagLGnP0VKoH/x37UgC
p5hvOXtPfYxWjT9uS32jdTbxzs5QpcadD1qs0dju+6jGqv1tw8hfj890NPFfqJNg
Is1VwYA96F4aAP6q4EGRUWMHpo/JmKVdQylY0QMcBiXM0HgjdEHBvXN2EUnzsQk+
ZlN61M1KKqlSXW7PBFRMLZFrwQte1LkzYnaDlVMAgidbCnVMl9N8JsjkBCA4zW5h
jwDyekd2BdvNlII27jUKfVmp8Z/hcmXdtYDPk8PGYCuD0BPZ6ePto5Z+o7CV3fcv
9YAZqyCBhBiKKMdIjXQ955CO3BCeVNON+O0/YVH38bU7sQq/UVZR0PBOnNcjbE2q
6s9WxCPU3e6NhFc0XzNLqS4CNi7sHowEa3OaWpmCaK2cO/nznLyfBVf/l3b2RXtL
BR7xf2HgiaXuf4A64hlf0/IrqEKRmRYFwRIYqlfQovslxry+HL8KFWmaQXvhcXc+
eACHYF+GlRWDOPc7bc66EJvs8/cpl1UQU8sDkpptDIEe8fDJ/WhNpEJF126qcMHk
MnByUDEOda+u+Hcb3BmP1EKZI3Y5mZJHL3wXx6f+emcSv2pyPD8W/K0gUDM1aQbz
o5bVRG3NfrMWiF3sWit7NwPIJBqo/hxFzXzOkXVHTHLRwMx3JW99DTtJv8C8AWn/
eS6CrIvBF8MGldpYsLDk2I+kgBKprxuHTNjvTeobC+ghQXi83wkt4KkQLNl2oG3z
ZU+tyXixHcwOoVWuSdCl3Ug581JWi5J7wJ3cqsLXBzz6WXzbPMwtnbyE8yW1yCg1
uHTj06I1ChDum8Qw5cJKa7Y3DeYrgEcIytYc5WNyoVVjt9xlFvin1OrYJRT6Qpe1
lJtW7J9ntKpI1Q4buELttVq0pooLX1WPcHAW2ycDlXUMT3yKDegwsKc02mb8hnlm
VXdWKw7l5JcHNjhIZ6JGy4m6xYdKvNZDi5shFdYSStY2xSpk7e1xbh8iUhK2NC5e
2vG9H11x9tg5pcC/07D11Cgzw2ujzM4g2riKCUChhEYUmFsayc11GMdaCLHadakA
4oL4MorUwBoB2KyE/yEEsm+CT67/sY8ERmAS5k3fTs20S69SUOXqUwgoke8uiqjm
LQr/Ult1VTi3pxO9/xyBGMfsfelRyJTb3A1ACjusRHxmyCBubRzQmSEz/5xFpw+Q
gJmX6TA3J3S8CVndgctxjNlpdiXacy/eolioLGRt0NCLaipnSIYW7f09Tx/Q6j4v
gQSLcDfYOAWSPe7vtmJNI4QXW+yVeOen4Vmfqoshoal2321zihHMy7uC7OuNYRnl
61rcXQjzbMw5tCK6Wi8/9h7955nCejSoZw3F5D9oON3v8mmHwu5dB9svhK9O6h1q
dur+cJkYC9Ue0ULEIl1JzfBKfFA+CuTNyZyIEYWY2C9EaF57XA4r6Q5Mcg5Efbhl
kbOzvgbH5tPywz344JBZKdATfYOstXjPfcgwyi/2YKOTPmTJ/JmM+v7vx7DXQhwA
wcrt/QYtE82cKGM40HKU0yfuZ3KmbkygPMHsUkjAcyQmhqzcGxNrmAcQJUK0j+8h
ImjBvvXUVq2WpR5f8jwS6j5TfqCKXlpGgOPBW87K7jWpfqPpMIFXKgKon+wq3vx4
6s7gWpdApX4fmuk00328BRoLgyXShAZqCERO2GNyus9LzINs/M7S7/CvR7PO9/EQ
2PfTPTXGar0ZQsCdzd5zEuZP3qaxUtB9x96Alh1j8eKp9KJa7SCXNtNCGg5zcNdE
UxLCrBFBoft8Ilji5O6DKgMQO95xWs4bRNTYLAhmEuwyNJ3bpzidMwMSFwvanOJv
pZ2aRgNThPy6a1EIbTtUUKQpp0o2lC3bvZBJwgQyOexeTecwKjzNIQBejPLBt2lF
7c126bqcCUr48iqfoQyVxhHdiQyZIhncI0ieVN0fhda6bPwdlcBjpcSOjm8ILoPU
MwZDJ09u0a0bOS5Tctu8ijhouX2olbyDN2tWkouEnoGj3T6DCZNkuE40AISh6bJ4
NQU43Au38r47fHvmV7Vj872RQOxeckIcsZ8soUNNVCW1rfS2v8f+JMHqylkBJlDf
Jt32xgKvtIcKyz6xlS5fZZEgfWwinF5bfNv0Y2zpnLVDbg+abdFmT+lh0Ft35TIY
cvK2BTop3yq9H2HEmOx47VZdE5WvRt132wZQf4DWnCDf0FzxqJtmr5PGs11RUOJP
V87Cl1nvLOcxjcduW1o21M1RSgZvaINyEDcJsvMF1RvP+GxHTiKAbEZJxt0G6e37
XsLuzxfSUewnmkvy/kpIlAmCMQzTRxe25UG4EBl85AAYWS5Po96FZaGlZq8BdLdf
9RG9vrQ7aNVnB5D6OOTQbg6igwInnoeoBr+hYX5SSwbepe2NgpBAXpsXtblKGdX0
guUQ851rj1LHnPKKNnbz3A5hqkP0vpH66h2kfTgVQ7St3SipGldA77U8QsL5dq56
f6pkZ/crlLZekmc2SP9aYqFeNABeuLXQfLQCtm3ZCOdcpI1sfLv548FuILrci5rf
QZ48j/Hsq50KB3Xeiv0UXaXhxsOrHskWb7lZjZHNToHIhWtcZVzFOvyQwOTJHoB2
3E2mUKnlXcTr4KRNnv4Xd9WutYFaV4c59UCk9JerkcBaSt/ItlcsOR5nx99ABbJq
VBKldtPYCu/j0OtlEc/QVZmkTq6COSBUIsnOe/1B1o95a625NyiaxnWDqo2bMVQb
lINHev/61DdRjbz81f/HHbEAgR87aXmclTZ2zCSIQV49AGoiyEH47u8G7ZFPjLc9
+6wg2VVTyJAvh4Ljp1HiF79VnF8dI5+SScHAZQX+vCc7SP3CcFfCDOloA0yUbVMr
pO8VaQ+K22PVxg9qoWGPYssaTbLldb3l+BSh9MiHId6yOVUfhVZHqPf2rSWnLlo1
I0b+Ljl3CazHlicouAiRcU+QALin/nvsZBEIb66tj660mLzNkLmvYmPs0t3qtiJd
7iMMJtV9eI+DsXQmm1wP0EpXXVZsKViqqUe9oR1GgVUvFEnZwfCSnYOrcaYgD16i
XrkOZYCggE1RC8kaoFopfqna/PL4bzahkZFN2FaYTSHnHNfuAFqbCAOIi6Nwsw81
n6MCb3N5kqZs9gMAT47aurBZbVAaI+qx6B9Ovf+0r8GHO1M+abktfF2nUGhel3gY
hgu7M/SjIHkD/mHJc17fW7Fh8XtrlQgTpUV8//eFdykqLL8+yLM56dNNzVgl6Mkd
wByhS7wYUbTjlvVHX/QktInnGTF0fMhsBspGQhtu16yj7gtQk6ebP5jmuUkfNaWI
d6fuY3AGVCrTc4GyU9pc0UOaMyGCqHzDJFDpbHKX5HRV9NuNMUlkFQZbwqpd5xf6
y8zWR2QWdVGpbvEFssoedGIq8WGnhlKZQeLd+9r6LUASXUHs7HcUk8WQMf8IYg5H
0qs9GIXVnftKAF8XukEDT9za4b5zq1UUpelEVBE1ui9RXlOGzgvSmsp93yMW6abm
tDe/qk0RSxAUJUdyYaLblsun2uVe+2Xr0Su2fPaq9uRIDqoenGud2zPypp1/uk6N
q7CeZjpE+kKfUAp1YUcXmNjqFvg2cZ6fXPVGniv4PwjOt1J3lbVbFdI0FHTQfdka
meb2x22qxU/WUvqtqXN0PjBPKGyyt/6HIn5ihfO/pGS7F7kuKz+pT70rIscfQb3/
zj43QPav6IXXN/h1RwDVSnOMthwsoJXcGG1X73R6vMhgN/mjo76qhmUwH+mNW+XH
S5H5yEEBi1pFfCTfsBsBh6pIJB/1wQSGUiDwOSsNz5aJoGnXX7oQ+cNUQyVS+pDe
ue1aOBNe9PyCd36Gp5bNDaWNdVM98cNS+seZKJELbvG4nXxpt/Bxz93FEcoViGuN
hF+AWCDZONOq4+hqQWsDE6WbMCv/ao8fsAMt9qfTXkGisEup+0kCKqCfWuDCfeTU
cJtVhWTjieThKg0mC//1ELThf7h7zl/kaq6vHJD9/mDQO7d7VgKA3UqAeqEIrHcl
v+CDk+x14OmhhvOuR8Y7Fcsd7+m0pwDwzewCMdcweBJQusr23HzARbw1ex7HNiV4
If5X7V8/zmQ6ABQV/BmkTszhyxb8WNZmTnz6/usrPYfRiBSwxp6lx6ASK0UxB+e1
UH8Z0DGVuC9lEaanGzs2V+E/CCo/VUo55tLUtwDqq10v+HdvjSrwIFkaUiaeW8mv
BZWrVfY6Bukni/otijWL9CfuhP0O49mJMf8YPqoZrx1UdNyKG/1FcRF/rUQr6Phk
Z3vOnNaPY/fH2qI8U7jBXrI0RvgpZKDviD0ajTehUciUDyTSnDNFhHtcaCv79ahG
RChV/C0lCwRNJ+I9EeqjSjk+OAHKnzytxWYV3vXnm9ENNEazgqcekSwwtroPKsr1
6EMGEn9iLKCKEbtjjX/ydkci49TV7cQDS3WtAcGE/FqWOkpImGkq5aRDgYyqM8Vz
JLcZau45TS8E02pJEfe2RWqTo6kbR0pBuwloRTTwCsxG4KuwozmGY03nrYr60jJC
Y8eRbCpF9oDvVnxFSQ6RzRkLm3clmgIftzSLMyiJ3wPTCzx7MmrBU8A6fUp6Ih1v
4jKdzmOrW2VWgXLpDgO5UnrPeYfWlwLupK3iiPCG8KOsGNU+sSkAHvTiDei2d6EQ
9KLd00dCrAv6A5+SpUx7BLjQMnipxa3zYy45IOWiB23PC83vIJmz6w3KiwSo+Ms9
y6VtBDuu7jR+ldh4rNc8wrLhIROayQKWeeJAmtTCePiuBl4qW6yAmvrRbMPDixSp
63d4TXmsPuhZzlT95RQLVj8JL1FzBxL/1+kNY942icQr3LufzfannlaFxgZl6khg
u497ZLTZltfFL4RNsQrkmnT96PKTYaYexfX47+/+KXE8rEnjpWC92IWrqZrxhlSo
YqpjMR2z42c2DK35TLW4/I0YqhYlp3Om/j/S9JiWpkw2z22Km3z/DZzWbpXT4IBE
hqUEnq0d7yfmvC2snyUo30I46rA30lpIw1oFZbwcttA=
`pragma protect end_protected

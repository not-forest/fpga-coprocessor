// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
K8lKxZPnHsvnzxLhIx6vFw41Dss5Nbl0oZ0lr/3cG7Vh9agDz68V8Eq8gKatnuiz
JZM5QXTQIEaXeORoiBwP3U6xSTFSmjc2wolGSo0FbPgDybFTc0G2GwPrr4iiF5Ui
kjyKV9jk+JBwwaVQMBqrgWqpmWF2bwEdExBggRpax+U=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 67568 )
`pragma protect data_block
006b1neyWSaoqXqdbn97VHIiSY4f3V3J2Sv58+LR50lqB1MIuVrUDy3JVIVnc2J7
L5K6IHtGig36Fk096I+KbjyTZznioJDlDC55qwfT4U4csq5MLScqdaDWOnCcK+hH
4sYh0AigR8sg1ns1mE57l8GJQvBRO3CZPuI3cC+DuaSPtfDIGJHAadHkl6fhyYST
n12LF0TLabW6fG11iDRLH1ruXox12IcdmtXP8ApjZ51ijU/LRbMHwwnSgzAg1gPw
6tV6oKfjpjFwusYbuFkb2D3/FtzNZz7ArAI0nAxm4EP1GhMkXVmR/iSoudZdpU2B
7T6CgoCYR22mhhSaz2iyghmvsATGT7j0dsHqKI2/dhjEZKkj0I3JgFe6sdPlikiR
ruSdWwrz3pIt2cBsy+85o8r9ZeKfnuERepvfI/0wXMT4JkqnbSBdEugkd+yXXziX
QSRN5IBpOg7ogMqTI4qDPuFejpWvQkQCXEAYcsoYqHaPDk8jSQfi3djFVp5ONGlJ
JDZmcs2snIrDh8GMHIoNFt6RFjIDhMOhVmdRsVZQToF64boH1DGjHcXNR/l3phri
0F2SD81QckxxotzrMC7UMNdmSbtnhHyft+MF3mGGPKf6aykV8b+nfSU3QmH4vQMP
hzPeZKUpS5wJ4chNcR4FUcDA+bbpFBo6+kJB0m3/axw/dm5G/1sVNB5xla+2WaPq
G1oxhEFRihHcu5p6EPVtE+QBycv1SAoWRK2T3EAYEYYi6m9rnZ8FK7CWbOoWJuPy
yiV9HInZg78Z5SOutRANy2h+ua1yUmmRlbxMQ2pGN9gW7WAOB+CTb4MYQjMoOdPn
tFD1PwPWPc8esZS5mksWCc5DSmFADMuDbPz6VZPicnQd5mf7t7dto1gs/OLNoiNT
jZQJjyTLsPj+os9Xy/OWqmdw9huQNSQkvKwRLU33LAKKR6RPPs6Tqgj46eplds58
NprPpTKXl3/CzmJyHPRCnrvwxv8/EH0Lz8t0gVKGqGTVjf+ik0cjgB3rJ/NaY6KM
oG7BBwzQXcmYl7hKfBH6NEimnZ7gSNhQRfauxV1kY06LX73PxJwL8n29L+b6HEey
SJNO+wIIAGh7ca36gPQzNPlNLmBMuaUzHQ90d7IAdKVFXG6evn+fQElW1Nid3daR
hOBbFtkq5SXM0B3G9ewNzfBrl0NFLgd6mC+hNIFEM7851dkOzE8tdxkxxOSTLnvg
sS4aom77eFqYIb7FvtuFSqmYFGleJyUCl7u4mns0he8rS7IASAO2RY/Gsazd0nh7
cfsuyhC0RyNqgGnVn0bB2DRe/E6Xu/NI3IjsDzGFQZnp3u+cW6RxX1gBDEgPwOz4
yXF/LGchDKXBekzBSiDrkaSygQDcZPB9EFLVxv36C7NQJAePyYe3U4sIA1nhSIaJ
KBxXbHgcwxTvxyGwu5lc9GDgm49KWHrH61gGCd6qCGqpXoE75HSuBkKGFTy7o8ud
h6vfbTr0vUx1mEe8rmj7mwbyKaBiqW8MMpAdki9FybOsavbb5fwpb9dvVoV7qnzS
5XgZO4Vlbk0LE29Mu0KrlP/6FgKr/o5QsfWn8jxqmXKvhIlkdMtA/0rxnfJdyHgx
wIwZ/1q79XccEOuPdpfZebOV8YqZRRL3lkIQPYPWBeHE9NXApNV6Md6Nh9DUqBRa
KyJMZHB+o6Ypsh91kolTXPe92Nvoup9pL7KM5Coa8hj74aMZ1pZZpWcuVira+6Us
ZLbjtqp9zBWXWB9h0IgPE+t4RSze1UKMO3VBC2PlqhjtXTsAKEu/lvXmqgm+0GK/
ZXYLJU18w6c1o4IvMIBxUkpYPKYRqBangmoJApWzdnvZZiSoTfIRCzQVxbWKHNmq
c4OgvsDVWDvG9GQJ2sFjRbEUwHIErOMe9lC+8ph7FqmP2Ej6gFPR8TXUj3SpvUbY
niSsgERk0PccIJjR5nlKfEREUVns1g27mOZ/Sq3BayyKwuMku4s1SAr+HtP5Vvkd
jOnIyoxFJq9G4tzina6Q+clLzJgiM9Sp6JPXt59lsgs4deJd2W2bsPeYOg5AGDXE
/oNcXYVBRAyUNe7gnfuTykJANp0wjpP3Wb/nT6PLUGtpQQyjqXelPEv0ApJ+18/D
G8io5+PVCxuKDI9WzBZW8YpB2XbehjNoPLhNPq/p03MFjHx9O8fMYm9+T6mNDhcz
n+jgnaKzwQrEAcpJ27+M9aII8b3BvJ/zSm7DxUqxPOAlqFJk/qOAMarcVi4DPxHP
35TfqjGpVfL2tnc7rSgZTpIsqI2cPfbTTL8/m4p9CHoWR42ToKnJoDnqTBFIWqPc
RRQAY/7HAvEGA+fhOke/wzziavL9Z0zyYDH0nkRxBjPmgd7DkASg0bUEI3mOEJ9O
uCUzH1pWpS7RDEstXzSbWHZTX//CJnt1OvdqCSF2liqMMM9URhOTfMgE3EJTMZiW
ZpE0IRuloP6oESSxjwba4RTvcF8n8X2Hd5/wApmo6Bvut+W2RQOm7jvbwrh6HCN3
BBtKr4Khx61T/f908yMht7vNaZQX/ZqoLIHxSZOXVWLER72RNRY29YlPPTTAsKnC
PLf6KW88Fm37TUr2YtMH1eEpTN+P5pgEbtmIPAsCIoBdoEkp/8DePOrwQlFsH+TO
OQM9WlBp3QIIBdMUbxUKiNYRiBmhqTiT6pzz0naC0139HJEzl1BsFXnNf7J2fMal
HNoSpRTHbV9yD1ZnBoeWMUjniPjP/LYQE0U5Uce8JJvcnk/2gx9qpc7b5fqZamMW
q3rV2ZpZ4lZ+tBOqaKaoNHU+GtcizQZG0UZNNin3/U37v1q21Jsq5UhpakvqATqJ
gCYnUT4O4Y4Me5/h6img7397ZZZrEzRGhcksOxzEj/qinLQ04tdpx8e5zGYLDnzC
eauUiCac56t3l9l7NqrWU/ucLD1qDy0mDf2/R4pjjJBioUcI3MJLJpCRAWWZsM1N
VXN7Bv/UqekPhjKq/Y+ektWuEmhdGPIuUC2wcvU83Xj3B4UDD0pV1JU80QSz4dCj
PAl72y7zPt3xaBiJtP8XWYLMuB5SXWtGEL1VSQCO6Ez+0sj6+flPiBfWs6Am8zTh
E1RnWuYAmFIrqxMomFRp89KeL5RytDrf57vJEepiPwco466qgGay0WWIIYeYKC8Z
jjz66JnMwkqNdh+8UVluaOiqMu8cx7UDUcdzqE/xuIIVmY+XhhwAqMKiM1EXBtMA
0cnvHEu4kFn/53jmnfztq+A5ud2bY1Woapz3X4jRtKVO0Q8Fbg/GDN987V+cM2VN
fls/kXruB3vTEwGN2KvIVwLGtX175mf8wRkE+MAvCj/kEqTTgRNzSVDW/X5NpSQG
hsRNAOUtHoqr1ni02XhDe10zJpare1U3/vHC331lh/iYYDTQaTPycwmhZLh9yLP1
5PmKDCOu4Q07/QtpyL2Y3pa3odRqlVhyjy6iMJtQwz8sz0LzGx5pRKSCTusLfv+b
treglxF4d4exAjUdvSrFmS08/ReebyiajYwio9ZAVTDV8VeNjr6ifqNvYPBkEkL6
O559kVzE9w1bfq80tKaO+TK1aNXqoMvVwqTk9LmrddQAqpRfeRgACLdAyjlAVHPI
BKLkkSnmQFiX5oQmJhTpXf1Z4/j651n5ez+PY8fgooECEyMZABpRgtLjPaDRdCgK
EwuYECJzwJS7TEPZihYcD3GlItueZkm1zF/QZ+IK9uRQnHeE5cVbUOzsjEB2M2s4
aSRpZgF/hwxlhXHCC84foLiV3IEpOcPwmg2EQp00qNWe3oPW9rJtFAOKap14LHew
Sl6p/o2pkPG3UcPCzg+eTDe6/wLyVR+7Uh+Vgk5lCHH7d5MV3qb906la8GCczokT
IFjQi4LtBfzCTbkuh/R5tKp4J+TllHdsNilc6Qksr0OdhODG6jryiYEytYHmU7zc
TWF4bVni7bQNyH4rcngvVxodSjl8zH+P+n3rN4egVlFhujmNWbyDIQ0+G9ntMl73
v0Dkjn2iZURPizGsy9z9UUa3rVwovxw9WHw5cAiI1+mSxipagIhteiB3S/jvWoT5
KBXQbJ7X1g5tlqRipecf4i00KfGzVEpAjzZIQEKxIl+VhvifwTncNTVe/oHS3avo
5TxZ0E+J1/JZG41f0GFlq+cWUQANwYbbGHD7z9CHymvhQWzg4gBEZWgrhJKeOpkT
eTls1S8/dtRIAbXikQqFK8ooPuPr3YK/0GSiZNZ3noFi+EkVZwQQz46poBTJ4yOR
e+7kfp81S7YQfdPxDc3n+ATdv2v7/WK7NR/Z3d/w8sGtdgrk+k1TB10uQ+67Mebg
NSUeGTfeL8Db/BsAQ6GK98NUbp5Gr7EKPTPEjPIupyNBVbgUO47zpfx+g1p4UGwL
l/R9zyp4Gup9r8nhURMwXa1tK63Y6n++mw753xC6pkvtTjVJCVFsDbZQWumI8Ail
+pphqys+k9l9zaEIZ+B1FSh1atjCAnhkZ3GPUeh7EEnFskLDpQcV89Pu6rScnRB4
c1+FT82PK7vDeEYWvDKehgxhthfSXyJl8eFA1OhFrjpjZUegHV87JpgcN2S6a/X9
aPqIZHAVFf4OJWMHqWUiudUtGkreS9udZ2y5r0BOpcP5HtcKeXUmdSs4QDPuo5pz
aZ3+BJMqlbu0S//n94RWDXjJc2419XQtlDn+viSJ5tjOcLwf5hjfL31+aY/cBrmj
mKYVlflIoit7fC313TjUegF/ZTNOzypXhw3yoNchn7X1f0gXKUwlAQRO4vDalFzq
HTI4vgBcwSZb4pOt9h2i4M91FENze6bBr7P7A314rZzpWeXWdRO1o6vVe88Z+48d
mlwq9MbX5Fgb8gCiGzoIrG4gWqTma031OkrNBy39zvHvIK90mFVLYJhfYi6j/5sO
NRGhFLc1MAhTJJfCwldn+tgScSU66RUT2Yfyi8hqMNEcNjYZbRS0PkeOr5Zmdd+o
M0Zy/jyaS6tscv2nBArAnBi1uGHO7Wkv+0Dw7E9XS1L0HqTlUptuH6KMRTwsPcc3
8rJiinVe3kGdPvOGJ9WngJQ8teZXFX1QOxwBaUhcm09GC5JGae4KlnqqdCZkfwVR
cFn2RDNFp/n8NjW1XOSz5cjo6q2vhJoWo2JTSdyZp65DzoT2ZxG8wTFEJRlgwXeZ
/65CeiF1Rx3/73cfwxc414MFraII0Sk8MW45uCArvofm8HntlZOQMI/sFQZHw7GU
+ITytO83KRx4gxLrCFXiXkkh2JUzutGSyYhMHOL04eFJPGcNt1cW5ZpBwhCBkwy6
dYe+ktrDTRdkYSemOjvXYmDZI+hScBJUxb1UL1HBf7smDrnkubl5SbAUbYcWKvmM
i8ylTMGJL9ux8zjgYUtSJwL2i0zzvSgyCIUxN5HCuq/rM6WR6nSdOfVogHRwRoG3
UlvDjSgh6s4hbgapVsCH2pu0A2BgCnXIahoVICrQNEsC9M9xeDJ4/wfX+hCqt3oH
1PwO5prKpI4nQqKW4papNkWQpK4ZhaImyyMgghws+ntAAb8kdzql2i7ETmKhR/IO
7hduKQU9s+umGbjTBymuk8S46kWGd16fYqyu5l/CCAIfKfrVy8sOqdLvwh6EAEvB
81QZFWMeH/rPWJPma0HTGzTK/yZYsHgx/V9ZkUohnk0scbUoD5Z58IvpyIicus0e
rIbFYvxxF1qbatsUP5jpBLE/hkdyEDqvFneWRMSd258ezNgnrst+ef97HDgSetaK
9hNFqZdir/DU2b5a+xFfdTjQm7BjNyVtOKp+iT70lQjU5L1/jo7eLNG5fPp668Ay
vvaqUy2yU/a3p6cIDvb/eWckm8CHJ6de1o3TBLrxyAnJihXwkdAnIdml9TOtEZ6A
9z382RCqXt/PBMhlFDW17k3zHdgChmqpsQJ2KiUOKzIcfqobuPDEZLT/tBvB4T5T
ezb+AoV+ZMj5/n+QoqmGSL/eWEDyaXJrZf8NkOJG0NC+WvZx3YLQ7c1Ipdxz+4ec
j3avKf8HvNdNGG2YC1RBRLRfRQolKQTjx24dwjl2fp66d42M6yqJbzZfpatbogus
o8KWvX/Bn27W0+Og5FdG9chnOExbVv+kxNfh5/OvfN9OlRj8BaUVVbBtxJXAiPz1
n3JNwdE2FzqrDjeqmIcdDL652NnNIR4fp59wVfzsr2YepxNRqLJkJWh80y0Lo3mk
JGarUJ/Z+WpczjaKUU7ag5qt8qGIUNGcPfr0qP4CPrO2Kip5KpJCSb4siNtpRjsK
EL8B7ywNP7TcVPettoQ0+Y+EUovd8Rfyj39hhBCc1d4rguagF/OshsrgONVXQYT3
XyqYEXHk/kCYoHHkTUNrzZ0ZEc4wwwZWisFhD2KM1RYYUg/f4vepHPzUB362CSzk
Bkb2BCq6oCkmpkJAn8QvmCRPkJYsmPQJ/I/5WTUv3D+CSJ8PBH99Rh56wO/gYFyK
uHwI4sqP1bBoK+6WmUzolLoV0YHFkcE+vytIUj/45seJYggxBm4q8LnOz/qPBB5Q
/PQSON6KrkyQmqaDeGzv9augVUeuru3HQCVX1bf6pWeO7UNjZqx8SY4h3Hd+GNSj
9J78QBzlcAtuxp73eYHJ00UpHqdegJ/TOT+Pu3nY1uRshbyt0K29FppsG15Cl2VF
hxgu/CvPqgh1s6Pc8K7nJSPKg3fMsxF2bwbM67TaNWyxgrOO4XPsyiTw96Bb4bAY
0lTxEmxUBbwnS8unhqq2dtBwq6cTbDhsIXJtJI+sLpuHgcpwtbdhhkonztD+HSZa
OM329xAIkJZT1g4vlBE2yGIJmxwbel/KD1NKB6FaN2ZNGqxWRNS6fpJSLkfm8mGO
3g7lCTFyVHc02hV7fHldBLanZnVrx22C/aOL3CBvI0qLam2pt8+axtCn42g9QPs6
ZjqJ/+i/otUey0dfnOq/kNKxXRQN24LF69Vo2qmqEo7RzIKnUJdkxnj24ZJDgIT+
n9EijM/y9vtksrBSeFdx0kZ0DAxrC3Safdu2fhn3piw2Z4q0c6kP0taXUMP3oFlV
9EV+pR/zDG2Gt0mZluQRT8j3uQwZQIyB8iZbG7GboEaE6GlCcJXo2461pmO9sR2j
NjfEDEyZ3ZLO6zkoiEBJ+cShTp1u+c8DpNFcmwS0G0rNt8v59tBKad/zRDNqTG9I
P7Q++o2rtXhv2/UMQTZ8zJouYcCOMThgvwVDrMILUdssiRsFE1fEdCy5rnM3GoT/
vqTj0mCQmrDb+NNf3xlYoJrUwrpEKLnBqXBfVX8j0uois8Mef8WAvgs82qzl50cF
5OlMJFUgCT7y06CY3bhAyyT2CID8jBzU2ICFegxr8SSOOoztDtHVM5DEwOdKFvaK
Xtftr6wvSd5r3OjQp+6R2wNrIi7XmzOxzyYKSqk2pbRCDRYX295QGp8NzhUay5Gb
GqoCApvKTwKI6A5N/A3sHpVyNYqQ5Fykz70Oa2ZULyiMSKuDA64t7wt6W+M67ji6
bE8KY6rSJieYNDjje7x2KuKffF3Dn/WG1A4MObMCU1cD3ljxdhDkluvnZf6CIfvC
DYRZy2V/hOPMDvcoC20reBguLxxVuOTfuebUFABCEvq05Xr4qA397ya4SDRbUaAx
YeMi/uJ+86auJ0ghHgPcUoUmaBdGbUvUSNBlsL/KEz6BJNJCB8YYBFqd5M9DpeTj
mxRaZi+1mduvo+20iZJJ7tIsq3DNp7Y7pnljKsvFf/z/B0ALggSwy1Y0DICMSl3D
lOaqx/wCJprYJe8D1DRWoKdHXRJgyU6E76QCeZz3X7aQ23JtjbOsCjxnM/AiRnhu
P7Lujack8ylJAFR/FPCLisFDmLWiUnKE8dNXUOLsGNFQxMkRXtKXS8UGXFvAsnmA
a4bsK+lTJgLPwGCbV4ONBQAEjvPvYYxkDf/QawkHyf0UrZ7MH9F6dBO1M549eb0L
MqeOp2uOMWFcAbktqgpoNu2gl2QWo7p0SeoQ3pWEFOea5iqhN4RKza+PPJAYboth
AqlHY+kKmeV9kqwDBYdgvGiFEm31xOHboqp/OS7WCL4/FU2uXQOElHzR50zdGMB6
BBpm1aWhNqEffech7Ya2zs7P5j58hM+NNbpJ2odXm4/8c9hTNhZ8gr6wScXbi9od
S+oXCUbZv4J5ep+hc3On7BpIZHj2957KMeaOfICkiWTcyBF8Ckqu3uYQ0JZU7RGR
BT4OBoOL/dhHKy0UVS9544dmWndzoc9KFbivk//Jf8OEAV9izq0Jn25/S9QM8I2X
sJ/kT0kp5H/aI1YyD+dajwMiWlgQ5dAq9tm35SBijPsA/5taXTHJqJjb2VFXSMgG
3OrmwapHtLBJXcwEPMaXmrPxW/b78axXWdfbTYQrgKJGdzb4CqILyd8UF2nQPZPE
8gW9WJHqyUXjsvg/K7nJTrFNVKj2uLCvV3NqGuVNA4bu+vkcaDM6iZPtzNWBmK34
Jy31LM/2HS7j593Lx9lmcA7Q4jSERlXb4B/ZlwWtfH+74AQy4I1SrHAgRvA85gBd
C4MxbnX4jFc+fdj6iQTaziU3IQ6Xajd3xu8QbQspgAtHcpVo6YZ8L5eAP0F4BNUB
+RyYZyA1XPD+ECxjkmfTSSIwFaOL4n0z7qF7KoDestAVGw0JJiLnUOukV1nGzw3+
hPxXiwUqvZJ5Sh01AGuPwCM2KGRiAf7IKRdqgj5NsmunHpg7s28F11QWLSIlkwNJ
ZicKVoGLCxP3H91qLhqU2LiG8lGEMRW+HDxUayQKc7/ZFcB570nxUR2jt4BFDvnx
k/9HqISis8Hvf6Hg2siNV4Xks1zuny4+X4v30QJmXWhjXnXctO/SZu2OBYQxKu1b
SvhzVLE99Ru18bhn9uiLINb7MdxNUFm83crEmCboYuKlkwMEyeP7CR1wwy06BrE0
ItNKw1piU2C9KoYYXzyGlJp5sOuvUdKPDQTeD/mW9jE3uT0zAODDXJ4VF4e7G9rY
tr0/+8hyV+wZe+Y8cpJprdGoQt4wFvVS4sDXtafHQfqbgzJ0K291meYrQVTsr8iL
ShFikBXhfJqAmFkb7zHOjIWSg22dc4dJmoXqQq80RAU8aLDbXRGjbWwBMcd/6P8g
2MXL0XQN1u5qY3LeKbDu2wzDKW8N6vB15JcYiXKTa5bhNZCi2hTkGzHi40CpHjz7
Gwz6wRMstpdHZ2j8BPUdMYk4mcdBfUcwkAnsq0OJdmXSlIvQZVvY9nH86q/BmW81
U5ZMauwEN5FqtbEPN4LN8x2PxsWANaVZaKuhz3m0ThOFiqtWdQ93TOGZeBxuuNQX
WusWSbovRfeEc/mZmHh6Op+fXCPv/plRFaMYiEu/YT48uvFD2V2wYkIcv9D1YN8V
B1YiH0nqbRbHTen6UFpS5FBA9BqBQvwmQJFhrZYEroyRVL3hppQozAOxU4Ie9YcW
InnAyc1hhbJXu76Erpf5mBawoSfDokUVxr4LwVgpPSDd+gdJZrp0QdY5CF8oFQZX
mUN9WpV05UhfKGP6es0JYQupqY4ZOImJ9WlZzVLfk/IsadhSMxzXdX32KPwM+lvk
uIeCu5a56r5vktzlofqc8iqYg8is6QsaekYsZbZGme23MlUdCIph7lXz2uSAWpl5
7mA0jYYElRDDg4vGnl3u1prG0/wA3TMUiZvk5Rri/hHPHXqQ9bYCiPIID2PsSqOj
DvZZIsydj7VumrcBUahYb2kCa2MU6Ku+M0hU/hDXU/TCDNQGw6LbSe7y9kD+7e55
yyDItU9XJKZ2dKaoiJ7infR6FgF1x/sv23chJEmN1o1rQCOiPBUqCA6f+PfI854e
9oHHVqipSV8qt7eXLyePcyKWjZCcDep0I6bJxTAUqPCkc4NP42gqTwp05+4jqX3u
uJBm8gLNauI1Y2DjC1sEJZkyLx+FFg+tvFY73JiW1thuL/XiBCM8B9yURemJWmrN
bRpnniNwa2C4uLsW5aSkhJ13lZNCL6JW0GzEa2X4HPHnxvWzIt9Ez3nxryndNk1n
HhOcsaT2jAwnYxJFIK8B0w85gQmet6nX0VlXXRAhcjitlS7szC+nVVIJPivbw7cM
qDtI/x4abW9GmZEbMRER8hp70dtSw+42cna8gSek0IIEaA4Fc0uy97sM4yIK+oCr
DflQ7FMbJhR5BQcCU80oU0OWDOjSw8HidzngEUvepsdCQAXo95y0J9dvXcVtEdWd
kVTELoB6dsPX/FJnHrua5vEHG0rKGNDcu2DyAAyXzfizdSsAcXOXAMpNP6hLNMW6
nGj0XvDA+3NHmZeVaw1lpS8uPubv12dFBRbDrDC7ty1e5jVXLC3R80il0V/Qu0jo
WcBM+ymZTKKJ0y8z3rhvfRqxQUlPJqDhil1ZGWfFWMgRcF7fqxDqyucwPsXiOTUW
ngJBkYKpoHUjvQR1ooIskl/EsV4N/MpwrNDl6eS3fNs8mGIO8hHLD3W4M7gY8Jto
7XI3c8bfapOaKhGSBV1/Ri4Md7KDh/LqC+0N52foJxcJInhQ+LEvDSkth4CiN/yE
1NJIk4gxLEY96F3NW5EotA66L3luYOFrc2VxU9On4bihUcSZtrdfiAryp+3MW9P/
t/97VGFeHZcaYjrP7qErk6gXDFKHuWcMXBiucG6dsXQjRALMNWvwkl7tPFmDWEZV
Jx5s1gK999IHWcrHhbT7pFXq7k2oPH3QIDxi04NPdEpOPZlnpeNgemkul6gOmZ0a
WMMuMPJqejmULyiCUeGfPkn2Bt+7VTXoaIJE32OGHwsWvZfDvlxRKo3Tp1ZPIfdE
LqhSIukFtF/a3C7rSyQYCrSr4GbIeHpb8QccrMi6xhGoHaMlTYAdpEwFJwv92qji
mEUd1g9HdGFFodLzNV4SiwG2e6ADhZZTHjP+dIW/NIMtsAWtyCbx4ivEjlo5WjzU
ee15DoVyMWHqyqqC1x/0ux8SqnXQirIw956O0V/srlaratcXShzdBH3PLfXXzjyH
DOS7UlHMhd5QF5yE7VgrOwfKS66WJkzbsrIRAqlkFCHWfs1SX6e6jDqDa74PLQsq
NkQ4KUTul7y0Kj/NPXtOBD6+raicBIwvv/PdP8Qz/n41Xlcciuqdb9mn4XYEBbPd
SBQXB8GvsRRuqKt80xgF3izX4s85FIchEM5s0+nmQIS4IM8h1tGGdzgusKRmC549
YXGME4XQl2r3E85OiF56PPjwIHML1ikVEdZIloD/P1IJhLIZcWXPwWCtyCTEIIdL
gi1ZsVeUxQyGzjPWb3J75VSoze31K9wtz1N5AeVW05ML2dlmdR4EaU6xuMCOQVPy
YX1OOwciIQqajy4eV/gmdyk9QaF4c94UN5ZxTltfSYZAw2dTYAbajvA9QcTWQc2x
8YOMg8eIAEyeq8GVnyatb20KgoxmorHBHF1Blrc4jyzcsJ4Ae5iRP7/Fq7N6J+xS
FFWNvKEXGubT4tLNlgPlvPQcdUvQOhJb4TsOpZmumnSr5w/i0MCxXvZly49FvDUE
nzvQywbBvmxhacLjyWgHecPY0KeNkfCgRbqLAn41YQaeRlIGnrolt1vnP58VmE+G
ld5/j3C6VTUv7keduIhnkczSiWr3BlhHOQsA41Xf2z3kgSoztTXhF1VgkeyHMKt1
nqddbJthUIqhLyzvFDt9erYeT2Qd3Atwy2lP4Q1PWyuln/+zQhh7cYBMbFwuTH2i
xtVrCdFXENE6JyY0NtJ40Dzmurit47xc5PXhTJZS7XDknC80pTarw8MSsm4JwKjn
u6cnrH9FJZHR8hZCNBrYI9uQga1BbV/aPxowJEXl+2KoxRrQxUSqhXbz7OoWBKP8
JFHyWSJe8hMEeK0iPCsEvrNnft0OwDhJXSaMGu302CYjEGNm5gsr7iyXOe6AvyCL
j95Q5g8tFKc74DBwfY9KPTOqvvhfM3yTdlwr59Djx/CXhTkBeJpvYp/vzelDhHhr
NlXIZTUeYpyM1dpnJtbEarZ//oc1ywewQeOw4+K1OFWi0LqJ0VxxUt76MXggIC3O
dZfayakqgZV0QpaS4zZb6lq8BBNo+P+50Bm5XyUy9JA54WkmEBP9o1wXF8ky1L/N
MKnWpf9U84xwLIDOPcwoPlMpNmaAkc8h33UASQ9pSPqsiKKeoKv6npir2TnOahIE
mpHH2cLTMxrmB5QWxnF1s4NsY/pIQBew5LY7gs0dPa6lM8CzQ66voW63x50fukYZ
TU++E4KEdC5I9GF1Ol15sKcqnLaxTp7dPnUFmXA/kvm71fhTRX5KeqYdCECt4vR4
n8XkqZfC43LctQmh4LlNKcugen6N9X0OK++tXtHrvAchbERTVWkorAdbukpyVIs0
IT43lBSWiLfI3g1kHG64I+EizZRkRQkeQAIrzkMg5lhv6+AmW2R+XiFc0SoaKtIp
2To2lNImXX2zsJYewTaz1PEJRvy05skxnGP1ztPyzP+spB0CJY12aA07ItvJyhV3
BTuEJ3EVQGtbNNuI4jyZeo/kawPCXRx/288n6NzaflmQIpOB9e6DVa7/pjKOe77x
qYmWurkpHiRj+W5y4DrqksB+Zlby7GzbHQKbkEvAavoBX6exxnImbvNbYpVkDPOr
D1xY25bAnNdIMbDqdJ8keOWF1fBxuzAYJ3LTYbYc50nLPqBysaa8WDs+9QYIT0Vk
viqGVW8kHchr3a0GxePxl1zANQoHGVapGt0oeJQSsmjo+3DlUV3QpViDpu3ekJ5D
ZJA8UIJUzZ3IzddI1S4nf44nMa3S89psElnfeYIbBjHre/DJqt5vNvl3CIqa3fmL
CUG9+XSSP0uzZ0HABtvEpeHlEgiZ1pEQKuQoPDl8COr/+jAvbTv2/6QQ2DPBqpwy
AK1ULNILFN1HP5EUzimoE9NKVgXoBczcrS2K7Vbval7vk5h5p8DAe67yiy5KAULh
rluLj6lreF33qwXmaK1b7J0tfXLh0jTLaGXmV8GInVGaneftG8JPz4+WBo2amohb
1yHPeJxvd90MSM0Gd1gXSGAXzJQf8bgzgD5zEdFF5US8cqe7CBGJRj4ml/Gg5Q3J
O3izW85rjWJUi+eWjxYvVtUg0zOitXArxUfUphuwJGFbtBrVAOTnqvtazdXpuVcX
NKMioO1m3KU8C3qI6TckWpY7ADUrVFMHxio1pqodu2JamWAfaja4k2oqmPMte+S7
CqFES/hqPtzr7fM1KKpmY1AjQaHI1NdpxX503AJ5Z8BMS2AFKofQJRS0zmdJ208f
7gV+pnmQUw+mxVtnWjkwtxa/FLFVObBz3a2Xmm5mwPQrgkPy4mx2jbW0ZBjA+II7
xMkeWAwJiG+M/aWDbMvANxAt/ML9MUCaWvWdQXd+Yo2dDGLijGNb6VkTasUfpVEC
5HThwM9hp3nKu3styOniTKx7rw52nA06LrFkEsRD8Jqc2LoVkNDvHwb6LF1xsf5L
trnlvrLkywzqYZOAlFDLnAO+1Za29i7yu4EL7Q3Y5A5rO5nzOKs8p8Zqm7bS2wFO
DE7EYfoLRq4OrN+uL2BII6b9MjiqNwx6cQiWMg8ZPbpTxW4Kbc8EvFbDxMAxsjjt
ei5yvpOIU7Jgkh4gaeEZj6AmMPPVqR9ppGzkhYjl6u1GoMZuXtP3MmhLMlIYRA2D
q2mCpST8rmELQ5SyICDlYY0xx0krpK/ku04KZy1Sq8mJ8wUXU5M4rN+1RPXTwM8K
PdRIAZDqWXIGRD2LlR0bhhOmB7Pn3GkanzQuSKfSHHcZs2HKK3RpSsqdMqgVsGum
kaeGCZ2IpYRzOW8e6eUZrU4FyVVaHbRd5zE/FOQ0a0Hqfuj30ez7/l4EnBvZEjOe
gq6Bf5f5KCEu+wtcyxNxxUWPfUQP/GUWaI1LrNnaIOh6st2brzD3wgFsprtmzpYv
HM4+TWhVvqnN+VgRR79mh23+LgltH6lbvdej3ZkAmJxK6BD25QkPIsMLqJhTQQ2T
zmm5mr315crKiBy1hcNm3+EDZYwFQOIuQroMA5lqKimu+q8th+0W+wmCWRY0Semd
S2pXHZao8oXqkVy4F0G3SgJBdNyTeMkTKbpyL/diy3HXiBgUKcj6WOvpFyx5kHH9
LSFk2rqLPcm53Uzaj93LpTja0IQukoCf0PkqBaDG/5t+03i6ThmnGfrL3fiV1yRQ
ouWgJAh1qlh10QxeV1NaqLltpvbk2BCxGfUeHz4iBxsyTLxxIHwA9FmUcDOGOHXr
eIBl4kSx8cCyyprxD0nIrfxR6rA+H+CpyGyk9OFsoD3/s4bGt5vf8TLa2ZiZo5V/
tHRpJ7N9zBR6zgcODrDuQ1wMypIOlNHbmEyc/hLBq7SRu8HkuF3depmJICyykwF3
BJnQwjagYhveAnWbWxgC05lG6Tq9DeGVHTdD18dtrisThr5y2q1zj9EFhYj/LPl8
xHUHJPyth+l/czi7gfz1ktP99SsjIxIN/8+baIUQZXQbYQmHxpXuLLsPB77zb08X
JL7qtdYzJJRwEVD7rbVsPunUqY2wEpwNDKJp4usFWg4YsYXFgMqZyXZiQh9+qqhh
bLxKE6icxsjm+p8itVfxMIczRW8Fhy/QEyDiw/ADo8WHt7N9YqwyherccrhWOR5M
kiFWBFh70scSjXIB/ja/DGQrHMMtV/S7SRDJqF0KcKs5seY3ls4Iq1w6TzN3ipBw
Z/SfzhU+fZuH3fQuCRe/yah3eBl3rPTtLIuW4bRN6NgByWf6y2TEos8Xyfj021Sv
nkz6re920nx0E0nuiu00LIYKoZ/T2reL30LUn5ZkXEskmmCbLwLqqvD2TK4vDZ9z
XlfbAvWoL7jcr2a4wZtNC3xIrWOyEhO2LD4fYGgCJE/azbq7sI0ZS3TsAsHfFGBe
sX5JhgCbvql4HdcxV6JriLPY6Wc5hqUl4FlwE8fdB4dmay9tyLSfSVdJtoC4c4C9
Gqxai0Lvu4ZbUcf6+xbBDiF4Chwx1hdnckCbuncbG1ZQZRm5UGRKwERnmE/wOIv7
IweMGcaVgwiVIyB2CW0bTHeHwiv7KnpwR7BkBcfxEUMA9flfPMuu6M6KhN+WSoY+
LdhhKqx7gxU+Rlk2ka4mlwiX0oJOIeuzmbWgRpdvQzaae3bH6UWLxFvwLAoFy672
UHa2sJXvU2vxq8vervXZPFv46y3FiUJCDLvagZFUF8D8jEZFlz0HjAk9r8grzUa9
h/wqicc3YbxmgKZu2Q/ekBJ8S5/PSA/fftVi3AQC4r8BEhshsp+FRQ+MXyNjxVYK
18AAqbFzlcHd6xtmeWRFZXoBgW5GowsM6JgbzRP9kXnzdH22OWTIIBZyyRLglO7R
sje865kCtKENAHD0WKW+bE5h7THwAO9GXybj5HDv4ZK811M81ef2IAI/3QdQEXcQ
hYw0igIwA7unsDLHImcJYIrx+ueW+PVG+1t3hKrlLvYD3RDxQwSvcnQgwBVvvLHE
1PAQ/MLJpFCjfPidimIm6QpdRnutC9WTBGCohb1BAqpg5vHJuCqYWq3OpXb2X7X9
aD6dN82Cz7eFx0zNGLHcsRUmhyZe2rMAwZyfs1HRBuKmdwZQUnf53JMxsjmgo5KG
9Cpj+oY3pS0AQfsnkD/yoS3BRfPfctS1pYv8Ni9kPmLSANKYdTPV0MR3P1k7x76J
K5zYK4ziTfIuKMZy1uOOm3NVfNR+Au6ef4AUg9tZ59eBERLbx1yjI7I8kKxrLdkC
Vj0y+iGYjMndVi/xiTjzWdQU2aThDsayJYqITqs8w0eaKmkJ5un+/ID93YBPvODG
QtXhtkq4b+DkQp+v1Wh2EnGwak8WtKSZKa1GGJLGnclsUHOFg6BKeWlOz0GBSP2d
ZY5NbGn1hb7cqkjkyc9GPCZQukBxJDBBYD20QkZqZrh0YgmkVZsrNgeJjpQAkb3u
3rHg3zxqaP2CIWddGdoRoeSBOjv1nZUqUEF4kwlhpP3D3jZxwuDcFHhrdAPFJ0fw
ZLqVJTdPpkAPs9EpntqEhzvDzKmUpAanveaRGZeINskFg76goLH4ODAI4eE6Vw+l
KJPHGNNtPQnJIJB4BTsBtxKRAT7d/iFVk1VjzmQ7xaGGS45KO9lAiMFvhZle7SLJ
qEG9D9nuU0K5R0UAKq7u3dAOAcdghHyg4QT8cLw9BfpGdgm4/dfuck+Dl2CXbQJI
GEte69XolrceIxLrzMDwiw4Wyz7hPwTR7zwpi0zn2Ft4B5bcgiGCxZ6AQSZn4iOs
SwlhXByNg6v9/errcg9Fj0y+7iuQopsLfXHl6H95RjqVw5hXFzpViJJrHyVq6CsH
j1C6OOZvZsfRTIc8hMmMKcL7IvjFYUSX8RvVcSTl1EHNsjBAM+4T/p0gRdB/9wgp
bj7ndTMGEc4X4UkONTMyQCt1sTMprqpKMAXqfJ52sT1ObAWXOZjUxJBVtCYde9LK
rOXf7xeKt0rIRiucgg1KPqp1iRuml75SoXTYPJByRj66H7fdp55NY2pkJQigSH3V
ugBDhfSIDLQFRdMTFUvtaQ2GnDTIXtLGvhTsHHy9rzVl6C+x7tk99QUyo2MI46L9
tPwEUkA9kUj931IL7wYUGdYYASjlBGQ6Ina5xgSUnkvwEAVKWb2guG6FYQ1PMT4S
pgOXfWlymSQ0EM/XlcoawAzca3Ov+p8xSfkBt/LxlXnM9pInhmUtgkL/v1qG69uf
j1CQkPiomjNi1UQ34PJP0bHI1vJYbSEhIHOx47O1n5DPeWaGFWne/+hK8RdRgieh
vh2uEnIDMnJNVg5E7yZ1oj6vSF31NHjIUsJynpVuzd1Gfm7La/z6xC/AkF3w7QfF
+snYF0WJP5ig0MxGNJ7+89tyhroxLw3U0Q4tTc7jO2lm0vNAPXh0K95VNwVZRs6V
L0c3UQEhvoQd77BmLiyM5pfQoMyMq1OgkKsTdA1ImLz12tMfmN6P2YHb7uGf3J7X
gHJRvyEN94lC+knNPnQ24u9yauGP1prvi+TK7CN5o75ed4l6eRoDc8DiQnrF4eG8
VfSm4RQxANEY+Ampb3gAtkyZ97MpAwfEtEIItZgc6pZk8PSNJqDtZbUvu0NcNgfJ
czMQsA6+1dDGipD9JERtxlFgrv1U1V7OVtl6gHXgO0I4nJMKoM2CGSXFE5PrEas1
1Ye1UORH3czmM3tZ1yuMsAIdZszom/0Q22wMxKCKZj28DPtl640U/GhgPRY4aNb2
THOiAqeMN7aDxYwG8EhaPm3EYOHnGz3v9IonvQORJkgmjpHYhLKKU2LXDMSfSsdr
wueEIVxxeoRpffKIZDPce3JZXpoIEAYTllPXCxy+BGuXzTb/JPjU/EZr5jUPtRQC
2zmiFvzES6DgWkJHZOpOlaitY3EmwagNizu6n1OT9gwvBJ7cLFRjQ0V6N78uLlHP
QGbSYdPULoESY6L7ZTGXBsP8tay/nNDPIzy/QJaLGxciMdEcRAmtQ34i0PqF44OL
sXUi49vFzBo7+uS/UAFvOp/bYjncW/YaH0U/df1rYCh1X694XvAMekQLuvNM1gCP
Lqh64/LpyvomIc0tXXRILbFItOETnyt/A3T0IWlFshKpVFhkr1/4z7lo52PB6Dwq
6dGW35ab9WjmT+32oMeBq9kcaw1p65lUChZwRzZe5ccJ+55Y2zzh8b8bWSyJlFpu
v6SDAJbCxiJpJHnQQealyaHOIy1KDT7lQ/xzKd+gT5MUxFDAk2pz0tJZarEBe0mz
JfOZ9ngBmQ/EjWz/4BXxQJ2DJckHqr6menW2DE2/eqKe+CMvAp12dk95GKZfOuud
MtMNWR+Kywmv0FIw5pbheMOg6/v7GdXHYSeiv7U7bzDpb98+ExMpxk/XpfMdvm1U
Twq1oPKVf3TPddPfDYEXTSMd4A75aZcvEsO4BYP+urAcWGpgzn/B27b8TARO9adb
tZf+axumnfSBDX2tTozMa/WZhD5d2sc7yCsOQ8DUGyzdJR64DUuX4Yjeby4lAeFe
6y77hhGOjAHYdiU6XJAV0G3XMUlvu+JkD0YSQ2ptBY4YuRID+8MwIn4b6u9VQVGr
JHao57xblf8mIlIdJBxohGpU5A1RBsAN/kBbJFz3SaLnnwCZKHDNoJZypj76VuW2
f5BreHiuRl3HUgg1QL+GSFup8e9RL5a9253HC6m6W/QwIxQFwGfXnauLYCkqruz4
4YU5rCBos9byGnl9ZYt8JywewIryc2ZKpFp2rxUE9FjVesv3KG5US3Vcr9A6YgkO
LslGLgSljbMnz2VqHveiC6weiGf2HBovUuvI/MEMG4ejQAIxJFZSUg7lQ7qEzA06
GJAyHewEkEXYAko5SiqnlDKaoUu8NjXXDaFaUk+xlgiqA6nvHQqk8YfMOF4epGG4
O1I606+9jeO2iYbzGwQLUwCjHumSkdTvRPdasOGbjA1OttZQliPAaIdN+8F6t7xW
o2XqQW9JPYOcr7sPtl29okh/7NkRLD/cLDhpqJZfIh7DtY7GrshK2EVB0mjw7SRz
KgUBxdoEb44QJG3wYmDkE7TnDAW4EiQhTX5B5PxD9qMba66OU6QcE8CaEh/Ff9tk
0Fm+aa9CuPWqDOzgIyLjlUdpuUmr4X0sYxEvujFqTssn9/wwjhHfATUIUsUsHKtg
VAhce9MP2G926yl2qvvnXsXPWZ7MjqywQQBwelDvZn476UJqN6I9mwzIF4GiTuE5
CZDLEfYG4A2EnxGdLyyMnNXbEhtkNDbfXtBQsF+wqz3dpE5PPxxptmMkeSBLNYui
OOkxoOOupUcRdxwpSWJ99pOkkHQD+pjDE9mqqV4ttfMAOvsUgaLDIJqsefcD6R3E
VfpdFyWfxYU4ct5pB7WpZ0LcCXOVsAfT+wvB+maAZAnWUIpHqVbkGhjwZTaMo/LL
HLCXrvXzKjdePNuZtHMQ1rWzqSs0x+8kxw+Hw5VvB5PYHitDD9UER1dCa0ZqxlXo
ijBUO3SbQLf0uJYptbQuTPsOmcs53lFqQij0LuJMKCnRG8jKPMeUbqeNz8q3Fufg
AMb4Ia1Wm9dC9bKrABeHnZGuUn5VwVuIzaO/fSC1GWuz6S2Hc7dk76Zlmf8wCYWv
+TeYuVqLHr1efdoXCUtVrNpZIm3/R77TePT0eDO5+JQrVD6Aomqorv5j7UXAW/x5
lJ+Ma3ON5B1wq4de3k2k1H88O5FMvintioy4nWARcFmVQoFPCSj0u3wcs+4Wev77
0U5ehz4UrU6eWwpho3SS5/ApfmLKkGJywa9R7NgEFStTqLbPWiwnkOIE2ab1EKIW
jOH55PM+qtjFvm737+EXxAABzPcmNpWB/9HUDf0DEilUprnl4Cqpd9YWro31H0rS
Ed6IgDwjlG5W/7hhhuDHw76VsuBVjOo3hEJ2RLPAY7pnVnEVKOiNNtKrnVsbbEzK
YHSy6Poo4wxf0AGnLGIxBvTz3ZpTvYmlv2lAbbpFVGir0fwG9J3l+BccCWOyeR/k
XJ/+JU8JJrEg1XUpjK9j5gZIIEdd4cebhulySW8EHpOoexSrwHYA/av8Z8YXmsKi
QOPb0nZe1xWxZ2LEnufouAcSMc4fV2O53MkUtYPs3L6Sr15p7gk5lpMraBtXrKR2
htFDjQaJsJvAjrSRfShWmUWUOElI91DTj5Z95BDg13b2frnjaSp9NZ0svEEfBBh2
Iyb9y5tIeotMLsqF9XWn8zmdOsMdAL6/DXp874uwTrtYgXvlkRTbuq0lIuLynstW
hcIam6B4D/ZG2BwWFAp6/Qj1TXfKP+4qRSfRFhaLLyuR6Yi+fvNIFyN+gMPu5x0p
ZStzEMvH2zGGA8LnW0voMoVMSiWn4/bxlaW6NTN9rS1iN50wd+eQzJ/EYQwm3bg0
PtItlEd08HHfmKZor792W03+GShjqV/oICF28GRSF79JYxvIN8IsfpW7WYTtIYe9
QcCEkORvlDqopAU7381cMVBqYPmT31kqK7UeUd6KjCRlDjvhsJMwyJB/RXYtW8v4
MUmNnnhoRMtTFzj/6Ti1YlFBp6p3CthENhRXQtgeBGzvEASPekd6wM2KBjD+/FcE
rKXxcyOvDtXmBjZBMng2J4me+vIK8xMhVell3EGjzUv/qAIVpy6DN+W1UdTe6uLB
3PTJFuEhMePHXrk5vxxeiNX2G5GaBV5cWYyPLSCXm7mjEqIu4S/++8Xi7r2vwlbZ
w+T9SGH+3R0SYpX6mWQnIaVNKpnE5XXn40qhffPRf6gpm3cUJ+BjWp2kP03sHE/m
RLaKtnsvSc9hFseIQx/aaEqYsBE4IuEDK8qJjXjujwBTKXA27HJuNt5Rtv6ck8GW
3twPRHkSbYOqVkkdC6FRoGnCWtGEXyjlOe+z3efNE6QDOCnmYRPZ2UGBa/96ggt6
2aZUHwCMtSKfam1AdqIWiNL+8jwKJoR0a/Xcg8MCaTOSpHOrzxOlDvhAoiudn2z+
Zhc8KBXzMWaaqziancS24BJdyCqyyTX4mNEgA4whv7Sde1G7VskYuU0xECcD5YV3
Qydxdva6zuCYJkx12mrvs3SAONddYb9xceYP3ZmoIKlfit6ywmEvYaq+xmVQ+EW4
TkmRHfw3K0qQLyGLYRy+HEY57mHse7/t+1w3Jw/rU2WjnU0RhTgA/UAZsum4N6Ue
K7vCf/GJw2HjpFXdgHEQiubHvapIHb4OwMmqE+HKlawbFgr7H1hslWt29TpcsWGj
D2s/FF8HxowbHYqex4KcA5EL0BoY9SedJ8P3qU+vxv3sGNfST3PajhgnpuwtHfY4
27hb/+X3mAVo5OOlcn8T4TRB1eKNUD+Yc/V7MghqyTnk9OX4YwDAA7zMw4gL67dc
pnhHXFO04L7B5c4f69Xu1F0VkSZcz1mkQGtMUZcLy9h3EQ2CpY7dJA7JtrFq/k87
HWWtyJHsmDTBztEHSP8fTqdoOJh0DuiGVThlrh9Wvai3xDrwsTfLR0Kj6XefIH/a
knaYi/5YP9WrWMP502SX4GAOSW6VlsMLerUnmo2uyJAvyterbW8/6Ut9fW2F1gOn
JIaAuaWFUSkTj8IIREZZHtBw99sybBvGiflporc1vKJJ0qpzWnEqwvpC2GflVwlH
9xbMkuwwmWTJDSpodUu1JX0Wr91n4UjNGBY6oobxabrwP8Ynck/uamJJpmH7ldOX
RybI7AerzGW9vp+Lj7ND17tH5kGpnupTHC4zFYB3inI0hcLmYoo20ELX1oGZPwEt
EhGw1K+nTXcB/a+p8N8Nf+k4tf7r+A7UW6Alga3/rwQVR/1GS3nFTKcjeThCAVJZ
tD41cUjtB9J0FyDOi+qc3zgAXHUt/x9AhdY0qLfdhySKlFtudpc4+vA5wShxmdTM
6YJqncOJW4i0PbOuHvJ4mHpYnDCK+cY5HbxVFLay1sWRtT1TSTGOYm1+Zo+Xg80u
ecw0ZiHfJiYK47S0VbjG7XEQuAGIuZYQtFhabvqS3H6h0ji2USVZvooePAHG68uO
s58at3ycSD/djPJleaBlULGHQc9V0voN8Hxd0SkUsINfgPRtW7LXjDq7TtffU9u7
2/kNYMhXVJ6RkGTGyT3oH58UPweVf+jXupo3CkbCw9iR7Wfi/kbDMq/GeP1fHZUy
5Fwscd76nIuiiLtT6M0VdMAkou09LsjUNsMsO2JHba9GQiMk7yRYN4hV/s3X7aPZ
7mC0wHmcrQk1peH6y9Kw5iI7QIxplcufk22AHi0mtV7V5fPr8DrHFxdSa1XmArkW
t55GunWUQmQbQoTqQ4syOsa9VDzB1QpcP0rf8aau24Uk8tqbEKht5LDV+GM6lxJx
pgOI6te8wX6YURz1M3Drt+chkkg960S4qIe5TyttVgeQXltM9WPWkw5EapnWARBw
bp6IWO5JpihH1EMZJPeMa/K4lfHOtbgphZwLMuTZn02M0GoK1qNYQGy9LqllLbks
XDXcm95wsyPYdn7ZJgA9aKzCaV61tkAJ/Bd+ZQBtTauimmvHx8v/oKEWKXVWT/az
6xNSM1JKyxCFDNPfAEsneMq+BlI8HuxfGw7g4pODES00GQ86wD83OTEUT/hz93Lk
ShdK6SuuzAAOglJllXW5di8DzFqvFjKXxl+VhdyHBRwxiC+9aIEMQ1+17rIveo4M
sBhImSHqL/PMB84iOMdTLof/W1pDRiFfxYWjvUk0IWk2d+mfFfyxTuvHLXMFaP6p
fX1BlPGEWj96xV2nKKceKey+8EEatQLnw1VAuNS3OomqRMTdX7YOq8RNJwDrHkHI
Vw7J2S9q+6Esf+Les9OxXk/9MmyxQKonIGrANgV+0KI3nYNaNCbPClcjY3sjTitH
eYeAVKc4OD/BPLbqWRAJ91kCnu/Ik8xms8DjS+mgWjwCBi1iBUyPrx00jUekBcVS
T16n1xPPpbNOevIquW0hNTatOjYKjf++fS8h3Z1OXy90QiNavfIFhPFFPV4iiabb
dF+soQl2UJ1oxUzS6NR2eHY+q3XCqB+GCioGKN838H2DIcBVdPHTk+hiZZ5GZ0Ey
6vB/QliclOKn4zP3oH7Ob2F8TtaNU47yIT1U7iMC7AbdwJyk6QZuZBaouQVf0McM
VqSOMaK19WS/HtklIgcefNTgHq8JIeOQGf8u76H39yKx5J6fJR0AZJXBnsGGjuT7
Bx5yBFmUieNXbB84FvWO+QqL6voEnnplnvmmCIioa7L79mdf08if4ReXHds9byRx
5TqpmPG7dYf5GJLZvkZ1RnCXV5yy1z89g02iuLcFLjY0i3xjc9guNyBhtplYOsnl
Q77/uUx4nUMbOt4LZyCH42MdvEWEl1EHpfesp+UkgnQbSN/QH6/GDdybf5jshJGH
DcfPKZUIDldwX6GUxWx5qhnsorDlB/P6R4fHd9z1Y9ZC3u9+Fkvhf+rrbzXCo03C
v4i6ZRnuPU2XBLngHxt+NmFeW9Z1MC2n2WlMIC7GrAcjqD5Yfo5ey6r/j6loaH6p
/Gy/iV48nwNOzy3eaHSDlPilZIslOwb9xEPK5fDiA2bFS8MlNuhAMwoGo2aOYMDf
IugLAhoL/uUDsYT7/h676PU2JxwtUE5qoeHBrWuhV5iZVWQJ20CbpaP0T/+rOrNJ
1akHXQ6G4cezMgDmteDCqc/DM2ib5hboIMObH+yGM6sPsFZimrooy0jUfZTF4Yal
/5NpgjNmPgEHTAUxVU/aPpQfl1PlkkycZEps9lKz2I8mKqY72hnHY0hGWSuBFego
OuxOnQZ2+ChOBZSZEbvVh7LlgJiGs1N0Vb9SkBaY1qBIg1BM07c6P5d1dh/8XWdD
LZiIkwHTTvf/sBARf+77Xe72taxhrEeDZF2bsPwxJJcyEhZ0LzT3czlUUOW9WFio
AckbcHLuVj/x6fRbFiDmdna46FLybmkpWxTHkcFgIqn0j1fKcpE4R+tFccau2/TM
EjFGTD1e4tGD4buSo+siHmXHZl86a1RTWwKdxrmjEbzQl8Ew2Xjg8X7xkRgqRmLk
E80x2KEXnms2GAxJVxief1ELx817daILY3q2Kx7fYA8gmXcZNneaEVmTdOb3Er2d
Uk1qU451RlQLAQRmabqt58URuHcQPd4CezoYmn1cM0q6gp2ps3Ean94n8G0Mwqpc
qivPsSflEdjyIlffsrFrN52/xmB2niFmmNLv9ezc7v72MIPU1Z/62CkvdsxobOdf
Ra6ZRf+kNDkn2/BZj3AFEp6/JL8beD4/T8UN9FDZK6MhxrS6ZTeohcUTo4Egb55Q
CSI6TLrVvfDQX5Xc7kM5B9FVvVGqaDcAOrcMjNecx3oiYn1bfCXNxq8ckhmEaxGc
Cg/0NScm8H8hvy+ikh+VcWZdZZQ9VzZuag8s6yCal44XMkEKLAaFCcnqlub6NuYz
7VKW++Wchae5haibKfCdE/yCWtzdwm+XgMqCiAA9PalDXh4C6ST19hwiaYV+OChy
bdVrJfcdZB71zDlHBmlcfeHXUHPX7PshqnxcAmaHdh5Cx4LG3qCs1dg5DJrW+20L
F/KLxrZsfFNZZjSJLhkIW4XDyeFYnvVHeSV0jbS5Ux/D6vnqXDCJfPnh/+JT5i9a
Sxdd/AGLueMtjdFLVt/U70cb2wdczBCQ3scGh+5cbuZC0OuSA6FJa+nHgmWEAKjJ
Kly1ucZWDNys4W9UgDGO/EpbWCUewFlYmd60hDuk9aPKRb9Xv40XXb/MOxa3lbHx
J4Lu75PerlT6eEF7sy4LXVuOOjPWY7VXJOV8K5ue4qgjz1i3UC3DYP4Yq1q7tFxW
3nwALkoyBOSzn89BHSNkjo2oM5wENQTcoG1K3fAfPeriznMeQWgVuCNwlhfnXZ2E
d7/HMIY8o2hdBQoa346gxnGOSN/UQ4D2IX7K7RMocmhBvukOhdXgVJdVgfL0oN7D
1wIopEvEoUeXa6MFsEBUpTcvUvV8yBxWq7yQISaWzf6WfWpOr5vwEHFKNFQwejNE
gzTTh8JMbQ1172DmK4ToN1nx0Z+xR+Sr3nJd7wiiI9fWiJG2UofNoncF65PsRcsT
SQH1+rGAYqec/PvGYTZUmYOG31BQyzkijYsRtlTiwTGIPDAP5yLYQZy0Y1FWgJp/
i1rVyWoDreK1+64r6/sNjOcvZvEgZAXq8aRVx9TmzD5xdAMGcdQ4muyc70wy+HAQ
1Khcsc/1eGXOsig8EkmbyQEN3tK3334rJsHkKgmV8j1qc2YoNuZs/fyx69B9tFL9
K6AA71ZR6f6oU36XaOQJGihCVAELPv7s2pVAv/WEShULUuu/UHbpm+KCyF7WOPbi
0+4y4yYkwJkMnHjWuzT6gprDk9mUgJaz/dg/Vmk+w5faOU423NHRU6ARKkvp/315
QN6GZtvp21jfeUeZraauB1uGEr8AanLzm2gA+vkb2EIwPPHI9DyFgQ4e2Ox7xywS
HajMQi7CHua42KI/kI+g7PcocC5Il421cidDmVOmmbbDLLv+Cq8JEjMmCJhz65tD
GLTXVrDpHo5pjvzCfZNiC5oCqB3v1MZiip1BGCtSVlS/NlrBDZGywD4kNWJwi+tD
9ookJeO8UqDu4zJySw3E+o1LJgw4UZSluglklWQk1bASFH1CwZC9fpQHA9bgyvva
iT1HWgsTnY8z4J0i6ywR/FMiC6lpFRMcuQpl+sdLKq7RmbymKIlotF7OkpJQpyQZ
3NoTdlTfIiEIRVTe/QUTTOMRq1HVoKTcwWhm3jLpLo/f2vdZDMZ6UPDdcVH2azmT
Qoc4rXp71G9MH4MmFyEC9gNqDS9vKKkgdv1Dm3t8PTICvcLQkb5r5JVzFS9fuvHx
DParGe6/CJkvdQHvtBSSkjgzDvX4sFyHYKEEn3SI7AMfhQaLqmNkwDDYASpf4PH9
ik20klenwK8rUmqjfqZ6dSbawRgP77BBwfS7ivX+j1dhq5GACEwjeRus1kKRB5r7
+rPM9WYPIsdPdWo4LA8Jn8uCO7irb1Fb+R7DvSGwbvnPj1S83ykpfg1KA7oSKcSm
RLxmcULGvU445CVs7aCo+mqgNqYAKcDKraiJGHD7yI0/6LHkEFIhfUE/vbVszb3O
IyvW4NDPrPVLfsKvWKoe2eW2YhYbBgJMuxUe029umHOXjUDdfa2Yc9atJeEvi15B
ArjwkW47o9XNRDB75GEzUAToFzddfdvNoyV78s71tpigYhLk/KWOsnh+/0xxOZpV
O35LfLhpTVZv5+GijyzKrxSF8xqc3WX4UY04QZkmnHqmfFQa6YCpyAh6cCnhdp19
MRmi4XOT93uTyL44yEFxsCkwgeYkGSKvSoOXPgCu2jAR3IrItGQr93OmKxpcost3
qHzr2qMZUeqSaU+Py8KALChWnFOIonneG95Qi3lM4YxRmMfWYV8hK6zcKeCETbDv
nvD4XB0Vvr+qJsqvp7f9o7SGtXiqaOpXTp6XSiXqhelq5U6oTIFU9YAxjeIug+j6
bFaDWGECBpbD6acpnCFMsseCGQov89Q02XKT30uJSrZwLK92TnDOa3Tg7ofH+kAQ
xtZc5u/OiiFtaOZI3B8sMGB0/kvf1d+by1NgXUOi8QwG+q4PVKwd00UwR0315Mhc
SeWMM6wRHUPRJmXuj7rSuW7UMVn7nmsXlmZ7M6ooJeKJNn2SGnjY0k3Te0mKSkuw
Y6/Kih2u2ImbzFI6MQF1KazPtmBXdlIY8WdJEPF4M0bnjyfLqhIU68UQrcTyhGfJ
dn2nEoB8imFzku8ieI9QjeuOV68IzKe+T64MsFYHKpzIvMMLjSjMCyZwNKerBw4B
TELw8jmLW0tp9TZUMVaxpSODn0/Lnvh7V2smgtF9ubbiKB/TP3Uadv16nF2hHBuk
GLwLBHoAOII7YTXwzE37b3QeNws7jyt0kAReydrIpBVsxCev/Tl0pnzeZE05O9EN
aqWkKV6jPUvcctjyO2nWAU0fitR10UAu5g0bUuuHBFikFBuyEWqctrl9aNYuWwrb
PLG5YG8DGzKBmMMHXJYMIjNvTYIE8MStOaMRRLT2ZG19pbEQW/Kb5dbDEOJp+2A7
uXHLK9GbLX8GWTrTsePeIgifYGFfhldFgLOwfPXOWkQ3MT60ZoCsJHzBzN1Nq/0f
R1GJBmgAjhv8ZdPhkRtzzTiabAj4v3sbWnIAws+bHtwGSP8hrYwVi3CYVjJz54Ja
pckPrTIPQ2HFJxuKEb0IhVlxK24uSitxCzapmsSormt6dRwEe7MbGJ2jtbf6SEbD
C6QjqMcx/v3iwL82TLYVGpoH0VuF8MXTH6W8hypleC+OTmHCck/Lp2QvpLaDWsNl
7UXx5Rq8t4Pnz2p4ajKNqk2Xwo2IEtmmecEc4/4iI25TwCuzG62AFX8jlY6HGPP2
t93/Ypdb6W+IsiDT+Rdfct9TU5yI2YB9WqFxqBGpqaJHOP/i2On+9RC06d+NftE0
3xcLyL3yM2vmL2DfUsRy2LUuFeywNpaG5azgDPnvsPA5gI+CmBv20F2gTKLea6bP
zaYDun+IoNJYunJd/zR/ru4RH1U3gC5kK1QBFCHGv4vnrz1u+dUM2fweH8OqVz/X
rUQDKAVSNB3EgUp729B1gga/Mv976DLrEpFHnR/ZeUr6GZYr2W/Da4vLxXOUqSE0
OtT6GxD6mmaorcFjazUT3fJTYX0cVQBpb0q6N/pzT61lVitWdGlWOMjsUhGjyaYY
Mk8x4PUIQR1J1NfzAYWMJAaPp5dnshrKmZ94t91SmVAebHrBKVUibpfxON1LlUNr
qti6T96MShmHiB6kbhFtSq/9/dBEi3e2Oxkd+zDP//Um9y5zE6Jxr4dSGhaJ+fRN
i4miB9njB2Dy6L+p0GEN3XosMSE7k4H8fn4fxQjHAIb72v/ZopG5rNLlTKysNwDT
HZS7H6HBstXznKZybEO7xBP4nL9qJtY+KsDXuhK6zVPd+bfr0c2WSCO7FOeocNUr
Y8/S/gR8bVnOgyurZn+8pc1aqlP8+Ux8Z0Qie8vUAIkXrbSszN3HTOSo4Ve8gnHC
xQbf9ZLnB3TUSZ5jL05zZJxdwUnDCGLOHT9LuLBr8jqjPrXo99ycFvGVhHJwDWSg
qYzTzmLfXNrlw6Qup0YCzVq7zjgxhYM95FTgvOIs2vO5fJvzahcEZx0mzL0a9W9r
p2xHwAOK6tiR4c/EZCsjijO+dow+HfDnJP/IVH61J/bYlX8oV5YiBaML/nBT8R4j
nr+/OCnr1NPRoVKNqUe4ahZGyNq+fGa1m0Dejnqm4gdTxAKVfTjJ/sEVufE0z8Bo
5hkwqT4eTSJXoBmndgK5bEp/WZ930OEktWz9mwYdYlXTBtZrqwW83D8gNw4i95tR
LxOEMl0m/1jzuIc0weQLD8Y8nmbsKCf5VFr0pl6qUKOysjb1gbRYs596nX6gLnaP
DhWbQNIn/hVtdJCE4R3ClK+V0jlvDKImgNq7ox5z4q0/zdcBqOf/M0HpdSPKSrmN
z5VC/TNkSyaeiEbTeqtR+4OJ5TvhpVwfZkHb/z9E9l6dE8l5TDuV2lx+PZRl7BFw
qBYeEcarbbTa0M2BlVWm78+ZpnQib4rZcX1KNiULlG7myfTrHckLm2KBZPp9nr2u
5Pvzes99mJyaThr7Xaygya4bATONCuRtDE9/ndd+UBldNWW4Y3SnPa2vs24CGfQp
5OEP1emwuWA/FKii94SS+9R1fOoFB7rAW58iFsioE32O7c3f/Pywnv0CRI7AZYej
QdyBlEgHDhYCqGDk8S5E7Iz9sbs7UYfAEUrX8DYsETITdg3aIbGPcOU2w/2NTRhH
MLcsOhZsvM1OC/PL+YvfUeBx9voIu7hTwGVaG3lrR497OkSTFYuKuoBgBL/ss7Qs
RgKED7Uv5USg44IfoN9cZEb2qImFjA2XRVUZ6c4hC0LJ1fuQ/KuYzqh2WYJbEp0M
Hs/7a6z50yCrQ3DgQ7kOdHboS4/0pIfjvs9rjL1oCpHU8wNL4yioVASaOj46xcsM
gXVf/3pFtwVbjt4cHQK5cypXAiz02cVvcmpGvg0E99BrxIXrf6otYvu+pi2eJo0I
1mCjuaaM9LQBfhkaNFbJCjZKuyVNDZRiqZIVQADBwkBDPUgLAnbMcNRpIS1CwRBx
k2cDV9g5zWjYbM8zbPhxkKfmCbXMvWKCbv0xLgUyNVF7ZZwj73YBLzT0PCLpwPre
G6Oixar2aPJAkQ3iEHBwDihA5zyrr7KKZuIaApEi3LJdmKYMvFe95/xlZJVGarGm
gKBSwPYU+bt/mnyRKA5iWBAVipzRj8qrZs13NhHd2M6kF+GM10c9jOF63kk+HciJ
NMc25xzIvUm1Ck4M+3AFgfJxjmsn6aCxqtLsLSktsdjTtc/sOjPPCb9PzL115+Qo
rW60S1SEBZytS1Il3mbHUe9m/r1FGe4xCi3AC6KtHUt+iFiOunKTDNobTJCJF0uO
YBm6VEPtnOxSoFOmCMmVL0PSn0AUl0mmaXk0R/mFJ9U2jAl/17fNAzzvcKGF7YJa
1/bOLZfwsJZhC5X4BMZ/yOBULhEkrn5kMIkwwqSgdEQKDpvr9rOVMyUjSlLVQT8t
nXL+wgs3KTcbGqL/PqfI4QRcAIB5mJEvNs99w96u1kbzdNzZMgQ7+epfeuwmsAOd
Bf16XYVAji98kVsxCY1JGVXuing27Z/Q3PGw9EV6kEOZjqK7EQBqmYgBp4CZIt1w
B5MD0JC5vCM8GGBQPho4zWnSimXBhyQqPxWcmyNjMv6gb9biRLJJTQcWQlUl0hNC
HoVhhXTX4wYElFkoq4Nv510xWYUX1uoezkVw0QbmKuLGK6H6AJ41HiYA25uaQS4E
3/qEKjMjkyxEZ70FzTnVFUoblyVwWP+ImZAe4Tx5XVZdNMNXy+yIu7VfjBqcGlgO
qAQ+1kLiurryEvzmn3OKhYXfm+5JDjyWsCYJwBc1pZzBmawySp2ix0sOVuokr9Lc
pq414Bmw+5nOf3B3bsMcKFSZ3W/nBzmk7c29LHVW48TYyxY3RcL1Aqvv+9Vm40YD
AbxyUgz+ysHEms/Wffwu046oFa+BIoVE+zdGRX1367DTsWt7WA4e7BRu2IP+iK0S
gS4jgXRq9aYK2lgXsPOCcDOAHu83cRbtntEUb4qt6g0H1Y/xZUsaLQQKDqzcnkaM
z8L1D64RYnNihuCYN4NbmfbgG/QsJrExcQYaCowm+K+zSUzJZ178kmS6ISm50F/o
e39wAbn19zsFgRKfAjFeGdzr/aHTIJd64zCBp7ZTOkBMx3YbtPA1A7bWbI5pzstJ
i3wPPXODv2Im2Fc5R+EIy91w3yLBT4VqVq0ipVpynG8uDkGSzGSL3iH7m80QQ69+
QXJTZsmiN395SZNHi5QeQCuDOYJpS3eGHXFZF+RpTgQ8lh+mLMGM5ZsNys80PPd6
5m+0g+UUWrdIRWbMxN6j8ujL5UAep+E3WFCbdOHoCJE1PqI5OxBAVOgv1DMelZ6X
tHVLBDMyPP+vXILCznhZjj+nTIzii4sJMPd61CI3ASMDgo71SdxbmoJf9vxQH/Ds
/Q5T7+wwOnr0gqi6q2N0EvZjSi47OhZKFUa2mR/ygDG6v2viCioLNViuPKrhkArc
v6IqVeyEeQeSG4neEUfo89HiG1JZegCa+P3s0VBUGl8Vw7d0UMG9eTTiCqnmGr2F
OpTBFahMkWK4Sg6QjVynCNSDI/++bIXp6PS3J3E3duhrZWtNZUlMy2Om8d3xKNvy
YJZToWb60wezAS3qfrqYixAk5X9bhJLXHfIz7d+f8ITi6X9FzcKjOMG8DAYVBfJC
2LNVbks9P6P+lS6i8ee16j9fymBvkRImF+9Q0Vki2DzNmbrYmAUPqwmVZeFYGC2S
5b2zvuTE9yTOS2WLUvXK/iyGo1vnrIyLpi5BWZn3i1BAlWgFasFFdHcGc+nZoG9t
n1jIsypssFezTl07Hgug8rNnCF1pKxGIPTJ5aUJG12KahrpjCzC6YeAWE6MwVXa1
wA5WKhUIqR1KMqMNl9de6GR7GW49bh1T11qxCNeU4CKtAT+ruy8iyh5ZJ6FGY8mP
9aO8HnYEskjeFIIP5ZoOJc72aefrmIXKuFALHcVEYPiTKa4SAHTXIXZ6RxmO+goi
e0VfrLBR46v00iEF6+0qmEw2T5qzEUITGK4qFikkLrNpsrfi3ahu4AmjAPLQFhg3
/rJfCApEXHNwei9hBf6K3w2AmQoHJ+Uz7Pqs6v590j3NrrnTOP+PF5yyF68bQUvE
+bjDjMveiwOmA8BiYcMQaBf7CQ1+/uMN2w35dbXIm6WzS0os0ocZVr2RUPlk/2Eb
YcEjny4Lm2XqC412/WxBAQWTowTk74NrgxbUFMCNnQMJuzQ8X2p/4FeUs71qrk0J
4KZLobdYUoTfCdbZ13y4Zuw67S0I6Ga2rdvwWidLLlynddEPszV79TnRZwieCziN
VsqHXkqD6qk9PxXfSq93DECpekD0Xfnli/MCiaXhtiUkqCUU4u8tSi+SrZ/HbK97
q2lMjpUWkDZ5WVJnlMyM5KZHs1v+F5zu/cqMN7bl04IGZD4Da0wIc0H6Bm0yItfc
3D5m1JSqsAG8fdEs0EIhJDYwShzINMslxazygCiGKrSsc+qg93CrAhKhybFwagkw
GeOCkxXez2QQw8ruPYlbzU84LTkTykhvmipsiev+H2Z6wZSsjUT+teAmjA7ZIOv3
JTvygUAXbL+0h+cPVFp83XoU3hP48rdk7lW4BtqEIErJM8UkEYXYiMVbT8/OBzNE
nWsVIq7J5Y3LzLjyPn6LmZokbFG/yhkFIQ10L1Zc9P9fzmehzmIQPnmNdDF6JHmG
5dz/FL8G3fQEGjzVp42jfbEUjbChLzPP5zsORaUxQeq0UOiaoFgs0Fbl9j1h0G3D
GEZsKHOX4R65l0WHWryZohGi6daWMkbNhcvknqKTcKSPEvcAXHVMHGSI1fzzXxtT
1YjmgNOryN17E3YEXqca+EqAW/qUmHskuqKHtjr33DwMwhGDkCC5TOwrkLT0dxnD
AWQXKnepYOP/zp3qg9VTn1MK6fR/pRGZTqKE+whhPmOgnub9Bw4/WWNv/clT+ulG
hPob8qXacQZwg+YAQOx3ot+CnUP/ZiOLZnxiwAIR1p/oLuz11GsQcLERedTEaOyN
+KoILxxIfMZRMBGRRMZ4qYWIXumW7xIvIoqUmkbYjR+yMjCXzwm8LeQUhQKM145b
f2dtpyqNVG+Csd65AYoZA/xgcYqRYgGSgaoy69fLQ4A/We4tN47y9UFjwNpjn0jr
Ttzm4/z3MFZphDLbZDHqgVoZ+aB7FWhQxtcHNiowp7A+EjVFYmCnrEIzkyzhZVi8
hk1z5ouUmnX6u2q+ejozRwHkwPstpwpeyNyepuL7sRUITBTmUfU1IBQtOZysS8Vn
mud0Jc7e9ib9LvP5+uCdjioTFe8gU/jJW0MfNaj0VDwJHtNC7k+mXKtBCl0P26qq
r5vOskuo6IDZ7DWWtAjy1VJvKqFVtmQcPsDNv0jquyw1nMOMKBjoKpxAzOpwROQL
S2CFI1g/4dFmI4bDu2CVk3oEMIzEX6ug778j6XuT3sCQTU6avUDEs27Oh71hhfGa
TOm9BpYOHyAJHC+q/kxGvUDbPnCucfkXKUZFTLkQMH3VgSCvnd4GtryMGZXT8Zhb
Xh3OuZxp9TFE9ngDaaWlAiJmYVrJ5hA6sAjw/IUj2Sc/u23jNyiEDM8JZGOPSDUJ
P8aW9RpxiVpqxnoH7W2Q9xSTJ3H44kha6W2B6pVI5FxsL6xG2UVtpxktWYC+6SMP
PqY3XExl8xQOW8y8KXorKdOkRpUMEez1zWpGi8+vWjDxiUzkokIGExpbuHpBSYSX
W9lrmey3GMALJnwTLFbnK3ULjaPcUJB0oPNjeLako6iyLWqpUtvYcc4F2ZBbwVC1
pSApqzPFLWm71OSMt6VXNc+VnirjnUZSMw5T4IVgPm577ethLCJG5LJrjDGUMUeT
ZZOsAnba7FnkSXU1OZHrn7IwCFHkqRmmmmyraRzNZ+6WMWU5pSaAM7wXzVGF+eTy
uo62+DawsCf4xOXH646gbAI4Nwzg4uSOcJw5BW3K8YPaNQGl1H+n7Ah6s86FIk/5
IK7Wy+bVlSHV0GCgRrnJnTppDsFCSdaV/hPcmTbxSxwvaMauKtOYeJX9CZAsCqXv
c9lj5fc4rw4FiIFB2i/KRvNdWH5q1LlGvAskAlXFS2+ol/uciwjr50Qnr3cDUr5D
PXWjz6afsK9TLMcFCFuP1oJ8oiVcEFpupHe4O8868yjwzz/tH+651/3WY9sE5P5D
PpK/6SW15GIEpWeC8uenS8FzyOmehvTlwlRN3RLJvcwq9Z6aFPA7cfslQh4Z2UAv
x9J1bF0uTfNUZnR+dhvOVM08KOxaZaTuVNnQAuSSPEF1l/3DJvR8L8UnsaihyUu+
xm2V1am+jBKm9i+1tF75ivr8F2o21TMBd5bPdrij+gxl/Pu2EZZatCDY1sbvVBXZ
0LEc3v2KT8zfrJd5KOkXOOVt92C6hD3reH2VSXHzbN0rWQBzjERktFi3Moe5qtid
9yjPjY/KB9VLAIfjubDtXndOQf+isFScBPCldzFdBEFqzjdLLMVSmhJxe3NxkTZI
Xsha602g6qhTUCg1Bu46wBFjM+PYyzYTAjbNgFoD8NQUpDx7oQwXzf71ejUKFAlK
HF2ypakTXmJ+0lJMn3B2aOX1hysL4Njb8X5RbIoxUN+fv9Hm4h1TiyXm/tRzLVZo
FlvjpCS57YT4qf3TkryU0OuqH4hXgqsK+GjQ/+InrW7N1DtmjJVl+dcM6UlYRdor
Y4cNzet9HZW5CED+hM/bgqffMZ8gRLXO2A23MjYfpVb/theDJjXmoyb/c4jV36cI
OvOCyuITuuHeChEhdsoAmf/gC3u61OAP5p958YBlh5J5KsLIzdiGUp36916RFrtq
d4rd86oG3aSAXRtPS9B5VjZW4W1orPRwzaMI6UavJ8CtakJAyqDR27mfDNqvZ/F0
Mf6h53CIaLb5f6Woqf6AzYP+ly4tTPhVvUD0IpWRtUjhB+UjQ1BlLU3a/DnkPhyJ
jcdri3u1TUlY5wa/sth9Ran/qsh3Gc0ntLTzDTp2PdzXL8Iwe9/huTsP7B37JXX5
Ohbn0Isc59CsTqjHj0hBgv6PcZMO6i3KeplV+ZmrZuhYV06N74FOJZ32Rm6nqgFe
jMlPgaUF7g+xswxAhIwvqmF8NZgCdFJSxTtZZZMnnp27Iqn6j38KFcn8v3brAbgV
Z4sJI6rLd3K4drah1dAUGf3T9pVuQjazvYZIPx8138VSFAEUzym/p118M56JVzKL
7Q4Ci08iqjb8Pi86gE6JxBoS3LF6SgUk2INQ88trBDO3yophtHigetFnd03FjatG
j7fDQBg6ON1Nxz1mU1aDW6wpdO3kihZLeqjl0U8ilOrfs++t2hhe9gQAuYC7lP4K
H1Fv6xg15ffq11HRuIyWUVJ0Xgr+xzJePdpUVdZEYhjTUx+bSwcCg2Q3oyDfzMuA
VAqdJmGB6afWP6RsQEsNugcKfZCQOg8gKvcMa1TwljJHeLrfyAXEd/TdLmtMPUPd
AYG685bjPvknOg0byQ9YAeHuJcuoNZbyp13jefBg/MWUf2srAKOmmTplHcWXpZe9
7YIkanPd6mlZYMVhKLyRY0Fs59zDeJN/OY0BPp1rheNPX0ZOztwPn65fUTUsAhJq
1foul6XEG5ttRU+z56UmigsPH9PJaKRRJ9NSJlkBoLZitWLtVe393pjPs6C2Sa9C
2EDgTrrZyenfVzjNoT3HyxbOh+sN4Bmlydc3YOxJLONbiaqZj06cenemQZP5LAuy
rFXbkuDPR6LUF1gckgYbRHz3R9RpixwtP6jj28u+9qYH6vTyWKs5v0aU097rOxI5
91V3WpgbF82Fd1zk1pXAClnBCgQ+5si//VNsJaXwXz6QIDXwPbONdLBIdekWQOJa
l+eXWzH6qvxS/M+89pVvxwtEaSZCgH1KkzdIHs5GL3Qu/n5onb4tOn4BPzipD8gs
UWiVAfMgj7DzFvXMRfLVAJjVZNY9tGGypXbz+/laRr8vXkSL5jC7/IkWttC3xfS1
tvK9H3l8DJT5YzsgXBI3fv3SRJN+Of2S6QgPciAZW5jnGjRCrygiYYJLweT0jUlg
1fQ7GFCe2g9e2ndjGtbIDBIJowXliB8Vt/hIRsmoaYAfgYjsxNMTQOFKB6Y+XgFZ
9eELwFG8uZyjt/3e4P6lO1nWBJNpXEnSlppo62kyzMms8X/cc7rNj3J/LH5R7BLU
FNd4UaUqrVw1WmfQaHblT/V9Ou4Ifxrx8pC3mmiXNo+ZLUs1aOd8cE/U3XSGJkKV
YG500JBoRh4z8owHknFVyhzJgcrfLBAFoGk0S2224fGVPfyl00gseYGc9UfIiSpZ
FDhA0F4CD0Nk6mBw01AqRvkOzMD0YessKz60pU7RCEBqSNMzVxhjX9FXM7J2pJvy
ZgMzH/f5Pk6Wxtace1x9Fr6mO2qPS579R96vxMREwNUg9VLJWxZPv76AJzT42q0g
bONzVY0FdiNvW+DxfxOUBruF+VPPlYp/R1694w/XQcF666ewvdl4JUvV9u9EL1kU
cbxvo1BB6FAWSjm9ELwlUirESSGlPBix78RlMjHkYmpBoHZUu3ijfrmoQ5Avv4i4
mdrxgTOYo/Djs0eYl1w0CkF58zKTKOPg4LRmzqc30OoYEWtk/NyJ7a2BhsrJ+lk1
521eXm0Ek1OWVirvy4EKezWoI+72p8yMFkMT8dzR3jJKDQpDVBZNO0EarvHoCYI2
l36o6XgIZdxgpI9E0QHCBrNwvBGBvJoW+JHhD8wb24YEPoHp/dQTy7BBOflt5TyC
hdv4p4/+Q79vljW7XMk23TAfmlQ939CIlGwl0MoIG2kKVSQaBt/1M2xmLqsn53wr
2pFDw73OsKXvrGs7R5llzz9cZtp2YxlHXNxnV/YVwXy54o8sd7q+tnXv2qbS24eB
26OcvOqteJdZpBQfKug+2n6JE3aSIKCqB7PlsxIQ7BeFFnEXyGQ/kH0cu3B+Bfsa
xxlazeP8ycXrM/fxCze4vgGuvusZkN8L5qW+EKydghaomAKoB0YhuBlqYxXiVfX9
M2HFP16agdeOxjrzmhrRIVKzyHsxIh8mIbPu9Ndm3fN6ur7d+IA1/jQOkUw2BtXn
SQI3yHnd5p22KiTco6y8MQgiQM1GYyCxKLraAXSW6gnRBQoyxQibKfA0j3481/A0
Z6xbWzRHkQV1Lmhd0DzHQ37XKH5Xrc721hlhXaZ6zU0r7ryqaRvtanIcb0Ms3NBk
tP0ke31PpdgywD4jVEeIUo+/YSVa4DH2/HG2FXfhgXjPsm0BtcDPi5/f3+6fE288
G92Q4ZwR1+yWx0OleEg4oob3Hhl2C7Cv9ZVLMt57elkrT7JImHcRXfc3Wv/rire5
9tpvqDv/v4xlpZnyJdLnObwgmUNN0fqnf+U355baYsbYZPizyrVZGjTpr+6iflvY
Jpr6cTKUhLZGz8pEW0+jR8OtadGcKuSUHti/1nGQlXIv6A42HspNCV5RfmzP6U4z
FTN2NitoR7MB3nYdLqGEezjRT8l3O8C/M3wwdE69Ob4YEEQSgvwd3TebPLNIVPXK
4sMEqUwVAwygEjWK5WhWLH/Q3zyV52/V5h7wmN5fUOYiawqzApdOM1vNvhaRCm2d
fb5O54p1E28n19UmsZTTMQjoRh2Jfsjt7QqO3+p4r+uDtnX/0KNFvvOB7vSlwDUo
GbXtM5e1G71TOQfZHq3uTbTJnyZaGe3lXM4xgV36n/IIKXPjTyshyx3BCxQIWjhK
qh4oAGZi2QyBAKTe/UaaTfPnXZPkWPSqIfCm4xAjDnKhDfCCWBt+K7GCcVdf8R3p
Vw1vI8oRNMIFMJbQ3zhptjCWUCm1OpJ4JmpnrTdSZIWAY2v6/I1AKsjvPaWrth+0
RTBDU488x7UNdao8wcstmL6BZc4ih3kgDQ0RtqwbaSVosfhGFXxNiqcMQhRs61Jd
jgyTKuDyrQfuGX0AuKYxAicl96PKSraW6//peFygPg6ZiflL47dMD23CjyOc6Shl
CKrKhiB6Hk7/1eDJ/V1qfrLReuHSbyZEYS0XlqyxMjkUZ7j+oPbRGj2oRIUiVnYR
U9EIuVN3Cxg2v2QnMEVfQ6wkU2Jnt0+JUSN+7O/8g7xPv3tIe1pwM3hi9nvCwx/R
CwMkYJ3UK8VVtTiSuwlEcC9mWRRa9ajCT8aDXJofClrZIxPnhI7UIu5XExhJV200
MiFtAU8+CApb1VIppqRCyqmqiQa0TJvelJBFVTIcB6+NUVd1RE5/07rpY8YrecBH
lvjbDsw/q4cuH8fB9JT8Ng/TvIN/Mn68zgIWAzxisSMNl3wCHsCg3snkSrM5uv7m
wbDOFtIOPNG+s6ZBtmBYgRXpWaJP4Y+o6W2CblR/bpp7qbJWFppgjhlmtnI34SWo
KKJahED656iFU/sa7aadnbQYVhL2TJD3bhKU0ym6Iamy7OWBcyhXWeyd7phvoaCp
dX6dOnOvY5OiSok/xFj06TMGJqGSqGLrkavhlOv5VYXAuavkPIT/iRKZfOvkbihc
uy3dbwrbcxQuRbpZ0IrEd5+vi3G/J3bWYvF2LuNrsV0HGHxiyRuOBGpZch+Y6+u+
6EtgUrbz8F2y396LpVviU4AuoFUS36Is4+qukOJ6VyiTv3oL0ZJUIol9kisHsT04
mtMJKY2iyNKgR5GyrgBlT5itCLX7kgLq5qnWUjBe04gOuipN5UlX28ZIBJVOoYTM
+/FQv1qufMY1Sx0b0QT0aiVWE6MnWO1m0OcdO7dYY1tboXyGo0saRk01u37xq6w3
8KUK606vEfvc/+twLS4qr0yKuclbUQ12/oSGeAWP3DwD8Xi5RDSc7y+aq/YKetRs
c6F7JG6i7smwFs5yZ+F2OZspR4zwX/IHh6XUe/9uzDU4Bn5rUnMwCBCPyk2XoJ6B
o7XA+WwYX97XIZTnhjKksXS9nGCuiUW9+Bo5eg6DN34IlyfJNU4ln8cP6vZ9bAPx
W7LLSkXl8RskNPWIGYLLn8wNH8u/v+s5mtdKoI1JcOo5D51CVk/vyeR6x3HKY1Dj
KIWZtnAXxEjyxdmwEyHgK4/9uaPT1ryXkvxa/QwmhFKLepfyz80rx3qLnDVGk1Me
XxZfZsNtUwuxj6TUQfkWYCJXpOCsfxa6AgHkCNuJjtRZXFaSt3o2AeYdq3DHJeND
lKn8CrnublE/JxSXa4E6tyTe1msvxIwKAbnl+usXVAiI5aj5TlXdeAT+IsgS+Y5b
8cFtwBF9Kmb5QNAo7SuQ0VrH0tPecuTYJRHTpdpUESMN8dcnkbz7QzcPtx6lLtv/
ZkhZEBnj5gbddH36RiIrtl8WkW8Nr5D1eeHS+g/STrYrE4w8eEa0N0n3Xhh8v8rZ
pSdlpznN2UGx6ag4b+Jmg4vqBeaCrsg15TYCGaEGYYxvZh+LS1PoxQCYchHkU1nR
u5n7zy83yNlv8fTS70QAcwXz/gXNOn3RUBD431WV1+ZEBsrpH2CwH4oMiKrIZP8x
IBbLZXXRxoC2vD0UwyrCFazML5l987unYHB36YZvKPUZ1xm8kThW0ImBz5FuBCgu
eUosTez9NH1kmTptfKgY845D9M+PW5mFQ3AQBEVCmXkK5ywPjtTWHD77FHaB1lW6
Q4CbpthCIHsQVVmb4TRv96SdC0Z1c/NuhkoEAMK1mm7gxmgNiLEeasLDdl+LB4J9
x7KPfQMUSHroPVl4SecKZDhUUnnU+67ocEu4uEXITpZITz3Uv01ucCrOf97toduI
erdCKoCSF06akVivVKfkvclEHQ5NXQs7/+X5EvFqYLtllQpT06j+D40msHGIy9VY
Hs812yfWA/G87wDR3uuDYIuCHTYZMesvxQ7aM8TEpmyjC6ReKEXine//RWo76My4
2pS60S/+dxnLXngMfMRK2tPBj7TJPN4L3nqwNuIjq/Ad+KbasKPEMr3LA9UkANMJ
hF/pX0A6rGd+uFPHBnLeJ+ucxWXiwQaY57r2e1tNQwVEjRgmVC9G620vCKXfE/0e
Ex0bOWPzFB/fIGqRKUMb5sGYvZtz0Wmtd06aEIY/YsItwznJ6FT3Q0pguOwIL8Jb
Ci+FFmbyXUwH7IF9nguZlE5xOvfmQ6UNP8FQbu65IBbhU/7v9IQVjPq/E66cV4L2
ux6WJZWfV2p+bQarNFu2MSO5NmKwmxtkXoSMCLdAWY4bcfF5vWXO2N9u4Vx5rpx7
VMtvmP9mu8c5phqr1gflv2L5RKv1HyDD9kArU+QfmB6WHBjX4feXrBlmIvIKsCVC
RdJsl2Nh2A+sMl/8sEm22vCtJsTu9Q5celPFDiWjanN5/jmeRhDBemkIGYcb5g11
vvKdPiLl8/bgXwlktJ1yUZR98rCWB6QMCXR6VRwj+RX8ZiKv5xkrDFY98/vMzNki
5fllrmN8tsSWFfAj2ETfT7S7OtA+Jxp/MdH3dudKjo+daXG0VtsBXv+mi/v9TgrS
znwB4vsA+cpb9Um1NLUWJdDgiKXqdsI4PsYHRi0YG+LRt8W63VmAFbisVlxO2gYt
SZPo4r3OqgDmHRYPI+LaNep70nJ0Tw5myeZqT+yQwpPxdSyCx9uKYKh0Yipe7pEh
/bl0/c/2HPq0p5AcqAVrAKvx03gXoHxonuVsjuukotPwYUxZ7BVz6jYb4gMkkiAL
WnA2gfub9CrEcir1zxIaloGrS8dn3Hy+f+9MpKXoC9kLaJF44TCQNKMJdXmjCsbx
FK2Xwm8DkVxK86Ib9+KWRt9yEQSRxZ6egxXRyNpgGQhFhsq1f8KQwl29svOx26KC
4WDLgC5F1JtrPMla+0UzCc+qL20SQ1n0iCHocENYafs+osW54J1LWWoB3g+w1u+3
w/r55GnqYliN1wqZ+//43rg9ZALlJWgJT7xw4a+lIEA5Wit4g4Wl4bt/WDgEmkgV
yvtWp3Pf7VXXsO3gAw80EwnbqCgwiKGA+LgVu7AK1lWUIIHG4H+OAxw1fmC9DHxu
8yfVMjz+nyxE6kxOZDdWLABLdw+1dkhpkjcoSegVYCwOZ+427VGEcyJ7i8XzpOd5
YmbXhcOHFpKAGS3dveRgqB/taSKCiW1dMTvU752waIR3eTVuR0CA42zxIKYF4cg1
kzRQwWL+ousJoat1e24NTWYKsrTsNWT0L8B7uRgSDb0wAIvgFQiugNFGaQFIN2RV
kUQOMkKTyed3fRuy/QA2THryTl8Wlze5YybnR0NBJU56xFla5ipheaiPMjHHC70n
P2EKQ1+FH81YfONTmd5jsVmy6uovoz6R2IM/SLaGDuj/r70bA0Aq5diO8ZMQM/y2
zpZzLPKR4Jwh3bIjo3TzwWTwxwufVpvPUREgRKCC100wXFATxK7VKtx8SwRUSDcZ
izOCqQBXPUWAB+vGLnnMbS6RHxl6JUV84D2oLB0ogUUBXMjZqMjmy9yRxqParxIV
b44w+Hi91e/SCHfLD4W3YUZehZYDrFN4bbe6RNPx3WHYGkcQS6w9Ge6ivSwWAxh7
lK/BeEZfFJEJL4x1Njm8vyEitooXOF6CQYzg6rqLxY36MBwrUwZzqlIXOWjNZNH0
KFMhAh4oA+K10m6T6NkJCHW458WoLXlheAyuBHS8MflSWYNu7xROCZD0/CgUw4/r
6eWCuAVvmxBYDhloaM236Stvwtwsx1Cn3Sn46nfoH0qkPf2bQxEHvxiRNQ+qi+Bk
yLp4OnOTOBAVOjkXAR3597o9bzGArZHU7YsWr/UzVFpb1SFTvWuh0BtLZSpo17e4
IBe/Cj21Nl3d8/GECCOs8NS2Li/Joa77O0ZK4Hz5H5uzW9ZxBJt1IkFxoTsnHG2G
tjXMqEhU3Fn5ZTngy8JDfvCKo+1J7FYeah37oX65PqaZjMbqk/AYgrLJ1CiGjKdK
FRJjpU4jf+900lRB8qgGptN1lr92B/yMwNAtC829dg5U/8yHdTal8hV6BwApyJd6
L9Ao9sZAyxMr+mxYvGMsAIyzzujWvY9Um7KFdAV2Sem44dT6j8pP8YFEE75WU+Up
vY31tXnN58vWCB++Tfb9hLWE5tG7pVUgBUeoPn4w3TMfZNpvL0NW5tY6nj2tO02B
mcGcCtdIb0ctc72Lrs6ETYulyaiVrLFABulph+RaMzzX6EPc1g9Qy1DLdj5s9qYm
U5gHnhmJgy5z5wiBsFG4lPck0NPuguVmgRpKLRP/8chYeQAU1e6XmiNF/WR2b77F
8nJnifqqDzSFYv9bEE9PkNBGgyxhNtD0qUIxSuuciIIuxVcVmF3Ol4bKf9czL1Dj
7NLmBCpCh/ZXJN0WWxjKadTYZLmZ2Wcm/7dpchG38hqTvaya9MQMIjQ7hHPUZkXw
uh+RUunoztYFd+KyxdxSMdLqbPbC7mY3peK9iDhXNnOAoyGx3r3blDlwDe6smvuJ
C/n+j1MckI40Dzeo31fSPOcYxFkI32qPWFGnJwf4E6OTa/ZTMxDF8HPKZIF3nfO9
aA3MVpBYjqArRS00q3LIiK9ae0zaromRtFpknAw+33yjk/9lSIQOBKgFdvN8hnFU
uIiNlblNNlq8HsyPjrU6ZGqjggvxU49l0hpwoXsirOyj73aXlsDuOq+SaJDV66DC
KgngCRr2RSWrkXDsMPG4x5JrvYO2ZsIXk+kcqFIST4+U9v1zBsbLZV3fC86LsWVl
s2xzXvmZhCLe7MqJgljioQBRv4EtskeBj9WOvoArNGDUkcmbtFQQ+tMlCAmGDz1L
Dn6TD7+p6aJ398w1kjOx64HkGUmMuDlBduHQgBxg9jvIZwdFA0tEFigSYHcdBGg7
jLNkCtYLpVD0BlOFeMHf/MK5EY0xxu/o8alXwMCWoJwfp8lzqKZZJXpAnIVGydR0
TwuyD8E9zlDKvkJvwAG1RFsGo2TMy0y5GJl7E6gjx+UD7vwKw8yfPqB4h/SNTXV9
b4FGGBmuJKokaskS9USk6XVZmMu0GE6HY8z8930azFa2Gz8oQac2+1xcanABz50y
npofuKtneUjYcStY6N7jnmviJt7CVAusKeScKBj+mdqnV/5Uw58dK7DdL81dyfgE
ODheABN8Lfjdz4f0xxQJzAftxpb8Xj2mFsmwMtnL6K4CpiTaRJ2cLsqLSWHugDD5
9QS7eUoFJi+7UsNHNL1ceaAcMCsynau0YvxsosGV6AB2cWCLO0+T4/xBymvc1Wc9
+8KWzhHpKVSTSI3AgbmaddvP2yy2SlYlwb39sb3vNR0qnCsF+a8EW8lBoRTChbG4
XOO3Ra6K1sO73ZcavnjTWQ3ewz6lRsmtWwGyaNHKJPG7qxgCbcpA/e/Yl9GBmOkX
rKpWzmLajzoQyiOYYaDm487IDuNz75++QI3WkjXKPpDhQnhfZqcaO3J5VlGmYlAr
20NN3VaytZjzV6HkZc+aV9ISe2GrpQztpNB01n+j9xhRGnBJ98FraKgJI6k5gGTO
EY3m2d64tY82X0UMofNeMHB/vgem9YisAPw4PXB1hqhdATgKRTYhYL/IwfbSzaB7
IBSHNRKmzYHL93/1hRoj1Cj6wNIPSMTAd3rTwojPQ67oCc7k6PYCX2Hr6QHAAsNY
m2YT0Gv9w9Xa2txWvzJneTEzn62IHQL525pUiiZOwkjniVxBEAHpa457vbpmo5Z6
Pn8J9Aqp+AIaNoaA/PSCGyVVIbury4E/OCPOAC2NBuYSDq7ugu4nr1eqnIo7vtRw
Ko1TV9f4zEQUg1SV1gaSlHEG67C1HLpN9MCZjJZxi8UH8F9n541OjMhuiLdYNi47
Puej1bA9LAyOYWtFlAzXTO+JGdr6elp6iq693L3cS5g6RW60+Ur1WfpH9lVSmVSp
qeK75whMQv4+fYVb28Xf1Vru8JLz2isPE5Lv4jcRVG07aeS9rNsiPFMPznnu9kV8
oL1fgxOcfmx1KCnnOnOKozf0CGOVAfFOAHHJX1ZO4mq6cwGJP/vhYnF/x5/QUOzc
/ie2r/OJw8OpqHCqhVrdZAOLXBaneoTmVw6Ro1SffjguM0lhRpefSNPz8R4/WBIk
FldaGJOePhxvTSJt9RQDxHwqeo01ko7lIo1KwI+UkZu436pA9P5wpsGadDRdZ9Ch
YryOTxKIkH8h8+V1qUPOrSqj7+d8c61yM3DniDoDs0IcOr0UAYbrZJTeHdUuxbg3
zHo7W1VPXnixcQd5TwPKi0+HiP7oPl2QE2bb9E84wdlFhEDvXnLGuEGCoy10Hzy6
8o4JLRUgHLY1AqWRzUCVY4yNi3TtmnbXfcY16Ut+o6uDhr7Rv64PHKUwtczsSw5j
HzdGAN6VWgaUIxUCj3px7IEGwKSCLx136iOzHg61rglfUpt/UdAv506SmtxerWe/
sdPdgOzS+G4xY7Vq8Y1gqAtRt7pUb/hDJE+viLAOEKGb7Un67gkhHaB7GlAd9lhs
l5yEfg+pMDDPw1F5EXuwgcgH3Hw28T7fgf/zItHzJsBRBYpdFelYa/MhIlwPpjQR
MAOUm2MhVfQ1M8/W5Dr9aVhQLJg/50ZnGI/jIrfTAvvhZzATWWdpdwzj1+DCILJS
6dnZFoasGJRgsq6sLpgexf9guapsNxuSmcOdbh1TE3RW0ida1wfOsqmiYF4olraE
AShhual/xTJYojK/8OabYAiJWEYsAOi9mL2OTezTt7nchPKYV6NXUpLex4Nh5eAH
AUXZlQK88xl2v8QYigAk1EJu329veXekwFL+lMsLKdHajOMGZVLXLD5HShAazLR1
OxUs8iVrCBBOXqTy8QuNbCpY5uu0A8vZgiwEW3PDwpY4/2OqM73FIKnXzT0xg739
+L4QHGvnDCckqqyQ4rgNmLPnwtFEv6b/8XuAh++EnXs48I47XcHitq+S2TDOqyWr
dd/ykojMSt5fg373DAGgGMYrvWBFMRrK379EwIftsCrT/od1DFvtlbeqi7s5wu38
tyGoYlgiJdj/n0ZiUSSz8BpMJX04ZgNH6JcVrd6U1KfPuttcsbyQH4U76w+VYBUE
+AYNMwszaJ2bc0xQkrm+NrnMyXy4A9BxkbPk1CRIdjk+WIuF37elyT0WinAxaQEJ
ScOISYUXrG8L9+RrUwzUbG1AYACevIW+GKfFCA0iSpcJTlvqghzQ4EQl8YLZAclT
NrhSx6yk8sTTKCAfrba1HZBXXmLj1eZ/d0uRucIkpwh4VJbzGTcjwwvlxSnb5nTa
wQf9JOT6xlkserzcbFP/oKawtIC7hsdvRUU3tUHHmNqzuxwPJysy2MMnDqIcylZK
vjxOZByIKm8bTZeSP3b4zCfEXuhlRBaBqnQTU4sgTpD0lN6zciotzRV9Ozrktzqv
B6sC29fkzaeaY7ozrIUYrz7PCbYrJTUd1idIsUtBkgFoQYYoUGlqBh7bwF3I5bzv
xCZJqVO01fDRS1aWdXmvyRwOYlgq+39bJJze8yzlv00FNG5s4OpXBpthBm0GM7Jk
XX0te5sp0uujsvlxdAlFyvELvpG5gx6DVoazrmVHkTbbv88zhZyFBF85x2Wr3Wcu
zW2s1kkjAf6a1w/8KiqdiVlUJgAQYY+VSo1RQU3Ebh4/fByIAaXlYJQ2L8Maqg3A
FvV8QoMK/vsfPYmDqQrQZzxoFyN1B8N+2Xc5LkJZRM7D+4OLJRdXTUZnWcxPNF4k
0z/LYOozdGO4rpSGvcEUvXIyYzUEHmGMvAvqsIedLwWwEXNvvyNQQiSBLTSBlzGN
1C3qDgoT29gAEhSyAInRRTcsHEytgt9VdSHpo3aXgpOTSJW72ROEOs0vf3+/RhDU
7qS2GNjAvjQwKS0xIorsGq2Onn7SAc34oLSrJ7A8cUkcgzEuanYjoNP36fE0zCrL
UKUIxJ+J29hkyZUy2ChIkmnpn3KQPXn9ItjXABurVUsiNMXPAxJGz8//kJfXz2tR
qDFCz36yuReegefAbY7XupFJLCMmDTJ6Ec8GX6MQkcWXqu745ZGkvNdQdieA6Ci3
Odxc5E63FrKhYbxIcOGRDlQ0wY3AY3polU7soUtI1gbs001S3vrhi2S8YsZBjT42
8cbOkd/5WbpivH9soGzm5FOD8U17/F4Wg/Qvvgej4griznRP3CQ/1566p6mcHToW
2t0ylS6UkPd+aO4abBdwwv94es/u4xoET8mZfsAYeBNYsId4FyXsfXuMaSjHafyF
KP334m6/LvPV/hGOVW/tnY/rtmCYduFP0nEL1VXatqq2RoDALHf0jFHxLQ6OvVeQ
NtJnvYek++Tl8R3HwGG7r3y5jKAEpcEIuxWaBQP1o0NG0r9ttvVSqBL9U27iSt5v
cItbXBphU1kINhiurdCdOetal+WR7T3REEJr0seG/JbBQsFUnSntKvdVMIhc2sXB
FJVf5VfsV3+x8H57HjP0QU22ri/zIHUZP6Oj2u6bTDSCoLfiXCQ6RgKsHQKKv81P
lEaYXMwn8eQ6XIBPzE1OV/rteiedcmppGaERmlN2HpdtCazgmyQptmv5tzq9ZWwQ
QBr6OScuKJqOgtVHHOU+yP6ZWGVN2r9l4MzPGwoOrj4b3XQ2nxwlXz95ZMoRCG1t
nlJMFG9cmjvDMDCGUNU6lgxWwCIx1Oq4rteZff4QqRQicoRE8NLw3y7NhHMV7swn
EC08fj9ueVuv/3lmabHmaSkuwxB+vm69s+GX1uITEc6Avt73g0GPiFYXmfOKQbA1
TdoCI2ttVcjnQK4zRlta4Hfl/ayRZ6A5MUSiRS0iT+XhfkkFFrk06Uy/DzNSf8me
pW1k16Pht+ewChOxj99R7YZLOoCmY27qV76fbUjx9MUh/T0gGKaiOGW8alwcnygW
qy9+Z8nHMRyPbuejG+b4P9qETG12zpKWlkSCNu9rPbArVKJ74/VuCGwy/NMvw4wK
bGk5dIy1hfF01nEO40Y64a8zlGWl1CvJRdjR9p2uj11TrsI3N+qAgfTAOiYSh1y6
imZZ2nr2DnvFrs1jJ5eFuLm99YOwvITdgeYaYvInLDYaHZaTHkFTigUQZs7JxR/e
hCVoO/L6yYDLh68WnGE5/DdbZFOgi8BY72p7W81Hi46vgFNx1fOH1tqSg/8sSk8E
onL18iTL0UpMx6c615o93pRQwV53anRtZwnfDkHGppCnbsrnkq9/7d1XczTs3PUO
lTugCgO+VGXNj+Zd73nENYYWjO56/SPVpsVDw2r12LmsCmf89A+T2JW59KpLN6e7
Ogv4BXAxavBSXMhrWFwixxdpaSc5IMXzXtDCQVG0bRtbArhqD/NxTJmmGOyKYLYa
1SIFZHuVXRVyKG2zPOn1jIJjhuLk/TluwuGL1UAdKcNVCN0vM77JrHn+7DNHJipo
A4mUP2twnMzcRSUkNhOn3pOdhPrmKpAfvE3yObP2qoF6BL3ljpalapNtxcoAMtJm
PzpRgvlQgTAfFjS/t7LfJU50fTuUs8AkFuTkNv5GgbPVWlHopriyQu3Bz7KTjdmO
lt9jzc5d+4LI+VR0+oOE7eUdGO6zizmBxFKMEQ7Km8aDJmiwI8KS7G9mw0hWTKjr
bQTttLv3FCGapnhx3kYEbwVpawMNHBNKbOv0YBlYLs5PXaGHYf+eNOXmwhdFQWSO
Nn7JrIjxtHh6rrKLYPAwfrB7wAGQBzofmz0eugDIfkxDAjGnj3oMjFwF8M14mFmf
U/yNRdSjpyqArjrKh7gS+I43G/sZr12yskFKRoVlRMAdU3ot4Ds8HG9CWUiLL5Fc
SKw5cu8VgIvCclrzGi8/E/12/keNLsGSL+q7dPDPEvqt3JsVvPiYDp48eOJRNV25
WooxmBAeBw/m74GGMLZI6dXnAStIZgCq/UtQPy6jTnXNKfx/Q1QmhFcfLh7Ln45s
J/J78OpawWoPH4wK/E8Fe9sX4DG+BGT60wJSJzX079+7nkJv60fuhk3K3v0Q5W47
ZfQiClR8RHRmOJxJxKzjDbafD8AgmFnoN6iVHpwjAVm2cc9sUXC5kVcPllQqUifh
AiM6OtOjH294G3ONvUrTSISnCyunJOr/Y+IKG3ArROnkkFsuvZo+1CoqW4UnFUX5
/PXYykZRXCtuqRy0EtosH0HFCGmFbd3w8e6SFiJCTVRs+f6mkC8MvIWpfYbwqSJA
gB6xQPurXemb+iRos1l7xwLrSXm860OGLFSARYXUNDwM4BbFv5hy+y/At4R0vuN4
TMY9UUsB63lVtYweByO8BpI1pfn7oizhsogx5nvnIkRf8pMYjgqNRgl3qTWgC9t/
PyDjsgcue7uDYnmVS5itgA3XGs8dXE7RRV5RYgDASsiwAC0VUgYUtA24Tr3186gf
cEL96LFZvNzjjTkgjNfRxp1zdDlG0rDHVVgE/4+USG/voNDHsxswxaase+kQ2Nzi
9ITH+vi0kyiSsfzD3bctUmD6V80oNwKwbQ0Z9R1mKY7vKhEcAXgG+AN1nru9xwSE
fW5gEwn9FlIlk2WHzGI6vpShPLb3qrybFZdA6/fOsc/z1kml9rfvAxD3texIdxex
BCSAeqOhRFRQ3k8Awq8vY6/CFaV/QQT9g4OrSq0fNrcU2MzA+znTVUOcoSJ+gDYB
waak7a6WMG941QDCKdMFBezQ/WHM8UFnYT/nEJiRAyjtgIgFY0C3lszeEvF+nJMo
dpg24uUNoMduHKyRozIADgMlbFT8Kwydd+Ce48zTz5qMDAdlk7RAjl2Fide9P5hK
OXmKdu7ZdTBjWxCjDbgKmITi+Yb05ALF8uSBA3rev5HcJnaVAveIJczny4ZIGo+J
rlEO5eTRcanMk2Iz6aviGXx0z3fl3lQUqhtzURlYUqmUtTKLiLjElzEwYN1et6kf
LltGwOFP7OvGHRlbJRN1ZkV8MQ9O1WHtDG76ZRr8H5c6HnIRFv8GDcxHxA1pR+x1
VOkbiAkc+qPIm8iaxg2TWiKgu+T3w+HD6kAb89QdYVGREJO5tE2TmnpZYm4OJfiS
QeMkQXE2TB2gMIXV3ytVB/o31diuBkf8n79obFn1ikXw4tDq9G4A9VXWgK1DTGoK
VYW++d+mVt/v5L0hpB8p37t1SuylZshSOApjP/SPj0ikufEXyZ3nTNTdJwHOf9P5
m93PRUPbw25Tek3SrBlfgOqewpA9wRMIGNie0MHX0CHnL58ILvVkdfZ65OHTzO8z
rWLGT4F/jEciPGOB6PTnp01ZfP7a6TooGVVSJ3/wYy9EIYwAF+yjPieZCK4mQ79e
+cN8ZaalOiRB3IypkllXx5r6ThVgrbm7sCnuzNddsi+9fHCzMemmkaN6VZyQC5Xv
i+1UoNaBoKB7NjU5MvOh3izRo/8NNYsBAIlW/zubL3g4PvuKO2IraWjfVOAg+ui8
Fm3HNGznZ+lEZl12aO3OkY4jEQx0o3f91hHB5ezGG18FpKKtXzWZ77h2YP2uik8o
SuEF7KSp6X7jEtW5KAmnR/UVDBsuFcoVSYbqrR6ZT7H9/ZGONuALBwjWj6hyD73l
PYpbMEEvv2dcfosP364t/fgQ/IuBU4qezigH0RiGeXNRPr7ij32vdQuE2leVGbiC
jp24AU4uL6ZFlFTKVX4NW8ZzADHwPAj7SlJaayh0Gsy4Bg2YQkuzAaBy36ZhHCKM
fpw1djuHQWPpgU4HYtWDwXfJGt0RKFgzI7a23YzUqIozozEa7ryYGt9BYAqPqr2i
xdBoQnx/d6Gq1OKqtj1znOgpOsG7JTcrsc3wBfIRFg4xathZFWjq1kj6bfJqX7Yp
DdJ5GK9m8UHVWQNx34IG88UX4poVe9ayHHYFiChQ4vnchOnccqj8Y7l2ZOCj1bAf
x8J0QfHFyyoi3KaMPegbLCcBrj8qeictvbH7EKLbkyhdnDNcKsKoE2NloHP5KCWE
8ILRRlhSVGBtc6GADO7dON7/Qr4l82wzW7eyYiulESZuSvLfORLEXINX18o8vbAD
LfCbUbx6opWqcxuOPetfVBb5X3r3RsjOFJQ06ctTTaQ/8WKXiv51aNJJHsnTboda
XGup/0aLG5WBOVruw+fp+RZ2TPKAthmUoEgeTodGLrxbHXQW1ayTqopJX8YQKsCJ
xdvM+k6ppK6gJUZq+1oMu6A+OyDzbzWg9Q9IhXxKNM8Rgw2SJ5IvTeLnUeUp6u/P
7TAdSkl9VRkW3AKPus9O9wg3YL6fc+L82JUBofCS/yv0nD6E5CGjjpIS+224l8Z0
2/rgsy30MffcVcUp+acEdOXuBh7MSUBewdwhqIPADqoUc42kn/59x0bVHeZrtrN5
Jc0YGNtpzLgliuJwtzQtd1bnDKjeHp6K51Yi6G5eyR3OLu/6/sK3TFUD0+4B8BRz
JeCpVdinbO2bptwKjyXTtPZ4SSyGaaTTst2sah3GCZHLHo8r0E3qkAou3TSVbVPL
qb+oek5K3O0wFSzWnb0zbSCo3u2hMJOwim2nVGyCmvmtNo6SNurOB/wTuY4RdcCI
AAu3MtFYgiWNLhzRFLbLkWL+wQTmyBMuAm0n56ezVRA+yAIzGyfHw70DLkBHG/P8
qqatpNn4qec0DkSzV28vTKauLtzYUcj7qtNY/CHl77vu1LmH8zVbBWQqkD6m5ylb
2/6WeSAv0/JnMT85H8XtvwgfrgMvPIHoS9P9n0k50XVe0rYiUKJ1/J4IT3drU+Yz
UO76Arg1yQPEb3/c6/dVBcnZAye8ON3gPITwwQ+O7pC5JNMvAvF5+2djz40cTKe1
cliJEGwIMT+f+CAMxTAlpRR+x/bSH4cDdEzHnTBHer9iqcnv6sEsjc4V1i27fdA8
eNT3h1Ojg+ptufEKe+FsQWZE3WpNcO37JlabBEhWBikxMDahjppTg63vHSfH2gd6
V4HLzI3YYP77cnWaLEGviEqYk653UUQU73QNpfxd0AVhJFJhA/OI0saUu/kv2cd4
DzK3VUkl1qxM3Wuz/FbGLt2LINQaURbjhzBsTrD1vW5+2MailyyPnt7t7jSIiGes
W/mCJ/qp++cGZE5B3o70Cx9kRTmFdOrV7mB9yrPAif8VPF71rutOmPCCt1vOrAPG
y2Rqw9ezVsGJAl7fyS/z4MA+zKI0NPW4HgVo0wR8SqIaCUw3N5PmGY/2TdXPJyz1
DBEJ5OvKU+5qCVbdpPBIJA7D90wHqtGhvGkH9LDNWyC2p3M7Q0Q9Yq3UsmdqaTEi
T+PAkd1GEU8VKe7KDGheGVDXBnaeCYNJzcgDGHFgMRpvUR7fXqrYtr+oBKtQ7OLv
Fm+7aQ1RTfB8GRu2Ez+FyAyHzooZ0BZpbVz8zaTUCeg39AmqgTJBPCGxPeiBDE68
gL81dXoI5N5X8FVQpETqOC+NoY2ztHLKcNE+EsCH1UG0iTWgMuXwHnk7aaFK0pmO
j1SShqr9+ImS1w0noXn/J0zjlG+c+GnxAlkYmW6pKGvvMmOz4aa5VIqJDK11/GOj
jGFV7vqFtDMbFE9ox1bd8rrec0HDAUcOngZPIOPiqkjT9ClNSiE7k6XhWKrAEyRg
0cMijAHG63goiSgCiL4cpNhSxLUnyX40mQId+zVpsFUd1JNglhHSqku3OPuzRiAi
4gt9QSKi9dtFpqc9QDWdP94rIMS9V+wUIdZf/A9hiKSOWFuP0aGfhK4ges8xVF+r
84C3M+JV9yfGb2uKpVh7TXa2cMAGKurYsJrxpmIN67Ocl6JLaIUxKn31ReVw+aB1
csPSr7lGwXkWO5HUBCqa0vIXZw+R0evrtMwr1Yr929nuPHbCB9K35jVf/Xc/n71z
5EiuXsD5LCK5EcQPO6z2tUS3vLIdVNGvN7q8Uy31h7SVI6MOPS25VoF2BUS6iROt
OVYRMzP9kYehZnuHZZU0zRBgR9Zdordas54ZQT5sLJvU378HAx3DSgfy4mvRA3XP
cQH1kXg9vDZID+Y+NMT7wLJzJd6vBFPMC2r7X+Trw+DgXvdyD7SQOlhbqnuCUo03
xzncm07U+YOPiUxfSRWpPLua2vQcvdfFxzy8Nbt2e/+2ZUn9xOty7L+ANTcYp4d8
MUuP0oATjB24pBh97Pgijwlf1S5yKPVr/7/bo/fr6i2X5lTP6VzombRNQ0mcIIzR
zXw27Fd4t5HXhOUeMWvuoj27HvMe0Li7hqrzT2NZjrOuLKHlcJAjZNqzW4Uqz8K7
VakQFOIcOk6ZTUk/Gt/NIqkM44LZNx8Zw7RtgI3rdzLoDp7st/fYqUaTtSt43mUj
j74Xgz5dL2fyXnDWIEBT+wnH5iZALxhDFqdhigvSFp7JbEjNJEhBgs1dgj+SnYrm
UPe5XvFPjsZhEq2/PJDBrwiqXQPKbSMWt1yKhMMLxoDsC6cMYWdnk9ZMuy/LKypj
QTj74+xj5O9NwB+0LoRB3D5nwDC71EBFltGhifwKfq6rTg3oK5cmI4udASezFdQr
QlPeB/gEZYNRV0S6iR8zEdkQSmSB9TKCJtxW37GX5oWGrQJDuo0LtlFWHy8Mdxui
V+lzeciK7zybD1gsOpPAMCHuSuEuZCiPJPWoAwqzLZ6jA/1ZPmf6MsDERCLl5xhh
ooP/sNTpW9d/jTPTbuHfsyosCcR8q2UnvmJWgD5JBmwDoqZ9BK//w5S6VPKLROWB
d5cdG+/M9XGWThTwJJYsnDxiPuQvHfp4tgLDFW5PE0bDetr3R4FN66UKShOUxetB
t06+Em1M37kEpKN67ejF00gAt3RD1v27VjLWU14kqFeq2V0UFeT53rZRGqEnkYkN
kui7EXZUHi9KuRHJu9y88pA77dPH2lDNmnXxL+9JhOGp6tfWtNTujv/L4Fgq7X9c
nTIyXtvRIBH8UvtkN/qSvVpdP48RP/kmD3xECGm70W/vU80htGeV9XgnMGY1Dh/H
UqlsxgIqvlzqGd66SyiGe67a8pVhFnpX4MiESkmg/1dJ0LlFbyZliMttvBRRmYEn
oqGlfLQowXj03m5b5e2Fo0qzB5/yW1lFlPCcsAraeKXxstu8IYByPdMZJUjNkN11
dxW+l55EV2dR9i0arskxUORVDy44KiVKFix0K0yxJiWTQ95PGm5E9hAMG7Gb3vKT
Bobi1m3CgFutI+afvkjiAK4C3zH+Byc/fMSfmdVtaTZbCFgb474HAo3RLITqetXT
TiCOX1XR44RLEhBqXLq0c52ZurlG6TPNGyCFwbX/6L/Nx2W96FuJNqofX367q4sB
oFUsETGlrbeVjrmLkk4Sw7Irb86M6ANkgSmEvzwQP8dkragkLjcKIvNLXi5QNGVV
ZA2qqwr3ucrwMhivVgErFEfb5/lSMX8F8dUExACVrRzqzNygasdV3I/Iw+llGHgK
Hp2VqTvPGjnbijTpOWsM2pKZFlyWpdt1W7/9FqyWxBzpwpuybwE6T5KJWP1jOTjo
UMquaER/gJrD5hzOOhjaj3uBci2H4/zlrfcMNys1r1CtTleahv254rCM+B7uXrgz
uZCRhGi8cHCwxrIeDIBpnxM/Te7z71HS/nxi/cELNW0XRD793hQ/25PJSiP4r86D
CmHzGoYWcrfIOvEBWQQCaidtpso0BZqfcbZHAdyVWfReKbsxQBS1Sz65lIEFKAYK
Llc93TYXt/FgFDlLJjcwgpx5G/8pplY5ILzvlj+biwnTtLU/eOWnidEZDA5sYILd
y+Wiod96dPeFvgLuePAG2+iz7gRVN4Xh3RxvizKm6c8FweJvMIEG2Op/z1dhLTd2
8KMmeWJMXvgl76p4LS2und68TGXzDx/vnj9hLvULWBFBV9DB1yowuQHbIG94T4+A
TosPKFBPiGmfmh6XBbArmmMenpy1WUufxDnfK/18GfiEBNAE4LaMeC3SzJEwFyfX
HEJml5kj1ZA785mLMIizwAo9yKC7t6M+o3OTdCwJJv4Xbw2adve91Q7i5Dm7rkcx
xEFX4qPvjYM+FbIB4ClnqbIXalvIBl0KAyFEPaXFmGy8mvw3LRv72NVBGHDFp/QW
lRxs/bcy/Q2K64dIDL7Dq1ACsrxZc7bB1G2ZwkD1X4YYo4DHdGaGNLOYkNv3pzVR
rjC5a3XRDf/rJCNa5IsdSi+5kKNxf8sNwYOaowSglyf+9j1BJW3XyPVLQEz6224k
PBGZ0bK5CPW30VJCEb4OqBbBs9Uzm8mVtKTp/3Rrbn6wyJV0qYVk3MfyXPHZB5jb
AJ+Kw5Uc1M6WnGxotig9UYyqZcPP9dXhg4dp2nBPXSlPKjL6sbB/2IBmr5B9pPOU
4HkXAallfFNPvmbom/aSGpAD6dSuvx5pSO2TDNm98TC2keL3suN+kSjbPJJGi66w
rhDjwZXmVjgO8zFwE4b9onvVAmwo6fFdCr/okWPcxZ0Q5y2wu60mU6UO6rpzC9WU
kJUo9K0nn4bjZFbgtKqHmG8fyZuPtJpF7SRZBmfU+VGIf3Kx/YUyRGmUoOqK6yOR
FH+Py9y5vhupnaYK6r4ijNMkO7Y0rymXfLTKxBCcaNL3Qz2zD2/8dvWWML/5ostn
XE5cHCJ3LPu3ADAwt+v//oN/8Y0j3cpuTWgbDPVSaWCPx10q1LnGF0XVXu4kO0GA
3mUnfO4SApc/2ioldNyd6h0xAyIsbvmpD8vx/G0TLLKeD6ilKhoriog272kjb0Vk
8VQUQojUkJXgAlGnkvIGSN0jDDngGb0kemHdaNDQz/fgpVEM1kCx3LMbJYDUgvYf
bHl3ATKrH+RgVPbdcMUZJZhnD/Nils03CbVfbaTBaZ9ozMLr++gxZ99Fno29yqVY
DqyQSgXrR16PuPgG3gSvCNkOztfWFsHtpceJLDdxeoHAuIig/8CyoA+ZL+SVIHTc
NTaLBtaIuysFkHMh2QrAu4m+3eRHvPGtRT3G7rowB0r5NiZt8qzQUvBpPn+WxiLv
7/VnkGqDO/vAFsURht67c4Ja1pgRdRDPInMp3niSqIOHTtNCoEo2XiBFIte7JtOg
5SN8NBnaJ2GNbUsRbW8FKD4SJIcyhQsrl4M60HEhazMoXxASLocQVsxwFOh1Ty1G
sZpSQCEIJRMQwwieSulnC/hI5unDVlEx35uCKKP3vHTNGCxUPX3y06OTe58z1o+g
/eM5WEdMS2RljXaVEMZw9eovYEBOTqKR/DAaOPjAOKMwaUfZEdS/SsHo0EnXF/uj
bHNXW7bltwkJKa9f/XgEIO5EJYjBDH8GxQdmKFfVqV54X3EA0qZmNspvMku8WIFG
I37c4IxOxUBzzQFqiqunhWeRU8xz3ddNQZ3uUzhTMjf5U+WL/1uBJcpzV/jrvX+2
xCu4j2ziqREynhhBHzNHX1JExIVSso4k9NgWSpgZiNd9cwyWuxzZCKkJNIIPXVcP
c5ilX708XBWWVMe/E4f9L9fnCGikeSqHgqx2lbyyOhSHKEsrNDrM2j67G9VoWKWk
qQuw2KYSTe9zSLBdzNDKvgJRpi/GoVA0bsZ615GVPZiv/L1p0uX33JSRUQoEQgwm
l1ZByUo/IwPS7jPVAksSbKAAetoBSYvJQbYqyimKmhCUTfuHRdBAqxwCNarTQwTQ
n6oTTP3Is3vHkKCdFRfFfxNaaQIxXINu1dqOSsY07JM+IWnDCNSPnKqi+DLmfwGO
L553zn8NpkAyRvM9WiUWwH6yvqrRUkxrkhO5ScBju7IAb7m4hdhLdDbVZujzTFc3
LkdVVGi11DDcDqRqGPOdVrARzmF9/LKt9ivKZXe9nXgv9P++o6cGIoQuTsq8dlKk
NgruWBtrTlyTHLcV/fXTlUlrrkULKv3XdMU9PzMr73rDPTyeC+dgD93lntgMF+f/
yp3YxD+ZA8crik05TUuqmiz2pwPR8GNGqhnJ10ZvFtCWX14x+c93bvp40AXqrNLZ
Hf7yisOJLCVdv0uWZYaStzbb/aCFja8PChFs8DQISdDq7BBhpg2BO2yVV6Xx5fAO
EtjnLzhFEO3XjesdpB4yBajhECUY7sJwl3AlQIAadkoOvzx6DZc9MTFbQDwIVsG8
e5rWitW+yXj2qCaOsrFgXw6uUXx9Jbod7bQ2I5KxOBZwapM8+fjj3tNOb+W+cRBe
2HmcYuYLK17xJE8/eoNd/vVcqiEqpBdokSpVecuid3rkVcFgWtu6FqBBOgAF9R5d
pOpFMiKKPRW/Kq9P/Gu4l+jYO03NNra8O9Ae35puja0bVnnp9IweA+9BJNPxyt6a
WVicbcKsjdmlBCMeUFd0WKw2mKkuIuAipCZBFy9xaLdVUXq0BKYzXTUnakecKA28
oBhqepfDj1iTua1XpHRpqKMDZ4kQQ29BvpTmOFLWx7OEZLZwBEsBZlwXFnWt4zA2
hJlDKxMI2OXpLXTIETNXfgcfxsdfSGvEeBtYKibOSvGmVlRQxRq4FoH3NC1LHiL5
Z7JRUtZgIM9sbYc518TYoYGymCkXSxd4P1VlQR3DtAzQipjUV6NjjenrCym4gbuI
eSE6nRFIjdoVllbRsM31PkGSxeGQ0EoqR6ugTDJLXjJWcMJH7Ntiw/PkZm53Nf7h
Pou54yQA2LaKdVd3bRKgLPK9eEYQQ7xnNtNFELAUZ4t0pepeMvJx+FQH3l/qekcT
ScRdAPFgBv2eecKErfoQoFLvLI6SWBTx5gYoniTG7+R5IOgTZ73P2WWMvVktvws3
8zTt81z3K4kJ6ctz2pQVOq9JZEEbC1C8I9kj7xuRU3j6bKm80hGxCSBaX/UubQDd
vYJq+gCc49VnH7vOwl7yo+GeTWgP+4P4UaloqrQ8mmI+voZCdffnGurscYQ0sdsJ
SLPivhrGHhdM91kR54dFZaTTu08Lqv+wsPxvBiLdj4FLtiOUhLPwi6OflPn0aT1d
hgjWqsZhGATwBYdNjkiA/g+iyDw3HR4F9Sho4KYc0HpvO0hK4DJJ6vSz+QIunm/9
Y0JmHbYw13Ii6xPMclc5YLEI5BOxxLDpeQ9sQz8QuI2UzYnfE70cSFGOutd7lHtp
Wl6rVcVsIBaG/GrcV/FwIKWbl1vUVrLrBLutno4rmnRB0XVFEldqyPunqwIqT/wV
H46h+5yCk6s7fM8EVIVMri8mWsv+sl+O1Lq0OGr/exW4crcvAhjjyf2Wpa8JvOqk
E+hLP5Z1tOj2TbLJ5jE46hX1GraKGkpBgE4tru/saiim5aLw7uEmxW2dXwa/kkWl
1s87PwXmtsxhSwhOrQ9jS/7nKM+2aqN1kQR1W+XCylEw2NlbakonvVNSR5x1ipCc
Rh3FIviWR5naLAD+Dd1yj+X8chGJJiD3f+jK9Dtn2ozUhoHn7/xzonbeIEjmErQ+
pwTJL6SJ+KscenMBpAVrIEXZjn5wstQ/YHkqYAB8LIHh11m8jBgp+5sm9U1yUsbO
BLf3EBsCA3H7O290lhi60W3xTmzMChBDGl4mU5dE8rs6JvDcFhofWdfqDXjZWque
MGFFmCS/vf7xOE8WFDdcidb9OjZWmCf8E277UaAi46wwIwJUVncHez4cNKDul29R
y5/wW2PGKwQpNJrH4cMsaoWuvE72VYq1qYfRbdZk4AaqHiLLxBgOzESqZ47OB/ye
6uDPAJpjkgduNKEmYtd3neR2jfz99ly7QOm7P3COacesugiDDVO50p8rRPHuXC1j
VDm09tplnlzRLAyDh+PDJTAQ2ibTcDjj8iH/JG/b8yVJxdOCGl+W3/ZQmMEyBqL+
7XhKFsCE6nt+3EvWN+t3n2Flx3qTX7QN3382ncZZTvQ996d9I/R2Hqt2U9k1Ybas
LyAe+dTxrvdoJWRRDUNXCCiR/XgeLshW3Gr8dG3xhhQREz38MMca2BKZw8Djia3C
ChTCVTxCDZQrkcRtBy0yfSRMsoto4fcOeSkAx58L9R3sGmQMN4S+ZkapM4CWnonh
L5G4tPhVWd9f6FF6btAdGvsRezJcy9yr6hoWBNg8C/69n9G98p1gzlRLaa6cNqQX
T4dTOH3l0p640ndhpeI5HYClb3kL0NCsKgBV3yu7TLgSKy8l7zZuXg8kpGPRAdWI
BJi2oRuMt6PhNbXd22bzl/0An/hN3ToHRRaNSYx86VwkHtII9vBSMpiPMZ0p2YJD
wEPHh9xEjBI6A7KPL8nqDS4Hf1lnNwP6G9VARM72Rk4qZ4Nmqi/+UPEHepP93GuM
OnYcSHKoK0QruVtBkXPJmsIqjacxEsOcgkq6L8hEqiZLGvFF/Qqe6AG7PMuU1qNb
HDPsya4cz/SLVBkHEkjvYdUu41drA3W2j29+YeaeKG14uNFDGKx3PL5maxOeUpA1
MMMTk+01BvUva/y4gwEgn16AylEzkVAaPxzOyG8i9vvWglySG0yAqdds7bclYgfw
CBSY3fiWeuYMAUDKk3n2V/cFBjUZof03V4lkwqIBr0o1IU68bKlOHgYdjKFVM8yb
IfPHYsuE+QwtyEDdXzLBgYI2czDIkmg2IEmAjTWbbXs7ek4E0zlBd3oc9AoHTdeF
2aqZwqyav5cJM3Eo/O5Suq7m+PVvL83KuvfzeLGHvOZGKkg7l/8Y3mySAwBaYPHo
zSU3HpP2uID08gqtqhy42o6Sgerezw4942WJI72qkE5vHEIM36AZTBPFaPxS83bh
uV2MiTChB2d+mcOQjwA9w3krLS6ZInPQzCkUXkrUKwFr0yuJoWX5c3us2YyoSDYh
iEaqdhBESj+op7a7D2qTFiH/076oMOhCM7WwS6wLXJmEX8LexJbGZoilX+BGqGXh
nwbaiQ4s2uaiL7s/G4C0RXBWxafiZPEF+hSwRbD0zpHT1OlNwJul6tsS5wjK/vMo
5ZldJu+mXC34DYItHF8W+xOwmeRgT7gqsn94FCwjBTzjZ6X2K9W4uIIc60QOIahC
MYuxqUYdHmRhPPQy2MgPP1lJbPaEtenZq9o2HU27TEB8IB9k+mB6jPfD9S666y96
TYRU5ff8QIhBtT5XE3wvkt6V9SclXyHSPLzcKowUoRRBx3vA1e3egaJmObugVDKk
coKIvGgDI6O/DaGB4ZAsCqpLufYaWd6Gcy2UTXykicZE+D8n0BFCPua+W/22GUgA
5zNqWDBWpvmb2JDIYWy3HjzzVvR8Oc/P2qqpyRt0WnzGDdDPH7XkhYFYSok7CSJ1
YalsVJ2jnTyXpS0r03ym9fo670C7IP6KCUsTtKtPEsx5SbIlxKG7fZP9Hu37jnVF
jJp0JUC3P7Xx3a4ZvqnN0BmZCL+FpgP0xEYwL3ukASGzaBPI28eQdpIDTnTJJGet
PUgHzTxfP1kvTxM6F+W5JUP9/5PYpd7Nn95VPdB0B/hg5dmwTBOhwcjoH1XtpzYQ
LTDQ+ktQM01A9SoxRujDTTEDanrKD94uOgW6PwnUjI1nhgNwG45fjfQGLnscLEPx
aOLA1yR63N7wO2Yu2HJnSCINbrYX0QEbPL4LUSCKFKeSbvTvGvZbRQfGaASeFVOk
4yylOUGeBhGyBEILP49qiz3zEQhzwRQgHHTC+67OdwgHiLnTs6LsoB3TtKul0qKw
FpoCwtVo7RjopOA+M5Gd8bXUmk0xV/JuIJ2kKmIpJ4gDGTuUmVXB1MNXfueX15bG
zkYI1tx/vfTDzZqg69uicRAeFij+2V/qXHbe0RVIkO4MAWyfyODvhONqXrm11hhy
WrTtsqI8y3Dk2tbQ9Mi5Vxrm49WS0p/y0GzfHw+Onm3GZSpcNs6MXIH6VXOlPleq
VSavZS/PxYyuIM3iyHNTz+oVHq/N4y9JcFrXHA3APwGfoYV1xJDo7QqvDte3oYVc
Dz1THzoQq0v2qBNXwJ+/XYF/RVAADV3ghhzZ/cZ4qG/717gfa7xb4L2hAVpPpCcG
rWR9L8Nsn9JXbPFiTnbGGu+YZLprPA6dc640GgSq0BAvj8KEduvEUCPPexIdNzvW
PPub96Kc2oJ+5XWoai2S84ocKeSs2lFafALAzkm1jyekfXMFdDuQ2vpqEwHnfJj/
xCVHDk/hWX8zE5T4SLhtY2hq50nCFi96NTbxCMLhdnrRhy5Mbo9NcJz0u1LpPSzF
rn4qqrI6c9ir/tnDqwtlzvZmZIRBniua9Y0DfOsfxvE8nzVfmtyVL65LCdJGdyI0
bv2pRPM9X3RdOZsV/9iQM3c3KkbsaBNafGgl/shU7nmlD6LMjnaqp7Z63s+hm243
ToIzf8n9ciGdjLLCxLRJNSbcPZkHr1LEePEXNzRu5fzlAkfS7M92aYwnQCQDuyrX
VA5VpgfMb2wcfaaPztH7LwJiXvBueG9tJs9zuX7ekUqNZfFrNTZio8bqsF67+kdN
UuBcGFfNysNpFioHtlguRC1U5o+vVse4sm0wbubDi/1OzeA4rZ2lUQSh1EAO8s11
aMp3dYGzgAKuNCT0MmI9JXLwhCxdCU4iiSGKfc70+hNL1PwpBhMUObxOCuRWy2KD
PysHdLDfsYAXETcfrKzr1FrjYd6djZoKIA7xZL4/I9KYvnd5dR8ncsHAXuUSftPh
7rxuhvJ5BXwz/4Wp6fY47aL3B7PGkd5LBu1PFeDm4imJXoaNBg2J7Y5osteyOSc5
xYMPd4inrTBwTG5hTcsrMGOhoYwhE6lY3Oxsm6Rs7SZK7yAKnpqR/BkGw1eAuIks
LVDmzjeo6jVQZhJw6zcEMfetdsiFpo9DlqMjt24WY4kIEG9gAirSpHhzt2V4hXde
F13MVVLSiYrVyaAsfZzA+yJ1iP21dQb7o7eg4a6dWz6jjMRFRF6W2UvA2pbfbExm
xXGxXWTIqJ/aTJ7/8hBVO9XEFTsOpLWVv6zLbXm9eKzgyZiTDLMdfVM3HcteKgGW
h78W+49uIKDW3X4MkS/GGOGkhdmjemgPoLKUL4e44hWlhE42cQZ7rnkr7dHX7LHz
HuA55puuvGc8oQgAS1sNss86xjE+OIoA0hbMNy4Lk9JxZkvP9dhD8dFw1VivwEWE
jlMOCgINH02zvdTCFI4N4SNdi/xQPlbBSwtQ4c3K/Czx31h88f0pCU07h2zs7nfC
/wnPGYaYi05/XdbuVCh6PtvnWg8bA7QXBrcwU0X5BdH5EUyc7t0VwPXDctLFq2qf
9bVpgaFBlCopcFuNaIbnB9UHbflI33QFayfBUpnCpOE2/s5Suk2bAcgqgMlQP9J4
3kfMDgvIQ5woN4SebnVkkV15Wqy3oRA+2jtzhQBplrcDCGd3PiHm47MMuO1071Un
+EoFPkR0najzUdTCro3xLWm+dgYVIlO5DGPbx+zfbqcnVRjQc+MsFQ0GlvM54YFu
gkgWDYLwMsaapfjtyr5C/JU2SJiE20o+XSAc9G7U05ucwwxxXMpaOBcs7es9OrOo
KhgRIcRE1vLQa7UkwHSvJUw0JUleGejuSpU/sgN+TNr/gc1sKdH/3zpUcpGPOc1e
HT1BduNY+p2Ew/9PDfUcU2MySb5b/r96Mv8NmWHjXUyjTmNORD0BkywYXCtFZCP2
QUE9OZYhv6wQg3D67azAqtEO+xtqcxXGT/ig6hgSGJJvPSxm2rqoU5jXMHz3659s
jAsLwJwMT69Om8LsiN8YKI8SsgDbBWpeP9pZE659cCbgJm/Kuuhgt7rZFZgrvDmM
0lsJ14nya/Hn0Y88gIolI0Y0BkBa/m3bbtMLbTQEHX17ru9nlqiE1XWMA2rgAnrN
mibqxUgDDRnBmSTVr03GSsUck0QpmuqrsfFtpQUpo6ZU7qNI1VtkpmDTMuljlKOC
rf6waSsqIem2jQ92MA8zVLwnd4wvwJ1TRJtFfBD2cqpqpTLr2AUeU6SEUnU22wOJ
7OjQKorxukAlMGGqQpKHEI0XBA+amx0v6EtqSJb7FizBDYr9Q5xsM0n69XNgrwXZ
TvXMTh3pyJBVLteDuWJCqRVcVsKwIzkL46oSXhy562TIxXMvd0q9nxDNZk8yDGZD
4FaI2I3AdtjccdFyZPB/ccYr2IEsnVOpeEKIyYe3PJyELqSvT1sMlBRDNEQAgZu5
e1ladvADu/sQNZrKF5eMX47HBGkQ0+6PoT9hDAhUqunmXI53X9TcNTNDcR8Z2UP9
Zfc8cfsNs0bjuvEBC/sd/AcDEeGxHwxUD/WaH76S+Iy2CGacePurOegC0VYupp9q
6S16mIdOtq57IIbcNHhVWgQZx8dgmTqXSCYYhq/bjdD4FiRym6qDhsAumVms9aVh
lleKnwc+NMrMcTHNaLh5b4RBQztiSqAOLYOtILgpfsvF4j6+HKV5GtWlBjdHYAYk
OBTKIqU2H20py8kBgiF9WGhoGzWYXka65SXCnRZbmUKVe62G86uA0ebzHdwU2mVL
Ub6qfDis2GjozlbV8X9VbAjEzbj8l3u279t+moCA9bkuuLjND3z42my9Qd7UgWfF
jsjpXxQbHHNDKGql7zB6lKjrjs5tIAbDMFFdGpcCq12y+y0nbUVEmhtrJeBwUNXh
bQByY016CntW08MC48XQrMixSGbJtsW06Q/04A3S9q0Lp18hA1FlF1FX4/Cuhz/l
dHzbBzSVI6la3HTtrpoeD+1CWU+IBmMuz9hV9xhHu+v18o19fac5GrnGmBztUOuk
aO+DzSGKdzy/nbOK+7KG/cxGUy9ZQ+RXC4jHNo9Yq6z3rBLwGfy5od4g/gJ6Jn4V
t+UEO/2KMriGpiPKUPw6SfG5fwrLfRqDWi1CL0K7WpzGXo7feCcHRu0MSmjN1sPr
sr1jFV12H+BudEuxR7pDGL7KwS/zCeNwFakPS0Qh4JK3jDuyoJowA9IcIPfjnuJw
ULQH1SpxQN2N6YOrjQayXrqWSFSbfz3L5FG5zrs9U2Yv52+8Tb03pGLumQGB01Fn
jYxx6CUy5Ldctt12gmx+3NTXUqXEMaMKBSE0MpefhdGr1Gl3mgZ9RBlDH6sUVIkk
pn49/jhHxo1YRFRP/hCg2eP3B9vW2pJpKjwOWLzKkO63PD5XtB7PboItJ2cPnl7w
DIc1NfxwW8oyMbvsTiEKNTNnn2oGe5bYPHgF79Lzd8yf3APrVXBsKMwmsYVXo4a2
Tfk7ECh5Qu0Dj2bVLEchRwdfxW3XBlJGq0MMGafT7W6TsQuPEb/X643QYpGvCdHx
TZ4BhpecYMNyEzzlYGsMdpwWYlvUEEcfFNdBjoPz1d9NedbfD/Iakaz124CEJv5p
wnMoe3kz9O6DgdBBZ8BYLOU9Narum9+vVBOfvxSV9G5Lqq/cy1wv3JrfwcD6AC4K
qyQ8rCWgSUXBWOwEKeCrkcV+qTHnBcNwPqVGMQ2HcA7LspGeQRScTRdKPibm9Pbw
Wdju0yRfKwLYACooY9/oYjOdGkk7ef2VB8AtvPt2SJKQp0oSwztciT2Ob39Gm6nf
A88xvndYb4KOT3q1WrmfEarBqRbyodeoCYRgVPRjLwWw8PpgKUBWLDjkgpximWXf
732ZVW7sSLsdrPcY7ViUv/KoG7XkI6JqcPfu3L+vqM7QwrfKzQx9QKadReoyudXx
ub1BnW2qO6G7RYN3z27bAOrf+S+6ICTiwf762Hi8Y9+OcIiESXHx8WQijMrc9+Df
MINjjsn6aFHAqLtK4mKyLe6BBXFmM6Zzm2nK3iZSgfA/1aDwaMgo4RgJjfblfAAh
tuRAxCnI8d4CM5/QRv605p87WonXJYiG0CKyDUMM6AkMXSg1b/iKpR3Sx+BX4g7P
Gt3GobVYrWSuerH8JCJ9kZ0l6doLopK1ibegpsHII5t68MZ2UyOMndHCW+m3aSBH
YQdOyzq5YyieUnX1jNdiACKlicRSXSFQo2bHjdEEh/HbQbz+7xpleJd1N2scSs7Q
zAr+Gzg2a3TjF3yL0JCLYXMyuflWdPbrUcFowX+lOYHifCuaJailohrv9/XDYs6u
/oqJubqMv3Ab6pTyhRVz29yOG1AgVKCDX5cRNa2cKs/K59b3rpwwnbSTiszUPWl7
Q9lLNBxjyviBaB6Q3mknW1SKVn/z+GlmpIDfFf3rCurZSMsQ0MhZfzN8+B2yb0ao
gZeqVvuWSeOOjrz5rcb+PzPP9ePamM9AkJ/6wudSJo5976ggJ43XI96bfxduRE4k
5/WgyK5RG0YWJ4QTaFZS8g5/ZnOTp9YEAWcdYwNlyJSlcRGhMK7ZV6ZrMtAjlc77
Q4SPIwDngJsCw90xeBsP9X34yc0Ixf6mzqFaQxC8HEkpsR4XUWx7GrdP+LZrcnvL
SgV+am87h9umZdMq9vgbEyopIgOTGFG6eDF7D7lakVOSct11f/D2TioIPI/cXqx2
158e+JZmLqL/xIkvlCdEyYnGHxIKtLGaqzaSXIFeUCRqMVNbqtRL4oi2KgdZbTfw
T/r7K8zSbNruOcEkXnJkJjhlqINoUHDRztNh+AWOQqdsifTmogGkFBq2Ax78jb/v
rffmuR8nEgcF0m9DsmwDrxOiHpxtoR7gH/nnInDUe99H4yYx9+kcNUGno4HR7jO5
Vv/r9Y+OMEGMpj5skSjCyeh/dZ2eGTELWYuEdp9HXPRasuqDb5NcgqwskGKz6PEf
PKQNC59V51sipH1hYuGQCy5XP8L8Ghcf6P3ypjzM8WL0BEZivSJQstJwFrTlZOTE
SM5nMDadgn+v1htO5pv4rPLd1T3V610FjlozQPD4zhDaVEtD12uooXSaUuwuPTfL
le56IwmDCtBo+3ApKKWohRndrF9Dox5X6iks/vhIp+YOpFX3Nn+8UTQIYR6vblKe
Q3l/NZ/2Nik1UJeAp0xzXI09dTtPoNn8IspjUI0Xk6wiuvAMB2INH1GAH94V9sCq
/FOEHZok6Lef/JJP5vW0qZGQXoZbWjqS4XLyHlQIaK2blAX69kZL5xZ3/agSKgN4
Jtjf79TigbLahYtmsf34Epw0kgW2Sz6mENXCsid+qhZsVGRcRPjQbhMQZYmzh+pM
LL4Ok1J6TqG5pzxhBUcYPYSoTtSyqj5nUzEyt7NjCJMlOZx9Zl7rCcCAsJblIYUL
aoD1ea+KU4fipt1PzH5uOCTtFzIojQNbi2KeJ7cGze+YnDzp5adI+kVsRoTDwlZK
nSrhI3fdoRMpM3TRYGK4UJhySwcnnEJ9OtSnliBOop2mYeUp21ECgSJge4OZPs3i
fRUdPY/96pkUmf1610ZrwloF1jdpRpWsGLKmo4bGcQDNNb7MxcmJdGxu8Nz+x8wu
XmE2mz2AG9zHoJP3Bv3swmeKas9/tGGZceGkUlmsUjjwbIVUlZqb6KB44bl/dkj+
uiYi43Somq4dCZaybkLg9xntLBilU6X2h2R5sfXM+ggwjwn6aRzXRUaf85cgzz/p
DEwE0yGK2b88AkNYjEUx+t+0ZMrFCrFlsXxUIS6k9z8K88rnQLNDVesWcNfQa0fR
FG78Aq2L9pZOBxE7g2F+i+pOIkwcW7V+KKTIZYmzHTN9BZzk5o9NuXCRGlm5jKc4
blyyyguWRzVrja9nGt4ocITeatiHJ5YrRBdRFL2pgY3n7zckebmllPmucmVT/3jK
0WNrCi4vNfLcWTC/Kcz2a/pyjqFIWV1I5nxOUUTJw93rO34kJUXKvPF51MGpxMdD
sb3Ia8t4aBjvAtcZZ/CSlNfsK7+lFnoBCeCGJQboc7Z/QVaTlHHXGTbu0K7tS0RD
vDZwZa2b8QJV8c0nGzPe3GUJqerzrG/sJyPvbXwTqJY/G8UpFBF/A1WsceYLik2b
HxMx4lYpVBj3YXN6N1MNydkk7hu/QiXUK7bPVkLauJxUvlRPzc8/akNm2X8pUek4
lpUCrB8qp9ull1jflLaaU8jEkfzZcJIT4OVnrw+bn/5Cvzo0SYqY/eJ81ELasfMq
Qt5URWdzNF74myq1M5JWedWDyUuJiHdUkMqe3a67vn5Dpu3AeHqByFkhj5QpQO6C
TRBGV+1IyohH0mjsAVvbseHTdCj7ED5cV2NcrVYnZCzLLsP5jipCyS8sxS7mJJOM
o3My4YB2yFpcnotLYPRTWY9RxSs7VilVFa2+V/Y9YEMj3XOsVF0sj7lHiQgFRCmk
ys+SXavGu2e2pxGCT/ecEgkJQfOCffS3RxC8veJOFYiDdLPRgON6yVzf8amGnBTk
s56lFqp2Uuu0lTncmYmTIRQeJt4BCeEInJdR+x2zm+Oa/qwET3IuG2uhRr1hX2lN
iIJf5hI7DIgINAe+108GuhpJi1fi7ZFAAMs+gw7psKrxVH21/6cYAXt428g+BtLR
SNy+DvtWnczkSWScE9Six3nKQJs10P+x2ia0NWw79SixDaG2LOQHU+VjVb4WEImG
RSIL7bE5Wta04NfUgKIC6hc0P8Vn0oxmyO5CZA2myo5RfPxh0JUpw/w90g4Bz1WL
dlAGKjF7/+SRFyBOjwcy/qGC6jdNmwwWYn15pAiVS8zu/VZSMEhDekNHcMNvn42+
XzHKFFNW6Pd8+IezJKlM48g+qIQCMkb15Ejqcp7QB6pXFMc09ojLpMEYN8p92YWq
jBv4XMt2HiUbl5YkCIqD5rd7jBILq6ZsiqmwOI5HgL4nH3shaIdpAUEhPRb5ritV
eOsyWsbmToXWwtxLMitLwmwngmLzVSmZXsJnEN7mAOUl12EI6kGRDZcND+t07QPU
3kZX6dUdYUAFv0PIObh7ZtezvIQ09omzwWIcpkLXce1GlbRNyTMcWUk/xttzaOv1
nIMw39ejDbVqv1nDjqJJLvRDpTKrQTtD6iqvXu2q7vSYlxynL0PrrxwE2xxlKElr
9GxikfZsAmhqUf/WDo6xxD6v2cPobOW5l7cmFSJeb/d677t1VkOeABv1xRyRBkSg
0ozXPtHeq2Jk6YLiZguv6uAOl4c1PoMnsSdl3lC2KbIUsuAm0Z6mp9Q3AvySRca4
xDho7wmgRfwoQhMr9C9REU6n0YV4+0wGUz3pz7MaqLSseEY/ifdqSMZ/YgziDV+K
ks7J+nl2fLAo2i+GC3Nr9mr6ze27jqZEbrEKeT+dbFZ4LCt6FjnMSEnXlp0pckF6
ZJjBIKO/vSSxDdRXSmakuecyd8IcuXKISPxAwwkusst2rZWbrIS4SEhEH0LE1nI+
vTxg7nFeJn0PH+irwZxGte9gNZ9a03u03Ux44TivtXzQ8SHk402VdgufMMJ4khiO
rj1j/AL4NwQZZPR+Xgqsp5x8Akt+a458mYarzkm7k+rykfnXoT1mNZbGsUTVS8Cc
znkV9UZsv76X4fItf+1bs2c3HrGSLau8m4h5od9o5d1uebvUkBnEDKiE7dzLlGMk
1SAASiNxpfm1rTexACUjgd34Fr94oOSlJZAilRE7weTYQkAHznEMyF2L31aw8/qD
ItXmno+Cg2gJ3vYazp81cNhek1ZdWtw2AsvnE53i5mghrcgPkcPcpTm9W4hsS3JY
+HAdmr65LVFDkeZhp81r0+YCrvoyIf393AWFuDngG4Ogv/mCV4iTFaKJVjNjzBkh
d7Bto3vst8m9imvL2HasjjVNWIbMZIvrhj44o9HHwHOFaihdWPBd4mwjrmj7PgPP
Clt47FdzEq52xpT3jWShrljKlNHaw/xjM7BuaehCEq3zXq8mvbmEiXk2oH2eCIf6
dmQHa49pHVUD7GYTv8Lo+O3E+C5wG9RD3WUzSLnnx4HZ7N9KBeEDDrbuk+w5O8Bn
JNXLbBF0Wy2MmapTEYj52zX0xFy4giOzbt+1L9WZ7rwVSvgKvJXCNqgGM4PN6D6x
KZAzp/qGdeCPHVNuKu5dXCwKQ0WT7cXs3pN7a+ow4gfu3vAiLoFPIUSR/ZRHVoaa
dmNvujXS9GnNgpzFys1ZzxydOsATv1YPhQPCC1vADId/sWRlTE53ToUySknDg1De
t7IO2kRFXN7sLtARhXAf7XQF5lqxS4QkSfiSp5BNkg+QIEaBE2rG0FOS2Tq6/7tv
GfxcSm/uG1nHN/LanRPyOx1HQgw2Lm0mMA6AOmvdSYaD2kvSJjDBVOrDJZ0WWmxT
M6qWDQ2BqjfWi79sa/bzp1lUvKYizLfgOyVNuZnBENiGsSoBbD6h8wlCrWJHZSLa
6Ce5nwEeekPcCNGdx9f5gsOqXnS0fNpmg+0O0+lLvOkgYxx924SCUXSgvtoJR5Pf
ENe4tNYJx1PIIVtaCLdRBcr34MFPlZXOFzJiKR2Jkmjj3jVTbhIodoOfw7q7S1Jw
GCBJ5eucavHJCRLkt84Bkbt17Jzuq7vIQKAFCOmp+2EDIQIUdD18Cw/CfDeUixJw
n+I3Kcr35p/X0+f4zn/I9sCSoG66PYE22AnZnL9siebIzlE6McD9Q3+EWm5qL2/G
ar4gfgh05iUCa87L5UJic89ABvngk+JBmizGkBPTFzt/sCrIWdcBHt9H1kQaorEm
z/xAML+qX2bl3R39pJi/w7y3lbDASB+MuKxF1ODBnc2PUWZrAE9J9FYgOX4Dih5g
gJ48DO2b+zSzHDg4rvkLPA4Eq2skq7V1Qengnyeq75cYHc1BHGw1sZVCMBliYnl3
I4F+Klv1sHsXPRPnELArME7u/+VBKHDLUkV4EqB1xPIzkrBkYlOks8cd/ul2b/Ds
BW6nHflMZJxu6F45EjTs8wcwXZtKsiuPi7Ux6sdew+eEsBOQH3bWOundHlmql1Fw
aev7ku6TTnQMS/nDSOhoMZi+v3hhy/4bowR+CKg6SJZe5xl4TS+sdc/2A5VT6Qyi
mWcoxewHu9PHeuu9FBIXmtSeq1ay3qF3qd1OrG4NPlrTTivm+aXPtaE0iT40eKaA
F/Jvb0AyNP2u74BVPluFk9Y2uJMexl9lu8VDrh5Bes76e8DOUzZQDo8TSXFrDv3d
UV7wiSF1WtEIkS54gFacLz76NRC7Waj0ow2RVjJYIFEzPZgIDFfBpBKbOlgj+hdJ
kI+uaBB1EUVioKDcxB7GjO7yW+MPLGUO9X3bBmsqpc39RngP+RZ/Gh6Z1HlGgO9D
aC0wRlxrCk9py9E/n+dgIA0EPdKhb1/arH1i+CZH+VLrsYo5v5lleSfdVPJ4opXD
PyoiLKkZKRgl56PC9zjrmBtLe4i1a48unHPEF8VjVEduGMR6HHynZHCs+xZ8gV2x
FNFAz7DmN9g/ujFCiGb8gyjotmbXm68sFoxuP3bECd7maQSjq5itaYxk9PPufvFo
x44ZXE6X5w243bHSQAVyzVEj3rqVjvvF6bieM7I2hVyT+GsOXIL7N5/XccE4LyE7
8oylJjjoLMq1kJdSQPmxDqiiTnP0n2ToBlMzwvwvXfpmM61lU5DLMVEKZHOG+fSQ
s/Byuf2ypAvi/w6QBMdj9mrYBcakZRu6JfLUD3avwyEAii3WsZZzhkNREPu9wdK9
zZ/une5288QxjUs6UHlxiDimQmy5QZwIqAqLHCJtTq0SLW/5X6kDmDaarA6oBW0O
aSBMSnPQIZ04OF7y23C5Ce/ml87gIsh0RnUomapA3dpPAL3cLnpqaP+Nn24UxNSD
3DPALU9OuyYqSkfQwpNzHbAC1nggNKy3VFwd08FHQ3YYwbwCmmovnYNTrR/IOKx7
0Ihn8O39WYi518NggmY2UyMBbFvAylgP3yUPtdNDwwVnlzgm9IJ9FK0QstWeYDzT
QiKldwZfXI9gw1nTtB9Xaq1254qzOkQQ3MCa3XUSJP8EqYiKoPK9xUxqGD17z3VD
QqQS+t2z4OiasGqcArwBHEc4hPgZPbOdhlIlXPBQr9LEOWn8zEiA3bzX9xsQ0L96
+/VDAf1pLgfZYms7TTjNwbZnBMsDHOlhNV9AiweBttrXT0LzbkLVlbt3UCiboZri
gRqGRo+FCtyaIX6EEdMBIJZdaZpBsjFVJLgjjdJYRaxuvNlc5IpMt1Kfbp/JnQrL
g6RRWaZex11fGcHOLv89mCGn6MICjMdaMKxkZ/0qc2G8X9K3WdjJurQKgPjt9ePA
yKQBia63Eunv9q7/z6JsDYpm5dLPa/4qZs+v28SFpuooBuFsqoit78GpT5VXzqCn
EBqb44DMWq8U/mIcTQSVNuNC2Qn6NiKRwUCKxYvlRwrW2qM87UEaiJuVXqoFMlSf
hWJOGDCBHkko6KOVasAPtJ08S2XCg4XyOY+wCFV1AAYfZm6mIiJrbWrC00MsLBCb
DGqZCZD15QnS7Tnsha2Hgj4KfFqBESF2WvS0hlhkxbvcQBpPuUDk5lhC66BcX4x7
D8kY3Ovm3KqwEXftOt+Co6nOWvZxipTAT104RpV0IP3UC2bKxTQoGeYZoht3fJ9u
y7FOwXIj6WKfB23Q1NMvY2rwkU5WNSdL/DxAajkjiZT30Mdg/hDP3Oh6Tnd+8VLK
SGvmuKFWrM4pnn6uJQ/DpKT0HwsmWpQNzcJ8fHxlFLfQFNwYwte0Y9opGtxgYiBe
i/nv8n4/WnhnLpakxKEIt6OZjYsd1wvKhDr/EnDgR4bVvkvG+BTdVRbSE+ke4KrW
XUvB5xRP2bnqHMrk55s7mOBvwCnxFj7UxIB2JRK7O3VN9xuIq2vn56cEAJiCe+fP
3zWsicY+d3e2cFvKqpZodn4+4KNB6CS/zxH1C7ADq68JoQ0f7rgh5Tmb45V3H/lH
EcoeLrQTJnW1JwpikAgbrYuoIk/vvqH4VGRI+GPug1xJMUDDoZq/wJSEpU+GGjgA
/3LvEqVvdrP8ndC173XsfIaxhgO8ErgPirjK4zLhZniW5QrKk+ZRqgWddtuD+/mh
yT5ZROp74APNAvSYlbHVIyY5soCxHXooe9qVyo4txN80RQ+lZnn1jnPOchwtPzIG
PY8hkMJIvf8Zj8D4kCwI/1N3C7KxIOGjdAsLW/JXuSMHLNGYmHFX+c9THpliWQvG
Z6Zgtj7QHWdiU2IeRwBkBPIp0c5a1L+/4LDKAgjHX6zihIJkR5dFTLaFf3lzyVos
Dv++z+Ezbl1/noODtfdfIIsCnQOOCFUHyfx8OeuoPmh+YsapSjXKbj4Lz+7VK/3B
uBMLkPKNlvQHTifQzQU2XpAJgpBcP96zZKU8p8Auxgz0H4hZEjeT7oudQVBDgqpO
QIw7hEEITULe3LoAVwXnpTMZjXNkzwQDrCc17yrpt1aHdtdJT+YAxdYOZqAKeFy+
5hB27mWnkTfENHIU2MfyCGHHbcbH8ZLPsXnW3FevYunO6zx4Ic6Q8RcHTeWTV1CV
04ysz2+BAMSsXAG9urkNAlkh+j03B3Y0EYKtlly2uCI2D/12NcgdP0tp0wJMNv13
dKzcMBy8QcE5Zaxm5DetrcGjHatFiTB7sRKhZcCa0BSV1ZqipfSDJqrXfWBK2vBo
I17M61nrWgFdSoWre1S0GtWrgbRoPplWHmh8+a0MZVjXhorCW0rNWMVJw9c1iIeg
9lTp2SP+opMElGeEVPUYvur8NNNbyX8l1VxinM9rK8GrHPALXBlJ0u9tGfrLsP26
ee5dXM+NtmJRacVDiAzQmkXFdVAjN4HqE3Tv3ffteOsTL10YOGvO6Lb8WYHqgdTD
4FZKCdF68MpHk7vPd0oeglhCPQ0wvhsTs/DZvaUO+lgng/fob1LiBSS/L3OshmHP
XMjaULuPlb6GN022z5pNffx4BsQrdfGPlQobxzs0+mOsWf3WagDolhudwEpDuXnx
c9czUgVowWI7I/LYyYH0nszeumDn5ttHMagER5Bb4OEpp+s/FzTNXrNTJFs4DIrg
vcp2wgNVfeRwIlFV9gnPwK+ORK6jijV5ZXMtsnoZRGHtWmatcmsfluz+1DjzxTZI
kX5yGqcXxPJCvJP1Sn9uYeXZ8ofsA4eYUEZ2/jyvopaegBO0NITb9O9WoA4R1nUJ
e6a4cuU0kziCi0lYf+Hkkn+9NdOz5Kh1gC1ub14yQy+DaPm+aVv0sfoNLaZcnVog
2Sje5wI61EW2xgEKeV0KSrV7nPgtMAkJYNgoyvbBDQwXR242aLC6f3QZ11qCUtRy
Mkf8HQEMDuSBvB235wWhXLTwC9cjhAj0UJehxhYStCzx7mSFMB2iknxGUXddrq4R
7a6jGYNfESGQEHyQQx95ce3O2tOtYtbf5DqBBRBt/cfHZqL9CZaAf4bE4HKGXu99
UaYQhYZP4DoWUsy/ol7KmBvQnv/MzlDPLJNvsBPX4bkgDbE6O9TpgY7SVIsWDeY8
JXbZNglkJxWlQC2khXj1PLS59YnqCVG7lIIGyKam90Ck3JP+f0KoE6Nn+Bs/RlJ3
HuQT5bIj9NwDzVQDK5nk++9EJ7CGwC36iXjiQViw51kgeE1WHhq2I8fXrEH42MgB
jLfyqSaEE0Hk4YtpZ1hkZaeEvZGvknfWmrmZ7EHK0u8y12avvIK8kE6Z7+nfvNV/
A53dhwyHPof/Nik+ERJTZcGW7FuLVaDTPd6rb5xBeQZgpqND7J0yz1AkiI0Azgf7
cQuRdCE11wcPSdkbUWnJrj2+RbXxFBcg14ACUP008l+HObv7nPpWggxCEkfc3IJC
Df73MShqPwYxwIFFPI53NdJa6uOhuwPbKO0crqjj6iNGhFI3ZW5gT5NTAJ2mo2eA
TucVeKHz8k/ZUtPmAWnIeUlhqMXTkkDYqtsKM8bn9+SUsd41sa3Pj6iZCXNoc3UI
RZYA416Q3Tgs+F+Vnkj0yuhb5rFQ9QaB+bzDx7GFhgO+GXfnTvLWiZ9bx2JhTORu
Oe+L+Dqs5jLBTmrN+Nsc/142vuqEI6bR80Egi6XU91vHZ39u0BQXne4NM6IAdhtl
2t8nCtCylchkDde5swFyDVdCCwXhG+LErlPFc8hfVLfgviBm4vY1hyQMEyjt+2T6
B1Vl7cGAFD4CzmwlO9vy6H+7ZHIujRN2+4aZlJ+TzTvOcxDHLkkr4n8IAEyucNCV
yTptaqcQfUc5IPvM8jwMWbQOUccG4hsrn9dli0H+9GPHrDle9QsjxLkcLAGaJ1TY
wCUxsfnULbZL8oJE9rXJr6ZyG/ydT4xO562bcwH15eu99MckO60UQdPs9XYGz7lb
io7kSBzWJuPIzxcaaeapg43h//7EGf2WFt9MY6fcugjU+5qevGRPIAs/7mCMfPit
q0U3NXEfUs0PPoyUJHOaGmfIkq3J5MQNNYQRWBYMX1CwslcP127UWuUNp/GJctI6
OpK7gvpY3d4Arox5c7WDGF9F9Grk8WgHQBxH55OKKKqL9fAZJZvfPFGtl1DeZRPy
W4Jb0mSt9mvOJJrJzSDhFU3pPz5aqspZMh3/FwlIQ0Ry0LuVFAooZK5P1Z4SLBHG
AMouiOVp37G9hct8QPvRiq+BGlaBa9sT0jOidhSlXxwZ8XNthuyZqD5rf2m9wBcc
+2cT7v0vXIvMX4e33rTU6xdClDstbdYW5K6EmBpHo48wrZ3+qzC+Qv/8T9l4BG/j
MCV27Xo+Xjhvyd1qso2FfnfUAdyfJ1esjUPRNBgAj7UDx1dhHYYenJbK7LKoT0g7
Hd5wA4aLg02hv5zoYwweoGzF+KUnCKOsm+2ayycm2JWSmrxTu/15MLBxfim7pXoO
8kYuqX/EKCs45S2XB79w3SOK+MIERrOrae90GkMBbm+gix2BqQWrl/BLxoLNI3Cd
mnkpvgENiTiK9Kzax67sPcY7F8MkQCB3ZE1bwDwusIlrqUbi3cNmKxKFBAwfiyS2
LoD5TbgMPbNWCFyE5GoqDPupgGrJbecVjm/lS0324GcmpvmKTSKACxz43mJVzvkR
PJMp7yqHcAEnA/V+sHMVlQuSvvZHOk0mp1CLFwbTF4VC3Akhyix3HEUspS4USH+D
kpLsEuETTpNLluBzppbyINXgIVVryqZIE5YmVFiF1co91oGCsYwZ4uovLcf+HuR3
P72zVChsEpdhzFYT5xoYS/5ErPlqCpCDDVs3abPNlSALgDIjMOpw3ihDqdlJSbYJ
geYAvE78t1P/6eAY8uh963Y4SvDmQPElnFWPpi7jRdFUNt6NM3SUOzDhb2a1n0If
9NnYHHwd0UkSDTNvWchHsex9Vx2T3Wsspl3nr8hb6oB1aRftQeMATQv8e5ME7lKp
uDOGqeRIsH7MZR0B4IoMkt3gFxoKvSihLJnVza9moHFmm/aFqKR84Z8aMvfHe3oZ
yXcZMDoz3OfH4UPhFcz4vcss6p50XQealTg9A9CerJ+j4YB27zvB2846sK9h0V5a
msCbEydZp0Nmv2myldtB4pm9q2e7sj1sBFyrt/dcR0GO+rSDpf9AHkoLGm/eNYav
/eTxJ1LRi2/4FBxs3ldcbA2R8xbv2DOfQt2HEyzU1JFiDi3054KeRBZtZ0ObRY/j
24N87amRjuuOnEWxK6wMUTwwQQLeF46c15JqwprflCu4DwqTmfMU275i6gkqox/e
fp+3KA5uy7azb436nntFTQj6wJCDBzqXLiWwaeosVu9z4es1+ccBzODYBXXC9auE
JBBwZPP3j+XPlp9toiLWcpkUQtd5ka5ubg88CQu8sI9TwEFwDFc25MYXWXnQ5xN/
l2ksgDsT24Q1SAlEptmwTnWs5Q3KFVHmefcgK2r9910rEvKczJoIK19/Eu1Gvs6/
pPB/3f/UvRSRjXxn7gd+EBIoDLC0Nvql6RhCzZJn/54rTM7kxk5WUN8wHry8csWN
Hl9m5PEgUHemPOaK8XEJ800qscpOKJBFxE0YxeUQD8cflkDnMb/RFg++1GTVGs52
/h1OrNlJl9xxBCbz8FgwuJlRhPVmFVNiw6kF0WelYKlayecpCktfkr2s5GX+2mRb
oprGan+h7pAsu1b9XrqUGTdEhVKzPff/szpufcJOJA323LxU6wyOdn+RQ7fMdQsZ
kQbugbk8JZNH0FHv0epan7bqaaEv+0dIuYqnnI/8xDGSalzPLD1T5sOEShceYYSK
WCCTJqJ2I/9a0wFM3Zg5v9gDgYfSwg5SKGSFga/wggZpZpXoxXbz0Dww4yKkv+t/
oxFEnJi9BAG9bwxNMvZ/qryJwUSUVQYCfv2fgLH1R9340PcR89hfwQl8M3i5lwCk
YQjHwuzbGWXaVoVXPD2q4mptSPdgZQsV+zI6i15rYXPSuheJBTb202Q7TFMbntYz
RYcIpPiS5csfZmjTld3ead7fq/cnLGEfI5JMu2KhPe7NK616ruB+0KDLqA4zTm/P
VyeJsIB4PIdcZ3YszK66/DAxi3LIjEe5p01KloDBqQZ4jTwZcnVHYhTBXG7uSHFv
ZgljEGh/CCGY3gN0PvE3sI+tLHX3P9hRmMw8CCGZU0JWah/r6SiTF8lXhfJY9Qui
VAMc6eJGiU4cKwSmd8BFl6BGKr/r0EraoKrA5UdMUbuxJmKgpDRcacdvwPhRa12j
K+w8YWaWfkfIa7n9hZIgzlp/7nyBuJbaDAjhKL2xJbRkIuohG8P50KSwe8qWG9TZ
WVQgUwo3RSAe172VWt4xN1eGhdy92d9lbwWHGskbOvui0RqAihJpoa3579fIUC4k
CbM8L8XiQtzOuxjpuEUbryv7OqCmRxZ8gbn9HZdeI6yfG0ypAwHeLSysYd6+CrZH
ySEGzaPpff42HMNVxs8NMwG/S5RWRkyi2nE8MPK9lRHj3R7pWvaRPPNaukfFqtZb
uZo47KJPIg6vHK94ShmFhZ0cp/gyg8ymu91uqsDPkHlOSd32KLg/CwSZiYTOAxs1
rLfjFRHKSe8Pf6PXUXCTBjHEgTHu5QVpIEIwEB/Zf3/jEZXUwC52zQCsz2mY6prm
d6eoXTfaYRQsYzKsJstJrD/z+nTcw+3CkfGiPHyPW+M+IcAwjqg155QO/9vyWvii
VTgVRFZ9SzU+TpZq2xfxBC+PeIVF3T0fWpnso6QEBj0kln8MtrCJEnj7YF6ug8yE
BQDcXu7DfbUS/BlrBQVKy11QE5EF6yRuuo814yh3z0LJlJxK1E1rMY9Irplhnq+J
J4kMVF7klQ8RdjauyMKeCnNxjRGLnmNKrIEqA67LFyQvNlEWY+zH5gzKBAoJBNSx
2ZSuM1PZrAg5NIleN7Bb/By6Amj0VQA36LJMjGA//MCAadSbOGelkJVVCah3ltYX
ttx4sIF9G+dmQAL0dq1NwUHdVrK1NUACoszc9tHJNYr8d5k9Y5jxw7xF0ILmIuiV
FbaKZU+7QPIbZXnvZCWIBSRsoV7HGK8Fgws2tXGRScanq0AJf8yFIVmWRTzCiQJJ
V7+YqcVtwOO94M12dF406QvLCioWImyhghfTsIictZk9r1uFenQ8Xpz9vYFIEA06
Q6+DX+fRfVg9iQd7d8WXSN5Hx3XsoaNkEuGozRtPHcp5Fwd618eumlv89XhwCoEt
FV5kLpt2wMQ0gof+H9X/9T2jDzIT19u0km6PBS2p2n8zuxUrcMCTpcb580FnbvRH
nGTsUiCYnMe9zG/zAunR5fucspYYqmUehA+SIX9NE9IH1bxp6K8RM/getpndA1hf
1uEVBV+8CSJPV8yYhLhCp8u/Cdk6YpN215GE8G0lzfy3YG7HBV8NoEEp5AMJJ2BD
UTy+KftIzOvKmOaapTsalphENpATWIty/ytZSQzoLRtAaLmebXlylyGqr1fnwA/K
DmhU1XrIqyXYFbyNN7Uj51ldWCdiG7cyO/0CG1xyalKT1p12FIwCnAOXVRUgJUQk
vO0bGPOI5TsrP+mHbrE6DLRciyG9tPZOHaoL4wqWZpVVr4htsMm7aJoqdMVzZhYN
L8qknNAq1p2VDvh223GjlvPmUoiSCFJ17HYX2t7A96gl+4hWjeT6wLHSubUwkTQ8
ex+E1FnSc5O46h843gDQ+8y7enyzcCsqFsA0Q6fE+cYRybqMDLrBVDMY09SEtsYo
IfDMKI2joUqULMaNJDfKqngI7xElOcL/4vMlgbF03NlVo0A4/iFiCCB4OC9TQrEo
Eeo9eGSnAdDcGRWlVpHY1X1CBl8AJv9Zd36QWx9LLnC+VvtM8bLNaVpI2BT3W5yR
El88blwfCpAWNyig5+oSa1trCDiGe3m7dFuIBWzO6oc7Wz3IjZ/si1k8yvxawyg9
1qXeVIP9EQxlYpbqfH2TlrokM+/0OQHGRgYjQ+n6fEZpTbgqs1Ye1B25I4yarnnq
BFbcoBI1GmwnymFNACYeoFN8QCq9d0uGqaxo7rkh604uB/YS1wOLFWIqMUa6k01z
iv0yRLlH5yKAynPYBz7D/dqgXIh3Akoxcwoe1/pN6k/Knz9tHTt+O2ay1l07GVvx
gIR1+foaf6udBDhhsVQBOyDevRyIOnsrx5ieZRC1Uru0fr6XkS+6AW7UC/xcqyzP
zMAxGyeCXzZCYnbXuGfHr6kwTjNyK4gYELDpBPLFUgGgxCx48aiKCN3G4+iXD6h1
+FPWHMTwVeejneqPQUnHvXoExEmftIjKnUqkb7tnSA/Xwas9FiaAfqtysSpyyvsI
9M0CQDiSSXKXA12WGkxU3CmsaxBvNhCuQbjUVpit2n9vKdIh9nycXc4eyj7xiXEA
fhe/iijzfhgXymOmasrgw+IW9yiKeyl/did+9QtHikJ8Y2nQ2cX873ChLKILBxvK
BenxHr15Q78u0iJGuGyEw/3T+uGFqoQbN+j8PeK8TeP/9TYXrlqUg7RdF6SDkLAj
S5k/rPQDuLORwmMPHmVfnG+03MNSvbovA1Dw/fzNBgmeGVGewIRn+LWcfJHIwUDR
kMOpRVQOlTPGSTiEonbwimFlhj7B1lfLMb/h2ajpCscNMK65L7EamfYROfEPFCnF
7ZSoumLJkNA3mVMGyYBphuQkm+t4ECqHEPAg+zYWpqcQkDVscWDgrwqchzNTA1v1
+9tp7iLmDFSkIdMSbc5m2br5aPSJKS3NG9Ss+cJpr9orYHYVTDkbpGZELGePKgak
l1YzZbARw3rcQD8NpFUz342VvpHWnoKpvidNkWooYdXB99LPnNBy/QfEBepRfBxN
nQ+aTF6YPpq4s5Gn4qQDR1WDkqBN5PkjxCNEsg8yMapAcgccPxM/pjinCT2kUzcg
Yy8RQH8CWwkfnAHwPxbkRhersHHyl2OIfwteQVC2oK5EvNTQckLl6PVYLdRwB1t0
0hCI8Q3bRaHBm62OY8ZwU1FVzrPGDZHhqXbJr9FILArjisERWLDhRq3rJH/fTNFD
hq7eGAiY6tFUXR0zurJCM/WOayYGQGwHLUnZHIzPdkWNoD9HNIOCBFmA23ZdBWVo
JGZTQUsirqyXc/Wk/ImDaZRp+byLrdfJRYqN/PfReEdHoT2JWFIN4OX68bZYa6Xf
jFEu3fSTqZSFoqDL2zNVTz02IKT7K3jlJ/Hm/aGYW/dflL4kvXMI93xjHiaML0W1
buWmzE99p8Csyn6AjSKY8CwJ4k1E9/70U8Kh7EV3KS83ZDeZj3Otp6SbRKpuhiCm
pSJrRaxwK+w3YT6F8YNjyz6+iZN6PFMkV0Wo/jtdzDDYmnGovRn90ryd6oJW+al5
k10u7bSaBka5HrTcxqIR5MuwEIjtRC5hscAObg+hrz2HZvw20Fg90N6+78AYWNhE
ZmrNc8WxBvS1f9XgbjVscFROCf6Bvcj4lRX7pfHDdK9bEVrP9AmHi0eN0i/amMb/
lXvPZOYWJOKYIfmxPnKZjee/jFXwHOyqMKTNqiujxmw+jKQQkmTgta24yoiieOEX
d2LcHXMD5IlKjaS/795k4305mjILYiLa8G1dfyRYzeC9dJvaijYVau3XS6t6WHuw
F0/1PaBJOj0BWE/o7QwKWTp6b5iADdF4WdvrXpvDaTW/YIx/gHoqVEIVv1SkQUT1
15FJxHyQIVgsFM4P5BRgHHo2Stba6b/U//C7z1UyS6JZ8NyWluvSC/oAQpfk4oso
9WTGQDoT7whF8wYPt8DzifSryRtOOM63RBykKKKAGEkBpXOxwfKOcDpmLeA6Kd72
efG0AyQZPaY/hDEEp7asJ5xBNOURYec4I7n3Cb+7mnHaoACI2zBJ9qd2IBWvOpBF
rf+2P0RXc3e+TGnM3nu2X6eZDX9LSz8NS5H/VcoNKTXwp6aktskV9ZQDuE8M1RJw
juIFSv1nN9QM6e8N0e/EgV3PrPo8c9K3oWtZLhDHbhOLKvFzSvd3fti5zdntWf45
Moc0nYGdYizmYQlWo2tT6ZD7MWunLlhN/x7uVUd9ribROitDPvVFWAgg0R0OaNeM
Q5ewkKvMssG41ilvjXAINcWgdKJ+hensX+Y+W/Mra660m60V0FB74TtKSARVb/5C
KbVHcooUXfygM0B55C7O3V0ew/fNZyLE9z0PRGCX0ExzGBnmfcgjNu9YwWUZufr7
nEioIbpkOvhwKKCVegG9/ZLRcclMKbrIu1rbfIRP+x20Z0s9QywK9OwwANyxmZoH
j5sY2Ze+uwLwhysGgO9/PVKl4KFJ7PmcHaIgb8cznQO5s1QCQCb+nIMNM7gYzTBD
pYHrGD0U0uDWtanHhQChLbya4j4296Ti80Slb0Aximew+YQTEN6VKoY1kd48awZA
CX/TlcNUidszbdCaAK+wWoqoaManmhNuBeM+VuZdi2SZyEPzPfGEs+Z6rsmVRHja
G6ZApYsfXLlkkqrOysYDiNXqkPWTzyd8segjZz7F4m60j6V0xwlX7YlTMfFjJ8l9
LfYeu4f6svKPiUQ5WowNwfzxN1wLoJaen8CEcEwqXRj97FIj135ZU6INlkQypPlg
Rs2XKX5t8IbrATWEKR/+5oSymo2JTR3Ts8LlWuF2ACGTZ8PSRBhY7tFgCQP6LeKz
e2afhH96dAkw0HGfq9tSTfU6laDqftHDrVCMRZoo0i0YinFGrSeGzGIrlisMo9H+
E/1y34eDXM3zOpxDFogqm1K4JnW1uxN22gQLsjxcXs/D55Q7T8fJCaEKAc+qiwrM
1jyVO6rM4ebo+rNM2TBJnfT9EMFKvCKHaep7rK9MCBvzsmw86AoONtDPBx1MtPMG
u0/QwHy0ewi/MAe8CfHhW4auH9FO3dqfi+QPI00pDnC6hhOpoWXKGvax+N4PTDCY
K5O7A0uxXTzP4Ul9nNJYVLaTMhNu+JVTQkWkkWCaBApa/0W2arvp1sBdeHr9ZKcj
wNZL9ANlJWssPsb9yOzl2wifBTf8OjlnbynZpuQHG+VRk+0yBYrxFnUu6eiQjj2g
m1SNz4w7DH4FNqLXg0NHJgdnh/BzqDvmb2M7Xf191Ilhtx5xWRmE4y0AUJtkWn5w
IigVVHYRyV7NTiJ9M2QLLUT4PBcW/ndo7yxrM2yghwY24yJ8mre3IwRlCzUnk6DL
7/5mwLDMASP0XwM/RflHquKdI+VbxIq+07C336iqNhg8x8NaHRUahOkZqltGWLbl
PFVJl/AqflJhwc61PdYFSkIKgkxHad5lO3zWXSc6Xem0P7iHbNdILKfLWkB2Z8Wy
dvRG3iV5R5BDvOXGUgC5u+BjsxUA7C2Jw/GVppAPrkhrvOnqP6vp0I6AAlKBmGRl
UeV61Uo8oaOp0x3XCvfWD8FnPGbnAmQZI0PHdFvj5hcLYEQK0BvPjdBwL2wbKfa9
k55RbMwoBwS0c6oJIKJClqAxyTOnEkQezxsoudJxZ6uJhn6AfebE4fL9ZxwE2y+Y
Wu0lksP3+uY3v4pmR1laDb2HS4kekVEL1uGnlLL3IZnBL6ESc1HCoVdEhhFaHKAl
CynRiI/rTLYbFt6sEhdKLy8wmeGRj7jg3K/G6rfNctErXAGnbq7HZZVFEuwwlfIo
F9d6hKeKTAwSVCc7p5bgwGvFFeV1eNX6BfD2c+OfIfkscyCiFCb5baXAXr4c4+mf
jPXnlZa/QtcGllMrtHINqrDZnn3RsAUMHRBnY6JU9nzovPntGgphXuZZMtJh7Prv
k91LrT8hZ/10NkHG+ksmttYQRZzHFv6wzyRhM9ZgOtj2dFdp0+VaHqQxARDfyYX0
B/6tTsy543WZakevB/Bws4Ho1AaDWfHuA5ddhhummGF6AnzNhj4YPTG4pT1d9iMS
a4sz5rh02xZPNe5Uun32KxCXphIouzKiXqkLW6Gbt35jAb0dw7b7WQZhJOp/kqO+
BMPRm1upfixYkmjO49iLH/xEvwz6mkJl2bvRzGfnde1SYTrFiW4dDBAjmjKros1M
jZLCRuBqPmHpixDImHSmL6XBvnk1EyXp8KW66XgGN0tZyotzyZeecDTT47jeIn9Q
JsOx+rR6YLFA0RWl7dOybdzWH5Zcms+aEudQn39QQtWK7uZCiqzzTk/jyzJXJReg
GZu0D2UekZCKMnM1G+eeQRLCDt/ZvJJcfqYHLomMZD7KHwrfIUSdHQbZ/uvq6hc6
HbwFDAigGSGlK2fwZZ7TdPtBACJsRxFAGPHodMdA3APYKTsudtLajoNuE8DNktVK
n61BUyMsKdXlHvBUT/wdkyd9r3qwOAHqMlmjqUh20o69ZHwNSAUGC7Adyg7Na9tk
XRovwvE8rzDOVdWPOVSTRwyCaWQ4mTi1tnNy3accSWZPaDZUPKwkMvKMyJ4uRaup
rn7v00KXaHX2KvEtJMRI1eNdnsoYiPRCJdxX8o7+tuZzOPx5j17vf7YB3JTGOOq2
9+Yyp1u5xa4edmq1Kjj7aS7c/F/djTz8FrE9bG9mJokOznLv4n/ZSJtZuHDkP70W
msiDsBdV245+PI/rqRu6O0OfDI1HTEBYrK/Bjj13C6/IU9lFpUlQrbvPupL+CseM
j2mhLjgdvLvRZPKOsUuLdd0Tf/NlxCdsD9kAoa1zGzBoBqwW7yiCZJSg296yAX21
eGnOe9GYo83p9WSKKA4URNUGuM0yOobDDT1g5vFnf27/hoeyEs9IhthrVqsc5hu5
THsu76fMXgiwgOcS2FhdBo/1Kq9GB2a4ZEyIzXdoDFxeaNLsMbaUpKrRozUo3hS3
Lr5BqKXk7uLZwu3L9eM+2vHoWLtUcmtvqTnxpjgMhsOXgdeJcRqYTexxrs2WcxUr
cDMm2Y/vz4V5iRLHVxzbh7TxNOnLIryHC++777qSIeFeTXB+W4ki2G5+rGOWVxuj
8DcJbqM5rZ7aN1kEWUZSvH16TACN3XuY8LXo+6K8ZTOv1DGiWYTRJ/XBljGTwm29
6u9Q0sNfnQuoDiBxD241UmtVIEjOfNOBWTWFA8r1WByF0t9JGHVncE88Qs+nWXbw
77atKPusERqnurgTEvSz26o3oNcrUIQeeeRMk4ou1dncN+egD8MBu/nrp50kcvdi
Hz2SQbXq2potkuD/wxBPOjGLIKZUu/bA2YyRWq9PtQe/5qOKijibKkgWl2M2/YZm
xjxUqBtyIGie308W+rPF/026wTFi8HMlIDaTldCj2krIYhdRag6YyLmrw9IrJJQf
p/ElqIJEn883gdcE3RDtl81etEES4nLPK7iLDNZIGZeGhZXSr7p09WRautLOqd2M
bz3meVzJpBTVgGLhlOHIhtcyvlfXCIiJRzVwEJrWhh4zT8mV2me5dsUmUbkfkLHV
nDmXCXUM7NJfiHKxnLuRY38apEebJ2Y3nQLPrcfyN/2rCw7FoTXXxxPOspWNbMel
bfD7sFNsFods3/tSLmpPPSiwxb979Ff9K/0k3aHz3ZzsS0peTv0B3RU+udX7jBGO
zRQC6c/xD6Oc6HGaUqAFh4VkGtmEIPVeayQonxgNjviyt9JU8MG6Vy/6NxCQJjRk
mAqOzoJLJN2c9deuyaz+VYm/fROK9UvXDxLZBr9q7wOHEAxKNNkRE4Jxuelsa3ZS
DwGl4PqbqBbhun/neWpxvC7sYxOreufJDc5D3o4EK08AZsNGM5jI/eRVGtGX9Ecv
8b8FlqW2+susuemKdG+4XoUyAkyq4P8xAjjtKAKi+zATb3BNfXv7ZvbjapbT/8eE
hqGyqjgofgL901QDP1azdO3/X9ITw/S88h2sjvsrPar1tHdDECM1wKA4b5+pVAoY
d02fBebM/tXrGdMix7AtbysJacmE/D1AQwTMCuQrEj6zlsAg9EiioN4zLt9pDFal
uhdhaXkQDR9S4k/nmSZrvzEUvedfYPFpNGABS9GLUww9levv9DRgKEA47lbYnL5e
VUShx9pHyEj2/5fJsmKlssYvDry/MZIqwYQ6v5U6m2nmpgLdhA/nUrOjcwuHvjw2
JbG0nbBKwNRVqHLSewGJoMdO39i5iS3w99/HllESjk1SHwX6zXR8C/jmSK2LwA8V
6PKlgXN9Ejqlt7kJL6hBZgeK2I13L0vCGjpArpHrVZohpH+A8MzM75MEs12Tvu6q
+z3aZaJkCLA5k2zGUWe8fsY4HkzETfDnO1bF4bN3uv+fkjMyjPQLU4VhcAr8/nyU
Vt5TM379TDnk+zXnbO2ZCcVYXgPf00/GejDy2QbO6fKF8KDx6uNRxDmIGILO2BRy
cDzRKKMyt7BZjOMt8uoo4Ed1DH4n8yV/FrmbMFVcA/r3FxGmAyPe+WQ/1QZfhfKe
lQ1Bmb4eseDhDM6oWes4YJ4xC7nwyuDYhBt7JWFXhbqTJYIa64edO94SGqX/N+9j
Po25aq6ZQu2oH/B/jNTd8Nzh1FEm1QOPI37mXO8PFVHY8U1g5ItWzeHxtJXlGEdO
akBnrKsxrWZEF+mK4XmDcgI+Gfom5j/A8R8WwiDjSuTgglEE0OI5K5wvxeFv7MOf
pFosMhCM3l/J6WwCL0G5j7IL41xvG0R2sWVZj4LWncZoworvzBmRo8D1uwvSC/Ty
Pw8p4CaRxb0ymEgWY0pcSk43ncobSmvxqjS8l9RcNZs0WRWy3Gy/3YVfm90MwbER
3eSpo7Qm1nOZP1j5NuY3UgaH32Zl+1Z0EneK22rs2rCFItdOANbneuQ/Kr+rxn5+
Vqhj1o/OpD80/nZzmhPtYXiYtYK3kGrGvVH482iYEFFzzvHw89L9nsz8m59L9y7j
AFkzGXtBw1NfzJqoZmiKeTqZtGc8wLu77U3X8Wgp942iTzPFo9RyKu0i0iX69VjZ
w9cfJ4bZeYYZTeEsmkpXu7Py6qeFYppLVFW8F1kltvKzoxhOiywXp/UsUSnmPzk8
4Qwji2cDsNkB0HgBBJSBQUwTzRV0u0g4fx8vynuUggb1joYQPySonWRWshrbVwZ7
GPI051KwRih2j+bx9axKfjnifmJ/BNJj23UxSA/xhbMJJDl3hu1ymi9v2dX5Q3r1
DLMHawGoHVcI1y7zev60RKvbfO2zPYHYsN8f8mHGCidyoXhwhzEV+uABMV81CdC1
adzKLGIW8m/PwJNNpCW76w5IaWb5pzcxmmKXWAHMajDCe2fSJNoy088+j0+A5qH0
pQdnwxynhHboTvXP6fm7/2/FwhZ7RAR36OOOZ1xFfNAOM8JrRd6QeiK2y73CErAC
tPcgd6QSgaq2c/gDnZi91V9ZWiCjwF5wO/QIuqTqu5fzK2HfeSMWY+mD6f+jM00M
5eLZjlb03qWbjEOtnHyV2PuZiR9hyWAUnMqXMJRrPbT0VRUd039OqkG529jiWkfI
hBsj4RevUjnzNooFsORjMvivcCEOb4U23n5lEGO3eRhcZiQ6DGYQMd+KjBQWqfYZ
V0A6RP5hU1DZzCvW3QnSzmlxRyBQ8jQlLIpuJC8R9BpD+LicmFw83cs9cynpAXPS
K+Ly7jmXQU1LTsxM8Tf9YdEWexhOyHxhmuVhduFF3oUS3q2eh1/OpYv5GJrjsxto
4csE1dqQRwejQdEOn80KM1bRWwzA/5bbtYz2fWpWvvyiyeOFJft1Pv0bf0pRiShY
kUtJK4DjqnU30XByVkvbMj8MlmZEZ5NS5hcvBCA3S4C6nVRYQJ0zL0GeZLM+i1VD
JrOtbZ26kFy58ahWMCBwYwo7oZGAdTISy5Hx9+1KOk8uObBnUCTNA3tbGKW1K3xK
jYCfjkEQ1kOe0fBB6ouVRq8324dnerkq4oWHyymEx1pSFEfBErpuGcBDhYKDzc57
OfgtVSZXqWdoOQrL5fBMPjMv735Sy70BPttipgDJYcQH7PkoTnk/VDMmEmC4OU60
EGN34ytj3v4MQTWyP0hYkoe/YpQe7PnMKWws5pgM3U/RvNKOhJagpjRMIXC4UFvW
ZNKANP7+/1HmXYh3hm4SmYRGaM3TiPuM+eOf27hXncTcfGSItaBQb9QnTiUtikOs
SNVJjACLnJfBkcBSESS+BMCss2kKjgcpsm4QE4BvtmGPHAsKl8UasRp4vKBTQ46A
0kbIF2qOuY8u+6bwJff8FWCADF76yE+vmc2Y+K1VPsX76Oft3RqeVfz+/Olpp2Hk
K/IWBaQwJZGAUxZiOXB7/0/2zyQciUQh1guK0gGqvf7eJCi/FXteURG7KWym9x9S
u7Lt2lVNsjfkqtO2tswR0tGqSmJCRha8P2DSRkytYyTsWdkB1x7sSOsjDK2/nyX7
kfmBl/PtAqJd9w3rSzmFDccp90sgDGUmimsNYxJdG0A/RQXrp1EvsTizcvv6j2iR
99IfoWcX0BK0TlZ5RHbd72SdceQj/F0nIjDdVV5WeIT4DBxfcmQ8GWbfUO81d2uS
tL8VAScx1moW2qEHjR1GM8YFSdSDd2EmdD0d7vjOFn9UillDju/F6TQwV2juFpcY
xUFPydI2NSBNYDOif/CErcnTBzBhUvEt54qsL319x1OsSMZv8Pp5UEztJyhH+uXQ
HOrzyfPNsLNlZkXqdqIt7L3IKI6lFTWUFZjonn8GAC7kM6ngaANTm4nny9BPmfwI
pibA/YFIjsIBlY1CzxvnomVLH5005WlWM5GK1Bq6Fdb0tDjk+hVqv1FNONRzWRAM
0XsSY6ocII0dKGktCUGn17ScgOC7jE81uNO3XzQA1Zrpv5/UaosoTW087U1O/jRG
HbyOtuuXknvj8y2HDvvI4aRfFLwNyhQGs8x1rSVl+A4efKqJXNkq8DU1n6Dg7+z+
8Rmoc3mim99yJ1SvyjrpvH9MoAXACkq+7BhgKJlFXygFgIyPKuc0K1nSph3bBKAR
U1XHSNyuRTYQUqi2yN9sFCE7Oq6tozbciwTJlVrpJup9G251rq47Zl+256r383P1
OCDfiq0UMGod71+/PVnuEx9pbFmRhNnfc2BVXc7Ejsbq7GPAQKuFNgpFL1mb5bid
GJivd1mONi5GHelOhuVyPBa8UQzeHcUb2+F7uDIVxpV1OydKuQlIPqGN5xM1CLnA
FP6lVo68ZlTpPq0VKDQs8HX/MDILzLfLar5nMIdkbiLx/fXmQxbJPp2/7xXfCx/E
8j3FlDq+LarA8u+v1SBel6xjQ7onzut8kgujlUos+pXzZ8JQAIXvKZ99C73impxu
mel06/sNKoFcO9jPPnVP7jPPova4rYB2xVocHLDX5DzeqYYqplvzi/P4qekIgAPd
U0BEx5ige594LzD+qSoC91dBBd0hpEvmIZX0hpzOHn9Mq7h7qk4ypgBhIbg3ql+f
S7ACuJi3eJAfsYbR2w/nTJ+iXgNMvmPF7BLfWUrY4cMbrVMI4eflpq6UfhIJaiBe
eMUjUhZtI2HNy0Ub2bR7l9RqQRG29NjQp5MJbm7nRknDCxh8jcRWPVwEfXY0Ihb0
kxV0Sfy7eib0TGuZJeNW+1RB9G7psD+ItWfu4IE1yf3+fQKHJKuKUZmCLIwD09uw
5FjnnbZVhBJt12MK+0XgT5x20sQmBeuHHiwNLMBYFgo7dd7ySaqo2XRq3qitCv/z
zDujWXfAUDh+3Ktm/bKlja+ybcIMTAZ6kYNB+l6KPAvDUiz5aIc8YW1j2n9IHNq2
1DAhmU7/BVvzq22NS9ukUWlU0YFhh6BDbMbG1zyU1WIOxT927UCXoFi+DJIhBHOJ
ox7U2vs/lwiaQ9aQnKfjHzExix5QTEiP47LjtUFEpoanZ9chbVr9IuLUHaJLCAeE
O4lY6MgdYm2+WaLw6QaRCHNLKE37tjx2zAoLM6QLM7fogtgt0JWf8nTpF4wVQpqw
kKgUoiRuHqsqwxgxW+v0WpgLWqG+3CSSvz17N3AyHWjFfW4WtOwBO8YJ0LBeDf05
klspAF5oM7+vIx4L3jdNwTW8jN7XEOOPKgx+o3eMtb9rLkKX1U3KAfhUos6Kgua4
zz1pLV7cVqGn7gigyVD7GiwfqLJh3SV1dduYNfByQyVnZNJTCad8OXQtLPk7vlJ9
WxpNDtAz//ujccGG9qlTjMp3kdRT8weBdB0D3jow/u0bWI5EGfOmnJKtKzHiZGAg
msh3rZj0Be4mnR4fzR0Wk/guNPSwBz028Dq/WPEg8Nt9t+2ivjhxQl23h3BbtABJ
cMcX76BBDlBCJk5wE3cm7duWkICf2a8Q72ANlvlukRAIpgZG2G7oFHspvE3CS5PA
1WoxKg0DCUWp/Vn1cQ9UxI1pj87RwWXPg3/IoMWFb0GBPeOzjo0X/MRhrBa5Ha4k
mDz4oCJwQKEsn0NeBqumh1O5O+VEr9gBBOCUyxIAyrsOJlAYPD6PzOJUS5qM66Sm
AgTIioeqE8vRL0KWUM3d7NqPewnFGFfvMnKepa7U6C7gUZCB3LIuFWRLs1Q/y11P
FfqZC3S6B+DFhOTGPaHOLpjvJ4L8csSmFJvdsT5R97pmaLxBcluXcR5AA3+uZux+
KlJ2kJivjK47TmjKas+9xHI/iYlVoLzrlpeaAHAF/ATlCwBC2V2KI3dFOPLT9FUo
LKVduKBNvW3ayYDiwrldrKOiVpPrSjt6XWV6Aq+U1TyH7nEluEYb/68i5uSxWIOL
Vju4V9rk4LIk7ZbrjD0RYgGLz5JHWT/0XGREVPh4g2qWBI8tLvqc2rf6Njy5pEfn
wyN3zCMvpXZKUfMeJyIIDOthktX2wpZgNA4yHo+DLSHAnG20X+aOwd8/y7w4XSqX
vXo5WA0b3kEq8Id/RVqtD1XPUu23Sy3wwwPJROgG92Ei/9nLVYgq0T2nKU5r1px8
ZaAFXvl5bTdKZTeKxPQOQul3J8rRbG8vvSRO/668o3BINmvJJIRyW+iS/p/sLRR3
1g1PGWhA08Za4kk7ivDExLFHa3IOlxvgi2AVuNzWiPK/OJxT8BI5zhJX3MoZPbzM
k8w+i6VWkNV0LMrDr7R8CVKRTJ4Dbi6D/oaeYisKJLMrMqmedSB8Qcr8DnR6Uo3s
mO9iRx4TDFNjVRyT2WBoExfzJmjWk/BWOA/v1F5zd+3YwX1dhRBzICxdEivU+JjH
hK4dj0cHYmaOXvwFXStkKjUv65+tyK/ROxJoGsB+poxH6eLNRpCz39ftxrwx4gUT
y3barm2xVsiD5isLZE5u6jsSToLyqnIRw5CXice2NH69r/gScGfj7GUVBc2/tSCu
yoeL9Fqno2me+QtiH0M+A5korsSF063Gt6V25YdSX6j4C/IYYbzJkiFltz79Y+I4
7m5dJg66YWu77AAhq7DqCzTUSZSG62QlH3o3+I3gNF/qkO6/quz8pqV7ogtNEbhE
0oA8vZjRxMA6mYH6K/LNqnI8F6P4k0F9vL8MN6FPuKEeNWKH6TKuJCkMKGJ+b4Tm
cK6qQtKzjL3YXl5XcLpa9OV6HPgqSn5sYW+KTF4GPwrVK2Ny2UsZ4WtBvVIG2MXp
RtEUVx0QFC885NX69auawuyBmITEetHS6t+YyIRR7Ct48TeQUOOJoaOEMZ9RP1Nn
oG1fSqRSVC9kjhAJkGEBJ9HdgQ07tCzWM03pOWi7pldfpI4Gee+36zfescKlRusC
qpntiN6FNQUF2DLzN9FdbzNUbR9SRJidJ/GzKy+C51GIyzMRyDz0vNtciWpI97uE
AxGhq7E1EuLJLszLAj1UX0+decwz20RbMj764yJk3rCsYw/NRbPFKa31A9FmItGx
Sj7RmQEmbD1fG6hVSrv1l0wzN1BePlx2mFdSCRJc+LIe8ID8dEl99Uhf5scWP/He
bh2FKxFy9MroCpjch7BZlFbSlsnSsh2qhqv3KCwr+vhta4/Puq0dPLTuuMXzgZTU
m5NG8FpUfJmA4e4kNOcjdHSA/WjGi0o3/GhQMR8uJLSYe15ZrMdnPe8uTlX7Rl+G
wKGWN5yTYviOFPeUi2k7IhWc5eAk2yeNdAQK6CVkqBp83Y1Uijqmp9kD1BSoWvhA
8EVY5DUR4868KozW8JdSEk8GpiXkYz9pX1EYHFpSLfO9qvL+epb2voHIfTsg5aNI
oOvUOFH2+1ReAxzjf61BjpJalE9SlfBVI86K5cWn1ntaPg9rcuy5rZhlT84WGOG0
3ERCPZMmdHqLyO9l/qd7vMs9X676ztPaTRMuS4YPGHQAyzWzt9zZc3d4mLwQRiwW
4qYHSyvahBTwyX1l5FbsGh9g2kid+98lgmNoGcZw6APZBJDJrKZkreVm9A8AstWX
aw74ztepSaWzddbKsLSM4aUOC6d27uEJ5IIQSlFK90OeliofYLTPDCmdRXF3wWNa
yA472ESk3FlGSWNW/FMHTcYzqV0H59oCcx3wJAGDB4So3VZY8D+p0yrLoGOOX9I2
EPXILmQCszYpwiikSbM7cEViXfctme+f7+BRDNa1EfCi69Yhddnlni3Pjl9EnicP
yjdd05a9oQOHKHccOAMC6omf6By4/+92W+484yxhFm5tvYGItj1emlsPcLKCjXC+
3DYPE8aD0LtGe+pE4NB2h3mXNmoWh4+R8meqLIlZ+W0r4dpGMa1PDam8+62j7Z8E
hGQe0HzuNULHsH2U79R/3rIPQdD6BGt9vSKwyws7SalehFclwwpU25w453MRt6qD
1b4ByWjqJ+/dhZBQY3FFIblSmFmWjxchHXY4IZVzIMHmE/b3DixAqsJPddqsYA3L
/K3B//L8cF6OQlm8jbSdel2IRfUUXgnKbhlBMjGACOJJpmNayy9X3C9q51/mv0qG
R9H5Zp53S0Kt0ZuF/jjego3fA7eQihmNrgZntT0g6n3tcy6/srjOjx5BtydU7pLJ
g3Xi8SAw3U1qQwdpP/bhSHhIlOd0/gCvBC/yy4iklJCFOF09YGIGlKfA/arQ8nf5
fj5jBT4tIKRNKZNZtrtt5lJbrZGJbLwR9vbqKTXg7v39K4qmqIIF/unYMdqJiLki
eC/1XjT7oMgoBaxUZxbS4XbP4lD7MlPQt9bicoMmu1yDgRsL0mAD3ifkYon+4V/K
wNGaWtoZ58jm1bWNNDx+5r2ZaNJRRGjwC/MVfUWUa2QN0TzlE/d7RzVHtIcioIP7
98gNtI2wM2gNIqUCk6vO5xreZkcjiRwFaq6KsJ7gifk2HbgC2izrRqy6TVZm2BUN
V4sufUePgZmyC/m4Bo+cjtZlyFIeCALVf+HFPOu4Iu3aURDHl2sJhTt2mIV2Hlkz
VLsFipIV+Ms9F5URGMOp1+XeNFEQkfm+sP6VfHfFpB/iPlaTDGesFtz6f+kt98Hv
tyx8zydh7L9HBwIBsqPBQpKG0GVfmC87rgoRqY9Dml2m382K0xW8uu7cOYB6V5XY
XeYogOZS7YB7EJUrpjCJddu1TN82tg2gDfuuwmZqQytjfWb4Z+yOd4mDmCvXxWXP
/XOQl1JiJvGlEJYwcwcgI0BqePPd9irphl54HJeLHHrAg5ktATx4YbSWzGfDcQyQ
+aHXbL6iwuABHQa5QPWduNbLIzOJjUkQkWJ7eU0OrgEMdo1hsjb+dTzh9+u11rMM
YElv1Pad7d7FG/zbVFbFkd2qXEMxIy1foaFMGV16LdLxgIf5zaMqjJvNiLfMbc27
A8DmO78W4IW9GLaKs1WGMTu/NC+Bkn0uFem2tIRdb+HMxJvkorqGho7kPx4etfob
NQ0nwppLLaRuh48OUf7NmrmftPDZOa09sRJjqadZ+aQgjqZgEO2WJvGpaGU/5e+g
faufCazf4853mkRMRYo0qH/ndNoilzLaoCWxScLCQIOhM0Kkg5bwEi0YBSP3e1jA
tmgbLqTbFQ8L2bOBB23dGw33+SSNMjlsL4xmJpG/THe+Uu4HUuHb8e1vblL7aGVL
DeNo20EfC1Z7wcXiik21UHEQWrhGGKQ0fGbFS6V/uaVMsc9VfIFWELe0ihgyJERZ
zFAEJrL0BrQz8+K8VNpkWUtQRlkcpTHPc7t/YZ7Dr/hxN1UTgu97mMRgE+qV9n2Q
EBlVN3N2Qsya+5zFAh2iPCS3MM3wPGDcOGteSfQyLMjMpdKHvTCWDORm2r1j+V/F
IS9NM8qSZ7dqEFAEOhDBzQmWnajfxcjOjAu7T3q4l3qlfqEEMhrAJSxfvgkCgqIs
JR1BW7qf829077G+UTIjVq7OIKZjC+B9Q9YMBC8yxHxL5JquYVPJ5Lo/rMh7KLRM
viyY7v48QTJ7+3yZ5UaEYI1Az2VrqEW+b98VAtpY8CHKSJUj30duH8QSWdkX+IVV
p4ABcjaHjc6DVd1a5IMUIRIGge2m4gvSJrwSAWfur7c93K6FCKUFJuFIg63KpwHq
Xe+PrxWWK7C1j7LAC2SGRWvUVtMKABwHCcZBzLChrmyMRs6s7/Q6LijFI/+h9W60
JqIfURhDBZJuUYdQk/SbzeNW5imdEbCAIVSYgK+3A3vV5l4fDXauEqNOHg09TwLU
7zeG4wQmmcBGacNqUcxf9gVR68z0PQhSTD4ncblKI5MVJQZBzqx1UDLEtmTnjdYA
MDp+Gq4pSoBKrJigCUjCvn8Qwi/dbZAIYh+hRXpQEPgqFcL3bEWCwS9GWPy7gxXy
rfltofs4jXAKPbYeZEebb36NVPxjc0Mopt6jAUvs3oZ5LgBW73i8D053bb2RaArb
9yXLhVm+cMsh+t9JuKh9kfiYAyaYc7dkYQvvc0pV2Yh6p9PStY54WnIAy2/KmuSG
URFvOISE+IrXnVwDqzceQSZFjUaOi9T1YW+P/RLLXvU9+Q0f8U1TDzfKNlobnrrR
YwOII5OExEVGvMHVilc5W+lS5b3rxvkoTulnRLj/zMnf/dACGscBHlXs2HheZlvF
o1N0bv+3aqExzXy0qRYTRH8pbC4J0YAvuXguWz1k2cdbD9kCEN2EMDdwyNK6dDsw
H/EqyMhtLEQ+l3XUAsaZEGlv0jVlz2UdJBJ1QkeNzi6UTE8NsrA9+xTRrnF7BtCW
nULlkA2bntZVkPYI/JDR7mBEuRiwC6caUY6o2s80GHwTJV7ulp0CRDChMFQShR+M
4+liobfMUADyxRMTONqT1ybBTEkogJ2Bsb88MGltYej0Se9qWpZYSf6gjCuZfyPm
MG9ynSjYw/EMwJoen3oBi7W7gxgmho0bjkTBJ+MfzC0NVy1TCc7wqieocsvdyHMq
HTcEIavxexDCd91aC7dtPprnxhWFojokrkFRijz+7tOx/BMoHKr4kz6I8Vh71rN2
7uo2DXNJUqiM4gSqbRHhMHYfIcJlGLzMGWlCInbD+chDbcKbT5axnTaupoLJNQEQ
JtVmNZud9iU6bPdgRdrt8huS769y8dnHE6zwG2fq6EQEZIaxF9cNmUU0ttPNmP7V
uWJuRwGbLvPClTXlLfDNaD7XQbs6DlzCNXUV/KnMgB8G1VSD9OloLmNv0fDHIIX3
0aR7vKT7wSbHfIbXCLavm5BiQj4ESFOr68EAPRtSROhN8Zek/lJNOhCaP65jdwol
AHCReTr/lXv5RFIlWIobjRVzJVPjKd7KjkCLuQ84qf/mnfy8PnOicnHI+222Zqvd
01toV+QfGdX6zTw3F7XWYngrZDkjBX6x5OYgfv5Viqg=

`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
MoB6pSPfFGkrhIKSUcowAbSBy0MdaEo/vC55Xq9cJ37rkOC0wQsn+VNLCkJZ2/8N
GtwD2yb8PmZ0dEjzrC9Jo+xPAxVSL6kbpzCgqU32rPXDoGzcua37imrIu2kpuiYh
7s8KkH81ijxUo3g3AsYnXV5xYoKt+nZxhtBeyrJxNwY=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 5440 )
`pragma protect data_block
sl7BRU6M7YnlEAfCRiRwBuPOdYhsK0gcBdyNAd8V8WlGHXuoMxNAFL2h70ISQHMg
FkYNboqBj9fVqJCM+Y/+QJYYligX9WuwbXWdTuVXZs+fHZgx76ddODInraN32XIl
7ZIrS2g3TQ7Gg5CVZScbse1FppamyZkZuou/mG0O2s1/FPbblYfXLBF8fofu9C2X
B0I93I3cjlsk4YRCvDdEwAiI77nO7ZYSM1NzR8qTHdAJ3sKj6aV7BjPsH3D2LY25
s16oZ3QF0xwatoZT08mIky4Jw2VnfHxiacVdNZ14ukmQQFu1pum03U2CR12GB+Bt
/iLnfaCksARtOCY1UMOx3m0AjY8wNDA1Drn93bNMgRhhykKDmsnT5l1Kgdrg2PwU
5zz9EeqTLXBTXAMMKEjdAq+f5U26tT2K46iKHIsWcdETkk+L84IQSE8VeMft+One
bz3qUa7MBUbZqcjN7VAet9H8bcuWDuoDjGicrL5PWpfAMdm7f3TDWsf2M+V7JaA8
i3m4x2PqBqMTUchj4fNzHE6NAqQCevyPep4KUCX4CfeOE51kerOjdDimtnHoXcXi
wEtOz143cbrH4YE8OiL5WBrY7SExclVlyHSZc0jN/5b+Unj4HwcpsnlEACZZwH0l
lyd+A1ITHmx7Q+aKVxC7Jyu3hS418I2WouMpREfz9qbigtaYfTOrZqQB2BFbc7ym
M43mzmSfoIA3eejhjDsYVXnjAwdVS+OFx6L/DBr3ssjZ2hqRorYyLgIPMo2/SqOg
DmXG+hdMbk5yzg5+eaO8LnQb49xcXIWxPy/26BZ8Rj09+yUSY4Fiuvsm93OAsaV6
kmzfEklujG+gk+h3aS80S/tPI6hgIIToVLjbUr+b14abwrcNRN53plPwosxLJAbb
6eG+e2DRYq9HlgQX3ACwoBYm2X3R0isgXisKVbgBpov1c6yz6wiN2nz6pRJsr2Ca
6+juXgRUpOLh+g7BraF1ylN7izdmSHmnwTLblO6be17Y/YlrvyRxYPtlCN6KOkla
lholosRV6PLOc65BgBXR9sP5xE2YALnpMsjSxHKzk6u7LW0fBPm+Z7ur0KojQdpW
/xI1O5PQH7tBPlsULRrBUM7IUYT9fe8jF8YKWsfVhZNiOMccixz5HaMyHKnMcdAT
BVHTPw5mr6I781s/KJLsmSfYjNHn6Vwb0rySUjwVLgmCjgHyZkcCHxBBL1X10T8E
k7v3NG31zgL4c7xfpnj6UD1t5nWzG9Py+TVlO2xdHRp8Ne5462qHCD5pmCYaho78
IM3FSVFX8Q8YlqrqpWaHaQC1YmFGFLoA6n+YfLgcVlVXz6h3JHdQfls+2rNKAQCt
QGGdqQGifiY9AhXIM3EaQpLNQNjRncbXpCGLGFxO4b6sOLnGMA8htzOSm+1MNx3Y
qyZuYE2ojuxFtHL1+S4Ts5bjwFJ2pNLeel0bTrR2zX/bSHeORBOBqwiviE5HA2OT
ZWFHH6Leozo/GALExiRkU8SJL7WDQiwpH78hg5sWfLg+9l4VjW8Wmg/Mq8uob3e2
NI84RPiCt9Vo+kjh3WnP0XNfUheAjh7P3y8kOJSXwdB4/eeDcFOm9Cx5SGrwzYUm
VbBhgKD5xAuN9vJCJdyXqCgL5GLKmvDPQrrDqSp7Klrq6A5E4UwJSCNj1zr1w+mW
TtqGFK3AfgSUxvTDM85li7IIPqpobrqXpeNNaZun3onDaRxfDiUTKqt+zqiLDCjJ
ejQh6GzhoKHEBNmUKsFJJeCssypoF4FGo4Ppi/Dqcb7dnM6m5XlmhsHzQMIV1plA
Iv+7bH75kVvPipTNvQJwaRCifIfUmEfYf7nue3TSPbV4LzKGt7NpdeX1ooTGFrJ6
ProZQL9oWmKC9m12+GAoOZzBXuEafyZD0YRwdr4rj0eRVxvxSl9m05pIaEnhWl/1
xRC0lWSSu+mvwZUj0a4tj6aEq7EkgrXY8qf6VrnFuT4jEeg+eJZqPBH5p8aFFx5p
SChoUyL4sSAad8FWTaqgxQPi8kZjgxdqCIv5A/nez89tHtZP3U+s8ywYnZHGrJ36
dMN+hqXIBshTIjI9bvi2YvyrQHtxOOoaZroy1PZNxuLaVf7A1WjdW5iQmeBE7Mlb
2VGAR928Z5zx1S39mvqSRbmtHXEq2TfpMdWE3hxbZXSY0XvdTlsKq9N4Auez0lGI
i+V6+bnIN76yDZRSDS7wF2R6ftAoTmaknxNbNw0XND3wGShGkLDYj5FCVVwDCv+i
L7nTON0wZ6x/Sy2/My24G3EkWhum4yoT33GWHfR8Wylnwok0zqL6HFjQhVK8cPDt
0KsMc+8J54hMYtGLJJkRChgsa2YAQ4/WzyUxMmVuZuZUHDqfvCnHbq9IluAbeqfo
PugD9UcxrlHzNzLaSoOYJAyp30cXB1tsv+ekmisDDRDxI5mbAl43dSfQ28tgAdcs
jkKOESJ4E5rZQeenZujnBSZO9iqFRXi4bdj43nRWHYosAy8S44AycvYUkjsd0TBP
/Rws/pcbxEDYko2FxbxsluY3Rh3wjssfLE/00e7qUEC2Aw+mKYMP44G0KvQT3Zwj
0xMPmC7LbQ+LnHQpxf+0FYZwSYOETedJQkzvKyYx+fxH0vccle8g0jC41GaHuvuf
woEJBRmwHXdb/nTLxdKZF+O0AoF0uJJKSMsK89yK+QIDoAqaulKlDwrxCgLeDS+M
QnM/z643DBaBB9eExhKLJoVN9J8sX6EquPFY+2zTr6AIDLr8a6BGjnGMhQS7hILx
jk529RWxUjSCMjsQwnLOlX9aPRIPtqear0NIHtSU3Qki77ZzxZZQ6VMDSkme8eBm
1rDvDjrRt0tlhAGni4pSEaXL2ODKQrsIwWAIO8nhktzVUG6akBYR7OdPcjXMTOqZ
Y97CQPtspUd8zsM4o47cB65aRzcBIaUGOepELg9bOZySmCr4U5Ibn8WfgosFAH0H
JXczfw0GoUnNM2O7Xm47aTEvZlxqA2SYzU//9tdXUHGZ2OUkzx9gA07PLdk+AqGM
gpKfI9jjX/nv70n4eOus/L8n5I6s3fkowtPI2jEjlibq6m+r26PYKlP81F+1Ivy5
g/3yZVKdYpK7sU5aVlO2UUV/nXTCQ5yjX/a9U6rl4PSzuH4P5uObmv+Ir8yI+2hs
eHZ74lFTsVoxs+Syw7+Z87RANw3lOdgb6esgqxIzRR7vH7/31kg6BxhyqE6LYdFC
Q6G/mixOv4eZpZDbka70u03QU5txzk8B2lsykK911QHgUVgKEUj0RULG/wRKHESf
dUFI+VEynr8s3l3XKCI+BVVPM1/X81b4T58Zt4VCU8MVhRBbGzkn70BWZ0BucgQH
YjtzVEnN7AucKtvRNTOBi6Wiyx3oMP9L07EEea72MaYeNtG5D/BfwQVHbsIzc8Tp
JX6XpTFOj67djLPT3hZJoQxc7Rrb8n5ouW1DB2wgMgYCbB2lXljBoEnLeLQP0Snl
UTQ/iovvPD179VvBMga9CWFqzYL+qF0j48c29rygsB8nSPR7cNriV1CTrA3eexIC
OVpn4XaNNsxmGPOG5bUXWW9ipp3fOwSck1oIwBYnR6zRqneZnoE3HCeFIZXMULQv
lK+m1ybkHCZNIKqcHUghMVLNNvtza93cQr7mswJADSLsCzCbaCZD45iSc/b/K6Vy
8ov0uj5uDypVw+9B3vcEihLUwBfpW6A/VuWFgxqbf8KkjUrVo2g5/LiJNCqqbdZo
H1EfL3+/Od3mld1jnw9g4VMvQWuUIXQ9Y1SYVpnk5IQ23V6NJb0TQQcbWcHu3hnI
6/8/ofyn/nyhna5M+DVr4nL6Q2imXlwdzW51hMqg2PDvdf9B53/4Jr4tdXH2PxUH
xWRY4cypUL/nB9Z8EQFJ0BlV37teFMbKgyasDX7zWlGy/2S2Z6FOQ3sx/jmyPNr3
n9rfE8utji0fY5xnBkymfpI1V2Q5oTc0nhV3rEebwP9FLc8eS6ITJlD8lIsnDF0E
qHPoln1SH590/kYz7HnVrjzYtQ+/GfyDFbWQmtk6uPccRxcLbfu6lAsMWY/Ta4RS
K7b6LEeUYmJSPA+b/rTc8YVYqlsj444N9GldtUUva1PYkHYIhHBZd3cazegrmPdB
MYpm4tcLogp1Iz0sDzehkEwzJ/flEthSXJEP66r9VVM0YlD4thqpb4cgQHWktB0H
dCm//Ky3zSCQAg6LezwkeCPTe9SWQP9u2C2rpcfB2N15VXwhkfep/G633cZKYrbC
fkVK37wJ+d5iRywx8zpoBE6ESsuARV9j34lr8vjTyeU9mI0EO42E+UohCFWndsrY
HjDymBfX2jQd4mlLJCp/2f53F01CnJ13Pd297z3yYZ3NQ/0qB4xLvB/jcslAPjHK
sUHPhmOYEIakinp7EU68ZCKLIbl05DeaFs4Ejh4QPm52F0JqkbcRZOnSKopW3+tq
vDw0OzqA2ONTNKxGU5NiXFq+rVfXkzmf8dwZ3PTK4b7D12rBB893d8ZJnlefiv9r
GXEGPcq4xHxiTD6i3sbgURUNv/cUtN0pfLPVqUDmuMzuV+cz7P1uV2FRVR5OgRXd
C6vxqLbW2Iyt2JiFseBJrItMNPFpBn0HTIslaUpwT7mxxq/Z9DxsmOTZsASBJRQq
Zl2pCA+EQ/DJxRgISddkQ0npKEJiQIKAG3CW6ZcTEeZy+5QhFhZPKab5PN6fSHVL
d+B8jbmvZsJlGPYCM/VspY5QSZHdo4kw4QQzV/MBeaAXhafk+m45F4aGjbmXauIH
QyGqiB8DfDKFGRJr3x208za1z5Ci2vAt9Gap3k8jiinJeyYbfqn+WZfEc7L6SuRv
i7Dpol3DnZ9y8gqC+tzNVxGqivdVwqegZdNY3N/v9jDetfBmC5OrBMV98QKkl+8M
KENKZjinksvsezHfONbGRM09Qzexo9nnTOi9J2eN+hCVkBvRtDt3dFwccWuolqCn
u/dwhwflWniqEd/sYa1/cKd0jt367f3PoDi54y+9aTpeCad0ea7z57MQ6isO00Lx
3JzmAn9JEDkw4gorXCVZ+UeToo25UYUw+HfZHSxmbjml4o5IwIl9EgQcuFWxEF5Y
vkBEXFI4wQsmMLsK3yd9N7dMz++0oZgpM+MIj8NxFHrFX2TIXNv0Z6Nhf1ftw9dc
zo3ytgaHexcl1UTe36IrmvQr8c/B3Rts+MWjW4ishI3SAymmfZNGEdos0yC4JWiS
9+w3/yo7CGLD/rZGjob2FEQI2N66PUytCEW9drsA/enx3FD3Ggjp8zwXgHQBuvuf
jiTURw5kPm0Rxp/9bDejO7mM2jvSE++md4qnn72qvFeRGNFxn2fdTGACdUTAXCa0
wtJf1jTlmT/PXiYp1uzu1iDytTeir2iTpL9DDWq+gTI94NebKRZFKzCHlqeSzgys
nZ0U0i8dAl0kuo9rKwxWJOlH9Hx6APk0wVVxPaAyKVqzqzCZbcWmbSJlA/1N26HW
ixqFe5ccsfdPlpPLT90FzPmMDNLnQq1NiOkG+Szy9Ig5J5t9iP7FO4neno1ip1JC
Uwr7faVaHcf+O974irEdln2uiL1ilJqT5Dww4FvVDlolPhArFeAz2xuKaQNHdW9+
U6XkICEq9c+ddpBb9hT7iWQIbsEYv56H481/jzYKnTa7kiBIhqOMBVcIlMrTfsrV
COds7Pl4tThmcxLJSWvrLC3DG2XgCzo4XE9oMNxDgRm8906i57pNB6rUbCrC2aVV
Y0I46C4P8LGbzIn73Z42s02Qi0SERdIG23dGN0VfwCPe6KGTBF3Z/EniQLKLXhZ+
EgwdFnJMFylQAfn4W7Mw73WhMjbh+yus8fo7h6YNFJdPRI5bkzKHek6S6b1mspeW
/QZkmy70rOP5PuJz8kYMVULrukvom+mQxO3k2gNW5WywqW9M/bu91y7BJyysTB6v
f/sDTFyCY5uhctJhUObzk86ZUUkBerGg74G2muOeTbEXiGIoJ10vKAOxVOS/gEq2
7dITehBgXCgCqNkz7C3+rjFdf4PRxKHY7z08F6WYW2sLI5KlpOsT5ou0d6U3ngd1
d6xN97wS4PLYVvaw1lgnIFzpet5avpFiYaRH6+lcbF3AdXsCwOBg2400QF28Ewvj
qLFBAUIlJdaDVkzWlCYk2G4luiKqSNtur4dcjFCqEtiD9lgnHNGXQ1OZJmhDLBcv
YyJfETjVJRr5OkdFUDq/B+9BSP7GHM58xkJXglB6IzaUJONWqHF5WIZPwUGStZSC
zSL90J8RV2ts+XYpaj2HZJV6hxpE+WJUUW4wFIFC+rn/SAaeFmYWqqCY6hWH1GS+
xEy+8g3Kh+JK4vo1R/IR5ZNJKuRYplGPOv1jDwkz9Hhp5hRxiETH4o755PbXq9pb
C+DlfTTJkpxrKhGRhbL+E1M3PoUTruVPtTjSQun5PutIIuypYnwEFYk2DvLwRpwO
YukuSrtocxOeY0UfSVUnuCKXADjn+p43GP5a7i2A+ECdKxFX2LuFLEsGmLIEn+kF
UMUl5yoJuKdAHSRRdfyTtBFnkMVZfog3MGtJU4cMXrCavFxTjBrSKAxmNV6cy9Yt
cCrg7bmbiKxeT8UsHE5Zbqd5DlA5tkwglACam2XiJRBEGVhxHo+J3MM7Doe1TIfJ
tldyZ8M2Tkl8aBxwlKmAq+qG9nGVF+/txNHgs94mwT4VDjcSwNs8cKH9p+hJ9Mp6
faGMqmacDxZulHUv5SitP471ZWkyaaFViBmOIiLKzetwFUk8QImSlgGaKvnk7KId
PqpF/y3AEWBDw7gzUZnNmXQnARn8Lj9jYxi3vr99eldA6CXG0O2Tp1rHIzRzqOu2
GkppeiCzofWJ/XM6NncFo7l+aV08ysbDE5ykoA1lTgBRxZdJ3DV2HNFVAtP1jv2e
Ick+k7lXwD6aBQuYxUhrY0jUjA8FGiSmYsJxkumi0QLK5iUe83DmUnRCLEN75MDe
oJc47z6gosS37GwRL4IeWn9MHpVMg3JJYps3IeABCuwmMYvrCjrkYtfErKOXQAHk
A0ZziOxBkYSXcj/Yt7bnBzOP+JEeQNNR7ejk8yuAoED+RBsmnY6bpbsbh9ZsbsF8
cCpS7Qz4EGgb63BhqyjGBX7ZBcNP3NSYVrJyHnkleJ3DOeyB1lE53yK6h1ke4uA1
u6jfJ/ur5AVrTjWHdwlnY38qWWdsqto+GZ7FY0EP+/kXk1ZmFBlpY23Hwa+am5zD
/ELJ1rk1MlBxIlbnUcS85sTF2rdB4za9kg++aSCbymoWMO0CMIbfHU3CKzUQid+o
TjaUmy7VQPWN/95mc+SM7Q==

`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
dxxu0sOLNyFuSLfjdPpNa4JsYEJW5xwEp19rKw97SQLQYKTsQUA/orUXprOEGF43
OIrmNCpmPihsA42VMpmuTtOfM/vpGX8uMoESbk88H3aKdU8ixzYeeYPXSWFJgZqr
XeN/wcOQlAevw7olr1O0z0la/0va0izYe7Lv3KrFmamLEpD8kZujQLhwPuISuO7C
y2vdgyQf4c1u/PHeICOQKnmgp0s252yw6cXdOdQ7VzRQIpb9OKec1D+F7ARyZ/k5
x5lFbupbegtCPdbdQtj1TNnfQzfiLqdsF+Wt/OwyEaKBtu9rnLVzI4tnPVqZ0nXA
oQeYv/K2yc00tyAktgc2TA==
//pragma protect end_key_block
//pragma protect digest_block
85yXTc5XFFVGeg8eBuRGnI5h9OI=
//pragma protect end_digest_block
//pragma protect data_block
JVH13VgkRQByghTsSRv6OybARq2kL28sAxMIbGXhSJKpBP7fFuLHkyy6tacpU3M2
2smcG1zNDUYjT0bKZ3Q+UN9UOSJnl5ZgQV0zd37QffiQzI7N7mfVDt+h4GOKMwrO
FSiMTVqS46nLRQpFFpKHOp0wxtB8My7+QyZQ8PxpeaCiVuxe1tnHMJTco/oevL4I
nT2gKenVW5Vh9bCH90f+szPVeQl5H2IZjB7mypQRalDRE7UMj6Rn1U8a+0LBbk3r
Wj9CPawqm14IAiFvGk421+SwzHatpC72+tzg7nd7inoWuwuMW8tkIqBr5GKPsGml
hIfy4MDovg3CFpr64PQzIrz2QDxcDD3WtMZOWLbs+0noVoKjKRgLobrbsrI62evN
IZZTC4SmPWyHEYu7FrrkDULvx9LBStGltZjZKjq56sxespjm7HwWaYYUkDV6UFsK
aqD0NI7dZa7MySirWCprYB+W5UMtMwjCfpd/HiLYZxB7aQZ45nhM5Oa/JB8mVOlt
iS8bSTzwr93PI1LhEFkzNzZDp8oLTiNkVfeq6t7diJ4D/xJWpWaQTEkej0SrmZLh
R6xtSOn9WIjtyij6MgR8pSphujb/wu1jUww5Wc8rs8nWiyEKOB6M/xmiSFR7pUo7
0p/8iSshwRd3RNEIIcF5zWXWZCGzuHcWd18EWlLY10RgbIGc6FnFLUkMYzoAGx+A
DsovCF25e9rax5d+irxHoOKbhlJgsqbTiGuh850KgfbXJEC/65zuvrKW0FYIYnIy
j7Ek61hKlvB48W/Y/ErSHMDo7RLkc+Tr/KNZDbCQarGKmdOs9Y37RvCiWJ7rEoms
GyHRtfC/WsSAjKEkuRnyMlfojvAyp+BWQftOwjpw3aOBwP2VV96NxC6ACOFXYTqj
nMNl7UHZU5Vo/2aAb/TlbPtYuVZz11i0nNMgDF1q3aGVX76nGRwc/zFUqWDraF+w
rNfFhEqmz4jHA4PnoiUwnyD9gGi3wfxtM55dW+g5kDpRqtpA2aUaF8rbPcD0BorX
kefakp9/gtVly5l4Rbc81RPQN7ko5g4XKEptlK/Htsld68lM8/gkA6SyNkzwFybG
bM67zn5tB+WuI3HP+a1jOB1yA90FeDQ7xIJrI/0Stg4a25DGSr/TlL9drzaQ2bsQ
D3FZ3+zv08/NgmGYmmSu28Y6uRrI6BM+BTzvoZAhDAr5kzY7GsrCFc/33DzypPxs
t/PZxYZ4c8Or1q6ctQ0+5FJLtc9hro24sJ6cbh/zdwunSjRz/4uOUfBYtT5ut2I9
TJGF80ZMBKghWB8TD/yDpWKKoRa3icKqdsAbT0iu2PUR18a7zYq8+vQwKuU8dqVN
DNLB/GHQXdaMhWlu4EY/obfqlWAqXZtOGs7RUGNg64eUYzYhuQFuTTdIsOV57Cvr
h0rgIdee5dOzB2nZ4dStmUEjMeJ3C4ouojBekXc3FKuU42GzoRAsHLvvKnQby8K2
iGfVldSWanyxGjIhuCfpTZ/B8dnSrSChcsTPvqmg2eg/0T1tOhEsg0FNcBn9PChW
O0xxLm0m7Pj75LlRyPEp93RKNtlsYYUF2A3jhYmFPhJ9L+UAi1o8MQuN1NaCk0Bv
HxYclhvauc61tUhYoWYfV7bVXb+1QW5S+tD0fseSTVgOyyujmA59cRPtxGjhNcEW
f5cjzpe9b1o4qdB+948UX9BbpT5OKLvPLRtRdwo2xXXQzrpWYmwOon+t8lvRUCmP
Hkhk7jPZy+Yn059a5lAy0oBPOQAGPWH8zMjR6loiu3pPscXRBbJh7Dhtfe+dEMsP
gn1juMSE//ZCFlBa8hQjmSxGbMsDNo7GgKqnCIBZqjLEdh8eY2e11WyXATHEo8HI
frFBNQBvNYrMOlItk2C+v/wFzSoaG3qFaYEkTcS/Giid2ONAY2DVCOJRi24vR3P7
k2P50wHNUPzIsua+z3qwjok6IaEt0iUWSSlsTf54lAZxEE/ofJ0OgxaY2S0DRTDK
pUjdfDvLsXnLwR7rXg8trfIJaRuHOwY6jLky+cbtElWyHh6McIZqsoK2y9B0dq6v
f7RfNKc0mx03h29JnlqSOtuU7HsOLc2slxdkFiEKtZwHyXvJjFeVlQnzNgpHELAk
buOiqzSPBNGf9DaMlhdXX3mGM6OZ9fFJdBf6f3EHOcgGogE4zDhgCxzMyK6g7hQc
V7LM6uFfWX6p17G79uaurwIEqmgpHJ7z2XwDCbDsFYfk1lN/uPXY+i2jxGOB1VA0
ls+XjWHfas/sNoOiHZEFEbE05CX+uTw2BxjDsshDNn1YlUmdhhFIwN3ThconiOo0
3l9z1U1n+oJUhCRf6R0iz3/sAxWUfNG2PPheGp9P9ToNN8z3oY7OX4iEyTZ40/Sd
GQTBGLNMRaWmkP+N/NEM9nxuscXjbmZXhvJLYz4yf0q7Y4PgXu7Q74cggN1MAqDi
w+pfLmAnv2OgYfNUTDqGnxZuo9SsgHxlFebR6clwfRsFOuPfV2jqzUIbAQ0KZOjd
DMQHCcmK/n6SuYi/4xZaC17INwSWgsN2JNFB4OaRHNWzKqSvmRSoin7FFcvVJScF
goOf9qtWdhHpk68RNThcg5rgROBe0bbqD4JgheBBr/Q2QqumQ5g0lzxtdrkEdu/t
tUcy9H72GvbHUe4FMkUJ+jzWdvuzqbJPzxZRXbbCq3EuBuNJ4bv0fi2/BwJbfgJe
GxDkOdsWlWcSrWH5DeXXfy+OojQv1041OsYjrSYF90qD4HLZeW083Q0Va0bvgbHU
WyKmhja5kwQ/UHtK3wdbBkZ7ziy7pc5vHxcSuM5w/fcszur18VZxdxDrtbFgoUJw
BtZed46gz75ejGeqvHYQ1xazxjiscl4V7ZMb89ebka1HhdiYJtwv3UG4UNh/nqj2
D8FXR0Nres5xv1zVD5cXpoUUphlaQ3e100t34+soNyLXB3XlH+mQF3hbMBsi337r
9I+uponwboLJbbYVNIlqpxnv6U3NcZRcfmb22cxfVZ4P4gjjMuTJaUQJ12TkoEGQ
1awB9JA4j49WDS7uLPEHHZzmE/ujB3UDXTlY5irpzOm6hJ95MJs0+OVMyFw4EAZb
Y3c9O/Zjn3uL44UOL9lao5BItMR9bX+kuMCbuNSbLGQUuoWCad5ivTErz4BBhN7d
4xTYF7end0KyTLaypPXT6Yd6tINq0bNXomnTvvNpKLHrx+A3LdjORTrJwSvEh8ES
4UhvNCmLHqYimdgZJVZwBa06aY8tjaM90wDIFGxYkpsPh7evtLd0mrjoCwLstMUg
GJBUgC3ndWrOCTlIAaQg3TBcp+8lby6loab4fn9U4GhLD9FYpvt6l2J9BcGzMQSQ
sOQ0S97S/RHhdm6aOBKt7w+yX6zsPsCL9h/hgzDnmzAqenlwn+Mp5oOU0pv1e7gf
reDET8mdh+syg4nkXfvhr9CK9LK3psdNNMYf8PoXyu5MRJWvXDQIvopTkU9+tsNu
yvmLaUunr8yjhWKik9xxO4FETi7Z6Zr4SFUMDYL4n8eyZxR/jKssq7kU0qpfQGMn
XaBoeYTkfI1xx130dxl0ieC7ZWAa0iTVk/YngqyCjqqhred+AZcPfqxZS1GximKr
Ban8G1AgntghvtIV/RG1ij3VSVAPRnnv3Lm/nG1QzcDNYBN5lNw8yr+g67JeL2Ab
vEJG4DzzRrLNaZBk9dfpOKgCmJkzIR5w8d8LWwZfPO/mq+Vb4rjws40EJ8vFiZmf
g5dhkGBySmyWoG70Yg8OevL6cQczQ3teohH/PDz7DZlQKBi0gkHX+Ztx1W4WZXq3
E7wrZzYQhkCKWg0/uauaLTpI1QjnCZ+E1SoSOTX6AAMU5f5z2OE3QO4Q27NSJZdo
3LIL6zMwOSR8N53CirtqD7ibKYQgmsziEgvTiLfnDNP8Zmm/dOcP2hSbaZyqHjK2
O9fEmoqe2IKy6XzCbbZnZbZ2uJ+jDlPtG5vZsLvvU3HuiKE3/SXveBlUih2urv5u
yIwlot+GSBTC10Qe0ZOIv89Q4ilKRYgG/r1zUYvmExD5fs7DVPMcEoLScb9jASl6
lw4eIyuCnYflQnYXjIJ0QLGPsHxBBPuiYG4Rzy42It870d6IUCUhAxu+XhqvktwW
Clh7DXDhf5ZDJTHV7cZd0XWJ0xJoKQU1OyeZk8K+7GXE2IT7ozoReawHqxHcCWpv
O5MOqjs6T43dr8xlEiOkcWRI+xpehp+SycpzH/ZDSwIwS1UZ9YNhjwmoMet4K04a
hEDjQwo9ZcYkBFog/N+17y26D4S/dZBOlw416w7j7RP5h7YD76K2sCSMFKrsxSJo
aoWDhp4H+Vo5YxivLVUYwhxpmuemEp35o7k/AWK2lDwi/tiDt1hTSggCcoHEoiq5
C+XmKQmAutWbO/H/u1lKjnJeUiSh+pC9ix91wlOln0MNvDtmiqG/g8Q8RLRt9MCO
e2WRZQ15OMAibC78Ipl9YXOreCYbr4Rv9fTTV6jWjYpn91gFzhQSawz2Hupz6h99
pPLXfB4YeexKpYcv20hnUaywSWxTGu6RB7yAETvRJoc4AWKeKcs6/ts+mRrv2OXP
aHFSov+h9/M4xLat+sWTcj27U8r4gMF/yH00ERwecQxk8al70a8vh6mMwKz2MbFT
jvxQ8zDTBBfSux/YIQzVErBvHmpzX9tgqrc3u6Q/Gh78x4xW9cqUODfcjEFZm+XA
hym3FApfjl0fB54m7QgQ/Dvlja7Y1LEfhwyKSpeBUeQak12td3AZVECqGajfDenf
eWMgo3YC5VsRCpI5rSW4GgGbjLlH76bXEixY05bORafBhRUHiTkWgwiwSN2fH4Yl
Ot6W8+eHn5SCNBKq9eR5wn1HZ0vQeh7+gwpfevNrpdcUrMLhCKP+618IXnEKAKhY
W75LDjn0+RHALzokgrtbfLsCPtITN0qWuakXkm7kRPiVwJO0GDTALUQrsNGWwHra
iPDdXWeSKguR+xuqI0TUBgBIi2RYuyTApEbHExH9w0ZjnIzZ8Iz+ygNbJr0FtJ0w
KMZwu1phsoMB1S6wEKLEubBfyOkwsxMC4CdOVblh6SJKpQ9AeEYzlg4h2MC2Ahzj
wcf9njms34sgmYySBIl92pS/dhzpcjuIgbYt1YEF+vlHtiY+GZ6liKt4o84yoh27
RD/1rluGF62+SifVCPdwLB9B2APJldc3c1EhroC9BfrZQEx9q46gJqZ/1FRMalwm
bPMDMshiSxYVlMqY7iPA57tn52wz0wiDj1jyEe2PsuLMj7OyPmrfKa4ADzSK8zcl
PmdzAwpor/v1phjqIHxDiPYdMyRl8ZCUu43O0OBDSiPbHlkKg9/rSZ8RUAqA5lmO
RR71x+eLAGDmLrewZT+yJAGFVPhj/luQQzCMWEiBM9oB7cnhj+yrT+FRYqZUnzvX
jaxMk17htswhMs4uftUyoOq7DDcI8K5abxfXXxIirYv/Y5NHII+gZvnEjbMTHrdG
3ml9DoQHlKy8qktKYUbKCOpYLM4YBdsAmbnUdlYhSCr6wfFA1t7XopbSjZrpOtLr
e7rkndTuTFzp1pG1s2ZqD0YYGlgmrXPS/k8I+uWZom5k/oqumBbEw/cJVS+AlnL4
mSCpQcBKOhPTg38DgaT3j0lpMlvSY+xvopbPmeFSF0rxAV0cUns/ggL0+/49rRKd
cu8NuB/wPWWobudMoHJXbdR9QPJtgt/ei3G8sbXRH71raprQDrQ3EK+9FUNTjK7H
RE7n81F7/InDS3blCUAxPi7ofNHGnBIUIFX3twHz0yOjhb73MIODa8MEYrAwIB+c
obCRAofkMa4mR9GmigJH44i2reHn6I0t34CjPIil71Jmz5hiYrYjQe4kqOFkNIII
Ukapzq9Us6CmFsyoSRE9f8Lnc46RDTzacKLtS9d/UcH5gvlgitFuxDCKv+0rVeBm
brxv+yZM8FPFTM4O842O3+sE/E5g30wKGM+Fi9nR+iiQYRhKINuS6ueLrUBqbBh8
pFAHp8Gd7tfQIuTIwBqNYrxOyownVCzhHP0A94WUdPRyEja2KTbkyJh4OcSgJ3dI
u3nL2P9IhqcpcPZay50SuKv83h6HPEewlHmwo2kmSpTUvbtt3lxsKoPH34ysnufo
kDFIJqpncdML2OGMHMacpWefUIUujeNbqfBpMjuL/UTTmUe/a9zEHs1mKDMcEW/0
mHDT0sMsf6/DY0ExVUj/NSfvVSvcnCQLtU7y+hRX2yCgtNvYTxCzEgUuhy3GoSB6
Ce6KsO87CxSpFx+nn3azuSFXLl3gJBWKumpbQqnVh69VsH8IKVgZ+VEmqwqdpCBH
8q6KDaFEvG+OwEO37nNn557INYz8k1rO1ZRJuN3fiPiq2eWyDvmhBlcqX0styBsh
AN2sX3KJNXcMH8uSHDlX/xbOY3C8piatCPl3G4UYdZvHRevJnLJxtd3r4nE+6o07
DoQkLprIX3lOmhdaSGmO4cy5JkN5mlrS9EMacgoW3QUcBEpGFK6ggTzt9GsfJhqm
ldscust1xvy/gbiRZQhBOiHxptXEsJrMkL3e9LRoy8v6Lrnd8nsi2QbrZVDEd5Fp
Yj+DlrOA8OZtG58bkj0gWBObFR1kiymFYjQpwl89FlQ+okOahWkHse+kap0TOC1q
Gdg4EW3Wxqf+at3lBX1LSjEPp3xkcNeIuIwIXx4nLtsGjFBmTMs4w9HiXiYyqFwL
0t6SCvf8p/Ql0MFuj6VK7e3GCzqNTH1JCSiB07ihemOhbzsw43CdgYKZEbGIjq7s
8UWmywYpKGdolttmRdliRpc+IGCRfXd9uKZPtUnzse+KWQW9WNC5co/yInnmfmhC
gCei9VoF5bFl8bocQ3to64hKbxjtXXQNyFIyR6pOhA5Aot7IkcrlOmapY6WQ15+y
vLsmqFesclyaZ1sGWemJ6CPxLgFZhVPAQvU9ZA27IVdYEFaCXItRpToD5hsT2YLR
YbucN2kUh/qeT2FaDZpED/+aVcPhi/47KFFKdt5DSRbM4U3tONYTePKSe6EhfXaR
wXKzPyC3dmeAwaA0hdHEpg+dd2QOtIP72f2vR1fmNl/0gEwCsqAg/xLzCZ35rnpi
kFsJcbe4N2n0HdgixMgfGsE/JO0ESXGyQKIjO+A9FtsAJzi1KrlWZ92qlmFRjkUi
lHYbsDrxnjmn0ADg8YSDgMniZhSBijnJIRtrJPXrk/vhezP7ocDCPlOqe+aqzjV/
+yqF/EnjYW5dhbIWJOWiuCX/Sjiy7MbFKsoTqj9x2cCL7l/dXoosUwWpE5b1WaVD
Xr9kfulr9pZ3f8HASdQEagfCSyWbDr+8Vr2+V8RvzzxsFaVPvnX5J7kSo41i7QWa
cjfRf2zQxMkhcNfjJFgxcA7TrppD0kiRt0sYwIkO/n3zKlC4HKmBdxol5LHvP1n9
iV3QIvur6llTZ/Gb7vyaCLstLga747dBSMpER9A68zagwWuBA2Rfk5IuGSVsqnT/
kM7EnRYHlVPdbx62DsCO7AQjb9525VyOpuvM8a2bvJwrooig9jGOqgyIbLPwVwPa
hLgJR2FmJOWmkEG6R3LWY4bmU7ihBY9whC+2op7+g/d5k9wCCwO9TDbJYhFXo5J7
I+l0rS/Oq5vhqroWst9SSMmTi6Cv49jSunYeq9WvgwztzwMD+KBmHVvVpxVWOWhn
gnAHIMYHbLxvL8eEMK7XIFYHj7C4efxHx52c7FCZYMcQdRVqTzxpRf0rQgR3luS1
hY1Hsn81RsPGr8BZPZLwcud3nTA+4uJtV3ANPuHNihBhuBD3HAtos8CXEABcXBHg
Zf2p8hQ6AFWHp2KrDS/V9bh2Xl+g+eDX+JjmpB8dsz0Jd6jNEt1xHNq4EKTC9xxG
uVlYnYh3AlvZax3LAoOV0tLXyhgMXRY19kA3lMZPFMVc+ocmxJTDsQa/IOeWroEV
7+bngyWVRv7nkwmxmDpCR9znr8lPhMJzPAZS7gIbrSpuPjx7j1bIQmrVF28OR0dC
RYLJ7Rv9rhcn8g4b+LhtfhcYawD75sNKGQw7OwcHXgCY4YuSHSQR/uZKssbGsjOB
JYe56xlhd+xbMxpOu0sl4jhQJBAURTZmgqgXYFCQS4fie9HHdqFUCu/E+FRUvwYg
f8CoEwnp+WASLhiUoddcNJDYaLOsniDFQzKHPHE3fqaCgW8z7YNw/WanR0hvVp3e
L8+JXnflQo3wgcnBCTpyQYh16UP8Xn62ol7nwxdkJuHulllDy1JSM84n1YN/8wY5
RlgotovjElo5NRVD2tENJdg7rOWsQ1P7cBroje8K0XOI7oUZ7/n+aHxU8Awo92lO
4/PcUKWtPev/ZEMpzlTe8yvu7KOcXOiRVaHwCZa7uhAc32g2+LoJiHjWW8JsT5yY
AlJjavzZxgMYhr22hfyLmzNnXIVur/94SxXEbv9uD6NaKvHGwcHD7+q0Dtro/zyZ
1gjT/DHM9CaRdL9683EK3rah3PjftGf037hIa4bhXkaJnYOQ1h1q2pk1tURRV/MR
ccMy7g9q1X44g2UEXh0UApaUVN1I39PL7QNVGJ8fZyUdgnJru2qkaB2wVg6yQk6w
XgQgfB0jiTsJ4KQFyexcv6bpuOYi2mFYOVb1BIF8HdALnDdeMSF8P8lqr5TE3jgx
KG1LxRmrgyADkxc0siAoihZdUR4DOa5frc0+tN3Qc5youPF8P5UYrpaIXp5ZFDIQ
h8z5ipFHctJnaGc5+DoVtPLN31BWxxWFPwLfWHDOo70VRasPWZ0D0YeRYQXabaxm
PvE8qlSoErCY0U9XmIjznbAmGajf5sUS3r8PZrFVKftnvvxQKp6mAWY3llz/DFMA
Lt2tZ0l5jeX2agWubQjdd3jE/3F7wrGICvf1akEAtLheSEDPlvsmI6K9fAUPQnmc
JCfGU9CvmfMmCHeg7LJtv/h3S5+M9h2HfMS0rQSjgDi9bz11tkK2hyaa1/JpZA47
e0uTPa/ZqCkKMa9ilMKdALqixMgmQZxW5Wkl6Jt/4vybOhXG//Z2GBTF2/2KvJHH
zos+nudobtCCJyCwbHYt62QLB+wvKVaKegq34A16mH/S63NGRPj70o7oO/j5HQKr
RIjJiiPYeU/5T/LNktLi4DOrL4EZHLsDhzEdjQ2BJXTF8eVjri3Zqdcx0qVugRBf
GqbuoQP03yE9YT6xbJAn74I6nrhNBeETSdfII2G2EWdd0FRPa8OirdoAmr9/25yd
MjNOdvU2l8WyaZUT5pdAFZ+DmVXdZjvgUzwCwxDqnvSAt7iBHyGxljikmX1FbxOr
5/fcGNciE0r8wl+vLqm4/Jdd8vOX8qX9QFf8eenoQ/D9CkBqDQnaXJMCiNwRtco1
4gjBVr0Is7Oq0gHGE+SMXk3ELVpb25fVvAC5h16ruUS4rs2Valbuly8a/HTSX8fP
JQIYGY8XOFYhD8FVdVPTkWI4z+tU8N+YVgVEaHnAj6yeKoqu1ldglvBLycPM5DXX
/1+1WZRlhu8TYHHcnEnVfh65O19iq8Vn/MQgjfv6odoIdhF+LI6KoeNs/xNGs7gt
63gkzZ6+fDh7qN89IviMKWgpRJ1IQXVkM88iSVOpiqjQBvRe0NRVO5yLisFY8Aa+
L7nzhJ7j6dAhgMtiBb58nc0vggMzd/XCSHxGQR4Qo6vBBuHBaTJtiZBJ8GI3furD
NUY33eBY+fmssAKwBU31kMO4rL6ST/w5xSvD0PsL+OI6f1rYnOduGDQaF9GKwHmv
TpSoopC0WzrcyzP3UCFuZcH8aPBsDEbe/u6aKppAN+hpEkPaZzXxuj/q68bXrB+j
FCankm1WCXmOmYYqO+dNJz/1nC+B4JGgqtXVAJqEJC8KpAhPZfYd7TGVdLd6A96m
ItMforEo09xCNirHHm/yzvO+IkrWI9wVOBSG+VcqjT+Dn+f987vdoqe5qiJtFuBJ
3mgLR39pPOEY/+W9s8mXyVzZPPot4dXBjisl++HHibYA0EeWGPyfXeT0BbJs6bWy
QT9lLLBnw9PIITpnThyUe2ykeJyf3wfUoQgzHcM3KRBe0n5DNRS+LW5h1uxi8m4T
3PntfG2fJXG7y8qKa/3J0G+EQnUcloOZmTPMfcPlnn9SXthNLgjmWuVGkp6ulpG6
vNR1cr0LlkFMZVfG8cJtcITM/D8f//h95LrkQnWWgB7/nZLLubiwYHRjPrDjRUq4
/gHLtSE6W1VJZCypC/Ir8NThgHI4jSWBMtBCdo/qtoYd7CtqUpTwjNFcYy5aMx/j
Qd4rwjFRInlbm4nRa2eloAlewaNPE60V5uRXGWbIn3XfwD+ibcDHvkW8IfZM29qC
/EFcmq+bHmvF/UzPJuJrP2VuysIvfKm30cm+g+dxo7YFuWRRFuQaUTrsAAJT/rMO
UA7pRtBuXFMll61zuZabZtdXHiC9FNM+1LCE/YbNXSXz09bysGuPjFsrA0TDRHyh
BFnRvCw2D2ckeA8M3Y8hm8jyFpLBp9Dt9zeglaXL1EP8AmTNhHQqrDm/DzRo9rdL
xDzJc4V0DOH8/djKYrqh50caROSECma+TKYjv/UkX1k/+UyEBjeYhdxTLqWVAHKf
PBNYADezz8xITcORGEU/6qoHa2Mjnk/lXGZpnG2+RHaRV+7ApEu2ZxAstk2WSZY5
ybCdpHb8d4KDESgysrNFmnt5xCdjoHyPqx4yUTRV8AisnyXI7WaEwFukjiw247P+
q+amGonBUW1e5ZvgXMKH3aJbPnaHRBtfhI/voLWKuUQWRcukaO+e4r8Hn+/MKieG
bauARaKwpMOyC+NZv6hSYT5+aTZGBJp8xQFuB66RQHTdfICkBpmEFr+R7P7tcz9E
mhpm+p4qpT6Sn7lqU5IW61O0OG/0BB8sAA+pQUNID+K0O0mQlEr3T6S76B+ctO0e
q6mwgLd6FGsbcFwqwj+dCfgBectOhIgAzF/2OV51nx6ADA51oea/vPFz4rMVZ6g3
x50KHKAUFpYYmUJUhgG7zI21x9RRdaGqHAucfA75aIK4PKjk6jCo42iQvjGllfuJ
Oc04ZxcGvZtTckYdo/btet08VlGMmd/QuKOVDGuvqjSaFyQnCqhAWkWthZvz+b3H
2VlUZijfcPTDbsKSvqjk7G+YYBekR48WSEHoyrRPH4UcMPsHWuQvnDzhKMjxZgWo
rrrbxm2f6Q5PviuaM377Y0spp4K4QdI2se9wFry/61jDXh2AJnvsk7Wz1YqnzMdp
TM1pASR17Z3l1esma5VG71ewCBdoTMz72+Cm7dSzs5rusAa9v4Z0XKPa9N9V5qm0
AdwHIlRYGaJ4EXWwBHeAiOu0Mw4kXJhJtzrV2LT7w0r8qy0V1T+M4Lotf96z9oOy
/2tVGEGefr1QHYQ9NPDLCSK+jzYWTq/JJEnVseon/xWhdg0EMekdrgYteTkLiXdv
XmrVluWu7+Iu0LnlQ3HjYbR8eMQea6YNudLqQ4WrYxs8Fu00gBV1XYINVqug+bS5
64TM0w2zxt9LirxU4aKhg2vyrVi4JSYsvGHSg7NPG3E11OuHpFu6EJYGYfZuYpcu
Jhn4IhE5IHbLFdcXwVtxIP2PSyuc7ImdO4ojHHG4l2tPlPvWWq1MPnY5bbLzky3U
aIkWmwuEHrQcCB3Ut2PiUXTdmIKT6XPTrn6a2L6Jl5y6YDQ6tE9xXs37SRqoPy77
zwq02y/QPYjbG0DT2DHr9AkF4Jxwjt5qRQtnq/vYjk6vO+1kg1j+cCOHt3aJHX0u
h4Swjj8LgfNaJoP6cWta8DG/f/JgAZqsByx4kvYip4PXSzaGtLtEMeTkvYHcgemo
Be34Rbm4XY4Ytm7AstxZPTRDFIXvQ8IzhsmY7+lplsVREHyTqs2k5B4oEXDs0L2B
uiDOhd1jvgHvK3aexv4RZN7/7pui2Pws7UmzeQJRA7RLePQXNjgD8oZk/slIxM23
j4iTQn6luxHIiH9QnM5v/nvcqtYe4JtATscHwdNWrJytU0wrSAyxnqjHEZPf2iYm
EnJQ5jE/AQZ3H7tbpu/0PSN7fWLoSEqfC6cPJCdUdndTjSZR+2qMtuGNr8AADS8u
Ze6uSfoxDIbODiKOGhz3idPW+ccABDdTmDkUbKM+AQfn6orenk7gnGHCgU+Q9SqM
d6oBdCGb5MhIz6X7p0zuxt99INmONfIfufdkB0G/XoeYV8pR6ktSqb1Wkma/UjmR
kwWAD2sxWYB9/+7rNy47EQrrOFeipIcJAPH+880ifFy+EvjFnmFOfo1D4q/3s9+n
JrmX7Zb3NbKaEWqIjMSFEp4ISujg1oemwo/xMt9nz0EBDJzf4+sK6H3TxVibM4S0
Q+zMD3ohPWtI0yUEsRjOgAFD5/D9BQNX1BU/nkmWEOSySKcuQ/VYTwaUzlEg6BNR
qfKviPSirukX0oIiBU8FwIZwt1jzaiR2T8f8kPztWKhM/57skDap4Fon6wSHFtD7
8DPZWg29kl3PCHTbnjE+kE0ETpaDNijPrOIaWa6888S62rjWtz8GI8AMkS6EZ9gO
6S+aCgv07+5lzrGEv4eBWcwVOrZJ0YQINXKcdnlwZtRFWnf4dGAKs50Cs7kyQoPq
fuf8Pm9rO/s1GwpuLKPjyXFze8ekhR85sCYp70I+p6dUM6EVZlrq8TJ4F4upm5nN
MA1q2NYRHyE20XjDLcm7shfjAweu6Pjn+mMhIQg6ItHEOyaIvCSdlfQoVbAM+zHt
9PLS24+UePVfanOOhOtLCBlQgD1InxZI0qaWJCooS9PT7cmbWHuckMR80HhTxlQE
+627T1yTW6Orx/x5ekjpj5EAF8flAB2FjJYCEnOUxnP7ompEKn+tn7QzE7p2wLfJ
pdbY3yPz0GA5q5LG/Vuu4us2Mbhi6RzHyNmMQ2AwgGHEeMoc1I7wwxeyoRyQZxIz
nVf99D7x9DMBDQfrat2jINfgH1YFUU43uyuhEGGQZo6W40dNmAH6SP1o1xQKTXFj
rTQ9XsbawrMmRpMAdyl4CZj7CSM0G5S1wB+0coe38ydyF7Oc/5R937Z41g+tclMW
Mc/gQKuesf7p+ZEvS9k5jqM9cfvEP7V6pz2nddB97AkHBUmqszBPITnbtYzN9r9o
YyVX2NXAsAPP6o5UsGObFViiHAiKRCgTyqjrs8V5DRS5bRQn6AUTI04+QNCNafYU
B+C9LtDBu6BFuJF42mgstBtpzhPLxmbxSXMOz6RriNNC0SPUIFvom0JcjgP/DeMF
dqwt5qdSZIbE3lrDia64J7FVZaT1plnSbabsv5e+g/bBEgUrwLMDFEHrZbEQFvri
EcVVdZQQtglnwk1DPKMBV7gQ82APF5Y/SVJfFQXHK1SZq9/+CaogYgqJ1SyuUwod
jC4XSOQsQ8MJHydOgG0HEUgJ6ixYJRZ+ReirL2JXPmVLY3jggsC6bX0v5k762cHj
r+5T2gRy4joVmwxY1/f0Y5fkkfQi9xIgbtjIrNUi5vrzRiaCI1ZjHv8MrtMaOvGL
2d5LLNIDL3z/VK8KPsZlKubHs0gp7l9pWh7B15B15C45ECc6HOd4nANvhMM+bWfF
fNv5hZaDGDGrl0CIPvFIzPt5rDYjau9qp0cWFYPZADC6zgOM6HoPhmrs5L1LyDUK
tokZ/VR1fGsexli7Vwtx6+LEC3Sr7G3kOpLaBJI5pX/9nQV5hSq/QGnvbw8oOq3b
HCyoMdb7gl6pv6v//j8+D6EnY4XOD+aJ6R2oLWm99d2M6ECZGm0SEMRY7VrEu55d
4vXod1rD+huq4HlsJFdNhK9kQ7Tfo5aqIZFsB8JHxeg6/0aNhWTkwBOGD36mBmgK
5U9IIl/xvXx+2tf2fAvgcQ9gvt+aFJPtzsAl7DmFriwQ1qw9seS4UY/cx8yWzJRb
8WWIE5hEFbeUwhtzjRrKFC03ik/m4UBOLjcuP4BGXUKye7eNlZ4LrtUQsdBxthlV
V1Zofazg+JCSDxIa7P2IlJYLf9ikkWHvyyhM6nd4OAzdzS1a8kokCzkvhliM1N7V
zIkH+qrmv5wThPLwjJ0r1GB/Oy5sYiMU7cCCHe1FVIUYOGm3yKtR54uyxwWu3LJs
nTYAQRx+q190WwAilnbc+Hm0YY412MofHT3zsX43mBzISeBRQASdu2iYM/YBbhRi
5nBqOwwYe3jNQ61MAz+dz2AzAiIpchKOL9BtEE/AbkotwE/JO3Rip6lxYbtIu2yp
bTmp/VKJCLPoIy3Ock5r3FIbfOBfWTTL5ahc9Ia0wE6uK9wLAne6p+2IflLL1xYr
fXClRLOPFxNQvJ81WasbLy+G1dEKJkxEZFO9Q4FqZCEai3zpJK4DUzpWVpEsiLCI
Uu8aosJvcIjUwzUXEHrOvGDSH9qlZ8l0WbFboK+neZx/yGb5Ffs7oOwqkqtTbQWX
agt2TEc1TRZepl0OB2y9n5LQk4IHb+W1yVxpCFp4SVSItOlfwhOaYPLZrU+z4AzW
1BTGDFU7u7eRdJxnkLiIQnHrdfB9WXW7Z4TCsSEfOnQsntAeYdiq+2387u95LWJk
Qz+hJGxMCWaHtkBhCWsaYmRsvyazkz+RABGrqh9dEChmhvR39FBehekAxrkyg8gf
J22UHotpO3qYt+O4ac/IDzDrQzHCdAmURzeLWcG4YQrG6d/BBwgdK6oSJJRss8tE
B0mtdc1tDb8MyvgPw3mA6OcKUuCCweOm01v6xj9gQ/n4jijpWA6iFm/1XdhaCqt8
hv2mbvsnK8bgjMe6LnmawPvm4bBMJ0Biho/h7/7GWC+/cY4UNVCVkAy5EQ7S09R/
DIM5fCgvFi+B80CdN6oH1zrILsCHBPiTXGP0HdR/hzEAW4O9X4iJSJ0RNFrvKWZ0
K8RH0gEYI8KCQkiCpcRZ4qtOjqF/xb1eMztg8eENSGJgVXtrWRD0kGZqk1hYPdfK
ORD+VOidrNRxaFqnjS+RuLKNbDn6soWx3Nr/bxU7ztxWUH05JV9EzxawwsxswV24
GZfe/+QS8XanjpE6G09PkuitEn4ysdKt3z8IeJAvtESitcxDX55cF9W/ey+htxTp
PE/wMYJ3sNsNHOCQ2YJwFs2+5RtYXXNRM4lCPpHymdJF8kmPd7Pdg5uFx6y8X3IH
CokQZcE2EAhfkzqW+qENRtWWcz7b5018w2vMTsRLwS5B0VkiEnrfFzwFsqgl/rfr
gKhtWyE9dJnjkmr0y8J8kTdKNywMHwsMcEnpej7E0wjOQqtGw/4psY/bJ+K56LkI
dETmrYTV92qCqgoS+2jGt4jgsMLzOsFcuT7RGtml6/Puh+A/gctY5YcpEeP54oH6
O5wCf7Y2Diqlb+q35EfijS363BCoZbC8nKR5LhFUUD3Zt2J8Znk0LVC0ikaY65ZC
Gd/5IQabPWiN229mtEPcJ5h8UCujEPqwHyvMKFWiF5VortN0bFLVJm72cTBdPtaH
Ut6NG/cCnE93ej7uy/IPWefYmr0f2hMDZADIJmbMnUpsVZ0RNzFTWpSy13cOOyX5
sAK/yA5x0NOqpTG0uvK0VHzbMqzGGgxJzlONS6DcII2SE130GQL41B+zFyleUnqe
9Xl7yhOSI5EdmSWDsV0Z87RSw5hCk2BtxxmkBl4rvtJTJgxQzWEhAgf8Md5etcWG
Osm46Dt0NhFAGv7TpwIG96LtO70ei1gr5uq1iV47EUmqNerBeshUh/EcMbtYhQnt
brRiPtd6A3nMOnkpXwq2Y0YDeyAUV9JX6xssI9lmnNr1uwMmz+rQOxz++K5GiKf9
1K6RJgGmHEOgg9d5QynZbywte7MgnfJiqBXVRalNOTkehhDvUz3oGIuPMwZWJGwz
xxL82cuUiWppyIiagpO9fNpjmhII6m6oErcCx6wxJlg3WxoJhyXeIW8fEBCs0ynk
SUN5/gXBKjFWMfgC++XaUc4KWNsN8HkzLs5x0jn8wjm/iRs6kT113nEpuaTjQRkS
qffgpoTc0dv6h69EkqAAfAgVg4aAJUVS66LAOQ20fgPXwxHLGEMo0F+/7mZYN77O
l4pfDyxW2feiXZFRpFbv2WLHyT7dSLFZf6ETXkvcb4olMSk0R9L3o/42/O8I7An/
np17IUsdlO0DFtHOUBh3Ywfjbe8iEOyPSPcQv4JQlVt/A6yjI9jMMPNGlKGTBvPQ
nDIH9PNFmCutXsFRz/ulATgrx9j5MSxj6T59LPfdpr2vluX/F5nPiEIa+fbBEl7C
eQmrEaQUAkcYNXiU4eMiZvdlsDYMSSYJMLCoXfa/O/FTzIJlpK+W8uJHXy24mccA
PNc4HaMMKstWxeo2n2x/zcXLQHN4MZWmTQ8O5aixP08aOmmH1eQinZD4YquKJM74
dQ2k66dLi4/zMXNQ4b1bbHzUilGoW+qbNc4rFemRMBmUHCssxUhgnsopcJcSUbUX
lQF90edKBMnkmY7sCXr3mnZl4iBeZgDRd9otIZC9s1bvkaXfwsATokW8yvMCH5tN
B6yKR9zwWW9lY2D/u5A5j5SPUFA5viAutYw2Rh5X5re0G1PUvv+yKiPFJJRs+U/A
uViG4fCWApwOnSQFgLs0hFKmmbDYTORV/aN1wyeI4PqdMvElT2AnGlp9B0s8wSIR
3OgRYiMsjF7HB9JbRDI6okN1FMdF/CR/nkk450QW5V+ccATonzd6iRfHmaE+UWvg
Y3W7SNKNaavt+Kx5rs+Tf2YnMovqeRxhGnqSRgOiieEZqM9f65LhfWn2JqQGMKq2
uRp+pz3xV+IQ8OS3DUauK1aS+ToRZJoI/oNdWuqe5kSy1ZoD30cMHJcnMcFUMliv
3ve1bcxyYUpYiogAIHWWEwQH3L6N/pszmjvEt44LEM4CR2lcwNSk29L/zIvS/IE4
pbCaCStOSQ80s2lqK+KQ+Sf3ZqKDXC3+SzDftarVHng9thipm0yDXedciyQCnWaa
eHbjBWLeCqX8FVKqUbz0VlkzBNSepqfwZvQnWWcMEIZlkAUFAnhgHEimMUw/wM0b
iizHATr8BmZfXh3tkbx8nMaCAGnMLLdjCA399FeFluVJOhz1zx0ShFH1JCskzVVL
Uxd1dXo/9T4HUQvjmMTKyto4brGsFtI/l9rHu7OrqMs29enMQSroDVYszGc+wFdC
JkP805oY7fbqpn2JNo0hLpCQ5lwBM50dCqUmjZsQtmv2PM/uNrBMi2X1zfwAzMNb
Z/m/j1CZZ1EbxUMI8pg9N6ItxKaFdoB+xu7CHwDueLmNs4CGf49K+GOBSm0JFIVC
QkD7z3fYT/NWyKyY3QHdO18JKbfx9N5T1h5x0bQq3elaE5Zk3iNGBgbyA2KzEwIf
NesFNCkZUaEwZl3Q/K5flipcERpbJ0AtFyVQDAgRciYvT8jiuiodlvP6gi0mveX6
TOqNF2rlu6rIuI9t51LABSZegdzivXsc/995/HS209V8T2nKrF8RpZgtfTSqhNQV
BMYsNaAp/TgaIMdEHKpMKC+5kjlTn5mhdjLqzRPMiCaXt2wSctKhuyk+1c0p9RU/
GdVx8aH5zJ+hTA0BgteQwKSO0ZY2f6IsHtsTr9O7OXzl7Rgcm1Z6BD+RbMzmTz8V
6Op8X4jYpTnOU7EksRobKxlLN3SUxcvZ9RBVITJBSfnhUnn6FnCLBdKBXNqfDrb2
8SNn664Hh8NsNxUXT5YjsXhKadNarGof9rMbWFZnL+aons46zt9mG1Ru8g5wWpiR
0JUfjFJXLkfydIAeR7BSmyR5DEAUYqn1yw+2e8s8M9SAmgO8MlzOLux+n0jPLdU4
QBHmjnbn0OtS7HS1waK5UdXSMmANVX4+8ew0eO9og4fF6WL2UrDYGJvwulrprP1T
kH2M9In43V3zflDcwdryQDTIfSe54bGPGKUy6Ocm3MkqKTbTN6JHKtTS0/JJUgTW
6cWwIwSBUO0Q4us6Tn7wfa50BdYPbNGyn/NdlkRLNs0JIndHfeYwVBxClHt4mOh3
tz5VU6i0BWCiwI2YeNtLoy0Og0nOERAxUvZveqKf/3FEBIYnqofiE9V3E+mvaaHK
QtbPLIR3ssMorpjuDIoEpxwr59G9tQa0OND95lTqaQeOjBf7wBwLahQ0obQVYshO
4rAqhtO4QT1cDQqsxrkIzucQY7nV4xjKyn9R+6bU2uSwf7BIkLVE7Pjkrm3xYFn9
DPU4+NHKEQCA3M3NMm+/VW+nHPyKI8HilRtU9AQNWNrgAaws0hp1c8LpQzdZg3jw
CIFOGX+OBSP/nONOTnIkhwIneSleyJ2PAeF9mP48CNt4Z3YEDkJplL9CKizTqnOV
vp6Ifje1LLwzvdgKF4K11W8pa2AZHyJTziScCzthFqGBma2jekgQGpI+3lnVcWO4
jiU6YGv4m+oxrMgD21JoMtFT1yIdpy0UZa5V8fbRVDtJrQoPvqYD1fSJoS5EBKmR
SaBXSXbSmjNBMu+aWquQsTVEcFcVCLjyy4ULr5+tea9RKRnwcwfJMXLlxZXnhqgJ
wh4j1iOpYjA/7Sth6yhTVVqTJxi78jF7HqbIpK72Ys9M3KpjvcfNgiCUp1OxG4RJ
FIbg3XjA84Rfr9ca9BeuA5i5vYBrdqM1NpRtG5hf9tauVckwuwpaGdUn0MPcBqQU
L6K2TzpJ/CDifxxJ9q2lOwGotaKbOIv2m9AIi+e0kho=
//pragma protect end_data_block
//pragma protect digest_block
odSE4KgVnNsnI0t5lpBKL2kwg9s=
//pragma protect end_digest_block
//pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
WeCw7UOnsVKGzKXormC9/TkJv2I7pKhNLYJkvo7Y5oKBtyVFFq6YjDC7V9X8eBKJ
iHtOpBdchzZdYFojAAcAOa7zdpHbb0hK1Q4PxFIDcGtgnbEtQP+sCaL3RvzWCYyY
/UOaz2+35DN2BylESyT6Le1glquAQ2C/DiMOoTlpQI0=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 8736 )
`pragma protect data_block
praIzJ+NA0GfqVN+AHROVCmQpOgE4oxZZIZIsV7ldXPh1tuAtgWLPEBwTQq2bsoT
m1kA9JXQhebAIbW0AbJlQ7Z9177dD6B9RLTY94x3udZ3w1d/2/as0kg81oNlvQiv
mX5FoIwYlJy2iGwvjyggLyjZg7JXynThnBifsWri/lb532sQJxD4s6oMTMWAjHnL
X3WugizXRar+nW9/gSNiiFmlKDuZA2Wi9eiawUqbOdx0MbnqEUohmglT36vmW7og
tmnDABMQlWhrRI+Wch+S2rknJlA1dnQWX8zyxx56x1ohO88Iv2AsOKBPM9O61xWW
FXnOTxKKlI48IY8fJnNuxnQvR5c3+yUDh/DE5XRpcaWmS+UQXdJ4i7pY5V+R3ONI
1nUOXe6SkTBkrk4F4vQ8sTAKphuoUSp4nFuyGQs5YRuTkkGvqZKXpe6pJ5OBSRk9
f5N96u5RDAiBCuwHw4QsScSS4QMWFKkncs0z2gbeJPHRVwlX0BhL99WeypfGaeu0
1/AZNkjrvxN9Q0E6nU5s+3mnaXxQr+spMsC663gjcNCB+rl4QzpKXN1nQKfN6twk
H/aDvQBAXUZQHO3SVUvxAClGAJu8k/WT0DW/PCQxnevXEoJUoC7b+AN5VWYuMDIt
L7TUokpJ22U1QCyhlOxG41WP7n20PUxilZF4n/5arJxgcb19eEC2oW4nzHnGwOk7
X3SdAvD4ZwY7vqUfqevuxTtpwoWWRZsOCqoLAL5fLfVXMNe09GYwINBWZhXQ48ib
rShesmkAuYava4CBbgigpXGHYd3Ra2PeOGUfZZPEPgp6IGVMrYXzAZfSEOi0ZSPd
xVVmznK4Bx/pygq4wgotCCAjPlUdItgicDG6c7PBf8s3WqOmWQkNxBjwx/2jyROn
UzcxqIMq1z0+6n8NRiCK1za1Ot+3x01wdW4TdU6v9NX3+xRd8Ifh9EEHsFmDldhu
4J2Os1ADjH0CmMQqKk+qnvLaHXh0KNmRWZLcBkEFZESrsPnJ4HpnsQv6Qs+cu+jL
swix5p94jCNa5kjeVPivcrzJTOwC26pfARkA9i9+5UX5758NyvFjKTv3K63PoOEO
Bp6TaTHVURx6OelDpjKRDl7GwpZISglu5JediVeYOC4Dmjrc4XCoubcVNPKpnZuY
Vi0qfyP5GR4ANHM7jbFAMD+pVUevHc3D677x5wCuA2FkVLOdObnji7+OrOMp2oR/
twicGwjbwOskvbqWxGixVz/3C0WoK8SPZocVXSxvHmPN7l2J8Xh+jadkQMDtZvCz
QBJYSGsJOj4hpsajDLQ3JpiXQr2HvdOazplvgorCO5C4dcGMWmyZqO4O/VQ977MY
/5lYT4R4P3oRF/mQysUdLq5MHB2irzok/nFKZlKExzExTVXWybrneKeEzngVjPtE
/EszAMBA4rBTK+lGnEFPg4x1xb4VgzDEP2dYxyOwM9A7ttmA96o0628XS/494t6q
0CbFd193cB7LvA15Nx+NHvkZRHJCmQp274WB1rifXPtW4Isa1EfekMVHoR+ovLn6
z3qGJQ+wOqktrZz81nY0l08FtA2uVdsCx3pYQkyljsb0ef9r2sWXfONUDjYHcWXd
I0gENyxCKddhdF/M549Rygp6W85n/mv97QHmBkBFDUXKnAwpj/sLNZdr0YaTpfOc
ZJEqYrH4BHy5+rY9pUrQkOTPlF7WQIVq5iuebBGAQi7IitzDwHEfqaHyPIyaf3LR
uQmDkww6mCvlQTkE96+mqBJBZhmmUReqE4GOeFRYrOKR2dsCxG/hrCNQKpyqACAZ
SW/XUVCiVLQrDmxuWgfoqxVnZv25lc3JXn1AnMxnwqVdtNvcEN7guej1FB6+jX0x
UCwlYbZncBLi6vLqB4nBmr2cFO1abcCXkhBzfd2pZ3rsWyJ/KMP3SHsXjwLWtodN
eQkfsPLx18cxPbCge3uiFHr5vFsLbBsSCHCcCnsivgwQHtlFGKbYtVUOfGUW3vpY
KLpdLYZ2pD0x9xPFteWHv/+f7+IM2ZBcuFp7eeU0MB8Y3iaGCYzC6mp1asfTbLjU
5tTz00j5lzUsZNh5W/J9nKAk9GyiLI+Y67YDAllxFVwQa8/ljHJ5pOb9Zxkd5nyc
2fGOBlKWubMKV7T/ayuVJfXko1m/MhR1iczY63jku5jJAmigNqAuSDRQ2RICJhFZ
KoHhtRvvIW7EkZmE7NtgnM8GGJZ1LoQxtqEUydDGDEdzi8GiaJ1fEqgJ9IwUDTdC
Fod+sAtIljYtF9rGyDxhwTmRGVdqxVh0rdl9wvyLyrbLwrk56cAVuL5m0OVSY0sZ
hIpmqJN6d1YL1a5uZYzDmkEXiDrZQRs7BZzwlGG1kAyfabxpUWIBiaUkIxeRgrSJ
eVtRrMIPGrNOLPNYDpCb4+9K5OtMxZWHbmpVm5ey0jpEzI0D8rJmdJcFNmJAbmB2
YSzLPAmIpvayoFD1b+KwhLssyiT5Gd6v3lVBHg0puew+TCElZdlAPkg2iu4CCjLC
LELSH/2dGC7mIHcPkuXwilqfCRDnuTcg6nj/G9KQ8WnMomjm/1MgfyfT2qlT0Yuo
DvVWGaS9Q0Nq8dvGg/vZx4ZIViWslHsD7ADQY07QbOgdRIUJ99Z0ArGq0CuYSMXO
Nh9Q5um+QWmXfUwVvnMbTFqnGvAOprp2pgm4lg6hXaF6/4W+T+DOOL/Y3BcM94zg
LdWo++fkKdPZ29gua6arr9d2z80wX5ZKq9m76UyRMhJkMbNj+6C24Hjrb8P/rjcg
+ZiQ5wWk0Qm/kgSmxqQbcNxkts3eKXT9i6P9I4XfY9MsUukWxyK2pxU7jhzhYDE8
s6X4gYcakRBkJZBv0DvlWLgG+qTf8kFsPXNOmT7M+0967WdVkxvVUmWy2Lu7qTJe
JWr6u8U8wUuS59cxGy2b8tQr/lpnVr7WQ3PffW97y8EMPJrE3+WLs8MzJ9qal00c
PbqEZnZXr47tLiPpboxtVdCiVz9X9LCp2AvzesUxddug4I5HmDOkbSx8+ZZiucaz
2I4Nn43U6Bfrtbwh4pjy7fMv6UVrBDeH8LOjkN3UGgW8k27K5ASkwT9IiHV9yXh4
H4nbTGYoJTPMxXMgoB37RbFgzEnqz5aa9BrgA4o0FA25u7jH11MfItlj3o9Sa91U
eyRpWce4DWN/rplEC88yTUW76iKQrh39eZzQjeu9CPrAo8mrgKnIR36pHUp9yPp/
eGnFq/5hKOacgMa6Tr/bsT0wTgrG4Y6owB0BhLwp94g0Dec1ofeCjXZUC9lNn4nl
Hp6aRyOhmnMySEjXJJfggGkNzU+Gi38aa2M/XIdFGfZwY1ktQY3oUgk8Z74mYj1o
z0e00V9YXsyX+nd/UrqwRW5j8QHrXxwyxN6FH3nzsIYp5qHQCcbgn/FQWg0j/XIY
1cvASNwgIjOZVFSgo5ZZsUco00emfnCW52uwa6gE59yxK2H7dxtCnmscvUvjEv+X
5/gI4ThRX4IuN9Ap5icSaJ8eISmmYfkMk2g2t2+Dxe8b7pC6Wv+9P+H4UX5sP0i1
Mz7b2mfazRmMNQFdRPIwl92CumwlvvG4HW+h3/adeNbArG4qtSXem36qJ30f43MX
QVyjiNTSo2rcmOoJUwPKzvpe7r+9bZIRqZ+Nxtr3bliAIJoeVZwXWTAARp0oVt74
LOC4KyMciwSTkp/HbQIOCO7ILn2am51Msm79N4mUJnTjhdjAJtyggFQVMzhjhQqA
5Er19mvzu0nXZClu80/mafgHlVoQ4eqo2Mf/RuTRXURVeEeAi0DS9UjbRWrXQ13G
oi+N/GoPS7oyLdSpwlmXBTRXYpwiht1wIWr0liHuSZpwPq6QUDaj0iMPtVpEIKhd
I+ic50P4gRh2JjZG3PE1XQe53NTFzhcKJOSCe1+p984p7qMIDTdB9cDuFQM+1sH/
69aP7Aj/dz31S11vgXdaLzZ1mwLYeRyYBzvxvUTCe38mxax4JmaIik4a0/EThatN
ZqQc1dTuBnYVNEbUh/dWyc2slRza3aRu/FU8sMuRCoZWuR7BjTVPfmuZjV5C4MEZ
ctCVdZTCly9lx9rid0+kI76DkvjSWgGdhu8z4Y3WjkFj2II8+Q7XyEWs3YM7q0yu
/dNYS1r1fDTxyxj1O6aGZT08ltCtzCIzOTtVEfMPVqy/ZV6SukOK3gZvDHUl2fV3
QpLQA7O6LTd4eDtmLhv3+Zl9FhoAxVnd4iD6hR95jV0j8WpGyWdGtP1gOWQSSd1Y
iloq3CLHL0L2Dvbf7K72C4C7gZcJE06vcExrlt74JzS+AZC27KlVkU2pKPUd8MTW
c5i4oe+2+/3NFoES6jaMkm1nJOhjdTW1VVCdEd5pEvryqLqWTpdB+rGsS7zyoPsu
pgEEKUCtK95XPniakKEHXtxdEKddJSrsF5p2AYFcs9udibIf3h0kybDubefp700g
JegGX0KRrW975wlyPu9JlBcTC2DCJDMlLuY0Qae3ObLJVJ9wzTZSiIadQDSiDswB
XXAyReXipkCZBqXomIs7m/90yp2XEJ2mjSw2NqtSy5GAgKKHS29q9xjDSV6qStXB
r1XosgDuxSFHQ3wESomNig5OJZ+DBvmPEhiqJb6OPPy0+wGcNcdsX47F2oXvPZa8
GKV97W7F4zaB8Nj2aULBKjtBx3Nb7eG2Yd0exPOJFn6ErraaKtn+e2XyQms8B1Kt
Fx1O8QrE/7rPAHE92VUPR2g5h5+MwvC/hgxzTj8IbtgUihq1+abVFL0nfO5ZBAc+
nfwD/7Sx4rISzjEUUc+bJw4fC+UDRcvtbe1uvnmarhgLsQXNvFfHZtD/5hMnDCRU
3jRdCCJzktZyFDDNm/aq3rYKNDBAgiFNefHsh8NlA99sCwSvlzA8Gej/My8FgOJv
9MQIdsfqrvEVu+vhervsHDYwMwE2YdNM45QKtPuLyrxrGS3Rr93jA/WIXp9R4lnD
s8a6dg0xgTe/U3fLKvj6WkwEsg6mk5fRzDj3dE6Uj492bTjywtEZIwNUQmrRMg7f
M4DclS/JOkOP4LyZbClkZB39bo+joylH5pdEcko6hGWqFElILK69nw34Xd6WNCIw
ITikLuXXDDh6fMtJHreEenwaO26txgKyTuciQj8MN1a3MEl+hlA2nUq1WyfmefIK
VaB4lUglFtfjhxeTpoaxC7hwogq6+SDnbCrrR2pA/uWbbqVjPFvH6gxe2IhxJYt2
SwgecnohnQrasWPFJ8qOF4QunVm4wBuV8PveTWDda8e5a66EXywJsAfi1sKopEc2
I6VpJbMAECzN67qANoLf3EnNDNmy+0cW7huBuJbvi1/GZbUuaE/ilHru4FZFU8c4
8UHgz2xqdZL+yAEE1SwPXfdRojIRlL/VIE2oIXg25m0N/m2yil4DKEpu6mo8YgBG
QrTOL0B38ky7ngU4S5B+6vIumyAjMi7AhxDZiNBl2eZH6MuaTJ9vbZg/H0CYwYDn
0rNiDr62SE3hRF8RazdYFZGwTMYgFfuov0/szDFZmV8QbZWNWxzKIJxb1BDy80jC
7inx5aho9VSTXWl8XMkL/QlsIuyW4i9dR0vKBT4hmm+qv40MavhFF5gc8eWiqMdn
9IlWaVymm4XdpAMfXS3PlNS9H0/SmUOP4LhnznpdeCHdjs3byFeuUC6gkmjAmI0G
BSML54/qjpYxhejpgx+ctdGJ9uVK2d6SDYzUuEDNjXZugkFkkd+15YJzkNSNWQ04
Cn8DzvpuJi5J1mdcYKd9qG0TDdn3k0sBKTscAqIcSjqkJlBphOlfsWnWAcZ7rZG4
UEpw+wf3FsC653jC8zsYRA22Sd9njAo2ZJuWy3gWvks7s47wsc1fUZDfMimP8GCz
u2mJUlsSK9XmNlj3NgakXf8CbHTjfCag6Dhfk90gzJ3iJdiVxF63OufU9g/PmaUf
nMu3JdKyc2w4Ilas1vWipyNJIvtuX229VWAXMfn/JZGU3tpLWITzygtXpTMR6l9N
V33U7yc5Lul34oh+pnpygH5k0EE4r6+YEJljcpDQg226AMFHzC1f9CQtsYZ3saPu
TYTRorkyrqIQJX99EjYiEAw1JvAiiyluCD9799+GmIdvC8FaHaI1gyOHEBx0nXy1
P38IDne2NGlz14Zc45ynZEFEgX93TO1DO6AA2h+MdvefM53gcEzv+y8RIFk2NmAJ
X8NiDkFezqLEsSgGXkuTDh5Vi/7h/LoSo3WIg3EqtAcuC9BvtNuatkRhLHFSWCxn
IVp1Oox0HRkMeF3DGOoGWlGdUX7dLPCoW2d8zp5yJl3JACTxli5j0vRsFLKdeGiL
knfdQzyotWW1tX+o4Dzz42nQ7Mt9A/eTSIRLdxfLuzcL++iBDP/JLNJ1TmoEkJbA
n5cLdhY186zsSRD1/1rC8eys2UixMGQ9J7dDoyrgx9TtKAbpbMo/iTt1raDjCLPR
p0wfxNRjSBVwn3lfMdUXZQhoS92S5Bv9YUrXCCDGD1G3MXJydL9DGdMNDdvbPF6t
KOhJ00Rm7uk2CtQTSvFks6oJuWx7JA1lvswuT0I7Ds64nOAG+W4cAqoSO1q55hkO
rAl44D7upS98U2G/UH70bhtBT9OH+sl7LsSL3MlQE8FuZnpAyhDTti9zyVc4preQ
nkw3eyOp+KmHAL76Dhw+5P22BjRIES9MpD6O0gtau2H7iOUZdRVVqPpEfrQTwr7c
huG3eHKP1SHph0b9UWvKHikgEHCnn/Msuw9OuAjtO+/b+hRRnfDCtMWHtXSuO60z
ZZwZ/ozPIxf4pL0QT7M1ZtmYI+mfFcxCtAdryCAAl47wRxJttdLcn2g3ujEtlAuL
idmqlk6rDKmqUZdJ4uVRYaFb6m/5PaqF3Y/050d3wpzFXLiBKVE/5quM45kDxcty
BeUiSjvuHJeUx1464//jHyfoeovwwrAKooaOr+VyB2Vl3P15lGAi8SMKYtXS15+d
qbhQmANbMSzPYavJszUJOR8VMnzMxuDvM+EqlENCH167nRc5epHUFXJRWsklJnZ4
J5V4M8h3NSRovYaHrec3oBjghLpgs2ifUHeObC7RgjD+6+lj9FFeWi2H80o/iiGw
NI2K1CTDXgbTpF/L+EvcjhsjGXJDztVt/8PTRqaKIdmtLk3Q0RB0DCSimoraObgI
dtE8D5zuXXFxGzxC3ORbYua51UwRskQcTg1kZ4y7CgH1siKa7bYgpB+TymVIxi3i
qJlNL6ky6xJOA3m1XQv8JV5RODSKtQmfAEjvDtti/ZIBFg5uxJpMXJyLfcxwoUJY
YY7K2oU+q6bYK/QzmsCCmsHPkIZFTTQE5BJC0mEpsySpW4qpd9xPei65ZuMLeMuA
EmCeiqb4VqMZ/pMRfsZrh1dPQy8WR5pBApZ/ufk/4MBsSeODlmcrRIRKP17ybuiK
RHVlpPhxSfTfhUGyl//XIQE75Wpk3EKgiUuCPGjnBwJFRX5+YoBMwnA2xb9EOvrT
+7JngIP+fzPmAYZf3M/fphX/F3UFTOVeXBkku/TC65RgOpvZ0N+/Bs1Dj0iI7ZoX
pMkElYJMm0LBu/gXbApNZib0aZALvRbGfNn/dHrUqd9JPH03hVAtxhqK87S9CFSe
BDv4qtUjMUXfGXNoL/d4fM1d5Gr0f3k8eWbnwAvn3gPtkcFAvIDQosITcCIkPcM/
jYD98ncxVkRi/apcl60wLmInJLNPv3KJedmVej+Laqaqcq2tNyRBPbyoWPgNFaSD
XU50ercfGYn9EiYK8Hz185elWgsw8lP2D/FBY0l52yGrMgMJZzUEmXDvfDkz6s7S
vRbUJz1WXbEfFTtvoqzN4l2lesHX1oNgMH+ysCngMUHBGhxv1ruBZp1xJTdbXn8b
Wm+IJXdj7BTGHwIg6Kld7wdAf2LzAycHgNu4iQh5VhFyiVWM9WSyOofz8w/L68MJ
XfeWtlbxQ9kMk78Tte6HeF7L5kFIR3NXQieqJDd/EQuifheXQ+wp6YbW2wpPpWur
0qGElwSuXUcXM4bZPyW2g9BEIHGM62Ee8hMJytOr75Nof4S67iWupur5Rop0tf0r
j/mzSb/McIshKysZ3fO6xAOTTuOYu+BNNZ3OwD516JQG743JG1M+XHLKe4zDI1Qr
rtyxIySQ4JbliffYv86hlQVW+A8MoNb2JAhiSVN+JnD2tGYG3DmGr2qc3/rF2lSi
CiSj90TcZaLeA0ZLqOJGGKFhPWDq84t9kZMQGaM8T0ErV3J4tajRH5eLDQwLd7c4
POHAXSUs+58Qas7L9j5GGwSBcrPqzk65tZRVW/eoR7ryt0dtPVOwSzBQD0R1M7zu
jd5/UFeWwkf5Qf4Nn9fW55xm31FP7FUwugLD66igZ+QSBjCp2lBlObFh7h4LojHz
j77zSenTZB91AEl46s64qZjri63RYxnOX12/qgz0nNQEdopvMFk75gPcQmzFewAS
MLUobMxPbtYoe45B7qSGPDSVZVedLfAxvTzN211HYyrZ9cHD2Ve61BtEcUsaH5wQ
LKA9S33jfn0DZF+A2KSr7OQvgUF/3JsVMT3LlCBPVQxlGnkJ4hXrfqJKs5KT95zG
abpo13eiBZQkw5Ch7339gD/Hh17mZPTdByuAH2F6F3j/RtyvDzH0zGW21zyVzG/5
jXfcRF/iOG+FUxkz3ACmTewH3ZzJbFPwU+b6EfGxqdJuPDlkZcyKg/tmyPtwH9a+
QXmBiktqi/DVPTF1LKd3iBVlGEiAyNYOZV0hSA8QT7SkFzq+XdaM+rmP59CLkGKk
OpwX52HxfC4O684sWs/qlHhn82C8Gl7dEGXoXfJHUOtEsepcv6vkqzxgMUrvtO1O
glIT1dUL2SImCibWrvg/r60BjF8VlJyiUmvcMg3HIST72Ik0ZbVKhvmX1zc2SlrU
C2uRQkN2fjMqiHTUjX0LW4c4x7a6P0NoJQ8wVn6P2qqspOFPv3hVIsZnMEDdH/4l
ElpaxJiOE2M3PVlDVr5Y85kumoXJulugQHFVt9Q20P1b7fz5yxqREdX4HMTTGrk9
VdfjPWa13C+8I6qbPlyDTYLl0BPJIpZ2ky9UjIdk4ptV4btLI7EkSm+0m2EWR+c+
I19xmn3JNGrNfjCkGLnKc5gnmaIEZJv28Sg0m6GpN+lB3BVB9Z/q8eiBURhMkWoe
qhgLxgnj7AHhpM61e8KDyuTAnp2Qo1lC38xE9457RQaVwdPDghCZJ6c9qn6nSEjE
/2ZwnPKXhBgIFHEoYXcjrVea27GTgeUqf/JJ5cpMsXJsA4ptf1QxNsKtcj50CSVr
XMih+p5+lStgxVgiRjU0OoiZdYpTqxbD/hzJfNf9ZrZBufiqQjaMAJmlg+8CpjLm
qJhds6d9UZeYan1dngz3cRdbSThxo00bFShGiEVMffhmftuHf+bvnMjBnM6caXdN
XIupPbaIGl3Z8S8hbDbL/unlyOU4PA35qufRJDqf3VpM5eXVhK1rYoK5dw7O6DXe
NoFYVa9oUvIuM/0I9gvJirCksz1VqPacSSneB5oOMo8hW3Or7VLrToNZMauNLSJ8
WxuOwYN0urXdmJr6wdUQSMv0Csq6zy7ZMSv58RtK7S82kGw53nfcpmZ71Yk/81k6
tqhvOkPos8XlotypfF0ON5H2GNNdnfuf4NUYvri90nepU+WHvwQatw9/Wlpv0gKL
/9V1THEUOW0Fh7q737KXN5bDwTH8MlVDhlLLkuLys8KdICYn0ChoUs7WwruNuDfp
MgCAvnmu6Uqt/wvtfs7kYaansHn7vjFJQseTVCvUQP4G3rCqYRsLTF2plthOFhgo
f5VZ4eof/e6S3QrJ2R88drnsggMrRjsPGbBYFnFWWVhslZPGU8aY0kTKgMKfFt4w
4fxuDMXQGy4GBDh26/Ucwr04bRks4/MJplu3H0o7Z9xghyJJUa2/jRrOtVdALlRi
+MQVjl1o1J+9q12DTtuoFNNzdSRHeDw55FtTuc+SXpJVE+6xLKQw1MxwlDGANTF/
tmq/CrOAgnIrkWeHV74Dfx8dSv7lQmLKpcGWAtM/5V0NEqIqZxKMyFqwTfl72ZzE
BuKoh7JpN0foEYssFMODkeOX/AarKsYANgVnjUd3PMMOhY3mfCBRzeAwXJ0UDz2G
0FsxCCdqBJ/sdOfdDI6uvWVTucw+3SUywgYBHhMymofwnLhFERgOK6kMcVUhoFqi
3d5a63WxCl6eAn5JGmjkIRrRNLFMBxmV7SupCmtesxmgH/PPZqGhjxGZX85q6X5A
OM1MBk1KWKrANCvA0xavhBrNZoWs/Q5ZbbIzc4sMqRjRcqF/Lrw394SVKfQQ/JRc
xG+1hcjXVXmnjUDzwvUz+H4rgi1fTj5/V+7NQKln2fWGqYHOFdoCTRFtZZLb/TT4
hVwcPFHYBJ2mHlenQFK6lbAcYhIxLE7oYwgRzsfFISWnqiWoednKyA2d9vpYiT0x
eUSQUqIlGAOJMLuJEtJ065bPHcaw8QGR4WG+IFRF5dVgNsIPqUoKwNGz1KCITf2Q
67x7ygszu7z07wywxzLyk/NZXUEh45h1fAZ4UnO3Fn5vzDqX9G5EoDBQIeaB5aoz
y+jb8pntQhMPPycViZtKsK60YMr7lIrWEN2dSDXjXzyZC6Ip9jKv1kFq+oeuurxP
x4/axYfPXZxMkg+oJkqw9mTYc3q11DfnzwGoHGsXxiXJHBtZn1egf7L7aPWXYvBb
BNW+g/8zkFGgOssolay8fMZpDZ9b2EcfCoCj0PADPfqpDzzwM/c7N2I++eWRm7Ts
1e1fNOC8Z7YDUHcPMAEu9h1ICYvQ9gteAglsPYxczCoVzGFOfEe6o7dgTjCmUvbP
Fo4NAfA7tyw5AWgIhXWWuLJs4sqGnaGiSJLakkC3qC/9dv2Zop81TseYC5OFN4GA
mPCt42G/yB8P0vYlia5zQxamK4aAzxCZRf2ZZHuBDjMSk077zsLTj4GUcpmAjjac
ztko/VCG1M2V4V/EqjLwhOMtMQ7KtjsLHr8JbRhquk/d5jV+fPMeA2bmu3b9cPHU
x/gCmi1f/uecfmGP1k4z23wTzxwQjnbtKF/gYwreQrlCleaQFbZ5fSRVuEWEcakm
eKIJJWsLzYH4iyZjsx+iQak3Jp775QmkHi3ag3GlZdOqVBBJ5t/VpCejvTQ6DeAH
2FZZLE9rw6YmvOrWIdXJMarXkY3mBh9UzsLy94WEik6/nExh2UcVlhDegn0QMP4x
baMB3dHvINFD148tH9GZL+8FyzPOLAQuVRudFtarhTz+S5mGeTmf4o5ajwPfU4ji
KLK5tiw9KxnezkBbwFz1ec4HDJQzAePV+bhfYLogohPk4JsM6n+sGkdBvoRQ+1gS
Wss+aRm6Haz/T3+TLhrylKO7TFjE78LiqjAcwjilvSt0TUwG8JrvI18oT2baORcl
z1ulmCg6kAbVSVYQ/KSxPh1LtQPQTBZX3jWhNioTgeHkWq6REDh1DuTPYz4bw6n1
RgFa/HylKp949kB2WTx8kltoT/HbtZYx/eCg9vlGvuuqyshawTYCrOzQtGl5zskA
mqK6b8JweEP2qOivUHy6xk0T6aNCqJNX0gwJuudKB0jcppi2EVyxtztlxdrPafgs
pALHzcRwSAOYAN+9tzIUzN71ha6LlpMyZcUgrOqAQM3zqwzBElT3W2PbXVf5ld5z
Fmj4tQiywxpAE9lhCmfMcNUsfhaTiO7uiQ7QbncE8C3ZkZVVdTM9k+2C0WN+rPxb

`pragma protect end_protected

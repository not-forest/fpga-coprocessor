`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
glG9IMYNO6eXJah61ckMGcSV0YPkvk8oMRkDMOIEE4J1FKPQ/2OfyqZA80C8Xj5a
BUJba91/rQjvxs0iMSkCwXI/XLsTngIG8eiAgSvv9X6KVzeeU+j8TJ0F0lWyBCey
NbflpzfTD3TXL9+5EJgZ1qJkOhy7emvupJ5Oz/eKYTo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15536)
BuiAKj/IMn5gMaUtWdxQ6riHjKi6hTwkheeM4K0lQi+kKOzs6WBO8v9eccSWZNuD
d9IBOFwXpBD9ULspPMxio35kitm7EVs8x6ssOx7z8tfYgJMtXjG5cfz2r6RLxkcY
Mb7aFgbRyv1y55+639uXET40xuu5VWXtrbMxT7B9P3ff0minHMjdEy70vxXOlBdw
cj+KFlWSDCrffIWVaqI7houvwoPI8pYHvjgc07gU7UnB5lgQzfBDCnNcxCyQHj4n
runrTm4it3wrPYdMhhoytq5Cbtw0MXiKZY7TkH8g213qKKGDj3yhFnzRS6UbnQWS
83MD+eKL7BOhW0QvExRNViYkfeDvvPUzpyIWYusOwjdAnCbZwhhFA5m0BpZ05585
l7ubDjTrStg2skD0TALYxN/MjZHz7tD+0sWHMFYqMbiXKOFu5bPZnD0dXnerGhWF
3DGb4uk0jJZAU6jCv2k3x0of54zZyM9GxQiZ2TGpNYEsTAot/SSDQ+DHEV9vUR4W
xkzzvaLlmzYsD169I4QPATkzQoxcyhrWiKMsb3IY+bczkXobK/TP9nuIjRtMXIlq
QqlLdcpCGZw+XEr8PnPCmFU6nnB8/IJcVjj6kbfvMeimPsRWPxGjg+HcfkCtnBdo
SO8C0V4hSiFBtL0491+qL1CEvO4q6HLzsgCUfByzJaaEgt44u89Mzj8OQodL/O5o
t9r98eWJfapI0hXfJN0VdTBc/+EkGXpSvEBC4vih1dygEP0RP+vzBa0Qwn+5+9mx
sj5Ovf06pg+78sN4J1+ECskjuOdkr+cebiQ4FJsTwqJizOVvNmiJXcIFHLmtHuWa
LJM3bejdIksv/MoTP7emjlVlAnZApq7r27uOAT/Qfo9BL7sulnV0rQaQWmgBn8qN
lVzPas1OdaZVvK8J3aXLuDFiFG+hr1eTcv4juHha4JGpBXBx3O7T+ms7rmKSCXWm
wR/RCEsHD6VDJ42CTU2MITKR/eSvhtiFw1cmhmwEFWepEiy+AqsFB5z9ENILnurV
PP92sMSQbowM2W8shbN3WVaaQWgUKIVIFX4BSf10JWWPNWGC6UtQNzI0tL9+pPqM
J1/HZpAngN9RxzVK/HNwn6crB0i+KimHMm4w4XBu8UaiKijrE2CejgTVNrNkcRIP
4RnCs+Y6VzwqAYtS1e87vKO4PQs4npUS2xth0mhRYfixBnmZ00sTKjC95S5M6QHi
1AM+IPfT4CfbVY8QGgkKqXRQXsLhThsTa+8f1HI7/BZkj6frNjwTvRzOIcXR7aV3
CwJXVDSBmf3dLLL57RWi5HI8rF2hgk2+RHAInBk5y8Y5f3u8hX1hrnxTuSwyztWi
cvj52rPXw4kd51rsSzYfcyFaq66T6OsTLdwm2VX7rGxtUViOsX9xqogfw11Aszz7
i6UFxPN7k+95iN7G7psI37Bo9vipqCANEypxGi/hZzhQmtFmEvrJ71eZkyL7pQP+
3q3KndXT5akNN65z4/QsWZQ2GcNlvJ9p5yhuOpCjTBgJqqUv1OFE2RgR+iDcrh+G
osfYPLzQR1DQvg/eOjPlp4H999DVGZpEFVm8QeW/6WEzXYUS/y7P5UkVtXR3meg6
63sEBEVKjJ9n5CmN2aaF8nHSA5VjDX2YBRzg+6AsOY08tZoiTqCDYIS8hfPgcRbs
P3/GkiP88cU6tUcvVAKmUyX6xwEZ4bY1MTUeNWyV4SPeDIsbsGGdo8a2MhJlNjuy
pyusuASf69VeSJ/vegwBP59FKk3AZZqsluUWIJumYZjonO7xihcBY1H3tqDQUBgf
NWtARY1SITHHAT4Bbt4aCKr16D7730xlgiNTodH8dQ3HoT3m0YL1UX07zMvyQJ8f
1lTMNmyzx7MjSPyuppoFb8Bxsc3PT34ECsgHnpk8czrXyTQMKYc9CgxtM1ai+Nx6
Hjrd6jgE/WKIaNVxifFl6G9sBX9Lhta0O0oG+16wTyEt/ryohMwVnZ96J+YG+yo0
c2uVGgCJz2hWDdbNmV8H/ifFWEWj0gVo3TwWUXuz52apWPjQgLKbxYy23qHMvHWy
3i7gSXvW200l/+ZmnwAOI5bVM6KxV4Q3sOrrtUjKk7KrGPpSocj43t/ZkvMABiL4
J8ploCTRqVjqijvtJplAOOcNu/Jxsc2HHEh9cTUhu1d0OwGT+kU7IRAJUKCNQ+a6
IhuM7PBnAWmey9yKpS67ANUxFj3beURZWsnBn0zc/PVb17JHB2Ai0I0wA4E/m8MR
dLn//E1fZwEzQ/eYC2ySZRepdSI8C/+uFlm5hjg4BUPTs4scA0BbGchqZtVVEK7x
/hepfBDSO4kfgP5W98aQCKsN8aNNktyV/BZFc1+Qr5XUeBQrdlIH9AwFfSYxxhqG
OhBpqFxiNuuWiE05L3hZSR0D8wUCF69dMa+uZXnAfV7mUZSeGimgapGcjZlP+kQt
0VUSKiArfknQr46Gt8/uLXN5tsKy6yOJ8OBxGIxXWjwleMUunr5FwEUPJT2pLZTl
N8L9ynY0PVB9uryHtzotNXWuQhQBlHPuZo57b0pFlADXkTQFX/Il2kMi24e/XfZR
D4XQO7rUEMfZbYSwoY4C7+FBOtM501siNcUrUkm72/y2Wm8x1F1MeqZqHiZnBosN
DQBbmzcFW7v94g+mBn6vNlVHgL7XP7s0S0ky3V+Qh4uZWDGbbkqhn+slD9PAqKuf
OunZwdCMBbmMQUGxMjoUDq/onhvubBpZ+jVqXouYx3C0xomOBr/PR7b7n19pamtJ
GrWx6Rz8uEMzKSxjZN/yPuHEAlxDwE1UYpI+u9JvxfwEeYpupSIJ7ZFp6SOjejPp
l3f1/jtr4gPNWl/9vSep4ROD7ZSEFhweOsr+ub9niLpTXFtoxAAECCbfioYBvgPv
zkZqX4T8LgdI92PkXrceZUWFuTXrzwF7POqg9RTJYBbgBb34JKmu697hf5K0u0Mw
/3r6d3wzEN9+8MN4tij8HCSMmOz2SjqVoOztxajc+0IQExK4FWcUa29t852+s6xK
pBv7F2mT12jiY6yG61euGgtGk2VwE6sn8uS2YCtyDFPZlcnMpbRLVqMLeappFOo9
Bt1NtjZEmm7aJ0fhyDHnwSviXkczy5HT41f5EqDqChVIH2PIRfBj+21lhUoOlmU8
qe4gsUhO3tkQfqAF/btkQtt2g9ghAjXxtp+Hg31Zl4Wls5QeL3yC3ULaM+Zo+6yM
d9tXPC2etvE/wKzbW/wHAlGB9WinYTGb2GBljtXXPVwBPnOJ7opqBxAiXZ0o/QQV
BsU97TRvSsqA6BPd/BxRmzXpzOc2r2JAlJQkoAs4Oo5VdHtnXINKfhl1X5pTVooh
WAK8ZYcF0Mk3xjd0dVNykXlVsuU4vXXZ6PSG/sbJ4Z3TFNLLvgjsd5R+p7XaUgeK
wja1Ohcb5cJ7WNbq4boFcVSxF6q39ACvVzOGxnixIp6WMmHf63X9bDuQXbxTR2Fm
Gjoi/f/N61AUjHRDkUQJ1D/Fwm70Jy9E7bm2msocifYFBICF02VMpWyUDsWqA6Bq
OzUOZIlVm8WBRQ8KgrSw5lGlBK8b3v3RpQtTU1bcTTRLW3JGywt9X2OTogjYpQnw
MtP7n/g6J0YM5K2H4yxPR7nRwg+mq7VA/zUacv0jkW6mbU3jnDlioPwRlPqFSoe6
YgmfHNfksfid/pWTgRDoFw47lnzyQQVCJhu1TQIXWPRYuxGcxhJJ9gSs+fWvS8Mc
8R5fiPuKJw8xrZLSm4pofA7AbojZ1rhU7HVbV7uLuIijQIPUqDtkNLqxps6B+eib
Rd5fGzGP4o3OExhd94PV/xgHKfGDFWYPLHFZfgKBFwQpeq/Cp1XblrJXcDnzwA3V
8pXFXmyxTrIXYmDEnRXEiaLgE1/+EnsjYjD29ife953xaDZCp5436fezMk5tP4wj
ULbLt8Ow0C8hlZ819l/B2PhkbYg57msqG5KtV9IJFqU/daAYxq3+7oS/uyr1Ph43
S8GTzRHl8YA1x+sgLQJynLv+zNBowB2f+EmX40aU5q4rFAKdhn7hNQCSkSaRRYVR
p+Bz1o6btr6GTH+IIvWpC/YuRtiklgAr8tKyKOwYPqy4RhpFfyYtGGnAeyNKMCMd
8s/nKIVdvENgEYwI1yKneL8Fx7j6FBq4SEjIyI4C0N/tDmvs9GsNy1G87ZqtXvzE
HpYiSVa1Ris9MjASE+2GPj2n83zq89y0h8oaVUmxZ4+7BDUm2K7Y4NXallo6YAx/
pvdFIN1nYZcdz9W/JxEZYbwR5vC0rG/tMPJzTHUoD6T1deqNRwX3VDHEmXzFjx/L
Bg9HDIdW+w4Q2LqUkqZBoFwloMYQQdyxO5CyGVUlciiaitqKqSzwHNmDfIl3ik1b
weutTq+miY8MPQ931EQxsXkld3pYCR78dwQhY4BxW26vzSfgszoQAcDW7g3YMWKF
3U9Bp3ZQw2ycFtQvR8kj4X1ruavpMp7KP50ruh/pJjYItNiAGPCtM0Ifd5bMYUnE
Zvkv24eSImrGspAcl8m3+JZ3SFwt50JvfwmsmVOUEY5IjxHcjQNQcd6zfhOk3Q+w
5uOrsTWpcviyI/KxWB2H+GIfUE9XtF1HsmcsHi+ktMuAZv2ar0UEc+9/irpgMOwN
8x8E4o+1pdUnTD2imjUzZreksr4Z4z8BsV9+n8do2SkH9J4PdtkhOms9eByEiC+n
VB7Mx0GaYrJiciQWOMRIHGKXouE0WKTIDhWuW0liqIijLcmP3FGFjn/+gworYmYY
8z+QxoD86xWKN1TK+xxDxpkehXw4Yin2mp4FRSZR/oYnozi+OLf0Or/rOaGBAJQh
sVlU05VSXLr61T/yZBqwsDHplsHGxp0FFbQ2XiKN3XxCM+EkUSMg/8rZiU1juWJ7
Y73KntyzkSjY9fqKUxSkCtnBvLyS0qvXhQriRM5htIPOvw3D2frO21pgFBZWqnl3
ONN2Q11FWgkVz2RJMlYqx+xV4Sg4EYjnvND6otBp/c95Hnou5TbN7dDqyUo69ZMC
lPegR9ez5kXNpPz+EJGSqM7GqV3PyFLTECqRn7WDoBS5PcFcgglhHeZXXzEpMEOp
1wUHh+lmDu6LCZT65+zkPm/qKiE6cDtZRSKS9tXL4Jb6IPYH9Ac36rhQMotXlS8g
7L7ngKOnWTn3QJ+d1sSySnsd6Gs+l64NDxsQEDI6wltx7v1KhNGCSaKE0+ljZqUE
qOJ2dFxq6nard2SaBW+WMbFgVi99Q5y3AfVAdnyWLiDLI4spsstpILEvbUdPsSzZ
NDz9LDkCYOo9kjqHLezOZg3TxKb+GjUUQNImgBpEzTLLdKnbBfVCVVV5yK1zw+b9
MXe3T0xpEcQ8Wj6xmQRgOEMFvlQ6ifd7jtVcLynVn0UbitNUFh9p37IU5WsvR+tw
xDu6J/TAY39x133lWzMO/vFNo+Igr5yWZUjntcD6p69eRzQrfXvmgwBCnMSgSxEZ
s4ZLgqtfUQMcSWApeUYz+1Q3r0eLIY1vQpUzX9RCG7AY+grQ3Uf402WeLBUOpXhT
6hToZiZWQDUHIN8dn0SJGBh5IM9FGiE/ZUkquZ3b1EP4R2LtyEboh5dD2F098+HA
AQuETRFMBN1KwxMEN2htDP7pZCBh1cq3/KYwRwzxmd3KddxPmN+B/WLEMHrN0lYc
qE/gsDL6PUjgQRIEZ2sVMfl0PvfyDKmBb/HFuFwAGJ52x9Qnjn7uyMxo5/yd6p6l
ULbhs6w+dnPotWSdOHcViw+zf3J5SFWfC0eegdk7LBnGNKwXYlmTrzk0f7jIEBrj
bLaSvRwkhbJsMlEzScKqhbAWg/2hWjNw7FwPc/w4NaUuIzrcLdeeFKczTcP3+qAD
EZXlWgT/tfvdLhCd9cvjU4xfSlnlHEn+GChAg2XrD2ywbUusAId+uYvLDqCNCz19
g8mAI/XmJnBS4tciFv4YSjyHMK271fwRsS4+yQ8hQMJ4ja9iySDwXS9VHZlFY/LM
4pcxZ67RIq52hZRM1DExD55ULnvQ3BmlxXFWAEa2kzSEpHlRQA+OYUQq5V/De05Q
DIWHuRE1lwSRm3imKsf5kvbhGVpCV0i0tfPyc+JiNuEqaKBkH8TgJenazcdWrOqm
URKVHup+7+4toJri0jEMJRORPbyShOEWwFMOk54sDHoafDc24NDnC2Re3Jlvbmgz
srbyvKDslwWNq9Ls5uFOH/b5rKr01sfkBLXRtDuX1YWm76WHDIuLZiy7Gd11WPDe
+0F8YTpqZTpz92/VCyq2LrIRge8zR+T1GoeymlsQZFfGgUaI5U+RtHebvht10wjt
iB9CcN0wiab6K6Pryqu6MTJ9lUKddfwWdgjx6FQb0H02CNPFZ/ZTneIoP7VgHiCY
vLKIAF6tzyYML2SwWJI+jMrlD2dLa1m5G43xTl9YBWAwluraGAs+xmdD8ET+Olz4
wntkN9WNwvkH7MN7/dyuoAaV/aThCs+9GozFFpG6DYzYZ0MGW/Y3NBnapmZR6ONh
3EhJQzPevuIFNQMYbk6MJFge4tqZ/ipcRkjQx0sOxjwgVyfxxAgUp21bo9EhQlsM
LW3m0deeq3ovXlhcuDQaMjC/isAnVoI1Tg5irNTe30mOEGo2yYMzVtFLrkXiDXei
z74k7RVYOMBvBtsasrbPBCCADPrY9tkakH0i35qVM01eDwiJKwlsmE6QKuyNXNsh
u9B6KdqzFDNTAHpwpC7TRyum41NTIwNRqZfiiY8y8cqRxlFWIxOJuoNYPEA/9Kq2
BiCxLVvs59TymMX+vtF57M8rxSTR3sBelAyd6G01W/t+TWAypS2qyn9jV2qY+/47
2Hw8Npdq6WveHM7uqjfuMJ7b0QP8c16oU0cZW8BJbzVKrlnR1hAEO2i90ugEBGjL
xIRT9liNBcoivf0PDfKZoJ9tLaah4JkHERV7DmeAScF2D903CZjX5+2UgjXbdey3
dPYj8jYagc7QoEWCM0YQCJFPjWaYjS1T2l7pxJUYqys7KvdAgQ35perZjm5rlhFV
6vc+4NNrgIxGEEwsokB1ZK3BzhmpJ3SfUbSFs0n+viuYaFx8MYnX1QUX+sE3W7h1
J/prUdCbc1gIPD8tAf+w1PjIGfRZJ9pgeiMdyOeNEA2fd0qOgF/QNauDwsp+MqW1
mCA7G3JiLoNTI/ikrDTeo0ERo0ZppcSSPW716jR9yIhGd4/IiVxbGmOpO0HaYHen
UvkcNbFmdDDmpl8fQASx75wGhJhPoeOBOfLt9Ma6z0fu7v2un73CLIgO0DFPgWV8
Ovruh4Tr9KlROLsR2DLjHFXR9Bi0ofnWQZSHZzjTPOhjlqEcXoSc86bUTjaXrduf
nqmsLyJFSvWgAAvzlsMYVun/6jVrTf+JL3qyXNNuepoOCqGor28uC581K9ZGFsmq
K7vfMu5xvmJwpLN/Nc8Bxb0HiOqTNnR91PzQDW0Nt9JklBB8RswFHdAh/Jw7Wdww
OsbIF1cF83205BGZn4u2d2IOXgwIHEteWg+IgLOphT5weJzE4F2NDe7N2hohUz4k
Id8lpSl34E/F0WF6h2pnm1DlJJyiTFswWUetq3NVLV6EYiDRWanAdJhej3NNPDad
eFFfYSZsdsWfyFrAbskEz9fC5DMUsPPid17fGWYk12R0YSa9KW+/LBSK38DeV5O3
Xi74B22GXZYPWOPuhVe6GNlFlBbOF+s78dHUTpuUF6sCFKb56C+JbS15AkPqLmQ+
h0VxF7MpLWQkSXJ/6CZKprtQRJZX0WAarT1H6nDy9i6m9vPYEL5WcY1qLmpUyVKe
Ctl9XUflVTslDGWz0SpUCkE2iydO7YyaucAuGyxhS2l+2Q+Ra0y5pORA1d7phKja
YRxdLncspnuOutwTxRrVQuP09xrBCdybsjMYkIrlvPSoJ5U1zkMyJXDg8sN838L+
/uuTpRvENLc+VBV7/MY++R4dyV7sVgwvuyZMXVfPjpI1EwDJzkBh2d/uFl92NyqH
wIUbn9iKo+wwt+xX3yweuCIu7fLTnRM5jHTdFaJ8igyKBWa8wjQ8+gTru35uwWBH
8vA3Ibz+LupbbHahmqdj4FHZVfcIp4xKYpQ5gMXa/rVCiQpNhDJRvBKVOxTKwOGg
hu8ebqcQM7QyALK8Q3+B7pUVQi51/k5dkScs7JEQ4RzNO5wHk64rURWfl5hkA+m5
fKr7rvCSUtvVwFlO5y0x5dMOpaTz/qWmyk78RDgf801qmtj0QtSGUCf+A5KmUxxV
9gpIcS5FYoDkA/eOEuWfxO7g2yyI0Am0s7/I/a7FjXxSKOe3TOSfiuSp6bvUi88Q
uMnu6eh2/apJpati1h1ig/KaBufrGk7pnwQTWfkbBJr1F0MgKwjBtA9BlrZJCwt9
CTiFlCjlYb6flNXAY1UPZHhxdMZ27gp9GPjNSTG28NR2zrfMIqflFMDMcHsmcYDi
HLY7P/vDmBFCUxRYoPbBXkrArfQU8zTSDa4b70NGHJKwNT40w7f5RikuTaWFi2Oo
hRGcxQlhX0CJy71t7Q6m1xnjMmBN30J+rEcf+bfH20La2rwDi8WfJ3ty6E6D990X
zWe9csSjT5CNOtPy0Ti45+azVent472Z5iHLRrS3Qf1EC7YGEhWCUz5D3Kz+LCJM
rrf2S8quW5w8zDnff5vP4u3mp7QqU6wxpa0L/4Oe+YjjVVrIfHwOJz+wPApinSv7
x+W8vOWZ3xsIABo96TQVFlnDmJRUN4Rj+qpQSrX3B6xTdAumD8MutOtB0SQ67Itn
uYvZNTZ5gTvl0i2TBm73oXS8EXxOzbwQeK2semGMQfRiZ+p/tGXkCK39zvhVsju8
6S7YOUt2DELLLuzTMp9Dla0HZ4KUSJVJgTnP5TK7dzkzQviuonK+Q1HhyWQgegZw
kZX7jSnMGo0Tu7yORgA4gQxeyttD5rcmYCWpN0AkU8pEMffDEufBH/1hXUpV4FlJ
nedBzHoEd/ZieJ1lHmbBb6CR9tPYNbtBDPJokD1OfbLRovWHjvbtTUJZ8TI1wx9j
0kGwVj2dq4ZP7j817GcZ6HHD+uHf0u7zjPYRzFOZwjxeZnp4EzQxbkfu2DX7idfr
iTtBmlieQy7ZSnF9iwbo2Ccvimzq3yv2MKdAHpbuCApxuPKr25+e57k6PMJzvwPM
XchMHb8v1YMrDqcVjYSz5YSTU9jcuShIMwp28z2uYS21xuR/Fwu+BxfgxJgVTBv5
9T7GlCarMa46nHhuj+TKpdC17PEieEaumFpbwHTnR5STOgdnzJI1LVKA7CcLpbw8
E0OhQerwvEIqwzwj3A0LbkN4FN49VUFeT34mMmhlMZXeUsJk9ZInalf9pWQpGBLF
bQD08PE1LOCO/xwzMRXiHBx5HUCFL3BY6MNfK+XPc7qn4baGb1jxxJsWe3EV9SPX
3iZOizD6zJeCgdNpxPLMweASlAbA2L53UdGgT1ih/DcdxmngF6joG8BR5CptR6an
mjSufLAGrB/bCJa36drpcG28ifpQjT76JuvwTx9xy4HpbaMvEW5oVExoebrz92Uc
dFfQ0uURTlX2cM4nEhs37MBA5IgXkLsH/drWCmDIb2Jl5eE5yFTKhx7PDplTVysT
1US1xJH4yGJErasNmHndYno0s3rja/ENKSxwPL/d78KhJooSseUSCCwu1fYVQHzj
o27pZ8xIri5jcgmqSvVoooG25y7n9Q5zdyuncdSPw9hk8miWyMWRRC4kXxu9JiZ7
h1Lc0na1TQCvGEusYjxZZ0lIf7iSwYPvZZhJ35RckO/qAJkLKf1duUmlmGuLhHRa
rbbMrOy+m6uiZvFF2fX0AESCGjDyCYwM4Lt6xsBhHhu63N9DVEZ2mJ9rCJtw5w55
H2qS5lLB8sCuAhjuWw0bkIg5LL4hjQeMgTqEJv5hK3BVFf8G1jArzwzax14nIm5b
t2d6NQIMijag6bZ7tvNds7dGj6/UNwDbM/h+U1n7hf1bnKA6mzV+gCucYStI7+3R
JA2sbQt9eby7wu3SnJPwNWJ5weV2m+FMrKpF/Lcs5KEZpZDxSQNgzp1mc15Mm4Ow
qLdH36OHGrAgugqNyV1iiRi0fndQLQUvyBipmZlLATHGgGYV3Zor5RjPA+UFA+7q
pShR0HRnhoPubSc2GnqoMYju98sz1QUnhlQ/2sLE4hAe1Qim4Cz1WkKj4k/JXsSR
3mb5oPCV9O48fJ3Y8p5MZ0AoEOHVgiDNpzIipALaiyY92i/zlHgG4UPlvMg6u3dM
Moh6QiI8dtIUmoyQ5/rOXDdrTrKpKxW6pZPelCWVIqZ46Trd7x6fSBqtfCKZGMl/
TNkrGdjCllMtUiVkTUaOMDBClHdch4VkGd6vyd/MGsowNELJqEZMJf4htCBYUeY1
0bcBneFK2/bswhFk/yc2M+UGoRF6U528iGmJsDsgY5IKX2rBuz6NftczgozMsiUP
lZjp/EEBDRubefXtTiEEL0xAVW4t9tFt7hhWq3PK2D7l2Jx6Np03KcIxzsxWqbyC
pi19SmkpbIYYVag9lGLEcc4GpsxWq0BhoYBgWXMLpPG0ZY8NJg54QWuljJO3t8x6
ePx7rDWHz1faIG1Di2pAvMTxUTA2qkKxvDjJ5+gsknXkkW4JMT38wJDpKopxrcgO
LEkU+OEG3sy2Pplrm2LqTWaEEg8wHPY2089yEzndrqLNF4nhYAoVlkHcN/429IzH
Yeb7lAIVO3/yPrz6KF6aoAOxmANeGdud3rRGZgrONUNLWGij3EGw0RnlyH+u/sV2
6JHOZkTbB3vgIVnfuO8qsZxP8vBT9OqsEqPuowG5qaOvkL4rVNgwoOULKyXeEGoq
SfGyXtgWX5NVSgWeesJuKZoZi6daSr9YOlnTicwtuh4PFKNnf5wyTkjTDJ2/vFvg
IkHo41PtMUEU6UIhiDMzSfvoY1ynfoqmTyayAeas03O5LcaTGuMDDF5DKy3QMI9g
D8Zm8suW9qeW4Ztmpc3JzxNST/9jvhQ96uK7L34eLlsej5JA6ba0oK6moYC8BKnW
VnHfytKFnO0SHU2UHwW9fNtQNZJSNezusUsaUdAbNKGqiP5eqM13fwCZB4UTfVdS
+wdW2OaYq+JXawtPNfCn6pvmtlK9lt5wjAlzDS9Dc7tlizO1IfEtFJnWp6QFpPoz
ATjGBV29138UFKFpm8BpVTc+fS2S0zTFWC2e/3RMW2tY51Nhr0BOlexHf3SXQwm7
3THelsL/7sx2fxGL/xs78uCEFldmfL1Jq9+OTZQ+CnQUP5FUKvTlb1H47Ai/FUh6
uKyH8TURQo4Sr/KEOpDmKkBuYRt4xgRw47vDq13KKc8wiPJKkD7waGvwrNrzB7K/
ue963pcahouevK0dZQn9uqn/18vv7iN36F1V+MQFMEIbJN6J5kXV+ocNZMnHvXKa
2VnZ4rPO4K5q4/pAp1ZMDBP2lH00LeL/VTeWfkD9ZAIdyDKsDYIQzrrbAUJJg8oI
NM/y8oLYw2JFBEsw90/xFJg4nNcG7IoK3nPdpIG0APjl+TdFLE1jhsjejN6GMVBv
pKNthwfk9bBg6mlhTSexhLBc9eQzhuRK5RNuPhRmR+S6qRxisBmzXBzYw1URxZ71
AruKF9sb09l93Tc3TJYuRtZ/Jqa2+fj2BXA3U9A861/Z5wvtDc8N6qQdoa5+J2qs
ExrMj9uBdoR/JdBhHAEIJrCcFYg36FjXuGbZOB6rvZPcXKabnNGZaG6rwfx7n1Ni
8bh/QVJcZT6GmAbBu5sHXl8Gtz5CuWFqIXGD4TRaTGqZjyKvS7+aVvt3U9y8r7q2
l6W37YCYYdN5v9Mz17p1xHh2dyXbjCbD84A1wGyEFHWmkAwsk/duTT/tS509nLaQ
zSHScQjSAHBUxbSdNhhyNgi4b3fnkvn/qW4cFQLGomEtwuFpjpNEKTOamA6G3PRf
lnwmHtD3YP7Q1aQI5+zlIOn9AGiStOpJGr8iimTv844khbJQE/acaCciiOCfY7IZ
yp/RCkWeTy5+ndIVx+UP8XYzaDgvYDuQ51p42KOJ0RVV83HGaUr+s2PMinmw0Afi
lt4a1B5DMZdR8R1k0HiczKVvY765QlqMgXNDNnoFMmfNwjmr0eAw57sCk3Grs+qL
AOomP8wLGGUQH48/MBVNjw3izlBTFFyt85Fa3fzGxIKYZ4Eex8JOkBC8Kf4XatqI
IS43t8afk7UU1djrneA7R9M0nzkJSTh13x3KZwaYTIWcfg9HmGYvajL90/+Ft8T2
zfOYIcJT3Onr9KuA7X5NELkgJtbve1lTlGZJRBEabXoWPfcBtRUPrpP3AAnew1Mh
VMGEzO2jR0vSlLGq4vsZ5h9a7ByqWJH3QcDAk19eXWami1KZY30MirMK7HZCE2lU
BV7DC03zd2B/Pby5qJxqTiI62+Xlv0JKdmcq9pgx842r69uoPfIv38cvLOHxLmOk
S/sm63rsDTjrXRDt+sJspLY5FP0w447J7qW8hJz/en0M7mbbMyB+MoXQADJijPSg
WasRu8apBkHaV7KBeFlnLJFOiUTXCy8iUhG2Cejsw8tdFDkYSl0FK9CLENHvc8sZ
NdKUsr7yMefb+gsUk6A6BfSMMpveGUPyUqbx4NTncDMUMYZ70OZpMTShNlFDwyuM
IWAi/tLVVHeDbLlio+WeRdn/XPB5yEE/7LO/tPbyDfBXbEY7C3ESZHhLlU835eox
26qFv0VuhLQaKalf5nGqaux5eqO3qDiXt2h3Pilj+biVMbc+fYqY9ef7/LjOuoWY
vSUN4C7qylhWmwcYeIjAspePuw3bVE05Yo98XaJn6J2oP0CVYmx13WckCuaZBjJp
EUQv5nZwRN3aT+oNS9prc14k9zAxu5eu1oLKkuIOlzpNRXvdDba/JaBnHr9eaXeB
6xrsJySgwaIB+ffsAUCnhbkiPNfgkkTIR9pIHg8deqjE3Z0bBw8YXelbqvXSGRIc
ke5gCS1y7w2VD+IIaR4927/T9TqANyLtnjg6/zmewJXYF600EyaJr1F3gp1USasl
m0SnjhxOqSZjEIgMm7g+dGlqLn41LRCQpGXlidXNkObdp01QgrbcbU4zKVRmEnWA
pndwa38SkcIuLmQHNsXICs0nlaS2iOFMIAht3RyvuNCQC1d56L1fWlzmKuJx31UV
herr+S/ow1FPtRofwy9RappUP3PJI88gNddedanu4uGhyjs0y5iUuYh3uDlu8ojT
yawIeaCkXwo71mKQw79C/xLeF4bE3CkFX3gq6bREaEFc3juUAL1FK+yq/utnJU9T
NeWtwcveH5oh/niQlBk9ks8cJyFRYAayw5HO34q8Zp+8pRnGDEl/mlmmT2j/Ya+E
y9Amtq9OZYh3XSxq03cAxSU7lLFyrRhll4jrOYktkSNBTRU2g6gxS6lxGuLrbN8Z
w5jMfU04cdmD6e6e2sLbuJtIJatLzmD+HmwoMI4BtXMA7V5p1PMXfCynOqdPkiGk
aDCJSOZnyxZJDLlSnO1jxUupI6G9xogOEYgZafRY7zRYMOM990h/5BM3/frjmxsc
yVqeN/0xmWAnWVlo4D+f0v37WuCYBi0rb2IR06zLDBNPKiJiKWzJyEfIj9Ta3dUA
emrPIPmGlG4stBsRLaG+l81iERyGk85jpsYWfGSXNDdpWLKJYRvkkEDk4iyrwRLZ
1IjqOVywNahQPH32eGbSNJ+h75Idi7Zxb327ZIGhtVgs44oyMp3kcykVj2PUxw+Z
8Lz/AMuR9zFpdWu3n/SddDT730VNquJsEqezSdz2D+eRIZibaJ6ZreDKq6dBW4Xr
ir0D9YDov0oZAajyEKZlQ8AMDVLl85meHM8L+e8z4N2qmdS3R8zVfuz/3tsSaN3X
UMAO0bM5gGlH0VbDP3PkhuHgx/wQKdSAvG2j7e8HZAEHfGl9No9AiuKW1l2EPSss
kWTXqmMp1RAOD4hEWupZ7gCMOvQH9ekJN7M7gAcsiNF6Ros1u4fuOBEmUK8M5BAK
xAilHvT/VnJzA03t2T3HSnFUpMRaO+bLrjDl5UG5mQF+Ri0ud+dsqMDSKz5QWMen
pgrVntNcJ2Q9rf2hVLpX8HkGLqvu7attV9Ajw9iV4DRYYB7CqFIm19jUsGNdB0lS
rNh+Lhpmn0Ur1yVjO0+xj65ixmEg0XeBM+8WZTFbZgKXXnyBKGV96tE6fiVJx/0Y
mj42RaoT1Z6vYXxj04/Esote0VNbLiHlZ2Cyh9fCYXuFQ84/43r7sb7rd7wm+WGb
5F7J9NuuAYQFH8Ast/7+flKBvi2a64Txz/wErBZDe1DGFJgQXEHAUd4vCvqG53mI
nRGMRnMYMG+MEzkt/4d6epQFWCI5pM3DHSPKtTEaP5HkSKkbNJiEztv7rI+sqUiF
z6fyIpqLrWlxr+8eS5s2AYV0kWHRWH937jpMMqjZMMC7DD9IK8UcgkkkeSLdSoiJ
B39GXA3686B8eNCMvRBi3kMam5aPAmGPSn4e0O5Tm+lk/UKZdLZcXBL+hojznjDm
uGtkLWcp7FjDPErRIqTfZ6d19ipar8dPkVfsYRmBAGw6eudcNZYTAfNaeY8NC0Ql
K0OzsuZnbc9nZslRfiRxqEpVPYU9N7uR9wCME+LwWsjsuMMjD66vSRxn30Wmg3eA
HKStnO6/7AZ+sNlBM5ANgikXKsSb1No4ikae0IApiTj35tjq3EK1KchxG/9IjpOv
40kyJMBov0mjewkS+FqURwvUC4qVTDz7s9vrmV/AbAANP+TJ9MppfVHfejmREAm3
UtxOBs8RJARgo5L6I3d7RQRgqxafupr4xB8r75VipOmrZsK/pnMx6KNBkc8CY96i
W8GEwJvyoeOgNPeWj/EuT0TTczeHI39/1vd5Ky9wHjSVRXzCHpfvIHwXjgOnp9XJ
H2oiv4gJFX/MqFIvX2sl5lB62d6po18Wm3dLVd4+UGkWUIIiy+URChYbNbyxMWSh
F72Xid24Bb7LNeMP19Tj7qIQKaEbF2LhGcUjZf9lHRheQ6ZLRbwsqmdlhyEPaJay
WC8UIcf/g1Ax5f5TLWEUcVMgm1wFQY8RIO4D4c+nInsdcDagJ16Q8DUfMbsxLXJe
UWeFNjnNK+jOXvsWLnay8Sk/UOHBKtc9izpdkey9fQm3tDGGpTSzRkRuh2IE7R+0
LttOGknnZj7b96WRvbfMLl7KjtPT3yFcL136mKDekup0iOqCqlcpaT6oN4egxpZ8
RRGOcwk2Oy/2IIUws8XsX2Z+z442xN6n4a1Zu/uNybMvrJlNW2oUHRCvmnojGZ32
UJsHC/yuWAeRfRZF/sKK0LdWLGGHaU4eV5bQwawZhD35A0b9E+QpqYB6y/9j2e1s
9+yMApT9dplix8PFVE3ZD3PuNrmnVZJx16lCXi23XcQYjSUCA+Vj5CeiqQNB4oHS
Jz/xzEpkrGdkHt27xHPWQKPZNFpsoWeq8g5rZvMhKAhV0f6vcPRqG9CkIbuiArmC
fX9xYiN9qG4PZBV7dIzyRbQd+ThuKU6VQapopUvHpmmY3roV3Y6nbn+su0q2urkt
nFLilyS1Z89zshPZODgR29ZAmArmZk/GDrY1PUMy2PaQndSSN3+6eAwVhgyta3xA
7icdpfLO/TAlk91MhDIx///ju1PFK5txpGBDGQ3AQZFGiJC5m/+WNAi0ihpdKOMK
Zg6aCeZY05ZeNEwL4rpNFqWi+dRd68jhft0kS9gg0rHpqlT8j9xGKYludSVEjvf8
iGIiwUFed9we9qXG+NWz6r7DupFAD3n05eEWLqupmfN/uHuPMOjYJs22PIny7XD1
PJeWGHGspSX4ys7TPyFBoA5NiPtKJZtH9rOcBAijnW5eHYGqACupvJpl4JvuB5nF
AhLV63ih7Ng18ZfSl38yGPneuMm/EvIi52phNSXXiFIL1Nzv6Bm2EtyiwSOVefQp
pXuhGgqcaLumsqag/vcdDsyqvAbXWcSbj3GQCRSJzGJNtBz5EVnaF1vI6C9c9AqH
jIKhvsoXyCZefo+8+peHWItRmMoYhHvGQJ6uhQ0/U7bwzH1K2OVyXBEFOe6S14iV
AeLm+jqNvWypj8INqnRXxnc5vriEueoS99ZQckfQh3odLMJyLyWRgIKwd44REMTI
h3aCV+G0uytV0gUnQ3giqnixnomI1iaP0TMFTuqx8g0X4vYOrYqP6dLeNtAjmJet
FjKpGZcQkm3xcoAZQda+XEj/9LXUORm8R7rGF/5aXrpzfP4hARupHFAmceOivuKq
Zf65PY0MXrynPefH6cC6kCI8InhF+p8u8rAPnRxdzD4FjwrMkDFMFsAXQQd4y7Kg
hfsC2DDhkFIizjUu9UxDwhPjUXx/Pti6ZtsPRgifoARJ+bRLijZO9sKZ/NB6Tk9T
ZhCeKFgtUE/hUaC4G2TkQhpKFnRB/ZC7b11pxhyxs1HD0IiFAqFN11fOUH4Vt7bX
N189sAYCxvrQ3E5DBck6gmOUBuzIKBxrvOI6ra3ChWYj/TETwCrXUJP0KpqOK5yn
giuXWmHdWdhWCkp+OOElFHrUKGqDd8vaKRC3GWSXxECWjrrojKDWLSMHX/gUoQvA
QcOJ3lP5Erd2i5+tZX/lawAhS32Ku8qG3PKp6gQ1TprOvWRYAXCA3ymvYXSVkYgd
PgV0gc63wlS7aC1e4y+VsZkO7WeT6x/w3WXIzBiZy3GJd9lLJXTaoECufpXJDcvr
hKqOnuDgWmhTu4k3efa8P5gmhC1JD5bHLesDA2PduBOAr/Hui+r0D6WC0MY1wMx/
3tGkXgafcwgwhgf9sKdwcZV0Ng8BvmRa5D5PlAkrtTlwyA5dhBH37iPOxsyJjtf7
Xq4tlDCvjZZ5WS20NRqkxBAjHh6pxZ4nFF67/IcR1cpWTf7Oq5/Ca773nFbu84v9
pCQR6Yjy1dnsX/gu2QwZ2SHqGgH7X178rfYnazUle58EfaYx7XuE7gireuHONd5W
8Qsstj/QcHJdLExSmgq0F8z0prpGsOelprWcFVcTThtyWYV0T8vlHdgnxHB6gGJ3
wGqKCA8BA2VUTQrzyQmSpHPJu5pQSvryTWScTHHsDM4cAyluWuIOhGChyUR56o18
l25IR7A2jApOH6L20mo7bqqNQQU8LPhp0wHq2c0d5jyIDKcVRa+WG1OjdQXcDowT
5wcgzPxv5jZNfWUe+6cCdYlsV1h0nkel9X+LV95OJRk+18+ebm9z751I9dcns5kJ
39vU7eND8s5ZGiiZxwr91MDGXB5HE1M82kC8lMoMcLzrTQDp7uHFJ8y1Ist1tbkI
uNYVGhtCs7TJ36F1ngRjEGLihQ/oXXXERpB/M2YTxXmszHeY3fDR0sGcTxWUv5ak
KOy49fE13QtYfn9v0ceCLJStGV8ThK7qPgGfnCoNOMQAz0SZeW3fosluRjsK8kLI
djITdk0tJINkopBHRfh6zTpiT2+X/czn33vgoQyNikKmMhzWv7d+BhXXDmJ25Gdc
baTQPwIdhmpbqMGVZCbRQQZStq9WlVpPfb4bTe/yUzxROc1etUIkOUZ0BYgoA/80
m8nM9/UdjB1S88Zn5f37TJBxXn/WuB0tbQLji7MJKNbKLOvlAF86PuqoaQPQYXmM
UHbewH8xHyAfzfB4uIVnhknRlALcpnIIoabpbUiE3UQ3XOHppVqqO+PKYhm5+hX0
BzbBXaBnGjEvKrBLeuFlx+rPaAsHUDzqQnC660MCjWCy3QriRBzope0uk0Vd8c1C
RltBqcSNIGFk+K87pp4ApZ29uaCPg5an8Sgcokam7pz9qs6Mcp1DQG3QkUHMy7uM
StdAKCeGD3QtVeFto7MTvzad2JMZw7LdkKqpNFESvNOipWfGlIqTG7xk2DBzw/E3
0lZ315GyZAWgVNAfz94SkfvOXAnnHBS+bjDA581VZZ4Pf0irZfA/LV3OINpAEVUh
oiAaHZGJobOGCBpC5wkPIPY/d4+wd0prhYyCVRPAIdpyKI0XjQqN+Nw1SgeD8OxS
sx0C/BshFo3/guUt87kru2Q6B0BUUDxvtOnlfVjQgrtfnzf/PG26bqIzB9dWBJMV
+wsaAbK9Qvo5KpPMPHOG2+f3YSs77mPrq3rw/wCAzzpnls1JMql8OSOtJiqSamng
HtqCrDNXXWkjl2BbbkYiqNdu5Dp7muq7n4/pZlb1N84Aie9pA/Vd/TlixMmlBP40
tNgWX8OMjL4/139xzMjlWQY9ZicIQLoMNq5AYBIc/4JDyHm+s3N4nYtrdIJE5K8Y
a2Kw+FAGo+UXSpx1vfzx9kKwKl8Ev0zLMZSvyTJyBJF+m5aAJHhoRlIBHPRXEkY9
PP7oO+Ia8lIv2CzKq5FM3waS6iqvzYhYe92jfzcju4/QYRbIssIFH+1bUVOz1ofb
GVuUzedU8XUnVIdWGSj5jrQ76DVQ+/NYd48NyCZ62l8J2eudodzfIZLpSo6EZ5iD
/yrKqi+uHCGzDbkU/0p988PPszwYp44PPnuE+XMrEz3ROwXWg046JJPkcr++KWzo
4diWqqMcDlIbUlA66qHqmw8VyPHsPcCxqhhwq1lLwxsOw6FkUppcDDDkGm+aWWoe
9H4EHDfcLku3blXR8oUFtDIJhAkcyd6UONy53DssaVybapB8Vb1tcqrfNePYore5
lYkg7mCY9mRdUsZtk0B0ZytD4x9WQGQswNABWtNSPflI/i2U4Wy+aT3rAF5naOUs
DA9qqlC9W3JoPUbBfr3NBdaHr6weZWuoCrF6KmXYOARYxV0KM2DvjInl0tgPpPIY
26gxVcgMV8G+fuOPmyZ0iFreE7UKQ/mAGk/mvrmASK/UFu2ZSypH5PWtEqxWFcax
8qCvhRTDaMB+MI4cxbofRXO8ReDH6mR4EcDfa/5756JZoHgmOXjhxrIXopTO0YYF
kATYu8X/QOK7vXN9Ft+mnb223WaMbi4I+69Vxaij5bvQ0GKFDADgEEAh2PrT8PiT
r0DU9o9dUW3iq/0lSHyrgQSLXBvA3tuShEBPqdaeY7iNrcO72BoC0hTxmb0Dr8ED
RY02dtWZwg3++F+l8R9XKPQCj0iLDdVIHcgVqdAJEdQOoT84h5O1akyHDKp3XMmE
OCgvDuP3zO+2y9Q2EYgrJ2iYx/C+58vWkIk6JQRUUPFheY4s9Lz7nD0yCWTkNvd9
Z8Wv2DFcg9VeMF2tkR557Moov/FJLv1NU9kYOyhbgy7GGfp6e95bRDiDzhGcttf9
dTO6mNmp0z7R1WuSJX/fd0gjtdeggo7Tl+LpnltwCqjGseKo9/6oq1eiTRNk5O8t
t5R1OTHInXDWNNPTgPiP0d4xH2TFeurHAT+YZZ4YGFY21Mn0A74/2ap46NCgoZPk
HgV9ujKFsxh8V3bt/eiZI0jrIi4DbvdHaDbaawMYYj74MNv29vSjymdjCmn3jSva
//+mkr/rcX3Jq7kFGx+gThwomHz0DzLnYo7QYmWwrL0vx8rXbmOH1bjiOg5MXFqp
trJ7xt8vxjGeq5TjtusY4sWbhBxat3ELveSHkxXNwJz7NSLqL2IWjIVs2mCdWsEs
N/tiRCw6k/UnNjkZw+kPpfe1I988FelQuoSsROdH+pf//e7srfJJ19xqR6ddwujR
c9wnAj72P8h+s7Iff3FWPGeOvfSiOyrJogASJA6B9q5xeFH/QObW+emYICxJYlco
R7XgcRaXvFYvdbtHixoIvNX/BqI5UZcA07R+p0Zexewt3H5vlLROXmPUMZ8yyUhX
cK4q1Qpl+KmvrY74muoARTffyt7TFhiKLU+U4djcKg3f8fpnYWW+cVN0aMw3Q9T+
XHbinlgxKYlRzYyDuhve+DcdDaggPFlQxxAsgjJ+QV4wSyzjyzqR1RZVp1R2qSys
a4JJNceoyYLG6l5NYsfsah64R0o7zkFYPcawFRMWmlhPpHhE0QBH7H8n9SK+J2B7
zAPhPY/JRkvvddXW65xeGGVNXIhyfWefvIATgl8ycxWntPRU/CrI3pHot+QmHa4N
AyUDJgqJ8NzK9vz9TbqPHJdqMNl4JbS/1k4cHCw9G/jlEsuEyTOEv3UWmhjB9Xla
RyWcfHDj0cAHGAfPbLLJNDOOUOk5jufP7vMoTXir4+nM7iQaWLo0ET6uGsipMgX9
Qyv3Mg2PTQscP+d+A4PgyqTMjGKWH0N9L7LnRhII1ZJvGfvyR8Iam4TbZhm8vusU
RDl+5XlW5FdabA/rHBYOxY8ZK6Rn2u4r/GJlzgJPUqiwanIv+sIHtPDdxCgprvcF
vMN3vtdrATOWG1g4cKNbI46Z9DPaik8Jz0fro3EOTi9XHXReM1HHx6XOCGT3f0jf
tL5WuiLEJUEk3cZVDeSSZSi5kW5fdVKp2vXVXqOk6iiOKTtQAtrdLqkBCJ/sxRb+
A2K+KmtHcBy5O0XVJ6I5Ah3Njdq0zOpGSWIedyP1Lo6DDCmcPNBFOx41NmjyLLtY
P8jG5yLYKNkhxwRGhE2ClOE+Ss+aN9lU0eRq8A11RnFFwEZnRtKOmZmbBGIbqit2
z/sLm7m8nfy3Sj+TmpTXqgi44vP/rkFYxDsFzFfIEKrwf7H7g3Qgy45ioX8rDHLm
OU0j10UwhJn7kHEExpa7vVuOtzoJtbFulvab/tiaMjCbtA03iq38LfBXf5DRPNnW
DBpH28/So1ruIoqWzMzKUZkNaN1mszXoOItR7vArvvFJT87p20Z4HfnI+XNYwePx
/yVUtiHR5DumxyvzdubFihWZ3ZxMqETP66dHRP1UYXgnp3JnBwu4J0MNnXvJuTpf
ZHVFPZfSYD/cs/GKUy5szkrqsW1QiP4+DGTcEDDCJvtLl+tgsqAp9+UXIvk0Mj8r
PlRc86hii01MSUOnjgW5TlEOARqJ9ANnuaeOoNxMu4s=
`pragma protect end_protected

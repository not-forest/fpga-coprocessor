// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
dAQBUmYa9LRLadjlhX9hdy5uzcRkLvmWixUyoGOgWlZfIFFww2C/lYwNvJl78BWa
9q/BlFKSWVbhwc4lIL4Smf22XkzweWf5i5C+S1RhcKIO1sGmIrUn0TQqdjvbxeeH
X601C6ssfdLNN2AbPprB9RJTC/OV1RJPmG5IVW/b/ROIHA2X9008kjFPyDIroprA
jLCKo78QXaeOetu1+r5mBGgIE53fQwH46hdUKrCxpWOWJlt9MII6EHyqisw9PSx3
UlH6xoPEg6qM6JOZw1BYKL4j4JK2OXTpXunipKVzTeUVQugjMRp9/qrDboZX3iGh
P6OCkO6axTlh2zKsb7BMqw==
//pragma protect end_key_block
//pragma protect digest_block
LiaOIuLMYQDZAb4CXffFe1xjA9s=
//pragma protect end_digest_block
//pragma protect data_block
OkcTbQAEth6pfDvXmJpUO9PU6JwXZnhFlvTFozuGy0lNhp9M7+DannWy6+jlYOdc
7SgKczJN8m1ROJX9hluLAz5qIy3UKaeGj0Rfd/UrQroTvGmzV0qovYFZQ3zUjicL
a1sTNf55j9MjcBytmaqgjBrd+SaHWPybm4EKhhRdhLOfQRcWvjZsi6TlNyxJWaMU
HOY6qBTbJ5pHuOmLzg7t2sOWC2kholsCDUCr8alcOELTqe7+vl3ArFG8peuzbulY
xxUkdhrb/e/MAGKs7DnECGK1kFiuf8Nh5zp9AdtxNnJPTKaUcL3A7nLHoJe9aEfg
OQsj1zpJwvUZ9XqFd3bUy2UhWA5W/SfPyBo9O8HgruCMbDwrt6jcsC/1BgI0KGO0
EWF7SfvQ5SCpX6D1zmLZLfNEgHdq/ZwRlAh6KU4/FKWvP5FPivKE6yOJfw11Vaxh
guYh8Jc179dedZL7d7wkofepH9q0JQ+Lp787ZOBFmaMsVPDKNO6779cCNsOQYtP3
b5O2bUVMuNv6dzJKGRtmSpL7ogncw1EvHV2g8UJ7wRfziKW5fu9bSLhLQ0QRnGnR
Kq/yG2+62T3Xb71jmrXH28HycDOQO2FTn+h8id6BMp5TOaDidqZe73T4m+ykrXYA
zCpz40hlfhAuSyTTI0fKAlxTGe3Nw6os+UM7zmLMNY8sqy5mUx29fqDjm1oyP6xI
2EOOqZ3eD5PwbdLehKbJNdzODorVDlIceWEk+ZHrMNUiuwF8j6CQDixHkgeXlv0V
nKEfXkK4LTXoEVu0F4qRO6BVMHr9pfZEZ8SRph8XEF3YSrsWWU4pDcwLl6gu8VyB
fE5E0NNHT0arL6Oumoy1WDn9Ne+smVgTP8VSV8hpHr/OQxsZreAw7J8y5c4YuEDN
rI88lXLTgcKBhEYIYYDodP3KLMhH4vXhccYYhH9WGlBLK7ITuL5m1h6+5zGXiwN/
ztfTIOUFwH0TYsJ/2offTMKFLra+L6p+jsEwpR/8z0FxKgoiknrhwZ+QVRYPvZXS
bdd7H/udU0PBv83XrVTaaoCPPrzQmVG5jG2V/3ucpogKXsNHPrJInqBCM95FshMd
43No9GAZEDisj52dw+ACdQ6U9wKclLanf6tFbV6Aa0ADHMj/KZDHWtHwjSrjkqa7
qsxdrjgeR/yoG+ws0RfR0BPgk1tAEkUsli0NpZcdm7fcTUQe+AGZiS43fYrzfM6q
v3/FT2i7SKbe+B+C8NqA/4udCJLHRmH2X03w9AgW8VGdUMlkcXKRisgQXR0woUiZ
gK+vJXMCCpy72JslMMdlWoziXdJaKc6OcwgGnBsl9nuDToa5vE3NOKbua9jeiCfO
3C97b4uqklgmbnO0KrkwXj1EddA8orAPgsBMiKN0sHsQWaGIYBOhNH1LPJ8vVf1X
W12So+dJFcTm3Jmd/B6V2zoctipCdrzwCyBaeE1s9l64jZCLj+q4SAflyxtRrte6
irXcUpu/2zq1TuDPgc5VLL16c4WjxKfNxKSfjmvqhebvnLGsmH3hHJ5q99VE+KAS
rGcFGX0Kwu6LZBN5DPcMlI1nDF6EMGfN9Msk9Y1+Oh3RO/USlifkzPUTlJ6Txeyk
vinfJsYVs3l9GVbVnD2VF8KJkHI1gPXPUCP7AYlsq1ZN9WP7mAPSP3dY8/Ddll+O
YMxYuo0OEeGdubVm0Gb+XKfcrC+aDCHXYE9gsUUu569nZWz5GFXQ5VgsLINugQxU
NGu5yGeenQMOylfuPcTfMkKdev7fy1Y9YA6Rikd5Cx5ESdkS2qv+scGwWVa44dsl
vM9Xf4WD6/j47DpdrCbrS1/itwYF20hwbcR6TK7x7+mh2ypphMMbqdiUpvrizxQl
CiOzesTVmZcAGJTSP5oMqgRP5OD5xh/+WUX/crl7VvdEyDhqV9RUNcI6YtpKEdPN
bpEenlbAho6LHaftnZn30yCemystLRwyPNHD3lhmqpSIYSRyUnncHnx8OGcEjKoW
pbTvig2saEw7qCSWN0zBefuewrV/AiyHNvdHXW0SsrxJuRXIzZHR2GqctOIGD9+A
gyNuulaOn4a7NNxbeisp2NKkdvD9woDka+mxf/wP5OZGvqQnv2s4KGuSClavT+SM
ClAB9oPkOIJkmMOnpyoKFzEOW5xxrAZk7L3HrERFxaspkgDQYFw6u/5E8pM4/sA6
XWpn0NXuNAYC2ltJqITxlpHi8H7I6rcUVqvsJ2zXX+RJfSr0l9KqHb7Q3Q1uTBqx
BOajqNfQ82Z74rrkocCqN4i89FCNki9MeBlcH3tv84l8ebwOBo2bs75i32SQNCcq
A3ZKFTP8xaQ92IHzYqfyMBVtCenIVupabOFDVWZ3YXj0OsTkVkq1FMmCUaPQDjBH
FQUhZNmzebaSPPQA1TGusQ4ZYiujEU/d+ZgodVebpVlKX2QnsitkRGc4NlrKbDMt
xxfKeSkLdfBGjyx23CsP3fnZERwCi43QgWBm9NUnonrq7gT2dYgtbdLMkl/y2pVR
jtHYljiWZzl54dix6OWmiDfkbW+6KhIxvZ72lJ3uRHHFepJ9g35JbIBfI/errSvI
J8ZOH2bS3LdwJlfhuOuxCf9NLQoq5xRIX5Gi3AoFuUuKm5RG0Rk/m3XfuzhgNH8h
0sXInkasGY4PbzpghYKzJCLsxAsK+alNghp6yD0cVWA5GGswDBj3ucfx8Q3v59hQ
CXM9tH/qr6SApZX0J9iDyapb1wcSG2Ub/LGAd7YQ1hGF7uo6tusOb2pcpjVp/9Y+
2GKtvBDVaHI99OQuPaUvEHPsnsWJlMRAvQGNi8T9MhWnSmf+NDuIdN660OLfgbeq
YPjNtjspBGrgPrF//NNEhdmq8Fm2HLyZ9a7G/iUVmI4ncE7hW0UYjei5BXJBmtzq
aFh8tby9pzxEII5VW+OloRZ2XVxB8MuUZz+Z5iQE3u2r/viSIAXRrKO36PUEcwDj
y+51yW1FqZAi7k8fFbDwjcY8PwHjwEq7mC2oIT6XotroAmkM91adl6cgayxOi88y
KJYpfOqbU6OlfFgLZCxy17XTFiH1DB+ALxyTf6a+SxKIgIPYu8U4vTVLUlBakq/w
ZAJksz/I8hepmlyiGstm6m+q47bOiA+DPOf63gH4d3h5kgRs1Cang89cV+3GYzMs
CBKEDDYulk2F2xEXPS/NftRpr7kcvjm/yOq5RkioSf79w0QSKi9PJHQyr/1zkDiR
xPqZHZPo5LmAZk4f4aE+ggufXAR6sbgME45roCeiI6VaY/E3aKOph4H5m6Cwi4aP
1LQNkdTiOcsik3Scyt2agOQEnEhDIVCdTy5EsM1SjtdwzKDwJYpVK1jxI2ftIO6V
KrHKWfbt+U/9UJ5bdXikAB05kwcSUMz4sHLZeXZCsq+C0J/C3ucIoT8XWM638uTs
xNn2UImNM/FVyyAY7SedeEC9vNw50aPVsAy1vKNbBowY2XOcfFZL1JBQnLnIm2AO
CrU6EkyzL/I/9BE/iF/exLLlfxLekKWNpV1sTXSiAebdYazeDFJmeC+RAlWBBzeP
+24VUNSj9MY5uPtVykar/IKRQgeJl650wJSRHSf8pbRDBcIVi4otC3u1zyDSLshx
rM4dlU8kxPXEz40xdMLxiH9skrAy1FdFEJMiOkBmnqApd0gD9fiHf06imaz7rLAz
soSIhJ4Nzs5FuEwiIR9bksZBnSadMFarW/AJAkdSIpg9NqprP0/bEXelta+eDcRm
LmvJOpWjpwxz7Keqv2fASEUhunsNBwvZcnE9gTVBoRcEiytIq+g5bnsDo/UsWwQs
PLZRAT10zsGBS/pjO7/avUgH7MYbjhgPret1wUtPx6zfs313fxRNlBVQOAOCGFV4
MCxFMxCNEhojC6rIoiyj//cvh7J8flz+uojgRMp13wb+OBaZPvVryFBRuvNydN8l
l6zSjECz0KomR+8ObOLKRqOUX/xopnvB8eATHacHkMnLFsU/OB1kmff6SvLCEuLS
ya9bbUDdCEmJleRubDOz0tJa4pQsnFLPDMe/2NIlROI04K5M+dpCjCDeYqnrysNk
m/yMZm5k7J5vhERdez5qo2NgAszSKNexIzzRouu8RYrvrJLJ0+hEe4IlVZEzM1Sf
0Bt8EBX8ZX0FrxYMjNKDIlxgNiMGNICXQdBapKes0wQtWgFANOjXK1nMQolTfjx6
z0CuitYtrYQs59cAdwy7eQcqRTiUDVA+3s+LqkFCQpmFOVQhYZ9g/rv+OZPTOnNd
eiYx7NxamwaXE6B+MaG4NkNKwudXnnFsh+w6dly6ij8fRSU5lwOK9DvDJrKb/u0K
YBoJ6TGy+hecwiomCCKQYLZZiELI/C9prOE3laisiBAbq+z6J28+wfcu7XK6s82B
81z2+k+9ZKbMBvO+KelHF/YMJBPecDg7O41RSBgzxJJ6eRWe1+9FXndge0tjsQmt
gPrSxJBjCJAfrVuplxLD1R29JxPdhXsow3qgTleKQNQA28Hl/9rW0df3c3FRFGZa
Q2wQrddIBd1z8qkTFvpEHU1YGl5xmCRRYETc2LPf2D6r4bUjgD3v1H5aYTJ4dHOY
5uz24KkPPlZzxmo75Mtb6r4G7c37yEl86jBmcY8K+YPJgVsX/PIRpNdreKGRhWx9
eJmkqUjQGdCRWjTL9WjPosTvw9iVJ7y/D8i92Kl7pndtXJoq41cMduQomm0MwbcY
bKaNVO/WDGIHb4yvGUviKd2wYlyOn2dv4dR2AE3nOTm6GwalUD0oUEgv4koWkGUv
Z13t9TQ1RxO5qRb7gXPx7WIB/h2AW98+s+cJdOz1QPabG1FDbupKgwpI2nXDo2x1
m08IcmDOSAfRHHBQcH3s4Cbq0Cp1rwlnAOJppCIsEw4Ad4pjgHIpoEvwB815Y64z
zRZdjGss61Hay5lbEsTbmtN9FOWOUv46vzYCRx/2mOjl7pFyV3EXcyy5z+rkxL8w
lgQJSVwhlJ25Wt3jSkXXW8kWLk2kQMIQlJwecJ9Qv++F3P0Xtj969olXAM1t67E2
QqYjuZPeRMY5r0lBhb+t7b/bGammkDAdYomP9YfQXc78vzN07tfLZLCWhyICrF3R
DChEd1SSCq7ZuBjiTjO0ZKL2yu6m3e75EHLQs08l73iz6im7zmVSW+cAtNsx0S9i
iCRnaQzq9tu/2NfzJVXUaZPQi3gCPA1CiUc5dWEKByk3v2b3lPyRndOknVeAnPK+
07qd+H1ojTMHjwgT3og6r5yNyM00oeGOjupehnA1Sgb7TRAPqUa22MXf3CC75tlJ
TFkl4QA6Pr9W8fF7s04CFzBFgNWZ674aH5Nkpj3XqrQ2Hr8yDxxq4I4Es9tKAQey
SDQuwiXb0wqaZk3FLeDCca+X/Qt7le1f3Y/FKBslbffgA3df6575OWphjYl9oF3X
xcSxRdS+WMMTPnn/uk8i9xTwpWR+nuZazJyNtL7OOvfJegdF1gwoQ+okdeZc9nwi
p19RZiMicbnOjglNIdyAWWxxQeQUZftL6CujgjSB8srdWozWHEoEAUVA2G0rAsot
NzJPVSIhoTHDVTtYvco7ONTXF811QAOCqwW+tG7bqNzlNFJpuRFAvmqV05saxke2
Qvy3+ZnAa4jyJdIa+J6p8Pl44w72yVMUNafyOvuGAOgSK/di8tmLMmgmiA7qnpxH
CDQV1egIxV1CD2Pzzqqie2GlwLvfXSHtdofcn2CD3DHmh1B6Y5zHZpa5lmlGRzzb
vG9d3L2oowAvYVrbC+zt0QzwPBOqgf0x0RAn0IkcimxzQYyTyTu5eUrRoHrLQIP2
kNcCJxAEEoHr0QDFKcmSUIKpcPEHY67F0mSCGnlTkfH0Wx2naQ7I0z1hdoeOXH4F
5sIUlUSt82PR3MywT8nyAMRozXGNRz6k/FpT3h3aNKU+S0oxVlkIJ4XoUP41i35B
cWz2zpiq6VkpzqwKCHjEm1NfGIO0PdXKvJRt5Em3sxztnvxmUFdwCaVzLsln5LOZ
cVENeyo+4RaeshfN5WBzb+m7LWLMBDzgPIDLJwk5pd7R+NjDTKq/S/d+fhVJM38i
ve2rCIAs2o2TVTH00NH2CG0Hm5zhl7/KbH7I59KWSyso8yfRvbCzuuhUBHQakdSk
rH49dD2d4U0lVsAyqmjTrwJmjkleq4MoN3IBpSQXKuSjIsswIgLyMcD8TfYC2zEx
eVs/VGRwgvTB6+fl1UJUSH3d2FXmzVTP18AFiPx4XHJPgLxJQh04kf3Xb4+oPTN6
VB27QDgp2N9WlqUF8QJf92Hi1T9noBW7vIGO7Z2bAKsj31EGG9QTv/rlS5gf/RkG
Lxt1N9ROV9awt7gKLEpY7duvO37KP2RP6yWxAAGGAuQ84C5dC4SgWxJzaVtYEcHk
eOE+7ndiuzOAEYZ0xuwRHvmHOmDn3+bl2Nb+FlISWaj1zQOxmX9UGz44nDeaDg8F
uobfKO/iHKDi4FZURq/NN+qvPdGSIR7toawI6tN4JbGWxWHwgRgOXlsXyBSgVG5a
3is4gKLrMhqcPtmPseoKYc+17FNWljWf/q7z1q/QK8phR2G9SixGKAeDRZytRR2Q
cTKCYKEw/R9Yhhrlvlq3OfI4GydgQ/sYHP/o8IhFBYtXFKIxhIsg+V/Tdsp9a90X
u1fNy5mflZflYR6qrQ9FBOsIw/nUwpWRTjJh+JZHXlE8/LlARjsPdT03vtAhN/DG
Np0LCFt+lhZ+bcl8xn6ATMVI7ewSg0OOxqMexNTx7M+oXpMhsCP11hBLLpoZnLb8
zji9MuFu2JiORVHGUnnbMuD6cloWmtfnpki5xg3BMno4DQ5EmOReGEORg83qSx5A
+O8lvOXIxPAolrk8i2qjMbiIZKGn8ebFbvvFtRe/UmBS9JsrO3MDtcimoQe1T9K3
cDAHev/3CIAsKHVJ14fdV6TeRRRccSXrhFI6dtVbWudaqvEM9T6CPW6XFCk0S/Q+
4HwA/GlgKtnFLEJ2Hq4gEHll8nNtO0WGrh4J+tngRi/yVdEkBqZ4v+cRY/J45Nkm
BxLPr8dXhvlwDykAU4nPorFeCUAGgfJvqqW2ca2fDV5c+eypR91MzJCODqcU2P5C
CVM1eDMw6sjMP+bPU/ZGyQJhTSbYzfVMve7gkkGYgREv4rIS65U2B8n9dvDCXTZE
UZF/2cQmQNWHtIp8aI9S0JUOgvKRE7nMIDLByhU3gUrRWJlhpwSy0nBVMFxryivc
c0lLtqFMCdmAXRCK/QNF3oXgR+s9jNFfN+EoE5oQFpG3HlcuChKHypGa1W1NDt+Y
n0AMtujc3b18UJOvsl1qX+307etOen+8gL6XTrq85qL2pkVaC1J3T1VxoB3MS+4x
k7W+2wWl+khbBWbL90Byd+WNQEa5+sOsRPTWcw1N7txQi3vhsBsGkt4JQt3W6lL3
TvnVZ4L4q1CLI1+g8oaXl+PJD2u4SCPoz6EIjkWeC34C3OhImUKL7Qa+F3AlWRZS
d0at6mEX1y0Qqrxt/8XssqIhqzWpzq4+XjBuD4rB3L9uLUETMi2WXNsXr9jp7fGj
uHduRwM42apBL3topeOy8Zjt31evcZUp3rGn2iDa/lu+uaJNU4EQXnlwemSU+A/e
WMSpaqBXyNqRdf7M1R8eWqI3rv9+idf2Uqj3bBd7kyh8Ay8BLGR1hbenLFhXG8ZL
3cqDbZoZkPTBsL3uqj20COiRQTZ36EpbyM/brQQnS1Z2EmrJ7zrzDxIpWKTJgIqW
EBzUUsGJ7CRPE2Aae4K2ApzvNFeZ9EHKDDbDSrv8RQH89c+XecU3JQLAWjSN+6pq
lfoMzBRNP3QqVxf77pfv/azzTnHYY/UqGlGeLe/1iPfZt8lDD7YfjncZ/WWF8Ewg
JsbfxH3eqVvdul7LpyH603frwHaoZZrBgPkrAA6tutPSTkQBiHZz0aPUdfvQSGP4
VfFhlPJBl1y0Em+rATWrnOwKALS4JhfeKobmCVP9r1tzi6B1N+kH98uB7vnuuzrZ
Gx+YcHbP6rWgy6toJ8Bq5cyFwKRkOncx9LzEqF1tor7/r/ZNNGis069175z01UQk
CeopPcafCQ9dtLKojC4VJq3hh7Ed6yZjkNerw1qKpXUpFwagUBagnBgC8YarO1jN
GCv0rarxdZRlhujkM+ujbXq7WTPG+uLlMQGEgz0OrUSNJ4UsrP0zUPeEhEjQ1BRx
L26IkkbXztnWQNm22r2nm+yLfEvot3rjuwqdNi8h9ZPbBgEDikv7RJNfhg7LWfRW
qSGsSOmwecPP/OOSa59SAkbXwgVsKtGQhChEnuavl6+ngaFZFDEohWVd6OWU9shf
XZc8EFpMrRW0+ot+6xOYMzIoOXeiknBw9DMCbT/93Pg8ihHcVMFRiQ4fjdiMzBa+
azhPjdc7/0O3A/k6lIOqwrpTDhTuxEwqLxh16bjw7DfqE0i2NkrjF/xsOzrsgzhS
AM81jN19ad39eNsg4jfVzsCVhZUSLy9/YSpj7D+PfqFY1dTyGtlnqhwPCY9O2NZg
nQwKA2uwAb+csM59w66Cp1u4Z3TO56NRly2PwKiO0j+QtO50i1MAzuFMs/btpeyw
rmFtsSpLxMXrETdcs9FMca6ZpvefkK/OT4yDNOJq6SfX4ffPeLomvKxwrUdjyFA3
24g0n7l1woT5IMn1soO7wxj4aIVzRQ6QT/d4KBgvDi3EiXwHRSxbBnefNn5zaPeU
mo0kny0T0lHIrIJff1r2PSYSGZxbJfCf4PNaFEUCh4eHlFupn078JcDDsSuuXRMn
QnBHUnCKja+sy+iadDsbXTvaHnnIRnbikmumxbcaqDwKnj1nERYKNiCQzHNHTBDB
hQRC6ZIEA/Eb72ZiZKRqzeBGwtHPA31DxAsMMcvd3IfKwoCd/gpcMxyNug8gWsDv
5AqanqsdC+pbPHGRJ7wCN4BsUHDy/DHUL6kdob9mI0MmqVMV4lhUaBzDvt931QX9
ms/i8j5286NoBeV+mUVI5dGml7bmOLuEkrAJ84VrsMZtyJXVRu6kSlbUTPxUjocj
n35DKW1D7K8qDm+AxpJW7E2iqx81eLdEnhLYDLyrZ2HPwwWrCst3TLRsRUs8IE08
+ydNWrsomhB4lEIBi1LG5AwkKk/VQaN/yw3h7PPCroNcJJ0ppnApqhqgyQR+cskb
bruxPkL9um2GnwGs4rrnF/8aztI5g/TydFIUcSbMCr15iT/8Kc/JRFIhpsB9rtzb
l3POsnGOe9c8ly8SVbzTAqzpvDMwN4L9ZKtJkZN9bNCRBa4KMKkrk+YgLIgcgpKR
jXHzqb2JSsVDJHRG00tp6robxyvvYEP/xn0KHucRIJHTsPRWZPTe7LkKdjfZEZzC
hZ8ElhedhbGJ71tKkG0D9USXeYLsX4xF89YXNmGcQkylS5n5WwPeb+Y4LWHjbXTO
Rc5mwO7Z449ZgPBcVvO2ZZxfZmQ+YnU0TIViIh1yEAiTWWlB79GjFjmF3FGI0qGQ
t4aLbwpurTjAtwVII4F/a6HOpl3BSvwfZfH0tmxsM2QfVl9ZrEGuY5qY5hb71R/D
e3onZKAVqK3szfYJHSvekQWD+gfA8c+4gPkOJ9Uc1sLZhU9lhpsIU2+Ms2k4kEFr
i2XXYeWN2Duk9Kbm9ArxLyqGFdheyWK0muoDg5UE2Zmj0nRHhareF2UFHjritrIY
H9Shf6UFPe5UIrkCZttqP//cXtuXzyHSVr6IyCghdiGagPEDjxHJ0rjFFidB1jqP
nvF4rw2efjW/Kqtw1tif8w0RBbZG+nhXLzXHASGngx2JdsbPcBbrdqOW+Xa68hqF
AEFHzEfy3IJRD9KGGSVVUTJ933UoPIuJW4S0EyavnixlKbbTijkaeBPQut44fyzw
Q7biuCtNPsREC3UZ2mFbrmdTNJkPMvmdczM7Mn9YyqfBHilfK25Yc7jf+ycrZty4
qXPcf6SQl/coHmE7qV4eO9V8awLUKC7htW61s44ahbodgcrG+9UXAnPP4UXs0R3I
CINR+JZ79HZJePjsy0dCv6yQPgnq0xY6roii2E9Gp/xVcHK0fF6FZSzrGohf1q8U
luDXRTgC4CfKj4O+O33pdN/of6hhDvcpB/ptYWJcHj87lc2Z3JYlIrm+1e0tsrc6
fxHxhweqGCBNNt0xIxwe5VYSDo1ZnNQ7QWpdfAbnE4j9yUQL7COWiGJLeWw5xWSn
cq8NTXSo1Ukzdn4rMZwjTzlMy8QNKuoln7mK+9LQbaycwK4sUzcLZ3Qmpw6AMBdT
AmEBzg9KJUMI0EbRteZ9ckcSxpBtEwfajT+PcTFO3fF/vxOKakrCyFh+LqsSnV08
1fVi/h2bdmfUX69wsD+eb1xko2O0a5x2nqoRZU8Yb0RfaBZRWqRSp3AAKduRzwTY
YOTJJjI3y6X+LhIiBgownwupNZixjLuWvrvwx9uxqaKB5tJ7IV39X7sjZa2Jf1E9
HeJQw8RWzcjrWhATKfxioJS9HUtty+J2mxmIvKl5Deck64oxcOfaYIhrK5y7H95A
OBuXLuhGmVf+FpmOSCQ9kPPMW6XkJ63zlpbsVJ2GMHjd0Kl/QLUDEP5bNgyQMAJc
xdT5riRSp+LxPQpvMAgA/vWDow4oznc91nRbRHATtYaqg1K+zT+nBdbgjQVBo4yX
9D+H3QOcCy39Iobs/wOe/wjvP7QC0Ln5otY2/nIGg71oE3zhXAtELi2bQDdQ5iNu
9pXEPp2lypPFDdmAG//vN6mqSVC+xQ1nAXW84qhiOa3vMThIZhl8NdyRh26iaJBt
+GUSpFOU9w2nGGiow4Ng6grGn+M9uzTWr/Vpx+WmnBLtGvu7pv54uzgcQMu6z2dG
TCNXvUcGnoghLqvoTVsbebr8GCo3f7SRyGvyoYSZSJ8Kvvkn5y0mQ39N9QfV9uW2
AP98ikNMh+RUp5CTRJZEJ4xxiUz0+gGK1Xc08hnV+vau9kRUvpn3U4DE+y8Ue+pT
VfEiJ4JbCs4WMUhQPdmBUXElO76o4Niz2gwBdGeTu1Cvb6zK3ePg63GBUfc3D6Rs
rXs7P3UD4ov+dTl3gdR1QE+aoax+Qs6LslONi8K5PgrIrQ43yhW67LSo1ZdiBAwV
VaMC8RS9O0FHtn8ZQp7eB67broZ1nKivGFtVg8mECnSVc4dSrZSckapOXgehRMUn
3b3nQ7uWgto/ZKkS9aTRv7TVAMQoMDmsX2HJpcntKUdCmAl2JFRKM8aV5o1IvUlv
nPXXv3DInKi+M8130E8/JhPHWTX3a4ZmHStQ793GpvLuF9agTLfVhchSxEY4PJsX
7BOL8BXm75REYNRThtfgtT755eXxx5eQr5yyDrzfQUcHHC0bLbMLMXdw00eb/njO
zva8iYlkUUWWqlVeKAivPL+lb8piwUZFUTne4ufhNuc4PHHcqKzOJv3YafKjMdsB
sO0q2+oNQQeJLasJX1Go/EQLqjz+y6znk79b4STnNc+jiFPLuP73OxbkpYd0uwPU
5Us7Jp9Quz3zJiRn+SaIKnIGRvFiQEHWAFJsegijHusgoQA0ZDYpW02g51OFZexc
GGhRLF8QltLV3dSTrBVTmh91Zfgs+gNYkwFGxGL1MbHYX0uAgzoB9OvoaM52QdRa
DFCNaU1BGEua2iEAueCT27rGH0pFH3Tikc9v5RnMAYqNPYPb4cJbXRWZfwpZyWOc
hmqRwu1wFll2Nasn2ptnS9OxDbIRuwv3IokWoGV03xlI0evusL0ks2b+Seac4+Fx
qy8Gcbep+FH3H/xGaJLmPZc2gsLGj9VsCauZ5rhrPE6Ve1LxqGnzqpYUURVJEupo
7l2hAgtWpZ+miIkjryTzpa82dFTnFEzqpzdY5OUe4Syf3g1flz5hOHpPPFu/MA40
dhj7oVzwu95ADpMzsmN/0zjAyunUwj9knSNt4wKp7BL0qyS0TyLrMZgz5YtDQYT5
xYfHAfBpYREGZIyTACURuPwse65ObTNVWWzQDrPpvTuQFOr873Efg30dvazasQOH
k4akrj47KYWfhAIaGN/5rT5cHVTs1mcw6w9IamS/Nntj7CmcpPNo/80qUiAWlw7V
+7ljSDseQht+9hoSEydnj2oBmekyxuPjSL+xQZGRPi3gGzbAgCWqYt+kBu27orVA
OJV3gDGC8JsItHZbLuVY+8OtA43AxqnTjVXTv5toeQS88CrhCxJDx0QDVAjJmJdT
XF9uGMgkcmWAmJhU/PgixSdysmSV9xO+rLeAZNbrVgp3+xv5cD/xxxDFmlKe3Q1S
SWFShkmpjj276GGb8SkQctavQY9vzmFqT7k+rZYA+zAKKc0uIFqCesCrZemNsgmG
WUfYGKi6uo6tcw/89dr8/qWpXKHLQDGJMRPE7gxPd4IjoBnF4D/Ry1UJRJA9D4PM
elt1iIK5b/4UGohizDoQ5y1W6O6O2cyaivc2akG/oqczzVRn5W7wilwM/Y7kI3Ov
hUtR+XfV65I5DBarR+Qm6+5AefMrcuA6HOcLeLUvpCV15x17b1SZYsD0tLrRpt0u
qSWg2v8vB/EzflqH4MReCLAcowcg+blt0z1s2pOrR7otHdOZ3N34HPxcoWy70GrA
G3CkjgWmHtC/1ZfNBTSfMj3kjBiX5SJVIrFZgmycvTMq1UpAyz/0fgz4Gvo1pyrm
M7q6eLn3H5Q6FpuOg+D2WVeCtuGWWnmbOb0YIrBgXuW01yxZezwgzhsIRIXmkNuA
LrqAr5zM02euaiJ2XNkbG6EqvM6fSVD9qRRGLJjTWRaksHbPEB8AiB2dcZcWTLN3
oluFsxvGoQ+moEaJiu7sb8cm8kYN+Db+g6PNhJ+41VTSHwZJymVppkLmth0Gc+83
s4oZYCOF9B9iP9a1LJdoOVJz20beUjIeWaH3KNZxrKdoi0+GCrj122mfApcf3SBB
Pt8psw6GPA09SIpmsE0VIMqC1/lZCvKuMHOMOm11yPEq4ExLYrDzhOVBlSV0q8GH
dlndNauejzoADi6iN0c96mNsnL9xXbJj5A7K02c7WxHVSaBC3W6aMNhe7MxIafoe
eqqlHlBMeOwHMlgAuwLBTbwAujiMuc1eWyYETKUIBFRxCCpTeMeYMd317HUtIilr
CPho+mPY465teCaJTqpaNUcepxAmSPsZxvK1QrSh3JBOKQjSq9bujwMuj4Jy8O3L
fwHb/Hki7YP2lPKLLCN0qoehsC2aL2IzU/WQGJzvmnbM5cZvkGudqc0qIAojddWz
isdwybNBKhkxCqf1yZaPDeHUT9zgew2S7V2s87LmONg+gk3JZc1yuxsqHvZ41Px5
bUlEOQsvHUqZKJejWc1pZhIY9hb5pVSTzv6GzdV7BnwLM2oj6ovC1PJfA4leQVmS
1nyHXD7oXS6rMf+RRhV0Fd7t3x2uoFJlORsenqf0ylkXp+Ru5vD1pFXPdWA/NJQ0
Ra0mIcdBM0Sj611d5rY5otCXrgY+ezuMb3BjF5trkPWbPfQflFh4QzgYEGCJv9PO
9nfYHN2GGrZGFOEgxOqYQYhngCyZ9Kto/vX2BncjyJkWVl5lN+jUerh7tJzKWyY+
TrnzpsnKIA4GEzzERZJLOQYWxu3QHTVNZwUvNmKNhX0ukrx4QHxFB07+r2HsrbJg
ta2Pt4pAlxK1tVL4zPaCMrrQIs+pP7YkGTvSanjIXc4XEflibghcBTuSvw3SNCUT
YxHBmC1CfFlnioXk4h53U4NLATo7lG+h5Ukf5mgNQw4TBYRQ7WWjNX2QIUqLo2Bt
HLFSNG/bEz98QYaX293+rpL/KHPhnv/kkq99S1oKCaw1tZ1CpY/MER93arVOwO+W
KByh+zIR5KoyjlvFdhpX3F2VT4ANg3veyNvvYN8hEzwzAQvUpxMgvwNS4+QTCEfy
D15Q8h3FzvdgeBkBjKPlm7jV/u7PF0Vjf2azCX6p7yBHjtJbxuhi7Zlfvi9XMpd5
r9Q/H67zVGxTlGWco9nt+G33u5mbH6hVZ51w/VsBbtHN+KMTYbhUfDIvNof8qA+U
Mtw/CFmvgNUa4TfHw5smRy4eI7hlK8SKGzrWCv7UxHiCVnU9lkWLF6lW04qGaId3
j8Ckm4ktq10KaDlNrkoFcYFgweao7gMFU+8hehnMbYBzf1p1fR9+cranTT5ZpFes
BKI1hqo6C6HETzjO4qY3yMv4lKArbCcp5D/+OUcocpEMUZyCsvHzSHT+ez8+kkfG
xJz54HrEzkwKsNYEGbHDLpsN32I3kpWb87pjfWGO0XWE+U0yNzy9S29oVhEa2os4
6/1GS/MvMTbqV8TQDQJX/yHclPFDJLWnKT1FPKm1laBwNvcxQJc3I6jUcs8Aacu9
mayPnhQKDSPMe7bwY9shlEuRZhftKYeBiDPbsQpMqqfWqiiZ+qAG7F56/zLdcdR2
XNQlqODzrZ6mMVwG3PANeA3pGIkbkyDbFHkczHq35Yr1MVbepmwRBE7cZxpevhbx
+hQq1A3pkqGFHDknwlZVU2OuAScJYmyd+DuPHfnzhs/538fyHrnaRNL6VDanrjzM
yqPLqMWL/47CBoNN9eMDGS8dMBADOBv0qjXpcHCucB0SIH9FvOJUkE6KMpL4SbK5
ZJNsBjPVTgEe47pFToWRzZiUN84p9OzoyJ0QFua//axOswXLWaACI5xHCLx4mt6A
Vr8fB4QbIcxjLFX5jjtorSwhcei+9hL1MK9hNJEVgk108W+wgJE8h9Sjf5Plih3j
QaEGkjFH8/0M/ZodJd+HCVV9uFaLzW+/J5uM85NSp9Stw+nsnv0nNdNZVHqg1SbT
YP9nJ2ucWz0T0lHcrfiWDJk4M09Nhzo0wyoI2QZOOJwpiyajPrCzNAIOpSKKfTMn
5SU0e9WEDpU7EplPRmSEmEN/2ko9yar7OrQ7YIE/P3sPhr/rWEKyxHonVPe0lpXo
G2PK/0oBxCfar4gvUQ0Hdy+FvMgVxZGRm4njjDiAtKggke8qv1jbqv0cVCkka752
Yu03aFy8qrIJTUFUfqABlow7y9/mdkvPL1Ga1PjmEgM299gNK0xtGax0yt2qr3Mx
88uiLnDdm97y11ttuqyYZHC91YHw7GeAGx2JU0BF/2Xmi2DhOZ3GWfCeeaP7QCiK
PBm7dV9xPh6TVE43BWgNJ2NMDqHH2i6F+k8jr81Vzy4NH488xpZtgZ+j12ADaT+J
AKyi3kb0zgV4Y5sdCL1l6kUiOgB+IB/0ohjca5f6lcMHQsx0QZx8dHpu3Ubq0HPI
3Nf4DYp6IGC9QCCq/n7ns67/d+2reaWT9yaKyq0QVh3AxeKhm3TC2FXyqaTwGmDK
uCHeavK7OUAYq3pK7o29gSpN2qPbFxVILHhyzXoCoshnaRGlDeLloe362QD3p/JI
WSU91lVEfZJ98xpnE4Gzb73kDCQ6mitSYx+MUZL9Z74fm2U9V6SlnV/Hwgm/JWXN
s+rfHR07mOKuaH3GqnuhEaC3TximROxtziswF2TTOwZ7ZY13O6rLTt/X1aUtvOaV
sIy2ySHC8AryyskNL8hxxjxp6BEWv99oykYZyH5rW+xphVYKU02b2dqWnsgSUhK8
QDumhNv55HM/vv6cazBZFUZKOUI/x+KOCQKYkMbAl44MRz6BpCWflnej2E6RZ3CK
p0LzDiqBeyn2yaZNhJmQLLcxjRbJ8kNF7kvTh/fnqeqpt0EcaOGlM+u/CB3mAOmZ
edmiLBgGvWIyt+iBX99yyV28YuF1CMPKXeylNt5oUSy9WCu8x9u7Vdu+DdPIxB8L
N61hl2hTN6DzPmWCwRueLA08JlspnjktaeoGoKd2pybJxk0tiobUDDs4ImwQbAWb
ymxWp/FVx6/bOhquPEr2EAGxZ0620Yk4oHaAmNr3ihZGb3SgcE2glR951XVWUXrt
dRGikt7KnGFddzMxO97cDgeXpV0z8nDup4RrQ5PDFNU=
//pragma protect end_data_block
//pragma protect digest_block
Gd29B8nsrKm7qDa85N8x+TaWeNg=
//pragma protect end_digest_block
//pragma protect end_protected

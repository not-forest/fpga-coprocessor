// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
rPmhv7Q5W29HZhULUj/tjtJqy+4CFocNHnCqRYbp6B3Jw9qseFIuy9cqg4LE1U6/HVFaq7SjADfM
85YdC6zf8bo6fgLN9OMiwkcoOqk7TUEKKgzls9GKw0aDaBaAa+NKBNYZDAa1eGMpArYH/0pA1ZHZ
q0yrckCK39Qg/y7LJ71ljRxil27Yw/woQ5tBtQjNusnrwrazhiYFvgtCCBhqmfvPd1IABl6mos/B
5gdP4PCc6clKdpHJ536lmETlX3cBsZ02bojzUCEwLWvoVwcZ10614NuBlspw0mRROgK2L88yB/NG
sllfsNxc9l1KUWasDDo4ymvAnHM2Z36fG8qRgw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 6560)
Aa4m7MdmWdTv+8XDC5gR7vB1egfmY+G5hZxUt6Xb5qpW3rbJ2Unl0scwQX5181L669Kzl8X+SFHq
Gd+tqEQB0jvxGAYDelWtfj6Y6vKSbVZFR6gVp/Qbk8h+sBn0o+nkeSWf7Aq/BqRhz1SWByL9yg4+
WYfF9MQJJPTrbXsllLNgoKswV0UUwQEWkEhJnXmbeAsUhEEYH+Gbm3pe0TG+KOA/qLQzkTgM+gnB
lyK5YJLlAhsmEqPZTleZgLAaVTw0BtwPmOM4DbnBAyEO4fWnNLzfAYsJcsZTygq9saEOCHFcGHC7
uTAxmDHEzRyvwcGXw7b6NyktVsa2ZtKTuzJ38yOO0uyvnk6UsHIQSaHx/LaZLAM4UxeRJ/bPJ+AN
Ujv1gKHCv5IsdaS0L5VIlpCk66LjTnnOrD0hRYsu3TVuj4QTwPO4oNZOeU4vOM3kIE8SHzuSNt28
Rst1wrI4Wno0Z+OU15p/GAZ7xWRwl9yyx6J98Fv/GWBdeCHXZC96TbEhu3fS+t4rhEMt3h6e4Q+e
kkxITKcxBp8b93tkOgdVWH/EsPScqNB68iOjzcyzamvW9uUo++V9PJqAuOBXE4V317PwAHBKXL9i
VGj6l19K8R0b7rZmn+DQujqHUXA1n3l5Ftf4gfhLj5k4cVFO96O5z1XDMOfhfQYdVud55RYyffw8
NbJgREoFrAPKK4bngPd27HEyPKPDeU3l9i9HaqxSX8b2KuaQOi8E1Dx7TzQ4yvoT5O5SbSLgXsoW
qCNjHapy6+6lggKYi5fA7jMj16xGKNiGYvT5v5amoErDkn0t0ttFBYqZ3vPLruo8i1BCWFbB/+8a
ftWbtI0/qA/sqG8ldme9db9bBrojT4xBHtGndc/uhk0yf/yF1yFB9xG2K9O4yV6qpn1+/cBIApAn
hzRsxruoABAEgpNqE2I2hAPVysQiuqM9pTqF/jKFwyN9aBh56Xt9EnUdDpc+3KxOMsN6HGggPO6j
ivG8cTwlo3PpPYnlydAVsydp0djzav+r8KY3zEFh1PTTNyShQl5chbCv++KBpb+gvpN2/PZrhELs
tOKclMrKBVXeLqpOXnHZ0BynTa3Rl3xUmTL6/5BvlOc8vwGmUISnS3vNgP1lSfcPBrcatGJtbJfW
KMPoS1H/gyz11wrR26JO30wsH2NLuClwC9jIR4DbrrVf9cAjAaDSR0LslGbM0hp3s8crXRdv67BP
cEQPNwRkEKvcHN4dz8zqfA76QtCpRkEgemUt3IjvZrAOLCZ/buqCcubmwSULm0F/ZS6zsvdOqJpL
h6xStB12BrnR3E4U3NfnCzUthcywCXizaN1hNymDSJPNfNJ36lO+er8lv8qhE2Sd77iu1diSugGT
FEa4vzfTDDD7BrkAwnyO7u4t6hRAVWrlHnAZ8tHbouZNslrWO19MKxqoJJiKfCr55GOXgZZxCfxi
G11VeVxozGbD1Abk+FKBrBLZqVHSC/rBtWCxUu55fAQwjfz/3h18Zc/1L/8pOTupG+21J5uPaC36
94UYrundvtJ0Z8kmYy2cAE3i46lRu5y66JWbJ51UNS+3PV2P6Qyt3PtHcl4kWx8U+oJKmkyihXQ/
D1wQMw9IoOzohJR6Ei3eRa+LmFDJG0yoXQLpqCWyXXfTIdSNkSkK7PSwTA2csfdXkwvl3m+eed23
6UkTGKqdyu3VWnh8KSStM60w1x//aKE4VhEOP1bPacIKhImEKDCkBW70bxmAnNAWouTyH75B3Ly1
c/+mxEGwro5/+00mE6DR07Fa64X8DvAb43yACLBJa6OJBi4TassuDR78MXWxVDnZJAKirpfHcgii
HNnBJ2RGrnX+B5Qd4MfXILY7asz8lf8tZjb/siNQ5u8uqleKYH9uzBwen5ZAzODP20+PFEkAn/q+
Ogrj2SS1P/mgxu3t+k8s+a62V28D2TKFlcP7nT2DjZ1nuYeb1jhDHfVJn6a95oH9pjYYR0m4txH7
W/3aW4I8JbYz7BkPXuQ7qEH97+DHhXkInup19A15R34NZnmtCu6vGRJ80MLExfFViWJnm4H76RQ/
lP7iY5igGaN1MtJA2nu99n/ByJGpBlC5ooudtaLQByGkLbcFsZPnrGamrWwbTgATTS8Bg6hvNaXW
hrtc8vI1bNRsZqmB4H5qOvGEzK2FaAGd4pli8feKRbMXMhzfZ63GNDK96opf9LWhY8m75BHmT3fb
qgG28yiXZFEfNDfvVZ3vlUMkSPw8YuTNuv50q00KNZsbeHgtOY4a5z637zt4NpdyPg/wxfO6JUyn
Cqua04Sq1IoJt87swR4Pu7AZITh+VDbZzrriEFG5vhcB5GmLayZHOcj0n2dXkmLiQGopWYzVa+6I
Y0Y+hxvPV2jnBcVcFhvYHhwt9ZeyDKHp8lV53yNNmPQHvCbh/WJtCLZrNM8vfc/ovtajiweVaReZ
oIBz5gDCBY2rlYQhNzonxM3cHyEJ3fYkcxySF6bOE8H/mAAJE9N/uADNdeCtlW6JdA2SUfw/k584
2jWToYxzSi7rYaEC7SdsAhAIxAppcz5Fbs05uEPlptOkq82fOzSZ184rGlml4LsOovwhGxpVvMi+
xHPW/F2h4c0L9ZrPuSLIyHAIAFUar00oDR8YxBFrC4SL4U056sWn0lF50WTl2aHtQnXkgMc1iQbl
FGHSOhgcHKkClppd1i1Ug/BQ1VRQ8Rmo8+locio0jCqUxq+QT2nk1JYudw3zkdNbKyFsEJEzIZWZ
fxyG2Wrm9uy6L4GOE14zIWGyHOqZZj2WlE7ESCaY+EE62Zz7dowPPf0ceJr3koNbTCyxnxowCGKz
0BbvnTLz5xOLEk3Bj5uqb1fkLxEbkqpSnPTl7ui/mufo+8FZMJoiw+QHHzFuuDM3rtpZpr8UvbY4
0kqFN9rfWbFK3lNwhw4sO/1NudQWHB3pV6HzxiciPBp8jltAMVX05PSPCsS/Rra2DUg49n+Q5BMa
xAjfsnazd30LHO8zFb6XoFTkQTafM0Kt4vUjS5zSvRlQh3Fuy31otINXqF/0NHODu8D9NK1Gb4VL
QhSI3CdbnOfkvYRKKC2xeir+gschiffdtjn8/uDy4uzTbjSdSRCqYoOtCJPQHtUuPHVJKXNt80+g
l9+CYdHxm16VGvtEYKzq2QVOdfUC+fmM9y9x7kFFb22WczXtDAa63gFmQ+UHFet7NZsrGtIgweiA
cp8MgMRcp/yEhDmulxLLo+1ahHSv4rlinFR2HwxWVACAl6f/CwECsh4tGycU1NLd3pebCcGodctm
6a2hq4qYVxobhTYqqPFEOKUJEwjXzRf/HT6BUpDRy7mdP0i7Kfr0+JsFccxdM80d8NNDUTkp0D8B
7s8+Lnx/NL9LyP4l9J812o26emuCmm795qXvIRF6o1zfZOOqOJW6ZUmBrtzIp8ejXHg4LU9q5ctA
LMMsRA9Rmt+t4vv4oYoe4SqpHf6vS1PxnixP+5xrLuU2Wq9NGRnoHK+O40CrMUjcGUOIelM2xr5D
CBr4R3nl6SJiYHTBd+uZC9xIHnHbuqLfCsCLA0PU3JIDxsKaR+t9tzlW/WZzSHMqpLo7C8NFgKJ+
y1eJVqkX5/XS6OJbAh8//o1+kzSbKajFyY9zwtZ/qOIJcqcnTt+w6UYvb4egwWQtrud+H7mc+Cm9
PmgpWm9E/kYpMUQqDf3lhNerwWttp2skn3s5AmnNe8G8FLu2InZ7Ci6rAiOPu3AFRWEOOcvmxEDo
ps0G8jiq81owC9R4o8LLKtp7xgQwGKsP8lvSm6j4i77++ow9SmYlh/xppYT+orrbQNIiDoKy86CP
JnB30ezuYxVOaQ41G7XjbPJG4t9nFNg1rWww0DZAt52LnNx76DRgdUJzAeYN7d81N5/VP3ZP+mIL
dl0N4ZNHLoDALS/C992g5Lj0drlnljolMizcVRFSaFLZW8NSwVSXZWg3kuc4q5flBNYf8QbGJI8T
pXfDaP7DT/KlK92G0k1kgrHum9yfUxB7inJHFcw+t8j9TddYPOW9qCsvq26hCgUq6HL1+u0qTWwT
EAYlXtQaRVgNqge2hagNhDRGunWiwD8hSGfgC6UjIYOnQfYWRfoo0RqNZJF8Eh1NAZSJ1oZhyzcP
rVLBJJmegIVSXuLCJK6z/41cCtXjmtDp/UyW66BvrG30TpRGojDoOc5bA5QoYXwQoSSOf3ilkAra
zOy4dzUvuiqqWuglHQt6aa+ztydfJUUEUAYzvEKejqHIHH15n5MDe9sodlk8v4yCDzVqQu82CiKe
AR8tmKfZ2Dhr9eq9uqqNWuxwOsRwM8JgFvYFVP6Xf3Z10vM6ri5E8OMVkz8H3ACA3jvTvUz2guCd
oqng+aS4AVBgP/IXgkIspMnjqXKkgBiDnUFXESuo70qnHM/kmyCv5+WGdHp5nrgC0yQw3/HwILfQ
KIUrHGtWIaKJZEJgY6VxVwiuQ+GXSW8GbJUZo/d2ECgyUEvg5dwzmx7QJBPfo00zK1+VZcsK7eEc
2iP68l8NVxBtbHmpivFaxsn8wHIWVCsoJFvp574sSSc17ge4LZ9amypUG8saK3kgJLK9sxlPSLgo
A3QmI0vNKt3PAl2ixJe0Viz/Xl2dpJoJa+CFpXB4ElYNwRBSSoue3JuQklkkl7T1qQOipJlJ3VLT
RUTm/t9nJaRTeCpEWf4xs4MUy0hK1ZvEDkbNOgIQ+F8lk4UlHXCg6JBbKout/08cW+dUgNJ5wOhb
Hbb9wVo4/VWBIyQ5JGeG2EFPKTs0aeqMNlEcbPRhVywoudA443VC/U2HMF81ATCjux8fsh3rl78h
s6bkgqAD2NyOwRIh3zn3vHun6tmr13FelhoG9arapq5D4kWBY314iaWe6yW/bEFAKFsfXvJO32Wy
Ih/BECbRRwl82Wy94FZvS0auPCHwUqLlh5eVGVPAIcmDz5Xbf7dUMBWJfYCu45ApLhqBrJESsjVS
uY0gwZ5hEXA2XrciKMpcJTgVDvpD0n+OI8KBaO7KciDWsLQ+5nc6h3bb6gm4TemOWhzQbIeAf2ex
EsESNUIfN5Jt++YcoDr2S3tyX2kCR/MVP/6LTldI0z9/M7d1W0v1v/wCW+e/jHWaV2QSqtuu6+vv
2rl1aFrPJINDO1IukAC+IV1NopDrymuYJblAJxEpnc0qPQQF6z4OT9Nlgj/qfnZ4N29MK9kXl3vl
OGQ7yvTTDhxqi8QbQLiA1eZ9nTRSX1eyROCTvA5SXZb+T0P5o+EkGdDlCm02z48tGAEK5+BxVHgH
4MivyYjj62K1ofKUR+gtg4gW+LZ/hwyUmWwhH3qsMxungppegeQsagPlZ11+isxdFedw1dHmTWdy
bKRoXLYSDsxqTvmah7kd7nV4/us6rdUG9hFAYPldWfJolm5/yLgnyGxtEc8mNl8RyCkQqMs9v1m2
P4WENO8xqmggdBVm1Vf622XwyB7RJ0LoASMHnKBxDHuXDJf1pzwpO92q9YgrZpXQZHBvnmAaavhn
GpmrzmwCMemn/yb15GaClrYC0VUYg9Sr6JOA74MttJyPKEQAAqiStNaH/TCUtSqIuu+xCH2Oy7P9
6qvhQzCoj48Ckv9UZKU3AYZSEl8UCQqTv5fnFGaq0vG1yf/dzPjh1AaNoR4XkdYPhb6wdTIXcY2d
wX3kTpL5pAb/ILWppo3pc7lAVeYss0FHXv+e/UngvWPw9lQmq0rpTknlqC1L0ahgWqE92RqG1ZQm
Ah2SAhB3IeWafZ13TQ0ncdedEPcD2NaWA9r9uydd6LqrP8Djpd+99e87dJUXb4XUA4qvAxDq6ftK
GGDIvlmZc0rHrPzxSGCVjbVMxW2bPuTyHlsp9MSYEdoDSKYHTGnvC95DPun0JKvLOXqdDpg3eJHF
SXxTpJ3LyN0iHOauRmTUascCAdh8sjTCLSKnwsxByYSxhlIAQiQQE97FhbppYFQNWx4TsG1wXMul
ZYq/osg7c32FH37G8rFwL9aJz5YfRWRp5fFo/9V50emtGhiRibPak+qhOO+4tMq7Nn29bWiS/+qt
d8+dAY0t+Brh21uE2PUrHxVF/xP7EfEuV6OTIPyJCwzf+v22V7ZXwJAu6vVv7/FiQ7LltSkEAJ2T
NX5yHg2wuz3jzgG4DqBPQbgBEGni9yhKjad0Dx38ZXcCSODDlzqIQ9P7hp3Wlgg7RRJIvFMTo+dN
5vB39USDkUlcOmAAeACTnP4eFk3Yab2pQnQRkCckCXb6vHNmRX22cPl0G4y+ekxri8L91bWZx6pd
og1wm7BtgYrXTMhAjimmXne89YyA4kG97wpLzUmGMY2EKBAzuHWT6AEb3z/fgpHWGLoCuu8fNhRw
b8+4gg07vziQTVkjHiwrQQCKIdAnYpvSNzVLdKz6dl8lRZu8QLT/ZxY0yCsUfNvf4V0cNpoU77aX
N3C9nkmlgxcckcKPADLVoaleUB+JQLfRyLn8ym5tioyKxz4NWNquUNdFvM28cW1h4wscB/fgtfNA
1gk0UPbQT8JtNPeelQSL05szKZleqDTBt2qXSEWyZV22xnvlriYpcheaTpKjolFnsqtYMygKmw/7
zIq4BgeXLdOwSMoCV7egOP9NoSs//0dL8PUYcDjScsJJFIAniNVIz6RdX7jSELA7fF1oolLXXjNS
4zCX14YukuW2zYC9Z6juClLqqMMbBiAjx95fpzPF4dkRWryOexqsqcRNBm0aMu2fY+7ihmK6ZUYO
ImqK/78RyoREWjTPC7MDEXX4jsYuyEjiARNbcsON8wjl4yFE2C+ZRI8SgsGGMJzeKWc7/RNf2xWY
mYKDb8pWBoFyA0QISYZSlsAVm1rdkIpfDLgQA+i+r/e+LWY+5sDcynOTK6SJgY2D9nWXLuCNekrj
fv1a0wR4hoyGd+F+Qmf/p0PX9epuvKocu5PfxrXpIEoKSu5KQFBmTTemcwV2R/tvD4/MCs+fIjlh
UPJW8AC0UMYh1uUH6zCIIFFjxZr9lFQc7PKXTA3SL4AeqHwybJiGpI/jnZHc/tKPiYrulS+Tf1Fx
Vyeka/ABYuKzeeMwOGaj9yHBxudiu7smYSSF8fmM2+0gXodqoqRx39gP3qXgvW6ZnxQFrsGeqGBx
Zgf9vUs+JZjgUUw33som90kfsnUnlNZr/vEzdGCy24cCipPJ6rEkGpyRXq8hpX6wgEZC1bII3T56
6lqnADbmgMQ+HGILOCnhpNt4TukGVqXGTGF7SzWw1rHnmA6QH2bQicIZlvelp2Y4PLI/0C3iLQ4g
UwREBPrD4/IlUrW4YSP+0RmenJDtVlpf2sJgSiFq90/yZnhurIIkKIekcWMgvTqjOymmoDnPJqG+
RWNupOE7xbHHlFS4BI5uF8g7+B8ChXZoiZVtAJi4q251LtOIp94TOO8o+pWVdTDkQ+WtLb4gUZfA
hjs9MVtee/WKwT4It67waKxCNsvF1nKRQHxuxWA8icqt66VdYwa1DYjFG6zMc5Hq8qKp4g7upufD
j59OJ49qXRAQ8gSip/0XXr/3mZMHzNyRWxKh5WrBNaLywmwIlvU17+qVkdbE7Ml9dyMdG7C1svVW
qF+I5/+uIn+mtvrP1zM7tYGYm2sRDUStN/6PKKTLm/UDgQLYjebqAvY1aItB4P5Gdo0qFbRKZbtn
4QKw5YajkGoBWJmQmT7IsdnhvJj3dR+5hSQtyvXJk5c2c91JwtG19//Ov2/wZpYLi6+EdMgjfH8i
5ibtHiGxvNgB0Iw0PzApif+TBrIKJ1uScM+33ZIm8rvD2PPbhX4o9oQuYAeFamqWhwcAKR49KBeJ
4NlFwlanCrp7in1lmofxiv7GDwnc3ZuiSBt46ER3qfFJy64pnGiQsg4IlZgMQy0+JldjdyrdSTSb
yaIazP0JAZffwcmJ0d5kJjKInU8wRwhbUWqGIQKnh6bSFnLR18GOLgINzM9t9qVQuINTWDGY3JNk
IJ9rmHIvLy+WKOZPoJki9aNDk3feYIGPUqyLSDEuHn/BA/OSe7gyYA16O4Q17jAtJwKW90tPcbic
7OFPWVGWcuUkPOWBMjg8Ig61az3/ibo/ZiZvVyrMrm64OI7Isku01DTa4vYp2qjPRaMZF0A9Kchz
3b9ZKKStjuW2LXZlagMuV9WKZTR1w7bkKbqcRIllPIWpzqtnu88cNOPEDuYn8D0GGJoUR/ovFDsI
qcf+CPJ9VbAyQvOFnRnb/FATTvvGYK0CPN4hH1W1aso2RF3sakqz4q1MLsvARZDTdfeiwH1+VRjx
rqDa3eaw9DXWNSf4b3u4JrkZmwscjyKFJvhdJlTxdsHVMwP6dqBhqHKpESYmEN1ZAY1hD/gqK7HD
ABq+nodD39V+L/l26ciDdqfd5zCJQlabTHGnsmRDA7cw6a4iIzxpEDmtjs5qXZYP25coy4jXNlBT
OUnfTnD5Uiv42hDS7NUmN5SBG7BswzcXsEs4FRI8OSalRarH59HpcjuWTOukbotyPRFzyZ4Vkiuw
e2WU10gElFb5aGlwccmckEY7d06BJIkNAnuck5NNc1brBrVtkrQva7Bb89bFx8R26SqnC8BwRhpY
Dzk8B6NevQaaY4GzaonmPipwnW/cOq6MiCN5CcTfQ7dliCQNhKvyVUZRSHsa7Qu0hP+WW7Wz1Cbb
8Kf2EKwZh8AE30vg5VfdMdzB+hRBTBdWnm9qOzExvhebtu+kge+Eff2fFR9KS2P9g0bK+iXzO2TV
cvgbqBM6wPas/deX4oxS7cvaZJi4AN6qxGJJcrWULuqF0Dz9oPH64fzyy9QcVqID81XuAh1FmUSm
dqpuk4A=
`pragma protect end_protected

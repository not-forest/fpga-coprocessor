// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
qlhuWIrkbGd7471Ndva+HEnHhOofVJZwmevIPJPKUOQljlsM3GNYmkwR2TlxhQkU
N5VJIsiQ12fnHUarx6cG8ATte1pafT8/WrhRDLGZ8hLVNdoRlvZ+lSQSGaMxCp3P
a24JJTkcgrvwjDEbuHCNxSI6TROGO4smBf0dNtF6AC7KTpnAPzYscnknO4bM2aHT
DosSNs3CmxCOhtALQTuuSKBscA9ZN6y1/sfRlLY6O1QVaMuprE6vrq+86HsIp2ae
uI2O92LEMA9XFe+LJNvksxvBWJyp9Kjb9pfBaGw9ZGaH/ynsS5Ca/VPAAelNDiM2
1L4R0OcVFwmBeUUTQNaN9A==
//pragma protect end_key_block
//pragma protect digest_block
qT5Qo4qznUUr2cCMYt0f0N8wDAE=
//pragma protect end_digest_block
//pragma protect data_block
pu/5mDH0id+h/ZqwX0qoXoDCcYRESJC1tNdddiqLDrbVSrrfzd44Ry3CVk4iYLdI
napFL4pKDIM/ysCF4InIOctJfMARp0wdCIofVowuN0X9149gXY1ETjdxAex8KJKb
o7VuIz7OxRzNipuMD5I8M/ls92X4AelVlWBGkABdAlreEL7jaQiCUYEV7nTpK4n6
MBhSGYsrvz7nVT1jkoOoYQ/zZU1RVpmbb1QTv5P8jrR8u2k2+4oqIhvNRSEgNcJe
YEPgsXowVPKLDkOGuB1wsZOxtcQrvDrXH+V6qBY7N81Kn4VeHanGGEa27/xG0Ae7
Up1DPOdyAsZ79WW3/0zCPwvfF3UEjzAUG5hgk9yan3qp+S+u8V2pJkmx0RmI1npr
pzo6zbiOHoHvipvKtkCalC7P1plAflD7h2HAIiL5+9R3gQqyl2Sj/0HPZpdCea8J
v7PvIrJ6scxtvdiPTnvN+cKccSEFdtlCzVQpHnZkUvTyKxwYgniqqqj6yd3/tylO
HAhkCw6p8ZSlj/k0HPYNRfg1BhJW8s0ANXYWuLDmI0n1mMcZloRee7WcnvT/hNc0
6o05KYQyBbvhUUcaoK14dGSgtUuopqayT08nNCccvhHMXNHoSFHGCUSh3Nt+/8Fl
akXqD74Hi1lVW1jmetrRIELiztfyveP5l7DSCDA/flP73DMJcuiTIiBeYgvixirH
jO1nxz+5ht34MdqX41PV9XhhgGVhFUtAOAy07A1EZ9GIT9E4eY1c6b1IAr+OjUYY
X6Bwd3sPkkCtAcqlXxj/rk6e1XsoxC1EJ1KpkXRsy/rI9gFyGRIGkwyAtSWo1zOr
9tN6Ls1itCckvO1QFJ5h9+D6vsIugara5iifhIjWeiwKkVkKMJKEGilAZQM4KGjW
PiJMLeffHlnubay8O6+zwkyOMQSSwcx3JDLP8/B6CzV6hLMVAoFgsOTLZik+ZiY2
ze3yxMSpiOgB4kJr1FE0x85NjOqLr+rlYQaTF+LxARpKPl1Vf75qMc9SPhVLidiu
NK6bVP9Wz+IsI8jwoQWLJhqWkdIsbU1RSd15TJXebHgfYmBzBJlmXfLCuXjwNIK1
P+lnIJE0WmVtQwcSnZnRZBPq4W7AHaNv4vctmypCBLGMAge6VAQmmB3Na5VK5sG2
Y6djanw0eZeXRk5apgCPRQT8KNnWEhI+OsyM6gYTBChbtwG7o1oTuJLfotK8KlK7
Ppi4FpRG780pGcU4QivpBsmzY6NeczvFViO+XVjIRtDZQHxEmUG5U3kQaGMeJjjK
O2610FTkoh8TgMI3kVWMjRsOz4CvgJP1gkpHBAayJjrkcqz9TdAjzRQasz9oVYt8
vnT3wB9JPY7IRq2UVhW5GemRF4sDJaBimzInMpggBmlCo44nrT5stmLIrWUEs4xp
ciaNOaXc/Ae/eIU7r0mIMT7hU1oA4aT1dgyWbHodkWU25DoEhgVp6OZtdSHRa89X
21WK5nSh2TeFYYEAlF6iqcF/nokKsnv1vs4VMStSjPvmnCdXOhBQy+8f8IMplHPd
ZdNU6JNAKQgA/WMWMaBakoQLz+MU7oujpgm38OqHw2W4iYoQ1DD2WV4M1euXPuf9
HJ89Km3tTorChIC8EYm1KZJHGBsau02hME3MowHhy0oXaMDOlCgGr9H3NP8IvPse
jSNC7XlBrLq2pp3CYdUq8yCzf2Xt1bkh7+4Dm+ebx4WqvTcMhkrK12JfYqrQnDwW
Nz6ikKIdy2Feb8646ODINXjg3Tj1kr60OKrn+Fu8JJUc/lr5r+XlQv9SV5iaaPe3
XiR9S+4LiETx2o5hztqaTVtc88Mzp9H1dTVR4t34cBSiTIccyBIzNn+8fCs160Ai
3JXBtayVDzR8BpA6MPdilFK3S4i6Y2ps7ZDRjUmshfXj8OqmYbW7NgVtQn6eH1Wb
KMPC0f9pdQYulETeJ+h65suRqrWF1Gyiu0jhCYIDjHe1briSpaD2547BZX0eq75K
xQeyV2tEzSEq9N2PmiBgYuQi1eI2gBTzoRmYiovJhrszEotZdsGs966LiCsYpxvd
fR/9ybcxWMD2eLT8HZpvJg3fnJYRqjJ1rRuOXAJIGKQJ0UNEl7AXosCMW759+Okk
Q97n4GMIwBL3aTRBjVu5L2vbagkoQ0cpPQ5lmY93x0ZxiP8BAKRV5YYaFUuH3FJH
v3P2tfwUtDRQq6q3e8ouEl3I95fe4XierIw3EFEina5a5NxyKi6eOUhEoYr+XjIL
esKj5PEWk/8/bAOcFq3KwAmMHA7eW7tPLdVg00JLGSEejcBezuh/IEyH7POziEmL
mu185uxIOWUUVmDBMIbgk6Lf/aqLuJgoBpzCIfWoGA0TbscpMSRhxnfUQGeLVtaE
jOZwvgpCRo5lwHfvY2M1Vzp6uycmkyeFC6tqIC2un9UMtD+yIVWSep3IiKT3IqzZ
ZsWzXnR5GURlKrJPkmArw9VmfH8RVJt0nrHxfDVl4uru2D+kw8LjNz+xd83jgBWU
wn7bgFsE3mm1DM0wuMa6Bbo04AD/H6CUBUqx7ONO1bKSIQ/oO2P+ea9oIQwTv0ko
pBVDL2hskCdJ/TdPyk/TfKyUXFIAAmv1lhXLWIPZDoK5S8UKVnzCSkpvBBh/ROep
2xssMkc7Y0Yqs9Z1N6tfdfoKNoxqNB1soVJ2bXcn5a1TbCjSIzgLy05QddMeu9AH
7SRg3a8tEqECfhtbwRpX/iUwFEM76MP1hM2e4J2pakpQwIuSzHAZErOZz0hnzROh
3yNXzZwh014GFNSRct7bd1jun3CegqWL6WdwZH9Ge+Apd+KpeBDNg4c/8bMfwOMM
c2G1iLFO52y3ljgZ3oqkguBVgChfLJpN4eLiug4gIT7mPirC4CIw99C2VYxJ8YWG
XMeeAG7UzbcYkwYLHtjS83np62fl/QfBRWv4YH+HBAof1RFQdfXdMBL/e3mTMyyb
9lYkd1EzsjYYz5u5deH1o90r2B3HjgtywDeVGdiHsjO3hseFY+v5TTtDHEiqTdwE
E2vuNs2cw4sRH+lJt6myzF3zxe18Tn6CZx4nt1opH4EEJTjMjsU/pk8vo4YQi4dT
ZKXJbO6HQd1KTlTxR+hb9XlN38XnZN7bRzO6xYuoEx7Yy4bO2hIyN2GS3bnomKKX
1lb0yofxa3XH6q2FkNimp1PGWtSF0i9bJstp8ELwW3vxfSsF6iVsYt7U3qmKMZCj
Pd4Pv6l0MB6DUfY15aTmQa4N05feSevM96ojn38F+HR9XQhfbKm2JAilZyJlECW+
b1dOrosly/yzalGwMpSN69ZCQzc7jt4BSeZs/h9IaDVmSymz3Nu3LdJD37bm8Y/w
/oKn7nk3Pqvr0MCoKBcitmfzHsvAwElmPCaQwfY6P5BqYsPvLUhvmoCrs9emXrad
cz2IQNtsOOvNYXoXo54YXPkR2Cyb56V8vduXv9OUKf41smUoC6kweB2pbBzLYDK5
w2naOk+2JDDCTHKbqFRJgSj/LbAVYxpHv/1DnIusseaSa11n24MlDewAo85IHCTZ
p8AR/CBFwWsi3AgmLMtJBTvsXombIMkd8AB2ywZdZZywFXJqiMsaFP94XELnvsNg
ZA323kif+DUShMIWNxQAu0Tiyo0Rmjpfy3rpzoAd8x53vhzf4wCD+wdNLutIwul9
9cfXKYIr91A7TE2fwVoqysRn8Jev6wn19y9zLOIiNfFk7qAyoDwrCw6JBgMRbyIt
sypwygvjl9tzd2Yce4DjLnRH9OrRBcSUsYCcfDRvkZHuWdVvRcEjKx2ZUpmXt2Bm
ZKg5P9yWA53aLzmnpZQiRGAgT/OFJYfHj5p72jC0q0HMvm9x/l/tqVZK+5wnauDY
BCQv9tyNmx8Q3UyWUR0/gqEcAUmCW93VV37JU/mAbI0/jYfGe7nkIUWJC/Z0kmLp
VONblvFFfL37CzUCAcK36yYFHgPlPoj8T6osYI++6W631zvKye/xeJs7LHW8WNy0
htPwaSHcapKVbrhDJwuQK0wqHdYREFb7ALgnMveF5VF4RRGe3r942mFTDumuRY9J
4bf5+5FcYecYAlaz4P7gJaDJtO/mgzAPU44WLMdWLFjQfzpqFUQ7hzI148SqrPv9
SFrPDuk7PBBHldTB8ru2Tw8p51dTZ2tE6L6DSey4U0hSsbwba2fd+fngZP+8t3aP
bwOEDTqhug7Uvwm8NRkYqngAoM5MQx+3x8QNXhrP8+wrZSLmLKrAA36fqudJBjT2
OwlVw1cNzYHpRScpP+l2HL2g384DeIJFBXRjwdf2dPAhb6Nbr8ciBAIvn2zdWByX
DpZ81t89wDmk/N1EHIOv/cNOTysXJFPopA1snS/QyM8ed2Szh5ssRFSX8jnv2HD8
nyasEdBoKQ2GIbFqZ6V1HX4jwO50iXs1RyD5VAJE3g09EeFYceh+er5nt4kC8+9I
XLzW976hVjeGr44/2szT5b+7wwAP53ophyhszivwF1TNhmqY1Pu/jcHueiVZDXCM
b18SIG6geG6Yv2Zyn+4/jOB3LwkurS1Qs+E3CAc7o3JKZWwLT84f8ZIq1iIrb1wh
MDv71zR5j0mXKnzV/tjdjWmgCYqmN1nxMc6UbE3EUXpfRzA/DIchYamMr52n8xbS
z97t7hrnnps3sfpaVkpsP657jqVdUGhq7SNrJlWaeWpWxBVODcfnIOlkZiAZBwui
Tec7sYCp6qu7oMRtqmFoPLnimNLSVbSugOBTJRtIZsYYfVLxixjM7mrQey3ANgVu
Qs2+8W/vyP0OdCACAqKpEO7/ZreEa2QX/ceB+aNNxqdPp/LZC2e8iUhvM1HNpU/X
ik6lEZafCIbuis7AvHZFOV0uM1HeRLrdx/V3iz+1TcPhTshg70WruBmeJ/nLlRJ/
GANHFYg84EEg4BK06lyBE4wIcLEar4KAzST3vJw9tUSyQtItbZXbjiV4sIQtEeXJ
8jjXpys6jx7qc8q3OQ0ivvMPsvbgwqnJdc0PnMo2XXBgYy1MM3cK67wlFqwqs7jA
j9Xm8fipq/yewCZXWaYl19pIkgJHU8bYJ0lFCaWUUUprGr4eQgNU02Z1LeDJmpQi
KFhvCH/yOOLxDbdoiNkelbwABm4i6Xgdn6tIqHtOwyreKWXVfwC3bhzMwyRNv3+u
Pd9YqWLPzo4bio9XDdoCvG4T9peOPHRNxp8NiAgkoE0XAyIy/GLplSFByhuUNTV4
0bfI+ZiE8JxthE+6ugmA9BKtOqNe9FukMq093CwQumedvJsZJjSoGYyjSX5BH5T2
1DfuuvW/NTWNr5VVSPSLS2Pyg6aRTGWkAlEV7NGP+qu6iMDFd+zGFEGcZ9WweUUG
nP8/5IZs3VsPYhGqQRn78qDbxBkKyYSSR9gBD2+NHDrFTfpbzFuchUJJKq3t9bXl
Rg60ZpnrCECfDM1Mpra5sUVOsI7+dAWvVbvnym6hNnIdU9STvmtjJWT/uDUiYL0o
fvKFr8EsEIzymkEuuYvD9NIUehrIgclUnGsOp9KXf4u4PwbKd5mgLzHtgG/99vf2
+QF0JFdbFTuFSIsaoQ4bYHIYRybkTVMLVSWFgxeaBMKc5cADQ/dHwWrFecehp393
339zZbJ50W9QcYK9WruDiZas6tJdrL8IZSLLkjUOwBVKC8iL8TjoNFY8fjOFqU+b
6f6rS8D69lZYxFrnltnQUzGUyJPznXG7/Ng74KzgkF8iz4Orug6zU52OCfpvPzCs
cEFbPPkBTe14iaePNsN5nkUwxuzWyjDD4V98XqeQcU7q0vc9adyMmRhdgBFtKCqP
ExaiCvWCWtk8xzRAuRf3Q80Hy7ngSl4Ezsx84mbneD17fBkkf5rZ/qmTkFhJ3uor
3ppOvdiWuII7WdiVnCyQQQkjtFzHWMGYS4MdxtzVt7oPShPBRaQRV92VfCo/wrO8
ZZcCpo5u1m87vGDQc3pEzaYLMuyP5+bHrTOcNXGCfqg+BPVT2VtDlBYSKfkH3tc/
T4WYn3xTNcDZb5ot8VpDPgXtEjSaE6whwI0mkNWn06MEOm/PUnW8Smf9m9j3wwPD
gxyAP3Z6Ydb0qk09b/TPGJZ/5BFjHtlQrTbrTGX3eM78byx8MDlU/1r9UqIsM3TL
6/RKdzNqGTf90hMjA94bqRg86CxBp1+SnGjmMK2rtrrdglqzmQ+o+tgpSIbYwhtV
dTItDqyuvNBj83caVlHfuWZX8vTy4NYs5IpyOpva8SFX+ecd3n8XfEnmCAHrXHP8
ZvwPzuOqK4kbzYHzAevVA28U9qtzyIIYPnEevCU+aYgGZi8kfg56s8EqTE8ACt14
laJR0IsElSHd/90IWxkUTejF2unXD1dhFW9uwdQXud3/nTzu2VRENSw9x1Fv8ZXq
9/QpEkaWJdADci/1yptYtENs32vvLtDlI8EBj93yGZlnDo3MR7rq+0JpJMmvlwIm
AZSCNM/BkuV6j2ryEzXcAbjpdV9CaPS8nED9XrKhTKjUabfMBvVEcNn4aqvdSqYm
dJRi4O9xVTq7ZfFLStt+2wU3qcTLJxM8LVfwHUnb5dyPjOJbfzTpCne5ZXE8XMg3
Egv+r0lZj4Kjri+sSUwY2J3OuoTyUv5pKyrSryRmN70HWUYxKw3G8zv7byHqSUS9
At19cTnd6dIEYts4XUotbU3HI5DVUPVTroo+pclOOy2j1dvY83T5T2xJ+OoVG64r
A0RuyFSr7tWBvJGPAVsowfMNp3rqbVE+LrrFk5LDbLdgjqXd1L1W+gp6vbzBGAZQ
mQQlqp7nSol+dyEzVCRzHFFPeIS3xYhHofBZSGHOfOSIbQeAPrL/3sSx3WpEAMvN
4DnkXA3koa3zkgh9y79JW/n2NS6aupnhGr+CBsznUOR5YQjadrVXzpsda2dk2u/L
WXhtHrYj6nSqX6qU73x8J4Wz9WKXiC8KhS56ikqamOKZo3fFfKjSobMLhpCaUVH/
ZJwnihQIW+i7w6Xzqgc7lNwkWbEkcZmK2BGArUDLv2j6rfj88Bu9OwB0DZOBWDJg
UW10pu8kZZs71W9kNF7i1DI+NbVivF/BszWjXnHl0AuabLgQ/rU+fCCtn4wQjFwF
Dl+rS0mKs4tyBTlzuMSfe9vtGC8Wbz7CUmf5mKTAU4J77B7nBNJZkZC495orWPFM
rD0Yqe1zKiVwO5A9zJF/NGDdNxRiKJRugseUhU9lhJBrl+Q+zEQ+zUs2bsw/k8RJ
RIZksY8Qt49gtEajpiIkKFHgMEcWo63KiFRa2X6RHVmQtzTiyuk6wT3u5/yKgZih
z+rfwqse1yIYKMC+82gyI3ttzD5HnMGpLHUjEtlD+iTStXstHrfnSXbMqY+PI6vF
OVm98hBR/ZHg083CLJRKEJZdr3e/Up306JfMflIDPjVLtsQ8F42lfMf++zEeMJcy
JohF5Dqifhg8dQGTUnBlgAPRIOWMcwTKNKQPvvq7Jkj8/gx+XTZrn7WSCGPmQr9T
Y3v4MrocY13hJ8ZvAPoRhvWIDyxilmApW5lkrw9NgB4/YE5wCW9ICln4ffz3LDSL
kvoEOmJzhZ9QYOym9empNUYWrtT8h0KMHQ+uAtUpxskaxXIZhxFY6/lAKOD6pH+h
wZFCffzs7T2vZR9FJy9K6pvwnGd+bqhC7timx7i2R+TTTwnh8csgge45S7OhKLoC
1ApID7OBf0D3lDQvRHEsCcJgppWOIPTuPC3j4YZvLN5LN0UvCwskeGAyM8fY8tQA
23rqr2jh2oRosWifEL3g9xxpxocHuw2l+rrU/LY/4se7aNMt/AVgJwAeY7qXQyZQ
iBmRIRaBgccg6+Y3ly1+SPk615WPkjerpMsGbxsUIkAGSeVWSTJ7CznuVVF6vq97
fRYrNKqvA5WynLQvPvgDfC19biGV2Xyh1ROk3/W7ZUNcLUWm7v3AXXDxP9f/eddS
ajjE1z95fvMW7Ve3bzXI8AWASXRFr14bqIa3jGKtnCOJ7aGcLd+TfKA/fPKPVw6U
9Lce2qYyQ1tfZGQBXS9rOnYWgdX/21b+6qIZJPeSWurm+s6deka6AFB0oolygY5j
ziOvmnbBi37SteZGwfBcaW5Cc4LGcOmTgr08C9oezD2RVBDVcNZSQZvHwR5OiPQb
uBxPm4kMX7aqdumMSFNweUuc3OsNhu8+0RTidVa76PuprBhcEX8ZswCMxzylcmdK
d6A9FxPy18YJpzwt+B2id24UMdNOh4Moc9PvwmRWjX8tnFbZ740EicLuDzY3jkDf
5NKdAwz+hMFvjYI9npjU1/aO3HALEg0z5Z1TaADl2d3NXaakEwWwuLrHFlnLe8L1
TMNBQBNIi0psYBlh6pTeWPq+yhbqNjriyUeOY6bJa4QDn1bEeGvH7HgA2o/mvJCZ
ZNf+fPCTMpjAVKbyajP5zjdP5cIikb3tq0Hh8v6k7/F5NNqoKYh70rIYP1MXciAJ
fuOmnimehH+xsScXhTL5ESpiXx4Yz87rj9cauWO45b/D5GjciCklhyqqsTbTXXXZ
yKOK985pZtcYDtr+Vz5Sw1GzujGlqN1lzXLKr7Y3DY+HpHdyBT+wjhPqPrAcgPT6
AfhzMlepXbz6rlb7o6JA2CH1e1M4tBhfpFeR3qEfalNuHtMVGmp1OG1Q7q+b8ho3
3RxIfWKELO+tk41mJ71XSgFUG68HkVA0DRAdn8quk+9cwEc5dSIlQov5naN1pY9a
yaWfO7VbqPoEG7kb9A1h5chwKznaMGl0bHE+4oXoEPjh1kVAMKWqN3TtOzWijm1+
TGM7TI/FMYkXTDrDg3CBvy7+lyj0LjG8gboNvbGgWWUuXhOzP6Xq62/NTUnjY/j1
8hq6hrWmi95qecEuoqc2+LOfto253RoaRsf/Wfvl1y7T7pa15HRxvHwF2sidWrJo
mH3TjCKuULcq3AMSDh7UmTkufgjt0Z3cvofGSg7ciiBX9u+wXteFku98CnD7FEo/
RLGs6ER+zagKq63N+dAGWRoPw8NjxQy+zCtBnWx7m1XjotJHRAeplvGw7Xc5Y50/
MlEOoFv/Y1L5pP5JEAK5HmpV7KyNhya/efyhKZdkh9imZoxNTFn9/9WoY3Aqv26F
2q8mhi5h9l6zxEuVC0MmwvgSaLatOMutQBXarXnBt7oMLKw9SaOWCkjUlq9LvTPq
PqFd0wRCU5/llMNB7NTJ3zl5jMIDPLFiQwBqLNL/y3xRXMUuYz+4gK9RWBeT2gpD
qz21+fszU8FD6RE77L16a3KJbndZJIQ6zcourLuXm6KxRyYU+qCjodBKQrfq5qLR
dMySQ6tcU3tJjl3FpPFdSAhj4Hz3bk9jCSzP+2zYH7SfvpuYla2CzNYcqBpvJqjP
u53WywYb067Dq0rFziaXd5CSI7R6F/WCQLo81WrhKZ/ZWpXXjoA1/hvR9YAQz/Sy
lnXR6G5wmkePqh3HtSZuhNcDe729tVnTtvH9dTEzHmHrggPJqCSbvYHBiEy+/Ynm
DY8x61DpJpxRjv/QNXGtQ+jzC+5oqTGoVdzm9J7yE8qpJsqR1Ft6f88KbwC75z7z
+0oUBZ+uA69khkXcAuJ9/+6+8OcFSGFnkiymKkhF8W7jHPEWueAD2K+yC15+xbtX
+vmqN9SDCB6E7gPxvG5/RxtNRC9g0ewyxzAdVyFu1i5Yxti+7L3kvOC+8Dq5nsUg
fxnu+/TpNgYSYGYLH7xOb0eSGRWxntzrsbnXGU2uzuoEFYhelGsA3j5iB19YoO9P
TAgsnyM6wFt85I4jOeZ84A==
//pragma protect end_data_block
//pragma protect digest_block
s8GL1pN1QTMgwm+p2tPeALgkb5A=
//pragma protect end_digest_block
//pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kLxrF4UFQgMaagu+VNS1QmyPh7wmbWamicg32fh5p9qGshbMRfgEdhxugT4oc5ds
2kDvCube5OgsnwQOgUPEiOsM231G/Vrtg+IE5xQI1a0kpvDdqfvwY8zYEHhgd+Ur
w89lvr+W8TWx7CR/Nd8SYuq418dJYTAaQe2koA2LWRY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15248)
35Ugf+BfQ4q/BnNIcmreJm52WUrJHnOKS1sW5O9y0H3+dfvnEVuGgTxnjAIQpYI8
+FgzVhjfMgf5LznjERMYqvlFzoXiaOge+DwQP7JkGHa6Paoah/X0Qe/ukeD2rRzo
sw3Y1Wh3EG8nNkm2Yb7BrRFBS8Q9TmbbEFSHCW+zowRBlnY8KeHUrIySXH26JiRS
xn7up6nv34tdyUvxfuX6inuOxzdiwdajlRoKRe+Z7iED+DUgWvCRjkBrcj9gyP2b
DdBqITwk8GZTcsJhE7RlPLWykwQVW8sORFx9XQxmIYtZpec9Ta5PjUcErRAESltc
Io8GbOhEaOAzlc+LDnVQazL7sx1SYuMX9VpNPK2r3eqECEoJA37V63lPlHg8nsIA
p7EedR1obEmKTi7e5LhpJw61Le0wU94ja74fpMCNc5uRoMtIFeYvTmlXbhCWTfvH
JbTGkOf3mhEovykwsWWK8FuEQZtQLUT3rBgJ06/cv+IbDjYECR0JYXrq/yHikCrX
80gepzf/0icpCRoMNnVuzxhOt/MdTTmkpF9a23TYrXb/7OYOMaVrpO7e0te4+VcU
owHJfe5J2pAEOJ+2uTClj/X9VajcOwkACjqRoZ/6l2ZLRS4tIdQryyEjrYPD18yI
RIlP3pmd6mFIoaxjj+sqeMS/pE1+CG6/29WB2oklGARJ7d7s8LAO3YEl7JDuwr+g
k4V9BD8GzAaipgxOORTOTfqMJpwNEkUJPnvQUOkmDeD3bexe2HslfcDqGMVLPEuz
4TR5+0TfYvtOoMai9PSBvlZ4SE8RgFD77yIzEKTcf9W+xUIMg7ZbIkXu7BDUHBuz
q1YG2v89WOqyyORq+qRM2M/ApujcWSMyvV85Umr1045uYQVmrOBzd14NDhw7cTDC
RdwzJBun6lBQDHM0fPFmkohYDThrU1Lvldso6Yev5MIHXezAkee2Uko7cAlQPR2C
sLqV/IiBDRBAIFlhEofnCgUKrc1K9mtGCWLQRp60QVV8fG5po0VllwfbWg2pksMN
q+HXBcHf3qQpjJkdXUF5a1L5UfWayJptp3M467F2/SbQDExnuceS2tAWjP3WoMVZ
PzblsvthZHev3zDA5d9+YK2Z8PmSHyxFg8GybLY/ysVgF41tL0TRXQRiD7VT5Gt9
3UgGZ62AJyG0mQ6vpwPCckFZoRgYiYGu8Cmm6sVNG7pOiPtMTwkOAlgd+n5fpMtJ
VFQxRcCdjcvEf8c8p9t1YiOieXFRRBouxf/mVTKbvUCMWYfaoPRgJShNB7r65olX
IUgvwBTn8lUZXpfBKLAzoa4nosTDiOQOhGIYrnmfCzM1b0RXwJGnWRzVIfxMxbrK
iPyuSEFfHSOwW0U1GxVjQrAzk2xeeIiZEhigbhZyt5aNcZ72WiqtxA5wINpKYOPz
ZymFAVnY9N8gnSZipOWywzGuzw54w46w1ESJh9pyq6uNcFx1JV7ZjxECaMf0Kk0+
0rE/odPxmk8k9DtjwEawhINpVDPvo7GzYiUxTzxE0MV5B1ei4EMSS9R1S6/qlvIl
jMnUxtTCDO1PPyR+cucixBw9SgGWh1mvSMNtlbv72qD4hdB7b5++L3WBqsnKWq7z
7k7t58+itmiPddnkk+UAMjlt73juHbDbKDIha3fIAwfhCibI34pKAGFl3qEigr0i
d6Xzd+abL3wGFDlh0o73iwyevWev+y0cKj+etnDnFOBcQFRUz53rgWPKZ3TeO1IH
VGU6zuBfcHF8C5VO9Dw4DiNrDTXQ7Eov5zoLT0WS3WsnXANveM2l0vceXtTmIYEn
tlCJhl2h4ke6K+uqMhiMLH5A/GUvoJJ2HnFE6rg1I4di40WSfPKal/QtttbcW8il
Dvs9Ux0OWrOFalIPspE54TP9IOedHzwribpW8K6Y+jkLfYHaeA6nFtn1SuYcZR8B
Gcw6AcDR5mscMNTAxT8CMrezoFoLH6k9pHteFNCYzVTdP6BnHrwXoc3XNcEpeNXR
YfULAM7jz2T70n52+AcTbsna0iP1n7KIjt5/ojhsKqKpqgeEehEs6GjWgitBm6Fw
t7WcEpuH1IzBY37CB0YDI7TQtlbIDeyWkPfoR0/tFdAkCZ4t1CsLRfzsxzcfmpfj
4ZJRtT/irvd5sg4ebgWgC0v1UK4dBuocj//aQwORW+QmLrcjbfPRgxH/I69LrLGr
TZ/wkA3oThWVzlEYzqCwYFdHb7Kqzvo2e0nSxCstfWsVXJKm6uHfTIHY2TXN1Pt3
i2D+UO/l08Ooh1PpCooY2uXGidsaMDeS1AEhncjYc9wfsBGBPZGGozUdjry2xDb1
UDyrE2A0PL12msOp7nRuBmvoLCdj7yy8s8qcypDuwZ9QS0kKezYIQ/+9qztkxMu9
pF+uW6CJCE7pR9USwBFaRVyglLF92CD5LeTMI2dMCJ119AcKr5SIppYh1RJmBAhb
Wc7CGJA7jC6NoLLpC4NA/xKOI8/CwO4Hc/ccV31asldaT+n6HQ7N8b5zlm5C9+tC
ISBoL9U1WTVWDRx/i7Le+aki7JC92OHAW/N3vJaTSH6koSD44jqlay9WqnO4tPK/
Z5t8L099SQ76DGmfH3L2TM/5E0S8yl4XIxZCfhC5bhWi89gHJSaiP3zwgmheHdJu
HLwf7ih24klCE7vBo2NXMYzuDmDH6ybDuesWCyKWVsXbZ9+ao1AalMBotIIorfu4
2jfMFeTYV4tFmRLbQICM4Bf/LGhKxzY8HJRc8l1ADltTQFdexKv1XCTlyluOEmHT
5BtcvN3dhbboQAnw9JPQ1UkhsDiqqMgmZ7zM5Uogn+yL/Rl/iJbE/B91SdFjaFxp
SHPLofHqYeTopW9oi2aSTIklHQ3E3/ZISuEiVNYcCQTnmukiwv9zGN2dK/pmf2LU
afNqaWM/LeukoIkykSXjmNne9UOYeIFIU5oiQrXJEU08zuibEU7Poc529wAgAokw
bmXdM2FNL71HIESmuMgzHYr+JlG5eV2KXwmgAmE5as96DPDJhAz6ZAdaOTCaAYPa
Lt3q+7kkaV+PqvjD1CeTFtSayoO7kXH2SkXX5w9op0CB/zV9l7HsuwwHL3RU3vS9
VuMJNCoAkCp0RH1NIebOexwbUe+tHVL7oISj88Gb/IAJqHeNMJq4vfpeqFVaQpim
JyerUW40UL5vdrCgpmVqcbY8J8bDmDJSaegWrA/zuExbYmEC9hVpZFEdwhe7XTQg
p+7Lc5t45b+sZb0UJ/K7TnYBvy/lIIg3gYC2PWYR15UY8jeFFZbf8r//HdaiSa1N
sl+6/TE/leueDKLxg3NOPhTRRsvDfVlB/esHLs/PoHUnM8dogaFtJUtSDcwf+g7Z
TXcO0MSJNdQR3GMRjzYkFI+fG00Qt2KMjGMcbV25F0JBqSvpSUNojQNQODhZloko
rCgc0bpSiORTrv0CIAVgU9JN2im57HyFzZGKEgqPLa0mThw81dRc58W+h06/MKTB
2Mczz4pIvbtHUfXicgGynePvEAl63Hnni9sv/xahM+zIJTy/auZWrTYshwPQONXt
rEIVIbt7MgFeGlTNC618jsL2r2oi50BIsLf0bCYHoaMzYEYUEfAD9WCAq+rIf2ia
3tMvHrm+8RXYzFeyFai9tWfjJK08wkYAZXCwGBpKrqC+H1502V1UF63hy2yg6R+V
/JH0rZcb3lp3Il1nG4zNGUmDUJp3OOmd3QCrBekdcVGbXium156c3p045VmZAz+V
iY+TucOz5vaTr4m5sm5tBIhrnmrumigIpo2vloPIS/X9FIgXqZuNkco4TKTBdFmG
rk90UyZaDSdmmf59pBrZO5YcID8WkpveIWw8S0uUMmeGP1mJv9TAK6C8QK1ue3Ri
KcMOykBQhOzdvOrHS+jkOTxOJr71RQUeVJ7BWjf43T3vjKxZ/CU7RMYjeSEWTe/U
HCNWAv08V/vtEVFLj3T+1obdB5I451Z/f+6RuGuMzLIaBsupwNKComA62krroZuY
0vRN8+BLgQQhRiEpl/PYt+WhJWALuYnwQDayVTjhHVm76KMdc0VNVXsSRjCDUC9w
4vvlDN/GUMPvgzS3KQ5sX+GBsQJEtBAWFzUNZ3ZoUQVRSSF5IkYBYOxpqk6Zce+d
ggywxll+4vfLYeCRsLZx7fSI2lsESkN1u6kCS/XWUC90xhzcdgfOs/KuR/JHhQGy
2Y1LltNKG4s5mtbXpggbIGI/EAIMv3PlQIPkNxaCGvsg4hTfdAXiLxDQBq5eJ3Wy
ckcRBmXqGh2GDiHIH6K8ND3RiRz4XeKA7Fp0ANwa4vCiQqLaJnb3wrwiQdSIM2iq
+X1sqPSqyoziG/qhKMhprsJ2tHUa+BUA7MzMjrSLhjmQxRrT43z7w4yaRRS69CGf
Di5AdzmPw1Yb7F6KYCzFvF60QNgLxuBnV+OEdlqxQIn/05E3BENhiTUMYNuNr/fi
/R41/lUl1ZbeNtv07aWWwlsaQJFIgM8MPaqeBYn3MbHFCrY/Re3RRVqvs92lhZvn
Yc77LYDTAv98VWvQq/j6HapKvuSJ9vmtI9dK19PBLy2tS2HIrCSWtSpW/xKlVTIF
/25IhxF8AnkLB0X/Gsks7n6bR7fhsfMaQLyJLycImZsJvsKF2z/QoYX3c8tDVGU9
wdKic99CwVXiQXA86vepaoMj2P1zZkKvpR9Rd6RoL6uduC1nz+hsP441f2zcmTnq
6Bg+j+vIDCPPXSXg1jk/nd7e8py7MzxVhNJKq/d1bEhrsVYU1vpfY075IoURHFwZ
cfgFcQT9ThyXKVlRYtu0VhtORbJOvERZiSTRAfI3kw38kdLoXulJhRsYah7sGYN6
8v7XO8vGM/K7FFDkEHjArm4pi7i194KN/okl+9sNv37sYOg/xccTpa3YsuRkYHwx
73JzmWyCHTWLdxsaL4v9Fo4SeU8gio35ssmB7qIhxFJz/2AoGhsz5gJf2YUqyfUd
NTucWxbyuAjWyku2IJ3AbrvTGHqXd9Yq6Tv9bONLO4BxIoORnxDUNFQAL+9ZtbhG
LJLDoXUw2EoYSu+oRjNRSOP4fQkKGkJ1M/rh8FKZneuXTbuuAhH5Qw8KScveTEc/
qZWbKG/N4x951Oj1AJfTO9AhCVkYA/4VAiONP75jD/UEzlULEpZb49ppyuRKL6Gq
yto5qgF9PWo9hNiQm5sc4W1vHvLxUqwNLWoOvycE2YJVNS4amj2pUZtPQEVPBowk
0TnRzT2ALNSHqiVaaSJMoAz4+Tg3fNZFjuHK5PtkqEqhnvGU/7ANDJgeuS13Hw0i
qgcOM+6VhTXpRBDeJ3r3/uj6ITVoxsT4ydVjcLP06BAvp94jbecrmlsz2B+FhWNh
8ZfiCDn8nLv6iqCyCFdyC6OSuA1/p/LOeCs92ewS96UtNdnGjL5Ezdnr+dmBNvO3
tctnfAr78iLabkgB45psxZ9Ps8HQ7MuSDDJ9qBHj5lj5sQMOXiqd4dvpXp1QjfXg
3EczIWfUvYAa70C80ii26Ho9C8tyic5V3VAE1akLGTI6sy80x/N1efQGxRVL/1BC
7d2XBFjUsdczDrUtMb08crMU4ZdhxdVgXuZDLgOEDggiK66+A9OgDtDiBG0h8UUT
dXvqSN5PGCgIX1IJquDW+ruj7o2W++mcOXpX7tEjxlr7NnGEPd1I6HP4H4mODCSz
3qCWhXi5OZHePQoZJutm7/fa35ByBFAeJDlV/SvCaLtGLbfWBffktmTzhygBlt5Q
C7K5kruFimOwWysI1pXHS0UFYQPjQElKWxkz4+L5SxRYYWvayr159/cJZ9myXU7B
eAHy80vC79/zYDwahb5/0hy8HNvOKOFucm31KCWtquLyTcQkyz3iFBPGLykdAMbE
SX5IDzb8/EWPrP79VUPmiC6+AHW3JWbJo51ubpLp/pYEnkXkiDdKckOnNuicDBZe
6Y3J/aoXUxQIdcIrIolJWZWNTPAqdU1yYzLhOKey0Zd8/EXYQ9bPt2bWvwN4tcXQ
Yox9Gg+v+h2Z5WATooSBa1DTIHqizwJcs9BZzf87fLCzcb8zrSjzaHDl6O6kwNRw
8PdUQAxWdfvmSamj8IPLYcf/aVyLwVPrxaFiZvh7NxLvF02vp7CZSb2T+zkTqtds
iyvOd6UKf+lLTJG9B1yNZKhuTQyyqWFdGoO8AmwlI9NHAiMp4PFjEMeaeyxeSo04
leNWQZVypSbGN+3suZ3XK24+MQofy3jg/gxRcuWH3iI7Klbr1ja2otXNzZWGDWJD
+3oBMX+HM/f75xPs66e0TtKmzRJYa27QzEBIR1xEiAlRL7/UiQ3kRP9fQfAgu1wE
0Qx2YfN/0saTI6Fefd3slARHIBuOLhIDjF6mnjOTkXBH4662O5cwV0ukNmaAQ4uE
wsOZuPvECOhJ6clw/SzozVlf2sOi9rfLSm+G+mNZsIfJWQylgr66bipaKV7i4pPL
InnxJ+m/+s64t2sgyWtiymLNj+L0nTbF5/ZFfOXBrrbcF855EovbBMinr5oURLW8
2huiz/RjxIrYXX7HSItFl5UwxGl4npPAQw8gQCPWV0Y7/caTXlGUgbbmRe3E0KtZ
CHFKkqVZ8na9PWWJ6CPwLE80bQSnNlJ6uJCwZ2F7GQC0x8djKfWzuFUv+dhPgHCR
BfpAQj1Xf+fIub3yNZOp1CNts0qzgeK7wlWNrhjWdmlqYw4PMbJPRL+vid6PJXaZ
ZOdmPXtEiJm5UkvTB4algADPMwW7iqkQWvv2O9zErAftVaZrAjCkrXHCBZI/Hyyv
5sfpoozGzw00GWpt9WCu8zofCcd/H2QhWlR6Fgeho9+9/aU9nXw0vNaVgoJBnw0z
ub+TzE/biFMZAkvxpABQgwAlRmpg23jX0OD8FRMZZ5wiQCmbV3wt/eUbIyCI7jQz
RTEXAGmX7qMPrU3MUGJ21DIbtlcvWz9d8y/5jfu8f2KxYxTnPv09fcSNgOwS+m36
3fbGSCWXdH4+AhMZ25CAw3jn6JoiMHNatq4rs4DWnj0xccWAP6eq6amqEP3gl/mu
2Z3dtRUE4Gv77Q+PLiFiPqkAUGkcEdGOudyjxJJmByPMFR4xm0V/ACwOMaqMAPfK
8LfZk02kWoryosvo5Q4rDZjHM8AbcRx2f3cQjFWllbzd5QTL+CcQD9gNOhR1zGuw
IG66mHYEsBiaWsAiNr8C4dcJFS9cJL1OmCns09eh9tWJShVVYWtwamgY0lVImWqH
ztgoZjJU0VabiuhIfr4UhYMG5hdJ+tvmqKBU2WO0u+i8PSdadt7IRieX1b/5AEMq
Qs3KUzs45fR4LA1yCgKDA/DCGVNL6iZxW4kVXr09o5RIiwzSEGO9pZVJGc9Ouaao
DB5DtZLP6fhzkfMmHPcFnu8fEDXP+4dbyGrFAWaPXElao+DpC+nHYXOzp76HhW7/
c8hrp2vOzEcMmcAGCY3ZIJcty44LYQSWNyk1D3xkU4YrbWwJEhS1jAFMeuDax7uy
jTOd0vOTjhjgLG9BW0kAcPdUDVIrHZVJ8sDgpj/EQxDDdDwqBYxNJK+wcNGf/Fep
3KOBJh4+O7iwL4wBXqJycllhKvVlmYJRMRwkpWvEysV3G0Cy37uFuHyBQGk3n8Ls
rBz20gHp2RCw2P06mIbDKExVPoRkZm+3tBEjnTfZ/IrKE+JBdfIFequxrVbkLRjB
aw8FXy3DByI3DgTCSnarPWBPMfRmBVW1uCxk7av6dxAd6Gdv219DAX18D6vXTm4y
PEvrrJvJU9QxIlQdrHA427QFQkdczVwJZsPKOx4OzYjpG+rlj8gVq/bhRSF0CSxp
d/YsK4tglpvVKNfTAX0/zsHBDVmmSXDYEEsuYzuSS0H6v/swNNONQCA5ouFPxtlH
MgE/fAJr55KaXNJ+3hq8V68xiteMbfrNCws1K6kwPJ4G0QS6U3dklGdcIuVbjtX3
3NQVFi3QvqkEAFBKi71Qg1rfxpB0hJQscLxYcHAkvLPa/UGRkWhtd5VgdWIaaZUZ
y4U8pnrZGJMauucKe82rNZ6j4HLlMv+DvdqssD9j/84LZAW2vl/ezMPnM40Obubi
YKz6ez/412YenIFnc8DcgrbQzlGN3fgCCdd5SF42+tEjdfnHQT75LmJU7A9+e7Ms
33AmDhm8nXDQQaVyGQWlUBRgJoLFGJUezKitllRJABfuh6z14ldB7Hvm3pN3F3L9
rObyvSVIi9uSL0fEy6HNypkjkqbt3gjTQJx3BNiIpf2ByLh3q7y/fpoMSIZE6E+1
Rbf/HQCsuWYouBRLQ/48zYyoskHJ6J6w9J1b+NX7k62v7YmupUUIbKWRU26S+QEd
1PDXwjPPkcmWyiy95Rrze2M2k8qKVL8RPzNXMeb61TBH55aONgf8JVPU+xJwK/6R
hL5hzJtXD4mbARMkNbAfDHUBTs7MLDrZ/Dq+O5pRPdntlMbgJVjRbWBatTSmVxdg
MoBEb5vBJsoIW+1v62up7SUcjcPxhek9Jk7gequqd1xmHx2b4j7ixEvsrpLpunmZ
egJe38rq19h2idBRRxarC7wwEmYH1VSmLgRsWb0vj6/6yaX/+k+DQ/j7AIgyd9LV
b7JqYpi/vJWXk/Yh+fVL7HeDVVVfA8COavuTfVRQFQ5JKjnCCErRx8f0yPpScDiT
5nqz+XkGSbydQHOl23qdamCYkLPWst/aqTiX2qJE/1ZXATgj53fx3VuXcSlmyvOQ
X9MASIki30zY6O95I2zyxZrCf2P9CwDv9NkC8S0wLhUor1B5eio58OG4ZyL7XQfU
oQnJGVPvYNJxB3uAinOopki5zk+Za3SjS6GOxIyqEqTLRvWGDIL7UqJXXp3VqkVE
T3dn1yB7BOdQ+etSGNpWkTeWMr6s+hXKWlL+o8xELa1OSrPBauUuTyCU3/QM18dt
seduxnbwq2VQyt6BDCHiQwyO5q1pdt4bqtI83qoCEdSHdoYQTRR/S1AiSxRdjNNw
YYLwlReRoX/MZAdhfhqYWPCz8Uaiwe7OLQrZNv2SgVgbC5M17x7djEoFNKAYDSmm
N/11W27hkEFCDUE3tNWs60EpQiDfZ9YM8mjYPv4qtr31eO171DWcHH0zQMFNsJij
2HWS13J7ObrNXvJvejuJDo3jJDz1ZecgZ7egmbVSlhtTPw80o6L4lyTjQKJOKoX0
bWfSjyxIOHsdgi2DLyugbUv9XwwR+C55UU+ZguvGhkLPBk8d7jM/b6KU84dQrTPk
HFrefq867xb6dGXkC1tv7Tn5He+bqFgYa3KX5gT6y+XC9q/Vg7x5DbE87Lt757z7
nyaNQTvwcAnOmoZJyW7xKePPNN8wyWb5vLkAgHhCg7kBbr9UzTucQmSwT+APNA+8
uXOy7r4iuJ3foWJ3mh/blz56ABO0zSQ28eYY6o2ddb29i7jnD4y3/ryFepc0mhxQ
npxJIR5LpYTelRahK++5IcYw918fXtF+XiofDf6b4eaa8Qh+q0BQb4fQs6soDRda
LbXlR6IDBCzsTrCYlBSUYaernGzNBaWup4BjpvQVwPoDoHEVHPaVmImrA10JIQZj
qPOpHqwXO5hQP81bmK/z+5wpww/feRU47XcVPfk6Db654DUfTxU/L2nUow8dFC9D
Q3Eq7rcYmvhBWXzzfBY/XfeuWvIBQwPgqCiea9Tdtqe+1RYq8sluLsIPs4c2BCaw
9X1Y9sTMIOl08EcRHGHoBIh4KhRQg928LN+4wa3VR+5LtgDHbYT1RZBciY1csVwj
rsrmHkRwzJLzqrFReyqlk7UvCZOvjrEmPPFxTBD4O56//fmL4FLxJxmgafErzG7J
bECra+9WpYAUUnnZDkgScIYJYAujJsqojpoMZ7bk5GIpsLgPcYPAaP8E3JB0Fj9k
KpvrGU9g2RXZA2ikN5yxqoT+BSZTefEhD8Esq6Ctedc2f2KqLmX+9PhA1Mv2h1bU
LUA2IzQbGJ5XMhWham3cudD95AMrqClySag/CakXsy0vQxK2JlicTZ+4l371ax6p
AEXboZVThvz6gkLOE/opYnavNGqMv/GKpma0Fim9HFH3NZCGg7JLn0xhsfJGjnbW
+Wfni3JCsfIDNdCMPbMOqKO/VxO+7YiivkDP4W7Lby/wellh/IJvot5eIuJkYPSA
Eu6u2DMObW/y+THxo5T4qAU5cCuNcABJK2nSvYAlz6/ALbVbqX9281TWyM8PWRCY
+/khlbPC28PRmZABs2mUGr8BWUiiedFwseXoEeAGnqN4OPIwmiuzngmxIaJiugly
CPAu/WpyCOLrVH/HHfqtYIGSJFaPCarAjw9qelODfIFRxSTiRvi1oqR+L4LJkKMz
iF/XsysSioCemDUJ5uQP4/TO1uZNGuF14vMHf1/zWYK6Zmot5E6x+rncCMjZ+t+P
MSL43QVsDFiae1hYpEy0i7Z7eqs/WHkRi63Hz+YQCzj2wH9Ics/0NlvQZB8lHhrQ
LT/U7hgiLZNl0yb1x1RtJaCrYzrvr35lUhSJmYOWuAmReDz/kwT6InAyKnlePU3s
vL5ObETR0g97vQBxk3hFIthdg4A+p8JxRZijb+3IWFt2t11ibRIlAdIaiD+QUlXi
wZezs1nIda4rWRIs09n98MbZgmU/puH2M2AFCT2aiWwptx5jauxqHHEr9JUA2Cgq
uQQT498uOQV6Ycnot0IBGtwO976UfkcAHbULes6LjedM9ME4r1HN5/GdEPDvgb6Z
w9XnIUrONvRn3dThjqBZxn+YPML8A6u/29UbkOySFmUwCoa6rDbLItvJZW2dR/WY
9i5FfeYXEjhv/O2tBYMERbkim1wg7QbIv/IkYdm4SWzp4gFSYYrKUyix3gJzNRZg
EU7Cfsc34RxNeyYORQBq83YsAJY2ShAkI8sfHuj+CRt2+ziEeWe2yxYWzxudRU/S
TGeSG3+JA5NXLw1152oqSVjq82BEbCrDxjsZMcVp1v47ZA8fpots/TDe46rDTJwN
8dNHJQwmMBGeJurvJj97kX+/AEZLJTcB6azi0XxhmVRwwCVqYVuLVLfzC5TAuOhF
rKprwpLmwY+OtHspzWSkxTIHurkrGPDfhErc4Z1xcz9NXPYtVk6SWkUtI4O8k7W/
GLBdCHZNolNbYgsWdXbPJK1+J69rCTcw5m3vmSAN2qoKKnsp5MbAcWJVDFnoOnXN
6OXI90HjjfHhY+vRKrQ7ht0lHn1PzDboFSHXs74FR4yGdBOTLTDNcpAsZZE4W6ZY
A/C3AM+u+ARrISLiPHarhIpgeeIVvL2GxAKjambIH2Nz4QbAzHzHCI/CS202p03A
pnoce80MUWfL7+BRIGbtrymDlXAONitw694D0AFNhQJPLq0gKWAihnYpmhZLjdpo
dXldHQrsFPBRFKyXeiL3otn/naPyztE6kOWG33UsTAUJHAyaKAywoY+2pYcYtB9c
HWc3oClMK2fX2JtMNvt3c2jDEgjT/tTsKBjVYn4GG3QfKXrd6yLfXvAa1wX+citg
FMi0S/pKc1F370qNDR5v8crK8E/OI7JuL0SVfnidbqS1gRdz+5+wPp2I1z61C7fr
CIt0t4Irj+s/RA8pLwigW8Sb4kopl3my6P5v+PvnT3RcU5uSWWUCh6otz8pBsckT
jK2IAHo/9l5o0yIpoKouZXd6aFkY0Qv3BTkscNNWFL0HQJ8cry4oCIhgm/kfyYuO
0G236bVMtuY9d0Ofi8eQocgXTEZ16Lcqjl0wCUezYvmdElR8as+zW3In4DgbQpD6
Xc5dPFHWi16Fk6PYjEYuWMvbTSQ3zYcymFkIHo+YzOPX7fs7XioQtW92nyEI0jGC
W7/MujPosOHxYcID4vz7MBeO7QXSX3qBkH9g6IMQecBeg1IMhUb4zt6bIQ4sSe0q
E1FAypaMHJcmSdJ3zGncU2foQm0ay7ctDci3lOOT+uPnSW8x+74V+xtr4IeBTarh
F2sMiDL+BS1lGB4mrNJE8CCr51tw+pHDbCRCHpnjMVBqjCclEmOWv/RDysFDWjff
XqACcM5SuLoXe4aZh/24hPlPW2jfDVWAG53xAUqYw6mN1zSpq4XW4BOG5kZDWXjF
N9gDaClcE/O+OcgHIC2m8DAqZ6rz0HK89n0gOLJDdkf6oJrOxs4ct2bpweMrhlnx
B9ytNlPOMgSG2HzFFhfkxFPCWp99j+Asops0UEEthOZfYtnf77/ex3v29wVeUDEq
ibeD6hBkro/KGzpcMVHnqAIsQXgScABjp5iKZc3DX8UC98qQV8W3lodDmkIyffD3
xmASArcSg+fnt5QlUb7ylwt95pjKFq2SLyk3QDp07lesvhjwUvSNOInJ58YzfIDU
FP4FTDj2W+x2XTELDG5J/zXIKw+cVeOED18moacn9oC9OEa11AhkszAyZO0V1Huj
6ue1opfHYRUBhZ3L1lhfuLARPFWRIxckvYnK77lqCAnCOBNz805lEN9yMYK1qatY
PlHxlbw1tZ4zk+M1QHMWq0ZE6nOz9QxkaYVBo1eMETN66AyBVlMoCmlPdldyFm2k
HF3vTsFvbsN0gd9KBRtf9aerVUw48WnL+oBf4s/5NV3uf6HjIFx/SVczjXwKUL87
Yp17xKn9Jiya6S97CKRqymS4/OVggWhFFjtgy020TRWYk/66W22tBRM96xuk9//h
A52xxaZsbDrP898flJd+ci6KU+rZHT3Dyqo5wpqSXUWA7wnuZhn4u3jUsbqy0SEg
Hw+0bp3MyKPafD0dnhEn4MH79pCzpxaoJV7lMMk7iHO5gZSACXqifR/Htol6Lcjw
KFWsILVC13FR1JyHLW9naDP9YHO7g6cy90wLMXHEQ/EDNVzk1Akm+of2jZEFihuV
8yuRCYsd/IC3qE8Vnay7WbBvx5FZ1j/0wR6nghPJT2TBUtEVWlE05VBt5ozgwU0G
izLcCOXGoTAlNuWqWY73A22eaI/6uabz/8rP7LdmNczsNwGq/aRiY3p3Wi+LLrav
rSHb4qibJSQ3jbbR5BHd6uXpd1ZG7zosND2TlGxAiLKndQDlOqINJPlCbtrJQUtr
jQOW6Xl9PBu6HuygRXb3xptaBnxP3rO4n20N6k+z+jkFmtNa4CE5FGGGMPBy703S
OWk30ClmC/1bKm2DJFsloF/Nev4sU7VLfucp6pES1Rle6G38LQTolspI3HNCHB5i
v5G5momnm9idTQ336ddf6iEMc02IabN60N6F6zBYG5P0/7DSOAONzngc3bVpHq4l
E7I+yhjWYSgDIlIHSuBTfEqFciZrxQ0lhyUmi9J8PXWH8BJTcAuuB3o99GOytqpE
wtF2pPIG/9/WDSu4UZP3M5boXBzufCb3stynTLH4FAcGsgYnfV3/UhKRNNqR/P2y
53bUSPr4vc8SL4k/qKpgecLCqOwy1bNEuwOIdD/Oig3ZNSG9LCZ33XguKCcbDSEK
8zX2ClUapoL9HzCI4HbZteSzHl2cZKKs6RUbumRzZLkTHEeko/pYaUbxZkGohxHE
DkmDdShaNODcVvnAV/7FaKZZEBtriXBi09Bhs5yJJQycXOy6K14oTSoMATWnjwwz
GVb11wETidfXwUjvO8d7WEAm6XcD+Kla0ZW6XAdBqysif/5A+tQEwcZ9wvzYS4S1
+LwXeBoHQz3/ry5RPxpEbMTRB3NyTAlUh9gjez9nlIIOpRwRN5JRa4Cm9zU8zcIb
esQMW+6IU91Xr0u6gj7cDqsxfaTG3p0vCX0LuS91IkTUsjxhaPMFYM9Caiapv8Zz
zdXN2FGU6y7AX0IsqEnQ1KTPpoOUVRT7SjJO4DzChnjbvCi93w7U7lpAqaivyfNp
oEC4mAP7nYlXkm8fnWIPnSyXcyT9DwwPCUAX/T7+qBD/s/L7b+6a3iRV7bsW98CO
+B2Fm4b36utzZTfXzYxPaQhpXR/5FLPjgZe0862pygeBAn49eLCg5B6LdAT7hCTh
TOkdoT2IdwiSYpF+JXCmh8NJJJhtbaV8EYRfqSkhSbZdvdTv9fNEBXV2JUsa4iPk
m42vzJT/VonLK18KzfqQnsSXQLgayddnLx0XuAlZUe77uG9XdVIlDIdmT/dOp1lY
MRzgQf72xxeGX59SMZoAeoNkkVzonEf9d26HYzZ3NpASyxUIbXhyuH36WJgnLbVu
CfqtHImYnViTDA3q4fEUxnHzNnSWVoHrU/1l69fBdAJ/Bf3qsgTCQ3OricuhlFhb
ZihM/0u3CeRoV1hiIflNT6rcq3IVrgR8AMbLXW0bLkhmqM7XQCl65N6rTW7DncwF
J/y8REbu8La+6XDYmU15rnYJZVEaqaudauUXY6SB8ID1A5zB11mmeCbUHgeZEjTS
jSxN4ZDwg+YcoJ/qfS/rxbvw0za84nsqlDKEybDiaSwhqXzHAju3pk2wgC0nJ3ko
dOhIFsbM9qy8LQ8GY4UXr6TDkXdU2f+2KY/zZIfnqJ58vCIFCmRdU9xjJoUFfyiO
Y8Ymi4EWqunx5fSp1DebGqBPxdKQ84v88fSLcRlB9PsSwXFxemf9DH1+FhKkuutw
QoeJzNrnI7Gwq7/prAVK4DtE33KfjPAWKzrNOadygclTesZ0d7slKIQ56bzHnE5q
SlF0UzHsdYS0bBqIx9TGCeBhkoY11uUNEG0w+ASx6a05FiHLzEkDhWvzAMPgjaP5
KbU3mLmhwfmcn2c+TvhIzNdpaI6jRgz14zr40J+12HM2hAVY+/S9bJMZMZrdf9PS
lCgOU+h+6CZ1Ap+xKb89E8huc6HcXLlzt8JNstJcT7kyO+e5mIgcsNF3ZpKVMwPD
l2Lz7rMHUVz/8wBR7tjUy3iM3Os/1RJB+N2Aay5AKyw0ThkdrHoG6S0ib1hD6f9L
qJ12JxdRsZgT1UawaD0CI7mYk617cS4CZAD0APLAbyluCfrOSYahxJf6tC86z+T4
EQIVKDTaxc2pMkLYAoJPKA9flqZSaakMsBGDGN/FLkAnmomFNMdLgcoZp+NFWlsp
vCiBkhQ+j4cCuNVvPxo/XuU7FDkM1B02jH1epp3q1BOR+BqGSBHMMfnGtTseezpF
malMSzAvUNBQcOWEUsJguDk9tA9gB5FtNdcy2jOETVgwCucvzsX6KBwFbEf5YlOZ
S6T6gCw88y8EvvtdYuV7Ntz1kP4Kj8KbGUYnBHfksOZEL/IG2/A0X/cfCLyp8KaZ
DKVjUnIAf5MNoZfmDxRDYiEpahMJLH6sVRgxPIw3oHHjgxUnzHSjgSnwx+2GXHlA
sL8uZzxGMOBHglwfb6+nrpBfWWG0xODAnxkMQ7LNybJvVNOAex+hIz17SiMJRTUi
XgEd+I2PbY5GAqJshUrmznri0jozN4lf/a2eshsxZudtxFNQmxY+sAsdvN3rUI15
tbsZxNKs119M78QGAB2iaJ3cmd+srEZlwr/4rZoaq3qblBubHgNVhO3LIsX0ouqz
2ccZzwFEZodBCtW1pb+xa5Kn0bPLw6ikQfF0mAKXnICKO5G7dQfZTX0sm47exVR4
dHGFgg7VAWqgtYYfTmqYxMGCp/Dyyt0z2b60dv8ZJZ6ZL2cXWIPBuXWHmFhxqPSN
LQIbuNyxG85NYL5+L0asfQZblUHkx1OQQ6J9asr1M5I8qsqNBIE7Gsb0kIiWoQAV
n8J5w+nMkZz7InJ5ifaRgOzOuNu7fUP+aor6HbRh1QDl3pACNk6gGR+PzhzTyqnH
fF8aryjkDxTIm126US4gYTgJZqwT+YJ8U4c8NKmoHkYElq9qrf99rob7O+9qSg13
+Lhe747q+0u0EUgXUMQLcUaySFls5ZgxMpAS4VCy1i59BxSrAQqaGV+D9zaCnZFs
RvSdcIYZdyLqQ8bDpqyLJ7DcXXn4qvVQ/akMb5NQ6Pl1pWTCul+U15a1kJ49yYYU
gAbDQeZy6ggbrB2GNR+jLE+3F6CUDOAmLu8BUykLVL6EcgNxDYSAFWRxnPd+9vxC
mfMrY2nmE52oJG8uNdgdA9F7d3noMeL5so1A/AuaOXt8BTMtGdiEWnbbmftRfJDw
TT/plf+4XDLYgcH7s5UTvOAwo65j/FKh8Ih7nkbp1Th9sA8kzq7me28aGYaKauHB
kv8bEjLFWP3fm/4YSyhGnZnJmFPpkQiayXgLvWhPzufIPbjc9f2NpHDXRUNsAgl6
JmjXMYTJh7N7So7TeronKrX7afCKwy89hPT5e6gLahEcxnD8/oylfADNTHoaceLp
/IEQaELWuOkwkrJpHdQSPgF2GwrVe3cAnhEIjO2KzCR1NVkYxj8KPHCl4jlB1TP7
qrHp8JYOsGHyZRMTJgl5FOVFyJZdzdg/kdBozMPoquesbnsl52vVZr/XPZwWmlYv
JEz5JYCc6ys5ZO1KxX4WiL04cb3XGOavDquthGKkXu9H5d4CzstLBjny4QQgA0Iu
o6rB2gqlDq5CuukuEl8sP5T0ObNLGm0i8mrklQo8Tdc5zKl/vEfWZzOgtp/Kk+JU
Wfts2UGABx6pZt+nnTpkkhR2YZ8+m6r2sHCB65yKPbd4/KGrUzWYAZ5Enm0PyDbX
8fbZ8NrItgd5eZN0wAr4pkRM2VskBpy8gFbllgeO0EzUql5ws9V8ouZKGa6k1QOB
iUVHQrCOzGmYhuLFyd9chvfjVL0LwjhcP7qE+zgD/BhopXHri68Ve/s8SPOB6NHl
goroilTwJbH9ScaPn5wKWHIHpVPrAHomKxmsLOUUjX1QgBxuRLfEh8Ky6Vz7K9iF
PNZ68wKc25MbrZwM7A+jz1kWl/C3ARZhYNDPr0fayrpuglbl/7QiudEtDlkO8Tef
J4FHIWfRG155MLpm2Ka0yPYKzfG0WRwb1Vl7E5Jtvaxyxj7S91FfKDMfa8ekNUuT
X+HREYXbyVGhMwiI9cUeHrSp9zxhzV0tHvGdjcW/vEmsiMqSCylqfHAtnO7uuXLR
7BWdoWW5FZ2HzKPsKsI6z7rU/4PznE5z9bHaDDYC5SZb4NX/9X4kz9CxzOezNV8w
n2WHDGNb8WkMyv7YHN5Cy7+idTnww84b7eM5sTzex0TbUBOhEBnNuVMwhqZgtCDw
XxjeBu0RxCxmoSnLeafZ5jntZV19HJUbJphQYesT4gO/SHYbxknHo0s3zv9d056z
eAKSKJqnlVZkrVHiU5ApMEq257Wj28xm4gBnJO7hOQqKyXm4xlmN6/DiGUD0OMfE
Oaot+D1cWl6fZ5EqHs3YqRv5VjQypfS5lxKj5j5UqcZAuG7Fl8c2Pk53Diz9iwTv
0YM02GfbDqWEq/HMiBvI8aix2zvBg2U+cMesMe5LOjhbz9FnoMKYnYUa0aAPZD5W
WPlSXgEZRjS0EZ2y0yc8ggQGKczkkOM+X3saq5MW4G7VxFkXLFR0m/ZdEomUxgS8
X6oXMrf0TE8XXb2c2Ph7r3PGYvfk861nX9hblay/Cv+kjVj0gssGfeHV5UdrWEBf
FIZf42wmZW7GEkcKUYyFhAtyHLN6Itv3c31Wn8CBm//dq4fKmb+fyKlQafGdsBLL
m2G4Ozu1NVFpzrKIBVfanHGuBV8eEzXExWNkJ7h89uAcA2M4T7meF3jqkgcyMEJX
z1Yi5/9lt5rY867s2MtNKU+JfFk+2V5tYdtvOUH1/OOz4ksdbES89nFp3UCk8x11
esi52hxUf5Sp3D5p94FTQaPbdUwmU4+rqvZjC2codEQxHt1OVyIwXXLO7QqKy4qW
Eopry0m/XkiYaH32Kc9bSGT5hlqSpwK0BAwTzrZSayLmSQmiDJS8/Es1mXJ05RvN
SAwfT8A5i6r6vjfVcWBwL2YWm1Ww07Apc3HVfn967wKVl+S0Mabntnahoj3ipqYl
5otUT7+GWBUn1PJ0uvwV1CYj5QjOz/WtvyXEEoYQzByUyRG/Jc83r+/WNn3/C2ND
B9AifEbhpdBKZYPoCEJBVSXj6uFihuxfh8cqWFYTudVqjmOWZYgjLH4z8QI0YDDW
j/1DqhxcSv1/8I/iMf7eP6a6MXagX3hwWt3y1VN9bo5x9J66p5xlvZHL1D3SJhbV
z2uvAVdXOTqE/GcLpn9PIBNfRYxPhKtM39HU2FnJzprr46SNAh0G4+F3H9rYJah7
YJ8StMb8biQ9uZzPxIl35c+81KJMWX5KkM25bCjInmltcz1/BEuYrcLqE9JE9MmP
I6U9EEqMb7lx6ZrLN6v7U8PND+vzq0LCoBGwt81rpqY/mlcVMyN5l3QU1NXZBkFA
m1U1NIuua1SubLcDXPDZdDUnb/4tfU6AD8LFqVgPRqg6cqEqB0tlXLLU3jHBArMi
y9hyMj7lLcqE3ja0j+9uNe+Nhz5hoEMmEk7p1xOfT+q9webSWgAo2vdi3e8/zeuy
jHNMpYCHTS2SHpyECr7oqG+/V5No/NmjOZMYdp9uU4MncJ1H4Cr6CIqgY8bNdqMq
X2wnRLMB8bwiTdxlGrPcm1EH65uoKI5BcKjl0eatoRGZEzowjMglrNB+KhujQUrK
w4SF4PdsPBtUMyPLiakr1FPi7M6PG/wVa7Nu5CuKRepOPtLWfJZ0Q0+tXFXwafR7
xazeHS2Cvo8xo5CdTfyatQoe1Cfx4zTHk2YL+dy/HXl08mrez0zjFY0QVm8hNhHf
cYlY7B7B6LRk/u/1BenzAi13lvP7xcMVWz70rrxl/hwAzEKGxzPnElrbvvZVGe3Y
wS3kYbtcT+LcNraM8iQN/3qjMoKVKzbiRaiSW5RjUqJ5pVl+AYeK7gT/ZiZ9a1RP
Q7+q7y7n0bQabuCzaGv3V0EqtwZYe165KhDghqQvK9k/fJkEQmuV+6ziryYFdPxb
mDH2mqLDxuag50uEvefBT5BScXhr2ke98gsC77UG4I4WJyBlwWpOOf2fdqUXVHvb
M2ZTQfC8EgAT3Yvf+qbhsuBLltlePJxmZIzqOPhQIDBf53niyvizkqDrqDgW7/Vu
InBgFs6v94MVtS9HmL0yxOopC+jo0npF0+gmcKPpaNddLjbLDTu9MIaImqajUTCi
FiN+iyQAx6xFSud6jUDbcncxTaKf0WQ1mBPn5aKGCf0+2pHD5f2pXsiCOyjrHpxb
NY7CGB95Nirx6/kSZ++8iGrx6I854/1Bxx0K84H08CNRr+So+o7a7BqC3XWkstqe
ArxwMJDJFNg/SYfn88nKM4gzhSIZ/qFxokLgKXNjzreG0IdBu7ys53+dZl9ZP34+
K6e2zV1xRRlkyfxn6H1R2wD2q1mZ8hVFgpu2+D/cFoZR7rvfsl0zcjlWFUB2ftMd
1KkBjuSHngNF3oLjF1MxMYJ7zueq40d6A7M6c4SDtvfr4LHQcHvoLbz3MwUpGKOn
r1jOyYNYf9f6ihN/531Jkof1vNPTh6LPa9dsjGutOzlKT3XsDgKSLowb9PFUuBol
vqdTNWKUD7+cj0kFP+prgZTCWlHw40DYKuxaapR5IBe+1ANegh7yovjYNm1EEPST
wr5WGr4YwApKvevXjV2NFS/slguvDvbrbPlar6vkl6Ya5nF+aX4IQ2artIxq0fYV
EQhBkVcJ6vdu9s2RSrqwOfrkB6w+Iv2U+j2B9Bit9XEDUYgUKqGG0048Ex4PT9KD
baEiWdzKcnVdj+XY1eCCksPDEm5TNSZoQKcm4YLSXTbAQMIDMoRQFZZkMv1xqF0w
a6LnVcKs/eWeO+P9cJozA1Q5q27c3pmFV5v5AnHmwZ8vCUy6mWzDCkEsiactcKmz
3zeAP8naPlTB+YIgBoUtokM3JrCqfnJHiRMoXopcb7q/AMxadcxlGif4I8SyFI6j
YFNOK3VhDjljVNN1eEfmrFgxCKW1rN4wnLFxRBsrZRLYLc/NPTyPCaMR7V63Fmpx
v2fUgOe1ydy2pkAw2IEivqK8Bgf8cQSzfppA4+YA4To1fT+pRNeAz85CCXs6P4si
PZjYEc9YjsrrZhEYYKAGcvGgZXHRrVDZeccTLF4TJRaznOXnMf1pobO3ppOjp0CS
a1vSwP2mv+sOjtlMrF/Lk235LFCqGJG07126bMB1nTj9E13bfvl+UAOpcNLefQVi
svZXey/qN7KGtUXB3cNVqHfAVL1pFmwSONeptqwhkoio00y7IshoXLP18WlVcQ6B
U34cdsjUEvIXtySI/s0Ksw5Nmd7UF5xEdp4ioOKR+x7A+ZeYn+DFzbZCVIvEwThR
MqaIG5tj2GlT+5jxBZgg3MrvSslbu9gDdFKNrEcnq+C9I5idl9SWFBrZaaxXFkoD
oUg1QlTvQkG9DhWIjusN3iDl13AaPJ0NyNBqas7Hb8IL2WNCiP9Z0KRLrKjiNTcP
tAHtMKQteoI1JZouXKpc2KoqeYQD/BatTsbxP5TszBZE3NQMwWHlOMW4pjcsTcLB
VTyusoI8r64VhOA+18GqqwYaDVWkuTJ69jcITUeR0KegXwkPkeO22DRhG9KYDz35
zAhP3+8eGWQV5mZBcnSfu+YOF4tqh4SAMKESTS63syQo72/Ogqlq8kuaItPv+1L7
taJzlybRItpBx66WeqoDSziUWeHzNGXgy02c7/VbW8A=
`pragma protect end_protected

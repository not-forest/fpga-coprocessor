// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
kfUnp1ZPjtMIJ4TZdHNeurkXGmKfAPBBhW+I6h406qJasnLlc7gZibAFBLqjsBrN
xxXc8XQezXkdUyq1LIo4E3vTH/ajqb1C/DiC7VPrPDyIBGTTEU/6qYNhYFrpMhJk
s/kJbl3qt2rmusfMWiYjnPd6vcC1tBnSvYqpbvaH76U=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 9216 )
`pragma protect data_block
pfckQwUTbyvc4dUsHpRiVDTHs14sWrbv6iS/XYlgS5b5vqGyofsmmkWbKZO+CPuc
q5KkJ0caDlzEWZK7FvueL86SPYhuAAzbkgeb5F+ex/13CqyvpS07H2YF8lglcvBQ
958N3RaOmd2n86lOEYX1BYAo/MSkALYmWsM5JjQ5bh1ZbqLrhD9VxwKgUsPiQvus
hfuiqyyC4rM3xlRXjFwUKoF9X9n+RbFkHvXwvx6ZDm0jxII3dtnzNtmsKEIRwqyC
AuJQ0PaPfCAMsj6ogdIhN9TZ7IMOIlH2loYwH133ceYAq5cx4ufIFNRL4b87r+cd
eSieZHoE6k1Y3l/dRTGYWK4YCQX/g2YWvlPtWKby6N0TRx+s8zjKzGn2o4f0+Ykt
C1UUWz2vFc8spPQZfrU+EPAJ3gr3tE+wmp4eY8P3RsV0bYgUB6Aog4HSaA3dSEzM
jHLvY4OYmcNxpjxi2Db8q4DHDtLAyxR7LE6UvMCYPC97IiUqv6Itr4bM1AOYdKts
ucekdW9NXBJ6JImHq/OlHn3zW9TmRWqpx5u/49PwRrFDXBtVl8Zw+uyjhJOZopo7
22R4LzgnXbzWPnecdjgZ0PvM0Ifi5Hq60sKuYOB5mUQsrwvUJfnl1a9C/eytOZHv
XHRSiFNhl2eu3Tsot01tiaZFmK6yFtzkCDrR9mjz5RIlDmq5Tq191lJ11LPBtN/k
DJwUje4BT5fO4/CLWQXHn+9e37HGBirRfuVX7GYaMyl2XJTEl3YzPSAORJgAPC8/
dshzG4ceQ+By8NDFZ5Ua8zr8CvCpbkB3aNLYMSncyut43WN9w8ieeRfu9BW5cMj8
PaS9imLuSJhaacr03FhnTbxG1JJgvdZVQP0aWJ5IcyETQTg9NJZwqRGZlBTvKKfG
/rpUuebWcV6K3zbizn7MlfsOo5UCzQpJIQ6vZJ/X9Nrvq1xMppz7wycnj310jdhS
ARDWaBRKiSPO9qoPdTpYaGzzWoiJExbbzLlaiVXEp8d34+Wfl0BTeRHIDnbI+yaJ
rwzZXMeDfeJnMBKQubYd3I8Olvw0Rhd1E6GMqHKiXVIMw3NppSUBk2H+44HGySyI
4EnqoR9ZeXnSiMAUz6s7/1ovY6HCQZ0NrJS6L4S7e21iaTGUruk/PLVJY2eIabKx
y4ztP32b9327FxN/cv77kc6/v21xM2ghCdOQAKBaTSDgrfc/rV/xoQh1TovRclVp
fQPybEW4Io20cda3eR2e4Vav5Li213O9DHFSC4AEtbckXV/u76HCGF4YfAfbC+PX
/erWQQQWgbqdlPrAl6sYn2NuILjMgQJO7Gvp9fFxBHGq2yzkQSI8Zl8O0HXyMjSP
cyV4bJSK6pCXcUBrfQ+Bzk8Us4auRuXdtzMaC+kaBQwDJUuzgmzSPEpqv++S5uA5
cj/zu8Y2URMpppYJDflsONr9BDtsoCl52q1QCd71jXeoO0dqyx2lYyp2DCTeppwr
L42aQuhQF+bs0cX12Kdv/vwIT+YaJ/PyRxd7k46J+sTqzKUPoGFkxZ5GXnm3j/jr
+ixEPCloeDLo+z8EU16odVlF7BliVhkREQW26RaH+tsGXB3tgQ4T0N3dhuUQQVVX
7b4YdfDkivm4YGU+jbkO0OOfjk/GACTC79CXB01DcgyXIkh82Rc66O8CeTPpj/vQ
r0oSEcFTQ5XoIcffL/IG/E1+bDWMjbga64d8K8bPXzNkitU2vQQWNFVB1uUsR+AY
S2eoCqrfjCIqlFe9Edc9P1vfKYDg1AgbLSgvJOnK1Pg3s0k+GUVaLegOhd2I6i9j
ERLybyC/jg2cgDVypOFcKhQwLosixnmc6VAkkrKELx//aZ+fPvx5HJgUwocRSEw7
/RjAmshilmq2wIyR7YjzbwX0ckwiKJg8UBUevd7HV6LHyn1Wi9XRlhchhH8A5nr7
XeAV6FAyzkV6+SY0QB9Ye82XXo+fg1aYQZtE3UAkVMw3xC4DL3WnEk86luRrYqyB
v6NQg79TCvoIHmfbg30aGek33plDVZZ+g2O1XXIVhS0+WYC5It7kNpD2+/foJeY8
ZCqUjptqAtymeuxzlCYfafAq/Ico3ydPHpXYiEzGT8PwubO+aZ7HtZhsWbCzrkzu
PZbsSsHF4+sCr3v0w9gH1wJFT0I9qYlHUjiySiqAv8hL8UkFntV5FfmC5uaG2TTc
8igfjBdxdxQjPrlvR8h37Ses/RCbfz3abWQw0jeGgznIiAO4SW/H/+3RmqBgwmYD
z1iUGEmtwMxW7qQkBnqIr3qFFjwWpD0GdmfiPEGptoL+CuZJuioXo2Vrb9vV+qUz
hxzPSuT74DsTn6VYF/WJEO3TsTcmc+nUqwFELpTr86BEGzEmcjW1XF6gKAaxAL4u
BAyeS+yPbjBLIGSXPVc91lVGuJcE4tt/3/HYg/UcZ2jQLhJ4IWYBpT4XzOqavfSW
r5TKHGFzwvVBnNiArxSu1nYRmn/wJo8/1FdcAKgUNoMd5yIXS/7lTuNYF0gU7Dny
VOVbTLHut1RvxjR86LyXn+wJfWO4nr1wEFFlyUMo04Mp3DOAjyCFU0yBZNWBt9Ge
JXfTL9gIzztmQZP1NVjVbfi9i7cVUxmGbRdg1oRbCng5gpaWuhSY5PcKXHeDnBYC
ATPDZ4VZ9k2X6EOLPGkJTBQ+Ouhjt+QL9IyYXRtfX7mQI6IqHPbHfaDA3mnMajgC
dKVlDMTb1dOebusZ3Ei6enlOC/lfXEiRQYz7F6/aN5lLeKmaXS8hGH5MedfdV/Zn
HVn6/JRlA67M/I61ISpo0tr40M9e5x01dEM9P7NQT3GruGbS/XdYEbYIvZazs5oo
kZdcQlqFPhEbG5UN7GOLv7dAcrtmUxcHgjEYKs/UoEHeI0OIG7umdJL19NL8VY/z
I1MmvsFqUDCzrzIwq3Iptk2Gn5Kr7+IRq3kWUU4QZbhu5RRAtGU2Qo/fchP8tNkZ
qdxFsUkYEusBkr77E/I67lSPWeDQlY1XLh2hIXsy9MJRk/GaggcLnhTQ7usNbSBh
5IocWI5PT21EcYeZIzlWO0cs7uHfgw1C0ga+6i8w3MdLMN+rLaA645lNiZ9uoaYY
mWQl5tTKJ49mrGStWqAZLX2+DRsdgNwg/omW3sFeevYtUn8K9Uwp+ykKdw7kQ0RT
nNjb/Hke9veEoaKFP5FSogB41mn0mc0btlBpgn2vy+Q4RQNQ+LvMUUZRMOfw+mvp
9gwOC9zSYmGUeoYqrekDk/ikJ9UPLqoQFxPWeACOUOyVKjwD2w1AjMVeNJ3Fdviw
9hqVZMZw5fQThXkZsJAxB75YQN3pR2CG+qjRjmEqRCPjDF58WCylcyVC8QP9vpKv
Ir3v1i5VuGspodnPCSKFJDh/tGKKXjyLzVvJCUlqePZPG/OUnEdtOlzPM/gIX9Cl
Sc7rEs1Ank/NrFTthjGDTk/Tx0pRAtkbxoC8JmabYz2WwAHKdulbpaScpyc/N4p5
AZPD3edDz6v3q09Bnv0D/EgJyP1SQGFvdaUZW+kLl/p728krijxl4xvwqj+OW1dw
LQxezu2pU6rcJaC1069LI28IzoJFrsprq3oBtl0DaqD2nd8dkCuTud/JfoZc87di
OYQyI2/9ZLIIuwMLzGl9eJsNfOfAxblPSWV/XmzvesbSyw2cRn4JTfd+cirJJtjn
Dpq23bpN6reVLLADGPEn4sMRWBXuW9RhbCkVsF440idxlE7+q6FRwlIK8020UaVu
aF8kc1Ffm18ORLquPqurbueoQFBWpSfgc5DL6CDLUFUL4DCj+RBYsPYmCoPUkkRn
VMVcnhWRYZRO4GCsTwVipxb6u7BUBYBb0b0JLin4m41z5Ea6LH/N6B6sUBtAf66q
OppNPfkmz7cEpZW1LNF9z4tYKCQIZT6Bh2FjFu1bfMeawLOrQXNb5rEDs8xmVRAi
X5r61k77nlL75SX1Q4SomTHf2OKHd8nSUl0FqRNOKs8m1ala7NuYwGk7uRWo2Dlv
Z7NnqGLymJm4WMnHhCYRQylbElzFizx/lGHIt4/YRAc5MgbF3Xf+Aj5KLQzi5yfM
+CX07oxhiq06OCFun4dtYKCurw/KKXsA6rI59Ah2+1S+1YD8j29VuLR5Fgf3LU0p
6cvyzym+cFoc0PlMAjSWlS0FB+vvPIPRCbvZcGBlW5PjFIE9yXvMYtUNkPUXbO75
JqRe6a32+S5qsCE4mLLoyFZtgKp62XphjTei/ENnBaTZcP6FKHE/BF2z+L4Zm6Ns
TEugZNY9unhCeQggmbzyFoMjOs6yzKkWcQp1odufMqEE9IMGRRXWO3L/C0zMdESn
/rY9I+zdVGNF+CvcoPMuB/1ixnae7P29b1RgoRo6WrRs/e1ig/eqBh5akn1FkIYb
p6TMcYOJY4x6G91YTG67Zbd7oaQ3TXdaVHjHLE97uIu7Y0tQMbxhckkB2qTIaMjK
zHlIyxDTZV8Z9H0AIWkfpcwYyH7VRkEPpmuD++Y+Z5fEcifepG31xFRp2/qw3MNj
1X+iTa+PHweBYki3eVTWCoJmya9GTOvucDT1pNYNWTyQHNfy9q+IuG880zDzXYln
V6pSlECb7wR3LQ1fgVc9I1NAOWZuTtDf8xIJscoeQHr/F5o8exLS9DgABWhQaStg
bI/9WMlV0S3AH4NMgTjGQ8A+mUz+TkIv2MUgfAww+eZltqLtC1e4iAcz5SY+8Gsh
3qHevTGWgQolJQSND7hx97VYruyvSuXklvRRu7JhHwBCj8/MO13yghZpX/AX1lp1
f5z0R7uHHnQ76K4Xu38FxHQ8ytImhhO0F9Bl8zDV4nZbxKDi2/mNvmYmXTXTjc9F
rVQCJkwGLlBwmugH7V3NncNU+ukvz7BgGXRF4UOi8eE//7P34pi89BoLxF+ALQLO
K8GpDs52WDN5rlLloCBVP9MHlTWAUB+p82vg+VXm9CGPqQBoYMlZzuPvYuCmikv/
1an1icfMhPwu0LDghQXsecZEEznXjTkZ+ekEGfonl5ErOQzGiEkWXOdEkSYYoOvI
Lc6W/QBFSt8Az6sB190aPBUPJsxnS28Bq/mpzEEz2/JoKEofnujoOsoKHKloLXpp
lGSTEZ8ysoqDN7elZd1FPdY9r/zX0r1JqPITK+oC9MMZUknieSbMbpNIODyyPX+0
GhQ2vyQQcmNlh8rIdSxWa8NTjyCZv0nJWdjdhQ7QLDPpRE7YsWf7pgE6JGqmnVZR
BwwJ8zLYGCPkJ0MBRHJYTLQlLvk1fBKXTZh1umovAAgf1VQiXnTzw2VLmwj0E/1Q
KjtkHOM9pjbEzL6QQR0DMAYl1l+OR4MlWqaOvRisXt9BeJ1q8teV9/v2O42y+GQd
ugEYxTDmbeiWTnvsNUhE9Nok2SJaQIoJ8hjPgNWgcyg8jIjjg24qDCkaEy5wdz5r
jFpVRhSO16MC9wDzromkcNI+oo2BLLs/OHf3tG4pyJGl1gfBy0XNlp3TU2jmqhv9
SogLIAlQ0PAODsu9OkWOcqK1bCPQgZX8iIWRK4wz+9y8FtdwpAs/jAiG7UzxEGji
VWqagbsL8ByzMWogrrRSr1wsHVcL6UBDlGPrOgBSqG3QHUx1plEQJo13JpOA6jb1
qGz8VkDClj13XEWYrUosaW5qKb5BBGVMxB8KquDGjp6bQjB998hJn2f74Azlm/vP
mNSOIUkSZ20S6ypjmggV5YplKAnkXWoiIBcz36o2riDjk/NE4pLOocv1Kj+AHQd4
rG1Wq4FcApqd+OKlUM7HpYgPTXOY4m92q2RvIZEUmd7Z9ROhl2E94AOwc2dkwjid
MrVw9z3dAYXRQ4Surk4RHDvo/owSsEBqWM30Yh9Np3cNigwRS9lt+Fg8SljcTODA
b8OG0OGDJwLqonJgWw/flzeLXUTa30g3dVhx5BSLqaTR5CLfk2h84f3uoKIRht+x
lfN/usZmD99c1TBXiFAJZuZtAwYgp5Mp7dskGCk53WWfQEB24okcYSOPGH/12kfV
SZ7rP/2aDUEW77lyGYYoSxeVnX22CRPZCObO2lJKXER+acrBH4//GX+egeOKDZ2o
0G6d1Y+7Xw6XObZp6PCs+AM+beIOszHPATogBAVdAqDqB04kRQcpP6POwUZZ7riJ
Eqw7N1ZFnF9ELvMMjVo8m6emWCOIDuvab96/AbNGho0wTywVO7R9/NTKktwosL25
IWFw/w+jELLLjkZOeCMsF8r7TshbGj9BpnMy7LKNTuuO/bh4kdDYKqcTmdmcDz8A
a2eQA5ThpLKMpq7rPXjG3MV2NvJ7thvZFFKBR3zWwWNHSeXgN/4jHxzisL+kpHv8
q2hHRMOnXyx0P5yO0UtBSNj+ySlGc64AVXDRLzpvjQK/nf/TNf1CCpqISe/nLKmI
oQGNVRGktleyJbF8mNAOIwSF0fPelMjOKEGNnfrXMZ4SfflLNV0+beXhbrWnvfkd
aWBBIx2Z7qwF8qZpLttVI942dE0E7QRRlKa7BNmsl2iRDnV8fZiRSJXKLJVcfn4Q
JQ6BjOO8/ouqBfzYsdDwjRfbH301ASpsKRFOmAxSPCZ6hx0cKehhdVqhmZx0HaR8
AD82u6tby9C/1ysSmc6XzS26DLvkGylZamfuQHyc2PWs7mpQGPfXtUDW/64XZIa5
4uQeqfM0JRtfjg/NOW7F7O7cSkluhppiTCx6WojZSNcw1o2nbmVZmY50XRQoQJ2k
SdbDhPf+V9guLRETRht11wE7GzLF4O/uutdNObckOkRC1ODilrLD8EpC8rB2MIcR
xYKvgUF6iCFMyYNn8i4u+VEzhL1miONWhtnSzVSAtdm6ot4yHBB5V633Jv8+iW6n
YPLptcK3rv9pDtgXjGgkyxEIvNAx8Uqb07hmK4oe3iG27dAAZoB1A7elJxxsxsJF
zPPVnAZJr/XvtcwTbz52d3unb1GpkDrdAV7sYM1Q0wghe+9aYjilNR+u0gLpxtmo
mUQC1lleORuBmlfCCR5/KbmzblduZqMopaee4/waqbEQRRSny63ExnOE1KSn0IGw
c1gnnxNhkQuNdb1UBvRV4m7Z7lzamC+86xJyaTw918XD/zd52lYrNg/MP3onYbij
TWIkWDrrYex1aajGe7S9x2ozoqN8sDWplszjrpWhL6YsT7CzphIA84QTdmCKMSJp
Wwg63ltMqHzKuqer7+GkoZjvC0OUsl7Xy1OTjUpUfvke6ULEu00fzN8BClg3TPj9
y12X6GfrwpBvPFt4Ab1dKh5yn6FoHtmOhq4cXU/RzcCkuxxHKON+OnJiqjF/00Uj
tXkHn8K94xtSO8L3uIguSeDKUIeTd86arUWlulRGWOgeQikHG6lynqaGRKNotg0v
6pIJscskqgWRmyOZiFfZspmIQnsH9HqVbR0xF/MTUGfige7X7hM+BrGrKbOkwNuB
D+HMB0rv00Dx49i2hpbGe5vnq2+WFjvYBYMCcExTXkpcJNtR+GpmwKxAQ4c6RxOx
9KbYeylzqMMASB1mnYG82WmqPyxc+qUi/zsWlNBoL4e5ExKeVVJ61bnPLs6p3EMy
RBAXL/J44VnEUfekChMSFUrcMs6+rPvrAlQEdJQuWDgsipSsnI3ZDw9itUtXHS9G
tSzqekJ9F/qnUyR5pRbYELEF2xj52VznKBK6A9YkcPq3thWPypy2Z9L0Zg+8UEnO
jiMpss2pg6H36XAyJiLIIOT+1pUO6V0unWfKzvPPeSGcGhYPD97xSLyVOx3+jiKg
RqWN/PsR8LQv2zqqu2r0J0HkivjlR+Ak3vDqdc/6rxoUE13cTneVhMqoVA21aMyF
4J+KTToeQDu2sD+eeTjuAfcCZmNd0W2rQb8QH8zsdN20tcI+XW8IYjVH4Pk6tvXG
4Dr00x38dVviE3LIQAT2q+iUnze4uLalastEsr5gBmEpThcoPcHvYR6tzfza/OYR
sS79e+Ykyx9K+4KXU00TtcEKxIvWP9nC/ro8sjkqT4v7l8Uxf71PmCsyvUnHSoQV
7GjG+mD3pjMUUUlopGlf+EwyWcDzgUTCadM7KKVEjSFFSJiZMmlu2MOPipv8reYZ
Y+/TRLIwa+9qR82CK68IDmRstOEy2iMyNczNgaLr4YaPSFXuG0JD06Vp/8tZQlup
ydRTxn7A30u5oL0tzAcjcPOgxhah06AUwaegCyzdWIrx6oAHTw+Zb7YvnkjhyGA3
DqfrOLoTL3KPYjXj31mVmO9oVvOxIP+hv0prNCJ9mr3bCxRsTsZUMAOEvBeil4PJ
uYcyz1MS/DYnvoRCWldO7KYBNwxDTEb6MgGtuKuy4oN5owtkG18bA30XpGvZaX3x
YdlG9vR+qrOT34AnHaaq4Fa22sMn1XwUdWo23mVLoGkJigCJCt14sTRQZUUwUw1a
QBcZJlbCZGtEfzp7rSxuIXUoDEy5Y7HsNBSRuvcHxe4Zt2ie8z8EGK3dRlGWwveT
uBIJm5plRlACn6wFcEyELBDjD/AgZXcFldwKpyWJGlKD5DLqXpAz3jvc86fA/eZ+
jk2Uet1XQE3l1cuTXget2+lEdaoI9Q4cHWEfumhhuA0I+D2c1zCkQg32YkOKZXhs
qoRciz1LY+d3289/EcCTxO9JEJx7VmvWmtDO7V6Plca4OKYDFEsU4KPcQpCT9jcQ
+xKkmfBVu3BcPs/SezNkYH0N0jY9R1wCBvHEEEfoDjG3r3xB0nv50VUP8QtAe9N9
bMRRiG6ZestdXqH9p7UrS4ckWk8Y0y370g9WbS3Dsg4ZJIuo6622POoIppNmwcnp
MrK8Pl7wSkmOM9Ja5K49TCbfNISvfgEJ/sTEsHtHETfQ8XrQyOWZKCcDEgsMxO0A
OYh1jsIlSnkXGhj8jJ7YpSz+cdGw7JyQeiEkP3MP3OY+ItptYqp7kgsy0vWmzOus
p//0SvlSLANCsFSw2/wjM8yJBqb1CFQDkFjEamk5/h7+RWfsr48CLC9A16OXp/Mz
UNRlSR+JmklVfA4kE6/9KbBvRePrsMQ33CJJHqNLDXOFSRZsjH01f1KuHKXupRZT
xh9VUu1UKd1A1YJBhr5EuJUJaepzgUx5dvw0okb3H0QAH4GFI8MbGkFyRnkbhI7y
biUJ6PTfMT+CRlDX42UjgoNW2IN5citJcjQULQwoPrtgOeKqUke7GZuwZ1yjXjsm
/HP5C1EGgslHl91TyYhZy3LUisN+x12d1OIuonbup0pkcSVxX/5ivdMW9VVhd3MS
cmvWEcmpq1RtpLZ5mkCcIUk+ZzZozI6jHuPqFQT4tBvpmyZUOu/YjDX/CK+GgeMY
aXq6KIhnnciO1n1UDtvymETid0ykUbHmCmfJXCuVd3AKKmSLbLMe7zDRqvdXABrj
HpTf/p8CQgJnRZTK2kEGEKA2EpoXctOFza4FobiDGZeu2Ofr6idZTJR21ZwumGGe
V4853NUbJc3/Fdr58JvUT+7Xr55lkoKPF6285oS0b3S8O6axIF+HCm+ZZ4npaYkU
6KdltO79EuVXjrGWGJJtnzPyPK3ltAS35XzeWm9B5tmfQd7nZmZOm8FmJ+c8zirC
heG7Nh6X0jYD7E0NYT9PDUAJnb5Hqjpe7uihcnu5PknF5x1BOYq3L8xts94gW1aU
iTAc2yqvcT3crjJAVxLhx32jCxOfXi30jvnqsYVJ8Jd4GcrVbb4fy3/9iiF20bSo
DxF68g26jS6yYdT1avvdCwLUALeWJDwxC9S47h3ew7Z+Q5xZQGIHEMScqm24qE43
wBe2C/PrV096ccGhmf/EsxuOySgfJa6AnAgmOF9PYLqqoIsSsW0YQRIs4ALVhxNx
riHuKPAAgpjZEFijs5CvLwPZj57iQOz0/Rh9KPHeln2aPsfcP9peDVwdUBOdcilV
S5kLdLdurESNZ/dwM6oL7lfx1Gz5VAi/iMNQDit2kuO0xomcGkAIioEAJvH0D3Ef
wxsxyjfHLEWV+QoVobgy9Prk5bXx4Y1LceQS7EKPlVLF44VDgMeE4/qe08uEqY0K
RlnH2qdwjTbnHPNQUS/L9pLoE+mZPBPShgcwCkKyCrZwfMXMoS6iRcYO1fbteAD0
asgLfT0cugUwRL6m/sfT/Ltu/LqG3QY5VB2a9OaQia62ljE3RZtMLbDVDJ36WwRE
a7rkbso8DG+Soxwz8y7lvT5u0rpHRPRhOvYWt23dYc32WPMWO9E9euhTdm+o7+Gu
8GQZBmmVEPQAQSRC8qq/72gaU4yo8X70ln8AQDL9TjMq4N/Z7CnZhNURDtEmKaE2
qWx760mKBqDjJmjCwuLD+8DWgpXBrik7N7D+ZM6cFxsWZjd6RwQx6CnzrhBAW6QA
nHjq1haTqOKR9QrK/VGvLuWpyivVtpSYm2D0k6r8xYpiCLrnsLzPcTqecAabrDuQ
Yo7bgziErdwGc7aSkWN6FXwQ/Vdd/nY3J05guclrPbzDdo9kw5QK1Y5wK0Ra9HzE
V3YHSHMR81V+ztgvC3Nk6hfR8o8SjoL4kYeeTIVrZOQFlZQmvUWBGVzLUQp1RI/n
Q501Fr9teCEbdvhU2rRwSVg1hzrqQzQYir7biZQCw3Fo7wH6PBL1AQuQEF1LJw/o
Kc+y0dFepKtA0CvRtP9pHP8Tp17FvSNUGL1NHjDXlqG54E8PEwQYiFKUvvTcCs99
IIw5EOjbUrBpqBuOJpm6BrNUoqheOG+Cl0meQAoQw5yihjqylcRxrB4AaFF2f1V4
eGY/ammaGH7GMveGAuY6tmQKI8RUOXa5fSC9kZtbkxeZ9EWLIlZ0IHnz/2wClu3k
OM7MavvFqJpROL6bnVuLpRyov7/RsIotiPcFmBv5qz3mzuCIp/+Vy6pP5Cq8yyVt
URb9Js6EPFz8GYvOpeIwts9t+usR41HJxLVsfA16WsVo3XnQ+/HCb/E6BVkvFx4J
yV0Z4EW0fDYju928llNCLnxjO/nDF+rTfL73MWmkOyLZHluVzXatuhznof+nifPQ
GFa4nhi+oOZHiroNzjJ++aF9fFmhbu3y8YWIR338JZqwJqQqkf09/TQ8YXLiUsAb
MeOPZHnMvdPOG8xxXojo/LSJulEXoiSR7Hp9lrFsR6QyldkniODyTaWsEarYeEEo
PfnRXfvXT1QE/jIDZyN7nMD5Mo6Is40HIUhSnws3nPb4ZLKUhis6XAL5GHoCb920
ZNvS9wzwK8bQBCOWVQmGkt/faYmAbpiSEKmrXUkzl2GVBIZ9Q8VfpCp6ZJ0gdh+Z
pd/Mw/rYK7c6rXTV6TMsWpU1+oI6s3fPaEiozyKFWuX+Qkd/pIKREnmAItCKIJOv
i+QbJCcov/qtVQqSBnKpEANX8bzB2ewLont5izPX6uBj1hh3HRropL0sBkH6so3S
Jup7dZoWR55B5RN9uOAerOvifqnayAKkpcC3sLs2zAiQWVQgPqAO25TId4Xw2z88
X7Nh040Dn4e+VNof8HbdqeRC1/FOUltSSLh5rNZjSEOkOJQ254XhoZZDbORZrk+R
P/xEtYhndAQCkMATS+GFt731rkKptdAkeQWXL4EX+zHMuDjEx5YDSS9AYKFcmPrw
frWlvyUGM5w54yfROGfFZBbCCmWC/P2AjpuhdRPHqynldPVad1aEYzL57U9pu+6T
iWewlsE4yLdEBpdpPfY3f1iMT5jJRyyuyXOUF+QfWlYNt40fJ7ms7I9DubEproAB
dEEs9UFaDG1wXRC0NvT1p6Mt+3m1HZegEz06cUakcfOxBu13y62D/5vua+uJjJIx
AoTzvGRVii9g/I+GBU3IIbrPlMdnjVWe3acDF7V3FKYbMJwyWtYKoHjovM4DpueY
f6D/7BkeI+80dq5At+K2wz/RPCRi/sn+TrTXdbJCUvC+xKYNAwF8Mw7cEMnxFf/W
BWbaFf7bIcakvhIUIri5p4HW2eHJ5+ifRFSkHyQv7lq7IEirmRl2Om3uSH2jlKXz
Sdq99ns/GVB043h2uU6pe2D8BJkoCje0b7DEbu2G+ovNuoDy8T39akST5yxhpHTL
sokEoiToamYVSRCTk2gFBATEE+DBWgqiLawxyFP1rwIY5yXip1WyB6pJsIRwlub5
IFzMXs9gl6zUnDVybgPHdef60jSmZ69biQJFhiOLk2b4+unpLLwGkIk5e2N2TRoV
0tWIYUHr932RBHNG6T+pv2Unpo+hqV0y2lqUZfx6ra/mZyxEZBFfhnFZ8iCYERx3
RtTJWGg5amFKxhegwxS8WDG+E2A8Ukvl9QGrS1sUkMqP/H7LZ+Im5/h0ix5uZC/4
ae20t9gt/9xzc+KFfl4R084lrzJdeHiyGB6SpfkQnSqWBefb5RdSn+c85klCIsYV
lQgSNObB54no4sH+BMDSuI7t3OCMDCHzHhJaB0lQcFanFqFNaT9cw8bWoxQj+aRa

`pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MKUHk394bJlctKuLEhR/4oQIbKR59xU6t+iWfrO8HOg+0bCdPnuNmg5Mcbzy+T7w
Du/XPQq6TbCQ9HINSHAJFsZ0df51cTBl+sHjr9pdTtklgdk7jTu7DV7J5DpU71PH
6VyxcfDFVApeoNBSXRq2M0yw3rgw27DlmQ6j/HMa2Ug=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13920)
+7Ayj+Lmlm8A8Hihv04Nz0fDxikk3vbSQfjTxVzjBy5+bt9m0nwpGBzHzZ2D/Ewi
7U3Pkv8huP9UaeXE+9EcG/GBDGrTravTvmvFRNGf8oXWenD3Q3/7F2q91kREHTvg
Gjjk+ekFvKnLYFePSHJrHrBxncOllVJvLkzVtTUw8dAgkJNS1BfgybyT9aFbyct6
xzm0BOPzbuXBfYza1Wn6R7jzYmSEKEVrwbe5OiOk9clrFz/CzU3N5U7PjThCxHc9
rudKhJDgZiwk/luFeKAVXdibcP2uwY8pnF1gBGqu6Bb8wtzxxVJh9g4Vf/qlDUEB
bllURCC0/cGIS/1AynThcxBpbXbrFoq0SUZouI6VY0jljagN/S0DHeAl+f7aRsFd
Pn1zjVyAJp9coqtXexhOT0b/lgT8PfMRzhaWvRn2hQ0MTEdBuieqBtdchNkC3TOo
ZxHtywvE0ONtfcvxZz4u3ehYzej+p/jrOsyOF1ws94v6ILrqfDUTVTBWmqUBNIA+
j2uoXctZKUyq4eX/FbfEHmLqsyq/6X512EH5ktAPvqHQD+JIuUGth2jY/0LuL/gV
veC6LOlBENecfSXYjePAkm5OJe7hsW+yLMbsqaRQMkItXI9+ts6UNxHoFnnSD0UB
G3LGACiCbZq9CEcXcoE12tFdZUNDDhVlwsGEmXhDoZXYskqY2/DPtk7boBOlddM0
SgYbuZlNuRY7x683y7IfCrKeE9OetTNDjRZKe+gwHfU+kWSa702clt0xFSbd5FC3
O8Qo4Uv7AygjGzwHYQqV0Nbf+KKTiq5Kf0JGTSj/cbyaNLePnJPXFDE9n2iQICaQ
1iQulOL1YzBZLitujGdh1Qryrb8b7RtkSCqKx1z4f9eQfnVeu4pm5NSnL9zwTB/B
TR0Tw/5QOQXiD0N9RYt2hUmRZ/1w9kZMid+S9tmz1LGgnbK9mgzJeNpnvdcKngVM
WcqUTn1slCylWo7VEyKXz6aYjFJKXwTewDkgCqQxnlKtTUI2VNoCANvj0xLLYvny
p6NK2pmIWQukuoAFJbGEWCezQIy0cb4QHLPaYPnLGO29SUbjZ1VnavyagMBPuH7E
UroDzN+Igz7ztzGPOOdhRfZfKxFd8fBXiDTycvSBKbOwhfvA0P9rqXUSWUsbU22V
o12CqXbaea4dOE7Va4EBkQlO5V73IIRdYITxyDyJ9EA1V9c8BMQEUdYaTw0HNz9Z
/F04TUhIMhdilsC2zYJxnmO53kpSyaATceFsW9qTpl3LjQbpzNp8W5oTxA6z0cW8
cEXA2VoA92zvp0hYFSyKhEqjvZ6ckid9QHnLHJEIhpBCFuMMmmbYm/nm0wkpxXZs
qJEqnsLfTantilE+ESZCbLcQIXEzFATZGN8womOPm9ze1tTYWaEoCLGcz05sqB62
uBPH8366uCxdQzu5HWuJFgnbTzTDAA5EyMWjaNwUmgMaL/tJkSr4ECh3vhbvVACC
hcEpmxr88N8+bs/un2pKuLxkX9LPBoGrCZEI4H8LHMRkQDREwHhPgQtfxtBreYwi
axP2T2O+ZLqAKesrbKeflv1aXdDDuCqmNhq5ltp5m4vZhUK+mbExoGnjw6Jlvpj+
s8ckZ2O8iKQaaj4aj1p4dnY3J3RUWc8/UNyYBPJtJOhfcGoIiS4LIC9ULvcs5r4E
uX2LdsmTXnOHnThgqowdbnPNi8NFeOIGJA2xrzOrTnwAY8I5mHAptoU2QlOA7xFq
K47FbqiVXH8iD0//wRILXnSOLRxRvUqluD/H8lJV1OZpnH/GUaiBd0WLqpfKClrE
RnoU3eKVQrGPtHZlo1HQJPmH/rvW3Gse+Cj7mM6DOGHphk4H6ZJ5YmfMCG26v9mn
BKHBbHg9YU8XqbhVmfT15kiIEdaBdBOT34oaadsDxorKKQxOa+lSCYNxz2cy5I0N
wcNayrF1VPwaYoQoGPNKGsK6sK8DRvHpYukHH5TA24EYXaPEjLAG92u/xg/XAa8y
wNFrcuCWRoHjooJ9h/McVrqJz+9qdnaB0vhpPVyDXfcnkN7VXeOEOILV0WCEOrE/
e8VuTkuJhIYOc/WDj4sa+Rk1rO5vRXlgEi7zYGgeNUJmVkP/wzBD9mQeXCF86x5O
S49mJ8/kREtb54Lg+ew1iSkrd13Mt7eB/3ob4ENkLhJeyNvz6ygsM26g8L0vut0z
/4Q4ecbjfxL+RO7S4kUrrwbkYB5A/2xQ6xt1sVF3z9varsgTlHLS/LwHfxaleApb
a+GhpilRZwSk4Jj9GW1tVwkbpHgwrEma2rXaE7em5MSq5Ip59mds41ALVph9VPqm
1lb5aNGS0hWd3D1Vkogy8cSWR9mFORpORprTrCgIyx2roclgNXEGKaatr2T/9BHW
+2wnAmpXHv2srmqNZKIma2uIGlfOcGaWvXm1KwK1nLqq4t4VC7sutCuT8H5utI0k
vOE9ST6tXWGBJoNuLMDX41UN39+5scjeZ6s5ldL41FwlSXbTp3bgkSelN0lFkWPL
iFa+AcL0SPyGZRMP5YjzJ3xa516BU4n+G52P3xjRMRmKCXF3/AVtBMn+6nmgDAFV
1mjJqGWPEvV2CGuQsKP/dLssdlXk4pxDou/dX+svOAF2ihxCrVe5SdULDTEUp+Wi
29nvubfQfrucAb8NnFf62SZWpO5/b9mAtKsjDdqdBt5mbq6gkOccPSSlhJC3rB07
g3fzIQyuzxIACCbFwRLRkicmqlLks2pc+IXoiYTmGCa1CDzXmlIjaHLCv4zlhQgV
zxHBmTwimLx4okiiRHpBJck0BNyIufQleXI1uVMZSJ6LqTL+H0O1yPxFzW1Px1A4
r3G03wyWQw6g5PiBt/D8+xUJJ9vEwDfciArvETwfbNOh4KdmpYnAWvenDoNGBtRJ
RdUEYpuAoQuxi17dfS+nx7f2BJcM8BG1byMeY4TWgWujYtgVOppEcKdGjNoWSipW
9UmXoFmH+7Zi58rZCSZqe/KLs0FMPO+54s4Osb769CBYL0MEUet6/GgTtdn42XGI
F7ShQQv8x0o35B+KNtn6p64pgL10pPml+O1nMs9mOk/9iBJaIsOWrt0V/0rcqOJe
SGpDnVOmdbH9ef+3+5YdCalg56mAmwrof+uCiIy/960o4Y7PcfXI3yEnqwb/OIya
kAfvxAZbt9omkdEJtGtzLh4kjY33SkOLWjvIr1kXyjdcUY/PHM2KjckkkMvJgea5
ZAiwIPEfwPoD1Y/nTcaO3CGRUnodBcv4MvLpgnouyfOLEkeP776sKS/wOj8BPj8T
B1ZG/pMNYump6silWBzSTuNCqXYcLMGvePet0iw5kkgitOBBGtkWUN2fozfwmMjz
g5Dd7K8SprpwqwTkleVPax6V6v9urVYRW9qtOKzEB1ttkx1LsulpDASLSetuTtBf
8SFdVnrGihuvCLp8vZn05mTQqOxNwHkOnau+3LgMilkIGVBUlQ1o8p5Ld9d/6nzr
UqPyEEw1p1Egfcuz29uIGlGMBM07b9fTdPMjvsFYqYIIf0vhUw7bMQyFp+wckEH1
/aZ6M7PCoYZg7nsPiTyGQzZ3RRi+ytkND/MaM77p4Z+6rFPHVXlrhTdPtfcp2I+b
BL6qLeq0KUYS7E6LR36jwm/q2I9h8WiUnq0SCFpWzFrauivGHiDqgJ3ww2k4EKTF
EoLYq3QbZtwjIW7m3EfrOCpFF/siwl1q0Ct7q7j2+aLQLDTnvfbaaKloz5oOz1UT
Fr2A3jWHZpHr2lYCf6kXxgHMA8Vdv+y3IBUZHwTy9DDsKVwHcniEDIDyyDUCaanu
KxkAN6s43OUgnEeT2pSVhFkq8xFLzG80BE9UdRdhiHx1m8ljeOrOERepCMDMrWcS
5nneoMLF/77WChRzMS3aDQCkDi0HdULKBikeRe2mkhbYr3dx57cZaMzuk/50lkXO
Nm6ewYL/B6ABI2J3fto21WdVznny4kfKvCEKxRe+GFSv6zwMxJKbKasX978wOYX8
oZ8AeuX7B13o1x8vGaOuiTzf+Dj6oRyZTpte+oDnTOMfTmAhY49B1xPRZYvIkN9v
pnKlYVPir1DatW52/FqrTu4PgD4rYOt99pSTZp7B31PZoJMdZJyvg31MiEyIA/1e
JHpchoQ5C0yFf/3ojOm4C9zX0uWuePUEY/zBRBxU0oWEuViCiiz5tBxov8sJLaXq
NFR9TWGoE3Cw1WbhiiuNk2EWilQayh2d4uSD9nGna2HdDb7jzf/R7BhO6rOJpt0f
JTXD/S6Zp7olwwdWLfrsav8rBHCQCW56LSpS3eM6Y5PMdZAfAEniizJrnlqujXHa
wrxWxazl/1bA8Wm1+fPPY4u44DQCtCHu7IYMyy42WUCvRp7lIdhaSSDhc434utET
tCCY7f7o/5WE/9GlN5VrLae0Fq3HLOEDvvrKJzKxaipC5VFhGajpI3p5rOhnuloQ
fYasb42kS3zeWO8mthxtuZAZE1BVhet/ahBWU4tsI6CewISMSoOx0sGMCrp82Mot
XhDWJE5VGvyXhA9tXelmHNN1mHM81LC2gxnk7RVj3Nw6VVBaCuzs/TJyfjxYIZE3
U24XOfhYp/f0Eav/9XQcIUrZ5ZtrIWXlsH79Ay9n/vc76wH/oF7Lae1La6jWqHu5
6TUHoun3HKF+Q4DYzVJzOsWaoctTVHUdVKZH96HE75zCThKFTAz1VNDqB5YQGDqQ
WDbEnEf1cRqm0KgEjiIJiddT6dAOKyHcS5N4YA0lU8fjxa+rrx8vYwRWVo/Ab1cK
ubljDf/lL0S+kMKzi2TPy7r1zv4+rrwEnCXPEZa4mnXe43epgpNsyEZVkPg7uMWX
Mj7kb+cXq7L29PZxQBYqwDPtNRAhL4DDIruU7/86ftYFSlD25b8sbDmKfSwaM0E2
CZHX0my2BDUhd61+su3Ilj7gAyOdL7BEdsM9mbMxJeljOOlaVKiAeR+sKMZIEQAw
D4xPZbKt8jDXt+vd1SHkksOsdlBATWaSsCoNW4NGdUHmgczbGAzbTMhCUUwcLf7D
uH/ILFbcFUdpDUXAdAVGXhbx1C1U2DmHIO7/Y6bI6/zxbpz8RkDIt58yg5NpRmty
TsF5w6y+Ge9zG5Cmy1HDo3fG5uTU7cza6ZRTw55e4CSrx7TGT0gwd4wSe5y+sW2o
gUzL4uBeqgibeabKeATVj9v+x3wj5EWkl5YPkrb8NK1ZV3WiBPiymDEWZMO4p8vs
bR13T9SJkuu6VcGiyXDLiim94WOwmTnWd7MyfaK0E1JQ/HTBm308ll34ATHoCD7T
Y/3dMChJjgtkLFSrDE+At6crqnBmF/Cf9qJrB/jQshbgEtKjhFKwI8FQ1mwTPdAE
1jTYBDWKOpPcHxk5fzPiLI6TVqXCaJaxBMF216ForLVw1S1cas8zeFrIK++S28io
vl++lT0GsLaIesT8hCpK1NlhOz7xiqRcUbH5OgnpoxP/AM+ir8guqs+F6pQubc5D
lepROZQGvw/SB15TMF6Y3gpaStBhJ9mSenw/aFEu9Rf7Lc7TkZJyynedRFhMU19V
5huZIZDZNPC38l4jn/AKa/3YttA5Y0q0Tk02VW4L7ZlStN8T6BuGgm1+fB3rkLtj
1S2wyZupDWijNOAjlKVHKlCX4ePcaTKbJE8sg66Djp9bKnAAiAQzvrQEgqXNKVT4
rgeY27lb9qfAioVVti+PKfUDsWPLAtsCNUCAux112uAjtTePMbE0JpUox623sAOy
bRIWF/pYaVtZvl+syl6mD2c4iTuw/rZuO48wn4e3+Pb/Ts3Mx9U4jjBwH0L5dAUV
qrl4filry/bT2Hq5IALOoRVM/nyDqDDtiXagl5Lx/AYZf3NZRYhem4K3iHSa6mlF
5DUhgg9DgkoLTQITgK3wDqgUgmDFUbITCPMdIA6GTe4rLZ2oaCXw4bVQX6N2zS/Y
2NV0LzdK+8hcsY/ltqY8i2DxttPrSNjP7ZK0VQ/0ULiru9Ka+aQYmIJWEE1F9dJg
FKaZHBMOsUBZy0gg0henOAKJgNM5YusUox5/M8kmmfPS34Nr7w1guqB1ulaPj4hm
PvhJ4fMxfoUpi4IomM4YssKKCvYuwBGsAASeLNAMMqlpahoEfxk2Fl6/YxSW6wkm
zbFyEjqOTUyvmvNrr1IoA69ylzqHFbBw3/EhPOfCPqdIPFs80WNd4rEbIF8stevp
f0zFjp29rIXjcOIITfXxeheDuJM93m27558j7aNegWxuQ/FbhPrWr6azd9lt4bn3
UkoUEeTqvP6DJb8BeadoQccymDSXcQAq4uYcz74mhArymb/d/gcn1QEcml+j8dEV
WoRwue6h5dEiS8l4ZdUH4XUvBVcHRWlw3xmXgK5NOvudFiA9eAnmo0wPpL8aIRXZ
IR4wqrwyuMnWd3cvMa8S/FgjPL2Q1GuNk9FmdH02OYIIOVF8qjvNSUwXNDunnYfX
/JIf1hPFJ7g4huCZmQbegYcjyxLkI6YRc2QN2Mlg6K1OOLMLg2dwWsVSpnFqYkqv
aLZ6WwpAPy3yGgPfauW/iVV12u1CV/C9ynyBJrupKxNNtCDVLP0khaR0saaK/JxG
jaDnd5W3qTAij0Jz6qn6EJtzk45RljVeY0+yDXZNgo99pn8qJxNOrWxIsYLhSDRs
+OuaaqRzR5Wqzho2EdiYbLrLU8hreBsUvTXkLm7jKiSodi2Y9S5Mv5TBLQHA5tHs
PWV6/nBDC15WCJ1ZOGAJVxmbtk6TNVEh2XFY9tzzSC03bV+KSQrDCdP60qIayDSV
8x/NTqt4qiTYDzq4tpstYeThyYL6CkSbPP4jjsffwu+t2POv5SbLxiop5nh7q8I/
AeecNzjimUz8biLVzux9IF2s2DigzcVPgbwLCMKBAoY7zeD1XbMpyNH/T9qpzfEk
aE8NZCNgL4BPNDpaAlByuR+e7edmO3KIMM9HX3uy2+Zm4cC/v/7jnlNfo5oiCxEz
LLUonRLCDQVNXhRWrOCyvrk+KN/jsoFw2c6pbr2kHyjgY7MmYTRlV9PuBg3yzYG+
yXFqyenNYxFC9ss+wjr69OmzQLbJqbZHrOk4jwQw23vdI1U54FogLm//R9QTGQxR
pUD4EfLFDA3f+xOdwrdjwC4eyh6nXMo3jTWGJRgEUpYYRkG1sa+lPVF4L9t8HgMk
YR6K9zaFQmy6q1IumZh8lbDh3LDUplnr8tRSf9IHPQqY3CBIzEzHimsCJ3Yb/mcK
EPLrOG7V0avm5Xc953PskUijiQWQh4n7xHZC4NsS4RlT6xSSlGojSm02lykNuqWZ
lpOTVJYo5zrZVpQ0lBIJ2rLNmEiIsQGxMpRij5usgN84smY55V+hl00pbXmcP4E+
vtbok+I09+7BlKOjDwH54CeW4IX8WE1LbO57HqPW+CyCOx8APA/yps/sQAVQliVN
ANLpV/P6gRxB7DKIQiCZfaPt6mAInRUCAoS9kPpI4cn8Gz/INyAzczKZCjVzTrTL
E8EIg7WxfIj7S+T1z+DIxSVH3VIZHOrpWDMYSb5STVkdq/R10meD0XMtv/NRHPKj
HvVEz4pRszBWr4yN2cJwyNMPQzvBQvBL31aMEYKPtwKsCXPibFr7NlsvTrtmVmpe
CjwAuAtfkh5lKmgLYp+nfbMmdmKJSvCRwno5hjzUDuRv37BbvpELcMIp/JbKmzvV
LQgZ4xp8E0gc9xC9ckKqo8hM0JSHg7FXE478e6NPJtXlFrWGp71woyn8MyNx7sHi
1UcjNuwWxDKV3t4T2BXRdq4o+fafoeJAMt5OC02pfyJdRIoza9G7Ix1/Zd+RvX5n
lyOHp/Lh4DaFGvF53zpUezstmjONBQnn35917HtNo+RS6QNnSzyfjz7DOCCNpTdu
GDl9/dRgubSbB8X9iHUAv9ui1NiqxFOqQvQWBnexkr591i3/pCJ9io3P3p08+xyy
usWHjoTl9HjduZsYg5LuEmdanXzQq9uBK0BTJTr/ROhvWCogfgXealE4AXBXiPLq
loXHvrBhc35yl8iXdj+y4N1Hh0ak5fOIS0RHHWDYubOk4g+cmeG6uR5IGuw3RgoY
+AbbR6TeEpyPNsCXxgywPR/gp1PVn6kbDJ8Pz1mmHm80bjT69jQlHK43gSc/dYlt
d/Og2sPvri2PD8Dc3sjy9OYc7NvqHeAEuYu2mfn8bilbm0ic80sLvdk+hFMkWCX9
7OQWCOrPknvKL9LPDhh2eCp5w8YaKNT3zc67TzrOboY9iOsXf9/TRmFpjkBMMqe8
xjLxDBsA8H6w0c0WpQA2IfF0ejb1YmiZCt0WNgwI8kQbK10sWZrE3VGJpZEYGt6x
ipAS6wlqHaj7KHoCIP1Jlw6VhEDxI/ewKGmr7Wwh5aplQ9HekMgJ9ZI5PREbQUWH
2p1uQfj/B9xGlzUfDGKMnGUvq1aFc9EoNy5TRNt7uHgsvgPjuwE/MidfGgezyKQy
RNrr+hsrragitil/B139Sua7VORlzcDYjR6EOOqbXT7ucAo8Ef9YX8TKWpbQk9J4
5QpVB57xXdK9de0qEOBDV4C1SypOSuZmSTt50o7F0gWAJDeaUv8PTIDC0L9Sontn
/tRpElzxvXA9BPSRtvvi/HrQlwAv5SaRTa43DRRXGScp/mi6JnFra86pcUaQhea8
GzLvdb5S92ep4pHtQpZhU/56R+UFzcOUg2yua2aJ+gVM1ZzwwHtf6EI8xuDOGRSq
+oh65jSSmOteHV8/EQIz22GhJdHZM8wioFDnHbDAd/8cZjCkOT2QrxGDNcDiGkDg
FgSNGtuZdGlPwm/SZEdOUDHh/bQKtPWRjI43R1vesSfAEkcvowTwoxiXjFRFmg2W
+8TMRyu6uX0ne8wkYTJbNVmH5DHgRsliGvjANI1BwUILykhJ4OKsnEcYgbA5MZvF
8WHPDuQAq4vr7nOHD/FtCb1zBkh6FYexoF91DWP+QZKAtYS5eAtYSdg9drRC+2pU
OLkGlfoCn6BXPZhfIXmYPP9/dDKbrzuK+NF5kNM6Bzftgz0kZ1cgyILFTOyVYAD7
591V2BC/ZibCAieoP3H6quGObZz+P3MSezV/yXgNVxvH9nOftiD7li+W1qbq8m2d
PS66+hhroBrIJQCjlyIoPn/EYipW9ust//YrfYvG5S7mg923o8wxiIdZzx+HNfq2
CUXZyBqq78Cq/7NCplZxCVr/vhHOdUK8stDQAPaacpiXReeTf17r0X4gUT24MQLd
w5zRRSnh2dpteP+eHtI+WCqQQ0jm1ITk3EDZ0EkoWFsJLzEQaEQUKKWwIF+SFAkh
EcCbEwQncJTdlANwo2t+mJIGevgeyRJ2sW6IV5Oco3chafN3SsllT6vcZdbHh5up
kiWFXQ5BqXYH8qN2axwC92rLUiBRD8Nk4XHRUpcbS6EODUw6HD6IYAROMeMqslTM
Sa7QCGaaH5xFxk6R4SPsM/lMcGU4g/SZVmh6goe/zU1mrJEEHHG6Fe19WKE2IX9I
veLaABL4uEiYfeCc+8+GdYuYxMEZVYBOe7GM8U0bXMBUd9MZqh4M3Lisk0kYYyPQ
w70pa9o/2+MEBFOI7a3cBIrTF0CVL4D0yEnXCTeWJKYD4VXp6fcYXGPInyXxc7L0
6FXFIm+/NtbyY/pjm1HzNx3wOTxXhTvX/EilqJKq7vBsv9dwUdvCpeYYpIIt0s++
J9VNs95iCzVgtECGW+zZr7PCdxQZIxfU0QtQ/vosNa0lXJYyJSoBKRbtE4fxv1Op
YD9i6ViaCKAbXEiknon+5wBFth2uoPKGF7LEJ2a7w/+5i3DxXRC/tmxOzwwo0mpA
eU+j0f6cN39XZ9i9CQSPQW/oK4QzCAS3Mzfm/oKNA3iWfWb4XMvVv0tMfq73uyGm
iu+iI6ydhXGcwr/uKBf3Nx9rQJJY9UuiN0pBo0NECN/vEdMCihplZ7zaYPOwWfb5
cpOIVqvt7NCXPC/aPldOvFQVD5//dvNmHmpB+ZHN7ybJtnqofLHY6tUCpB3SCzS9
4MWPJQPk6ay614gt87QqLhhZVMxpaZFhY1srCDVvMdlkOWDq5T136Xu6J8zHCg1e
2dEyQOSzm/i4k7VF4vf4iXtbP82AyzMXeLlUCQWwj3hHQZgSjjmlBo9/et94eyj/
cniFs1LoLycKJ6hvFgB3muv/gUsV9G3wzCfRm3VIlbdQXOhdwfKzbJzRA9l9xO0z
SkzTK0G4pcygaMOxXZvfrXJVOS6qfemNfZazcI7q3SbIH0OYgJqcdhQnt6ZR/ntu
ZQ185qE/EyNukP2eHs7HC+YQ6uRF5j/imLRIwVy/8THsA7k+Bq7wyvGOEmhkXHbQ
vOfpBeK+HHsldRizNyBXIeCjylkKr57QazEI09XyNn0YZ/4hOn4jNsZ9A1ixZoEy
d+99h2ProFOTbWhL5pHGtHWzteqCKPQKhLrp7T2zFSwBi6znTjKPOMTev3WOTv88
QOxIMjN7vSMJB75UulPWAUy1kqcVymOF6yVwAyIuFfKfQ6hAF5ouwcPs3ONSeEre
xZFBPlTiioHX9L6rUY/JFmFMSt/Uyn5UCUv3Eh1d3TjyGyVtFq1oQqtTy5bswdGi
CHho4hPUrUv2xPAWfZYLrcvBiCSUdyU5Eo0Vamm1UAPRnpXbw0Ieroyx0RRlXmHg
+8Wb09EB1viZnAh9l0b2OapOKUymBzzXiQrQRa9YZfxXQTQpfsKFe0upHLYtD5Z4
dXRINNubsVE3mv9WJlq+AfmNBjB94pxqXq/r+mKgleMRhc6249D9/AFgaxBWYrwP
NHfh5gn7P4QiU0OpDbXsDtHfplcByJD33Es8c/ZKnmkMZ7Qo5QpGWWMDbBSH506x
AJabMEO3B/Npf7HTYg/Ls1l/AnE7dDsu5Bpt6CNVS2H/CD61ULcW1XsCpecb/Blv
3EcSzou4Q3zwgY5GLhfLOUh1gF2EhaYUISjtk0McU9Xnia26sspHbcP0l40jNM99
4IOTYGa4whOSUnH3ZXp0VrXaNuht0cqSyhKGf9htSDpyUlcaW5EQPy/H6sUdk+Zo
Qn1VyMno1+VkJsJNW4TdxQEUoTS2dICYoW5y84ECoErAtw9Mhh0xoYWnZdOGkHzo
5RFbL+sZvmTF9zK2KEqYMZ9iVM/oFbkFKajMctX2vYOp9YaS8jM8MVn52wz6S7iz
SITd1E8gmvzdC9PCAs7l+cxOlVLgr/W1jEgQ6F4v3tYGC7N+Cf2WRT8Du37uQrm4
0zZCM02A88WPVOxhGq+q6Zxa3XZUJ5GxM/XWbRKEt/3n964sbZHADhwhyGgufNE5
j9RaKBiZki9H41MeDos0HEa0JufvCgeZFMkG6RZxXfeS1Te1zOKGtHtfIhhqyuuf
7PrmPlc+MubM8HU4N8WU+w2wcfEeHGY0NSh+aYsSicq+EA+u+LuEo4DmVP7XB0K3
GthdEmAMbqm04C/bhrEGXjRtiVSSs+hqV7X+/UCe/UfxKo94iMMai0Oqd3ox7BCs
og9/mUYe+nbTGujznWGIfFNT8XGZ7v+uRVZrzwOw+U/jCBc0LLtEjxMpAzBh6QQ1
xYKHakaGqj/JZN0S9ZLCKbD1KNM5lRCHieYsWTpr7rd/DDO2yO2Tb4+NmkAeD7hy
JmqAdIs12tUxs5bGxjdCmWqDYfoRr9nHAKygPd6WAoZ7dB4sEwKsRC37kjtxRbUk
ALwYiNaRDLiB3lMA+hCHdrc30eVZwOAM2xHnkyjL9i4G0y/PLAaAuHlYbIgFtIM/
jtRqflyg1d+8wevb+2d6D922NRLwnekJzQn8vSCmui2HjVHzWEzJIaNV8b81Okr2
mq1MnIU4iF59sa397OfUeleGfsx/IOPia/3LTkMUG5cgSUb51GFr0yX4HAh7lJZW
v5a0S1JGYI5P+uo5PI/+ozL/QFUM66PWbCS9KjCwkLmXhYXkP0UZT0/aFeRk+FYF
QNgYQhlMojsN+H+mpfpZ17M3gGfT2mAgSyJG4Isb4CH2w9CDUlFte3IUf6lDbPEw
aOvyjxgkwozibNnrQNSCJAwJU+UzHLgj+Fcxx5c1nS/4s+6zeUF+RbmFULbi0T3x
MMMk+2GZ3W7AEul/wU0O+YScNniAPp4syTisX2sePyHDq9kztpHq0Y/hIYI2FvY1
8rY4bmGaJI2wKgv408jbCm5aPCCaonhdG9LEI8GJq4zra5oXEAq4DVUdgl9hLgN0
VTMjP8Gf2jih2JPVhZz8RpFvE+QXbPOEnDVc91GYvKLSqbsYe3VQ2wL/fqMy/YSz
PC5x7sT75EUr5NEevqUwTGtVxYdOKlIrIiN4ldmllNoInzCIlXUlI6RR7kJ84J6f
lD2kavwJcPF+zeUZYTYagwclyfdSZy3+7VSUNJfe+TrQZEMRvpOuXXx5myXJZODh
Z8vdZT0Uca3RyYSiOL5BXwe+2BOm5sV0KYkNQ/NixbFF+2r7X33kJtbiuDqOFJEN
NrXOAn+GvYxWHnDiTfzKRUTxs5FHc1J9VOilXsiqWus3SFNnbQAnwVzM+PG/cNR7
ZZ9S+gjc0/q3rQ3HZN7tdHb7CN4Zb8V5cek1rJkK/9yx/54NDuh0XhJl/3hhP9XR
MNOz8bhSqzgpF42XS8cIFOAT+PNMxuIuaQlV86HJqOE8djECt3agyHR5VeT2WVQ6
aWwhovklfxa62xitJxCPe1fH2qPw8nPbNXC49rIDD9zXcKQ0TakxKW1Az4vXbrhV
KHFlHFh6lE2vVUWseU9KU0fPjGF40PvTbQdWIB8cK4wEQbiNkj6oFLTyDyKThKs0
JOh92RMkOVYed/jkqtU1GSbAMhvdBZ6CFErEhni3U7pPTfYm2vZ38DqGC7VfWZIE
q7VhcWw3KhehibXWhIILQVj+Pt5CUqkboSSkmCniN7L7O54Ccrz3spmmtQIduGk/
7/T2xY1tx5h/WkdYWhCstIgCjjxWqDZryztCKZbdcZl+f8yWc0oX3eGTnTluVf4J
VOqUUmOWO8JXGof0/Rks/ow5Shq97mz2SWnPq2SV3mSUWMhB/qIDVJVI3pdZBohE
w9XSPGxyqVhBEmMKjm6ETLrzmmPiLBS/jkPd30E0POwxMVaWik1L46whhzYe4/tM
Zqh7PSYWQP3WbDUAm+woFD2Ei1namhDgF4DeH9HrP5gxvlX5RkXqX5UzqkH0KnAF
HdwPaketHlp75oTE8nX9CIZH29IHx6KZoqtBQ5GlS0qaSVwn0msappeChlhbejHF
5K5qTM+S19WanS4Jlu2jeMj4bnJD6uGpYLBeeKCoRbPk5ib6OP/uDp7u8zYMG5iN
9CYwg7kw2jQJq3Eu3f7GOmKP+gdhoyxjxh8T2XmorgSUdYN3kEr5KH7qkl9jJ+4S
Tlu36gYcOAjFZ0HL93ba5XC4W0R1UOLFKguOp1VeYQ4Evn4AQ/dV8U2MnbQeLSsn
w9I7j2g/A05yf4UdQJTexSgynmNLx2NMSGTGMVzdz0bpU4cXLvYjI+KFUNypP7Iq
D3tEHkNuRw3QrsPIyWSCEBdrmEBN9242RepVJOdZrxVB3oVkRYwlwsTnrcHkQCYg
XpsrhCwKy6JQFAKG5saDcOGVEegl6ZX1YdsYHAyx18l13ZdQGx5acb0RuM2B3PyS
fwZMeAnUCxHkTVNTtJKd/itES+IE9xpS/oLlDNLcXXzgx+1U5QQXoNahqot3DkIt
NzIq8atqmb2epiuz3y+3l2belHNWzEQXykqM2HBfcncQG44IDlvYwlwkwMlhXLtb
klT3wZC7Oap2+8ydxXVb78a9PFNLrWQMTqSi5ReazGlqdt+Ut1rJzq+6XR7ZC2qW
SPY+mewN8ejiXbcwQxaIoekxjTVzabCbXApP58S3z1IcdK2MGCtQVC3JV6WHppkK
PkeGE3vmny200ipRArMkBCXgK07otaQ4FkPSd8kUaljrXz15IiXA6T8i/6Xc0Fvi
dq4OCAtoeInaxAs9JvfRATcif/bAU6iQ+Jl4FNMTeZd2CaJp/RyJ3EXuzFuPt0od
/W88tg4JboM0+UW2cIzmEusmMvjbhnkt+NOba3GrU05mQ3CGbF4iq6pgOLf0kS66
tzIYS+zrf7n+hRmdYPIrhL7h3fE8vnnA8Zc30F6G7BJSwAW/K65q67W0XnrFFSQv
rMFJxu5EzVx81uCehSowJXvGFNjVA796pNyZNzRjXWD3Bcstd4KjJ4QYAhZXFTGF
Xbax55QT33hmjv0oeEU5iuyRepTPKXu6rvUGjHgwsSJmdhSk3TYSfcepDldaTPdC
8mvrIO9B8+LcNLBKZSaFqAT/zuhvvOG0wo2JCamBT15fJtHn8Up0HfvTWVuu80TI
lDm4YM3zpmTx1xHH/aeg7PRIjtuJlXf5H87wCyz7uRxs6UWDiUtRlbHu1+wUjqoB
sPQORlwrRrM4MvmdftGw00mFFhEKIq5OIRxIZSpQsc3YuUCDItPNf/29S0KG0zXc
H14amGn553V+6GLs6h9Wxky5cpw2c5NlPX0HceApwAcLetIjrzeXQb+vrnKEEwAx
2oKpEOQhMBoOYHjNypaGpIedKYdlDrCF7KgB0TBa79bgP7axVtntzSJh8jz4HZ//
0w7av+Qg9mX2ManU2cx2YSPrZx9YNGebLKGlHcVovJX03Wb2EzRKAud/AI47crJZ
vkJX2mpMrSK3XbNM5OByZI0o9ggiRoqVQo206Haq3jO3Ph77s718LfjiJ3IfXg6j
1ATKhjdGug/k/N1/zlJDGtbStoYXffQOdrK6Ij1I8vtdtemFZ9a+o4NrC6fLntat
tiQ1LzJ7apuQjHNpjrbOv/XHkXYpP2bbqzux91/wkWqaXsnJIVccG3ejBj1LQk4d
J2z9fQ5pX95qfn8lEMynmDH1DB3h69r8TPxi+n6QnhFijMuczqw3MSu++XaSB5Zz
R0cfdDWl8zXreSLETXMPdtAkFaYWZRwmV0A9bngLlOY1c6y+OmVYAIqrC1CSderS
IbuRaWM1ZKpmU+hlLTDbMtHdzu/vWK2eTZW0kF9IvOvvJdX+wV968EQ744dXgnJY
ZQ03gBZfFh2DZNfxVvxrOqZjojFUhttb24KmgETtIfwggNtKm8Sx6UwlRFIdzqNC
5phlSnHTzpHz0qgrir6kh1OcTlvncTlKKid1ReNuypkP40pbfJlNkYu+JpC7PgBz
sWYAH/D0S5GIT/nTsT0f1garW29REJOOrxn0NPDdM/4+5917M+PZeWDIemU66TAH
5eNFch5rc6jdjKB4RzbxXaX1ZYynDCqfkGTLrmMuyc+3Ns7rS9uRUgpkIePOozmv
scoNGTu9x0URTeNsgz5qHHNx70CyoMkmFRYrEDUDTdksLiqKqW5alhb4fvL5R8uH
2EVbshMMw3a/a9WlSCwrjgVyrfTy4OFGiFJIc3vRLNq+uLvMDQGqUop5I7KVyP04
tnKaigapuewo9D6GNoU+v0AqOpJaXYvuZl/iwqQFwOsDHvfP9xxs2ij9oN1f9ArJ
A66sDRAUu8TO0GDh+R0DcqkkvZs28SRRkig5pvmUAZO6DFp9xAZuYKy4GHvkU1+w
C0mC8WHHkr7iN0Oqb+aTGn1wN6cBAuZNzVsTngco2ugDI66cyamu/11YD0zhp7EV
zhNa5Wlex5qascLxEW8PfQRgrLEF6fxoIv5UdLZsSxDYzYRBUnL/L4KBzopVZsqn
UvJD4XyBu50fbhUqWN9Q88I1G9YamEDJc412PkusnxWn7QfDP6MPnErnwMm8eHFE
rpRnlF9SvP4Cwr+IxqQmRdViCmk8k/Kj9EGjjYeM0w0ONFzKPBg/Q+ud1rSy8N4x
X4VT+UFxIDVokytlhBxV/UgckVgN33+ILsVnWMF4+Qy/XLw3wBpX7n3oxm1Q3nWi
ponNMavGGBlKIgSyZ6HU+dnSNY6Jy1ZzY4QPAyuzjpoCSUyMWjznQ44GrZWlmDwu
thLeYPuWj6GiQLs2CJToBphGDovs8baV26ZC0lEaaAzHYhvYd8YqPxzA2UwXhMf3
KK5+/mz2Ii5b5nSYqhvhWHVUB8x/ZbpGEWLxiBygAS9VVu1/G1J5RPJYys18+GQf
Xmm85w+OtoypvPkjdDpgRWpM9Iv6FzLlbJHierFfY6XcXQVKX9TRDkwpITWQR9zu
O/0G+mY2dliQckf749LaHVH8AR5t1AVNphj8uAtNPR0kskqN99grxko03sIHBDNq
dfjOLk0ke2b673qTuHqKH0B8vCT3iIabkYwO++PyDY+ZVN+/tayHzZd31sfwgrSP
wnU54yYj9FNYXVaoENIseyhLHwWcT+Js00BpuPmBtq3B023VoNiMqvcbUky0BuLd
9Kd4da9kG0p1dLxWmEtTWuhMM6FscCGr04A0sc7wEe0lhDhRgHsPY8egiYpzoBem
P46vv+KlWkAQIVE/V8vt3ciQIobwJvbSw3wiHQ4Ybdgig/nwdvv20u6t/6vvEPb8
rNjfDUxPmAibHaoJQZeyNrAPnIrWsCK9DcaoWf+F8y7vW328JSPN1lqSE9pco8a4
u0Cvte/oCrzCLXgj5lt1vVpysfQHjxdfvuxVxIvJkFo880kjg6+h2SFdJjHWq86O
rmAm0Bs4gUfKPuTitEO6IRWnUidF0VWKr3MtGDarTPVQq/0Jd6QqVhezstmbaoyh
wPMJuYWYa3SoAxvl2NiMiwbZ1R8qx7/3NgNQYeZ3B4E+9n116xAKhfZTI5XiCoQU
JGEBHD1+Ysi3whE3KwgAzwnYESm3ZJfqOT9LXweKmiphwJxtRPpipXBeGEK6LkVi
QIPFc04Q+CjFhbiBqBa6CLeaQa4k8pxh8JL+vH1w3bvaxeUgdBFFKTIIIu2RcSj8
zyjv+uet/yFx+X+PsUzw2iUeyU6CoTxzIQCkQqKWQytwKeE+r/R9d7IHFNogAEF6
xC1bROl8qkw3TDjOw/aVhG/EHiA9jRIq1pT6foqFpBdh5KKkXRYZ/jmFofEOc0E8
wwMKuTqI4aoUDkUUM3pPdG/HEvxnfdOQpgnfuEGNDh8kmFTmh0DXHmZWap6xoWYe
oawi3SylX3KL57zmYWOKfKogtYsEijR3yiZMu0yI/gKT5/U1PG0Qh0jGsXJKDrzs
1Q3Uww46UOANN0Et5+XoOuMO1DFqTJb3ZuBqOX1oJinWxDdNxFWWOEjjC+kuXthd
lGw9sbk+0lkHMLR5jhFKWMPmGqj+7WMNSsnwhUAzh68DLeLF/wOpDoWmQ0n1ErXg
7cH1gK5gFMMi77unrKgm+zrNcaZbao1ApuhpUCnP6HV1Jf+v8K5teWpjRzieSzIH
Q0b8gfX3gWpr+hTk/YVyDDSbnF/eQ5aFNqrRXrYXQdAO6IsCyM6TgC0+Jigv+d/a
GpsqX08p9iOBcDXUJRU9L9huuzxvHRp+YIcBAuz0A/KZmsnrQwzVRC6ZqJQbp0L0
Tib8vYbzcl4iH7ttSIvfCKv+FWoh/nld7UxSpss8YmaMEdD4o1xAsXgS9J5dIjpZ
kDTJdD536DAUxJM3vZdmEHpKzofwEGwGtY5aDoraarLBq1vJJcoiFf2QIsDaEBzW
GDbWHctY7FRBEN8/qLY+r9ib8/c+dz0Pp3cbimseT449W7L8hH/30kSpUUKyjlVO
nLTx9VcZl4sVGRDVtLg835Ak8dTEFIIihWHSIxxrWAX/juwLifhKvX6T6B2SHEY/
T3cABrnzFzUgoeVRkoUdxVNfyVKdidsF2eUFwO8Xg1RYFBYvWbDZCZZLF4X5APh6
ChIdPp4fwMlB3vC9I5qawI06rJnK3MRcRrlCpUWDHXnj17vCfYJAx/M1WJ9M+Tx8
+ir4z5qZFtGHmn1LW0W+WHNlUSooPbn0VPyzbq3auqP7fZWjnguNi+YKfcshNZUD
eX3tsM4wjf9kQhM1FqZLX4dhwPn0nVmeHpA2DlTgjUCng7hbGGnKOfzgS0oiulAm
eUmenz6pT+3qLPsFsPtaLGb7+AF5uM5KSrJM9O/RTLkYebvp/cTPbhSV2NUVDIpS
5X0iFe74KKBtDh0gH1alGlKKKpC58heEfpn6fJZ4u9SETPltEcXsFD9bsFWddtlA
WNpwjxi4V7XfAOB0TumVwbMg55vxto+WySpfM3g7uajdtugOaYx0DP/omkooAow4
daCkiUczEWaBsc0ILRzz19p9ysFINMiFR7WGkNstXo7tYndnM1KpVI/bnExIB1hk
PmxUEPF4asuj8GLA9F6OhXm9UlnqFZYNm+jnh8tEeetwMuL4q3h8Ym+ran+ekfEx
KLZHe6QtU1eZcCTj2ThSIsyLOuA+4e1R+RHYnHej5U9ttm6ZccGyhv5KGl6Hhqgc
zrcdVJBBE5q0MXUhMGE83CW2YcpUcsPkk2buTeAt3jW/4FvxeWULHMN33bSL1mwP
s5uOjE7kKORzEoO6z3AoijnWOB8t/mG/uCSewcTkrC0KPwbep3CjFrPj28arRzq1
ngVQ9Da1k5qBKdcElZOtwHOxvEy4Ko3bph93iz2Tx/QNMwGSBfOFg2phiFeZgL8X
wMWBsk34FWOHNTXq4qavOd8h2uJ57/uaux0jBZhGG1bZtYk1Zum7oY4ERye2z+4l
f2trI50+fpav5hgTb+MkJzh6ULZqMVbiNfXitERafZpb2CvyZ69+eAgBMlmtfnGS
ZAS1DJW2JhR8y9k68HqbjaX12mYVK1j+uq0j6GyGPf4Wleu3peg7xU2FpYHuyzB2
`pragma protect end_protected

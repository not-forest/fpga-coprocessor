`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GqproU1E5ZUfwFfr0cy51gCS279Z0KEeBNfJRFsDtFjgEYnTE7o1zyD5kxxIAcfv
i0+8aG0E9zsRoR/UJGzPWrt+uPeL28+MBU6csdFXq4I+OKMPLpIMyInpIdvCzRtN
a3+YV+DrWoHTI5r0g18bHdifC1Kha+fi5wOVJSjrRUo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9792)
A6MIGoRTxfY3sIZJ446fiAhO6lHfxIBomBmMWuNLn3+859vugyz9SVk2SBu+Q0SO
K8p0mQN7JxbJxKkPmqiKFiQ+tJ2UsTc1kSnljp6NRMzVrMnlzOG9VwiQ0R1coULa
H+sGvYl9vii+Ugxpv3fG0MhhyXdz8cz6cqnoxT0wdsznD06OuEkIW+93q+w6aZ3L
AXmz/6THkmtvI+MSC4iRgbOQi7SDsHJ+Upb09Bb5DOKnt0SXQkJ8KW97EtAreyWk
k/I7X0urprUEiPaRRYY2DtP4GO2TEsSeW3Ykwso+CYYHbleBDesQgSOyh6fjVx3E
TCAVcGDBN4awIvpjXN0tSwgdCjzvL4ni3k1sKs9lhBV5cbwjIJVgzA6uAI/HNY8t
9EYyMKeGXgCVWIKI0+o3T3mYyVanpKqjWR0hTTINJXqX2hVjmQAMEkaPr1qc4W+W
Z4lp97G4evSnRXTaNrnbsDFErg5rGr046yFHuTGYiAHyiInR3pu0GUGCuPUqTLzw
3sQ5PVv1QlBT3Kl/qS79f8aisthEtEm+jznlaGN5IqID0TvZP5tVjbhjrgWaE4fz
3dALvEyXUSsPhWvMrOs/ptlUORjg1HoVWKcRwVwss6obNBmstFLK7OhxPInSji0o
bbzeGSdl/tJvu/AEEhkwdSLILmzT5wiXEL4bFOxiROpGrihfVe2dJ4+CaRsrXLCx
ovBAxvFhgnAQYYQdLJkhk05a7Bt3X+ZxafLdDTAqCEM7YcZ5n8Ib152URMvwGmpF
zpqwy66qNa+lqFWiPSFf5A+Lh9NLGMPWdU9Bzqf/9IO/UD3D5HKBVDyM7Httl9KM
e6g0FvwBogfnwOqcUYiryK3tx5LdAT6erDKvL1rCnxzuFgfTrnBgvCfoU80jT5e2
Z7OxotxaKsae8kOd60lR5KnuHIg2Fp2DQ1NQfv5ItcYCLu9FSdxVsPT3l8yyqE+o
XJGeAXcageOwr9tfgiC1fNiQScU/2VGOLFPid0NdPNcORwl+GtKWMRNk1x1Kr9JB
RRjmsEB8oC7+IDZ+tOlXsEmgA2GW9NwOchM0e9cVlQVPvB1YzQRu5YeeUXUL6clv
CQevWoiBojH83cK/dcNcR39hEnPnermubxs7jfTNi4DnDgEKW7aoE8Yr4ywYtQ+w
AgWDbiALBNTcTqjQYD+2SlY0zq8ZIPsRcjPoM4cGCGbWCk7p3THLF3YhGx/QWjT9
9VevnxlCSHoHoDkXjy0sigi2bvWkDWUUx7CIw5ZZmqaIpIVqL2IxcGS5aaOKIT7d
TuaPkVVIfMOz96vTfP/WReiPLULDaIS5g3E+04kpuAkcuXS1RBn4VULfKLbQWJ2k
8LKXHzAmaEW69vDQfukbFrDS494ZhOCQF/UlTslmdBY4I++K1dvND0drl6j+Stwf
XSXZp8b9WFO4aMm8AtBaBPUGr//QavrHcFb+Zxrn1fsAo7bgwKSqOp+ah7j/U1Dz
V+jzRTEVhrUS0R397mRpBXa1BQ3icwgwdsleQYUlw220IVZVCsxU6TsNyB/D1eWH
NKJtkpB6M73aNbWKX55EC5iAhrA8C4Ldw2o6hIfHXqPUfbeJ7EDhLnW5FqMzF+PU
2RABHO0pCjjKvtSfgKvEQkGfTHKlfmPu8m9rYS/rGtgESuIGP6bhxhFytA6ow4Y/
5sx1s4FxO5fkZ1UtkXvbpHd5PdgcztTkOptUzF5AMGr1ebnDIfJvM4MEH95X+Rm8
ObSHWFJA5jMKaN2K8w84tpdZxlOs+oKpew5CitETJaFxquHW1i78iStyQkS6u/PK
FA4MkAmeAioDme5brXWNHb3j5PUnNEjZ2EKXhY62g4uMudWpYnoUIXQN+0dujE2f
8CiHBgAFqvP+w5WF6a2NXnwH+thQPyeL8mrUrQCn98d2IHxQI9vXJUQhJh90S4te
Zq3Rxb+mZ8a5Vqa8ikPpYATRv04fA4R/DIOspadxxN0Na+wXOzoJCgP/bYwRpyLp
mVbi+MNlq0DexNrB5h7/JEDJE/pTWUjI4tcrfYTfm69nhoK668NySidjc7UltEqp
CrjVnNK612SY7RMsBJNkRxsbCfs70Qu+Kfk2FInzZhCNlkZTCTMlxFU2fQQtyeFH
dIZ+uEnwuM8BslprYEzc4wNcwRoNgPgBALkf/LbYmf4t51Heb65DFmC+P31wHaRt
26t86605mE/itYeKU050at1i8f3/wkTXImIeD1NFZtnzZ+h3CGm0yV5YYrFocfed
u3PyFEaG/FuORdOC7KXP0G9vtaWdd4RgE558VdXewfz8ei7oA7R7DdnwFnHgiHLE
HKXRp3SQnvbelDXGoBDjAzO5nwlG4zdbihWO1mDL3x9qfmnzwknA+vWp2bO2AsTC
zXsFMaTaeQtvBJY13oUb4m4XRW+jRjGq0mdBhwFUGReDAW53jVm3KNxuw48A5VUf
VM3AJmQ18t38GKIfEw/XyzvQmWim2GzRgHq3bWsQEO5EQTOBRqzzOb04kBtyf26q
RwqmR8uRWY/fV0yWmfG+cWbYX4cHkT6lsik6rf+dHFDOxy4wRYI47USCNmCn6EVg
23W8Y4PKG6yJAZqd4U9e3a+YTObQwpwnu2qbvjYsQtc8s6QElBexMHxK9EvovR17
CWciYXY47+uiEQASvGqKQn0DsH0n6csBhscWqjtODldvn/5uqGXcW/HLbiWR4Ctg
NGIppUJfi3P85G8ZIKd9oqBiOEMRPLmocsoD1Y5btCGjOSjcuRSCTjI02L21I2TL
ajUks41fiyByzrzsWavqFiOHENF+q6fT5Clo1b7hCF81kT84cEzC03wgAulTzMkC
4NOa2h+OT1FNRKBliFDktm2IR7UAQaBI1n4NUBTrG44W7WX1Bs/kCJDn+5mb0IPt
MBfRDsVglSKTRepeGrC15aMJxbhvSDKU4hujqekgJ/o4iofiZTojduLKy4eEt4Yl
47dCst3u87Py10aMsxD2HgWkCl/kjdaaj2gk1jRm/TyIirvyKJldmEDXfKjVavOW
5oXkDicOGY40cK6gspTMKHYSRvYBznecZ+u/PSzTtHAonbV4ZNZD6uBGoMw/Hg73
dgn7ntilB3S1297Z4oV42IpQEiyNQmvnzhWEQnvrj6UX2VwKoJHnxlWVijgC2joJ
7EVORV/JaNeMdc6KL9R8511Z1ptGS5FscOGqq84sTaqz6/e0wsgTLnSfM+44OK5K
IFdwQwUW5vYOu+6L26aQqljJ2V2ifX/FCC0kKhVKizNt9vhiV2PO122ji48N4p78
be0jTqQw/NZulH9XL4eq0KeXNGoNV9SmFed37VI+oSFDMTDH0RmM+ge4nh6MSAWF
n6z+aQORn6kgfT5MM1COGaMcuem8e/YXIJQuGdRcxQqCIRYjHvfR4G+o60TVU0IX
Fy4d2m6HtuNl7/g0Z26fwH3veP7d4xlEwGS2HdCAKR7q/r/8O1TUgKFs/EMRnIC1
z/36u+OieFSCyQ2DstS0SxEludpV1S+T8QFjwGSSAV6jGjwT+gc94KPpX3/zXjHB
Wt98xb1G6ETG56btwzLtuF91Yo+zi2/FS0yzHeKE6R5h6ekIJMe7Unv3Sxe2JAsD
Q1hBNDrP2SucDQ8KUOeS/g/3l/EQM5Xl0kb/2JK6uJrwlESGj/7Irg2SD9Nl2fnv
1IXGe5KRHx7iVFxj+JOobImef9sQ0inUoAv0J7XgpzcXjdYsOua2TVVZLzaWSb2s
J7arOX2fak8/vbEKUkCwiMU8rTNLUHysRwaznXM4C+0mMDXPU6v1jhQkB2Mp3kpV
v9SVwdg15bQSlfPVIuDc9IB2Z5d0nGQ+Zao+y4pUTE0Y3NJmBZ/xfC+/8clCFghD
pCuWwEhCcltGh0na764SlBKnyhift+Xjl/GrL0ZHHkxRsfap9ZpZehJDXlIH9L5e
EvONmLf+iqcsaeksSnSrbFm0C3WcMDtN5ZKDB1UlNxLR+L46eQo3h0vGSpIxASdB
9MfYfGKF08axb4gRFEYXlRXIx9/8iaYLGeHQZSuGjY9EYL8xxsdGWfOZhMwxtA/F
20K8te4+9a/5NL7+my4XRGUMKfPcn4qnmeS1D6rSpZJQNx2F5Qhgw3sFmjYkumeE
CJ2qCyQPbq6YatjTWDzuwtIcbs0HOjf4L+HBm/ivvEwECuBwVPTTFqG/ON+Xam4q
qKb9L0HSwqE3aE7j62XQHguKnSKiqLhvNC24l4ARNAo2bRkp045Btf0p1lOlPm2n
fSZphB9QuR07nTOrRKxHUv/IkE5lR/Sin6Z07W2J5jYCHwzzjqZGsBR3UTCNfdSZ
mW78Z4+Jiei9wQ2gMjOTKRKLaKupYDa6dSB9mIrmU2clNdQZLszqhlqUQdsfWNqQ
fBhj+Yl+F8o34KSXjjubBJdLeiySIOpJdqI9FfH34+XLRUF8U1Cj4g9G1WeijJzV
ruMBhPBZXgnVRydccClXKk7TQ0b9M/NoQD6KRl5o6e4OeE7h5Zgt95Rw/hxxL7S2
q9amhN1wNFY0RV8Jclk4Q5yr7sFoshP5L4PAXo8r8n7SNzredZKqaK6yvYvd+d9M
bYDUXl4DY6VPMmjbs1RFL1wCPb2QjWaU/tc6ISMrb6IIlVDZ6gI+vELpqlvfXfKw
JG4CDfLql5eouOUl8vot5g37s9aRNUtJylB9r5wgSVpVsJ/uuwzsyLeQD56WXlN8
Mu+xJLPBejFXsrZOTlieEXLA3KirwGqdovYFLMeKNT8HwazILb0VlqYW1yVLbtTh
1HhS7Z6dgZj59sW1MnmyPTPRf8qgynXMUU18rk9tEQ9yCw51Hqs7Q6Ci4/Q6h/X3
jDUoowl1jcP69QtcCM7reIorYNjmHLchp1jH299T1VU3v3xZ1LnQ7267H8flkW6u
5OWS4tL1KGUoQoQP8DDY91mrrieCo7ot35hpkZktsshxzRPOsOFZJKt847X6f4Hx
0Z1qlYGsBIftzBUz4BaJpWU/6wWvuKWLnBzrHxhQt9Nv9bn9EzYo+fiEO0d7xSt0
vlIYEFgjJDssoxQGCECPiNB2sLqRulTDqICqLj8sb78MgjXAu1Rf+RFMf2205WP/
gfUqCiSYk961eLnntRs0mF94Pqe0rnZFAR0yvPgVxgpeRi1lm/rEbpDB2nmx/sx4
T89EVBtI9nfJeI3gFHKXiQQNyYNhtZuuQNYWo/f/BVc/yCxWKZyPyduDXcoGiGyP
l13GzfVljIb6MUDkfmy1pRxziwZSIXnczLzvv0c6CCDEMjKCt+mpTNR1w0YV2biY
iTvu9j/gG9BKzpjCZB2QV57Qf0WUa1tKqrphhUqBNWU4FypiXSRSAXyZACccicFt
j8XnPbJClyZUt9FJh1GK2WAxfcgiZIcYylW0xyLVl6pBTZBsWP6rOeU7GIznBaDD
vqdx/mcZs3ZXav4cq4VobUiD60QA0X/0kLh2Nf2GKPSnDJ+WMHy4Tqlua+KhELhv
sDOuChUd7Le+RqD1k8SiJD8d9EZSsjV/B0nCCQa/eil3E/bzrAXnywlVgzAO7QIB
R5nnaWG97kHqV0tYrYCMZkkSVSrfCi7z2wHr9a30xYU9/NJL6BFZhxcEF5HJvTQr
Y8sSON4GI8FfFjuGV8LhKwoPW2fv4usCLI87cwafK/67RmJwADUxBPt0OkcrEZcA
8ZJg6k5ODbYyzxc8DILJg6/s6/MoQs/+z7W/gUm3YFfjv1jZ2xceA7jP27Lm9AKq
ivEVEOSbFIURQB+8P+VkhBrU9YQ4JaI/IYmPHaZOiKee8MLuGsKrX9TBCn4gRfcN
wloWbRh90KgdR8qvhDqu+DN4iVZPDFTMT/9gnUKL5bKBtr738AUTBfUkLZpsIOA8
/Ax+z0bMARRWNm4dwFQhf6jIK3TMluTziVwBa2i2jZbDBdjwKe3xg5OT4ZiNbeXu
2Yo+JtAbfMWMtf7AOSAY3/MH7tqQS8HngQbkqCvLnmEMol73D+U+7O51TFFOQFm1
YXmXIe+TAozVa77ehAMd0VQO6bSuMWjXxnCYNY78n+7phhYaAV0MyGVfx9OyOOex
kYB1j+st578GcmxqDyB4W9qbM5O6B0j8P7RY9RpGKrRn5IOQqjNyVRmOs2slj0au
KcGgfeqyCgaSHEw+UBztapDDI7pnNENAjSOwPHKqtkuXPtPEgUJ7wd/Ue3DzTnMp
VmRl0AZH5oxh6d9arkpUzkE/TVJN6dCT33yJvndocu1MqNmHyOl+5J1Eo+wJD8vT
8QhUSxeLTY6s9rOqh2qgfH0YIkgKwYxUkY6tVjxkEPRWozPUZyCHs7Gzql7D6pBv
DBictAXCjHN4IPa6y6qfAkaVRWYg+mhUc3isP5tjzlKaAjctOD47++759RJdfCdb
+N7R/cyAxaqW3Yux0DVNz5H3oxvfAuJRAcVzy9QAlZ000mnPG3AHFRLtpPPEqGou
W/BjQ78aAccuTiudpgeLI2TLUICQWvgrqabrDu3vzbb3t+LsXYK0IHUUEG0MUl6d
/ITQt2my6i/ccFb+S4HzdYlMFQ86XR4hOvdbz30eLXSgLWISbpPEtro5i3UkFCZt
3l0cJxuQXSqCT0l3Z9+V8UV6mA3a4pfT66R/wPT1UCq4ekIGd2Oqvw/IL6OPo/iY
TLCRKIiCaKhVoLJHZlLYyvE57SuXdGL0YOFn3oNLvcxGzPMxIIV7gPqM4mguMwKl
PXo+t5k5qC/I/lNoXKxFODYt0Hsd1ZXyvM3X13cL+4dw+dbu7+e1Q091uU84yTG9
Ouk4iZdG4f3zcwfR0jQz28wvLeihyNiRfT9Wik0jhYERqYQ4Xv/OFF8JD5RbiwJf
EpoUsqMJbZDOzGUjEOwIGO+jJJqNBPWZWv7UQhZpJyfS1EEMKzNke/MmmqoCQH2g
DTv71TAXLN1NFGmdmVON4nfUgsev5nxGtdknKB/z0hb1KrrZtR0KCm6y101YNOLZ
fLhIBRaUQa5qytFqboIc++pQiMmKjztHHczw0VLSXv4oINiZAM9rdJXtHSaYaTO4
HuJkWR5J3OeFaTETgi0yAhlgfPJYAEgVnkYNnzun0O7tEWVXS8AoX+m/4SuAKc1/
iJK7CppmZZyFvyvNqmnrVweilHfUt3bQKXxbSpsK9XJaKkn/IHyFQpx31teGW7Mj
u4V70FTAnMpd8zC8huJUJMVsdxK2NybL7i5aiUMvFqrnGEbpsBBwjjRuYIVCrC2Y
oCRVcTiqluw8+ySuNC60HY92NyosQtk2C20XjZPWfZgiYM9QPHSJApsb+LqLJsVQ
zhnhw+Ue/kTZe3rX4F15gFMaog8R39BKHwZ5Jb/AiizZ9JumTrFT9d7ozkrhbZyA
YSYrY5nmEXNPMknOzXi0dHlnk+dhCRmLsxbLSLffrGhn5fwz5pXyS0lIq/vIEyD/
z2nYEx/ZxKzIg+rmGhRzWSh/GpT+pmldk0jWD1sMZXx7EKlB1YzEALBf0NjDeMID
dMoETBw/taZtlEqRNL7sCfOgF5KIEpWExueVqhtzWNxWXPbvapIHrfH/pe0HZHX7
Q40TIgxaTJWFXvDrXBZ04ElwSUuONeZrSjS/qksLz44G6dIqY++1lTvTzRLSPjbi
ctFDzbKWiQtnjCv4afOwroWy2FEre87DVXOMDvLb3ZsoKGo2nf5Obc3ztZu/dkoF
TsGrAryl+enFhc3aV73moVk3fLOIWm/BGMgxp9Vkr90TQz3e6ynguDDFHM0BuZba
BuqWGzE84vp5ZErXI76I67+f7jd6YmiJ0fyo8vgpECpeNizJHOTTS+5ki5MWxi+O
53tBkB/A86r6VD6T7MhsFQD8MpyDaKVpvs5HqftuM32QUnxKojWRvWdejBQ7LP1F
Op5R8c4MTgafZbvXdmGGcpmyVwkfN0/Mqzr/z+ObNNy6lUPZSkacdJqNffRThDEG
d0D87UuT6X7WX6V0XKAWlHMJc+D3usKHx11Q9047pkbC8FccQzbeXRSANWp9/kVf
WGQ5Jf2h7vydS+Mjqh1nkIPn6IYxIcI7Ouhu2Hh5PINR+qWM83PnqVPzHhRl4ITh
GEyKnT7Hed9ek97JNAr103ptRorqONEOINvkUnrpWVFV8jSY9d3voDbqYdyPIDH2
lVGIrRe+XFtj2PwXHcj6C1KUzRNutb0Ynnz/UJMdC+w66BuvaSrog2fx0gAm9Og+
0NRnT5G0I6veoCkH7aXm4RFPT6cC6i06dMhCzknNxF2LBU9ChTRbiH323QdvyKpz
vml6aCe+auiU+f6CbxKbqD9wQCQvUupUmQCdo1xnurgjNupvzBPMFVD8JNPgbBXb
eYNZTgzppAv2dtCOnY/6TGGjwzEV8zzoyWuymQyXrPquY0glkQFMap0womDKXqps
IHwwSXfq3PDYzUg2ssKMYWifHCBVgQKq7XgafExuV2XTUoYq8e4ZI1W0+P/G6JX+
VLAmCQTGNGE5X7u7QXy/NQ4wtCYB3QdpPY2PMiuyGEM7Qxuw/a+kJwB3lFn3V1rg
wTNcsFEGo7jKXNnLHOAlermOuvQpEUXPufVBeqfyeOtB8fg20APDJ0Vm+9Y9FNAq
SOto+A7/Ev/O07BtLLcFThwO6lodXA/LbFWLVJMhF3DY5hCIVuHxEyUrTbLoOGNC
Oea1abw7deEq8WTBVhXmPaKvQgQbNRYX4Us3Xl4QVk3EQt2l4J5RcaXs5t4at5bC
TbKcabwSUS3NsuQRu+0Z8Mtk+qcmuQCoF+yn4jnkx85441T57YfbDXE2kz/tL2G1
6k2jwOtUq4BMcXC+roSpsBkQcYlEYuJRRCgGD1bBaKZ19gr92f0+KXomV23hwTCS
sd6J7HosJCl7PTCHit8EoP0FByJyhko2VHYAgk5FghW0RIccgRDtnOojYzm6hcVj
Xj/+KoYFC7ugvEHWoDJzCwZcZxpNdSNvUA4/sWM6tYwqS0pBK7hzavCujdVlKNiv
MTQbZB1FXNdEgBCrtgF32cy3QumCLlpcCkCFtPMbxWIu7T1twjsgJ+cFZZBLh6WQ
ah0lkG6GYmhY2acgHCz8fxIxoTh/HW1tdZ3Z92fZ2y/g0RZbAhr0klRsvp80cEKg
FRXTglukM1h9ULf1nAxDpLmRwumwjPGfEJTyhn5p/Nh+oYI5pqL9EK8K+ph2FiVq
YPKRqq1ZYkc7jxzXU1hGYIQruw2w4c+GTbxp5iKwJ+zsgvfi5k7cmBi3Yhl6uFyt
X4uQTM5mTJ1O/1uaOfRpPOrhMvRurhK4ltlxY0MofFJstn17ag6tAk5y8pLsjNIU
R9HGFDSxTCuNPwOleWTKYkKgSfGOzuzaFAnoiUt+3srPmuWRz6JdPZEgZfC502P4
eyJK9WjsKf493E8aKB/Yuyr+Dou0aClT2okn1kPeimQTwWyxIcnF8k9Gu+MpQTiA
5cHuruHU7XesLAgsAHZaojpFgBOTwo1BrhvE+0yWisVAemVVoTyOBxzht3nu7mey
rHx6HZzJ+HczTUzxzCFsy/QoyHrFlggSufi7fVJjNY3pvhB52e7PiHMVZFfCml19
SWpIzSPLsLeWrZon+pY2yDMFuxxZ7anJU2qQ5N98RDOXtL/iaJ7LqY67laPXA0hO
33c83JD7DalYVGj5dmRdXPNR9cgQem2UBwoGANXfrRjLkdr8uX3Xh2w+8Segly4L
YnWI/+k0SoULYI3QRowuFR0+46Frw6+BUsELuJNd60DqruhYioPC/MvqO1RE6Z/c
3S3jf7Gat8fwGtR2vG858kYCqeBXRiI/FN0xl11XMZ/7wOT57eyrBGjGmMH1QllK
/kJ2HaRRF3O2SvyOhksl/lIgpcl6tjA5XlXV7G9dicj29p9GtzDENCoGfwwgsJI2
HdscES5tuL7VXCpu8SK1Cp0X2oYPyf3soPc8TFARbCUa2CXm5n5Glif24+dSq/cT
4TUUwB1TYMfgr2qQedgtQ2CTcKpBA11PcKdfQBWa16R85ZU5Yl1xzIvuUOwiHWvp
tScBtkyghELmCvyxn+Y9nw7K7eoMqDVi9ZXVn3xHxMr4IDJLazmzIM1h1fupjHcq
wdbe2/nfRUkCvLi3lcSJFIXrv8IZ/t6Zj7PIYEOpUk3riHIu/uQifr/FOG3tFKrz
TFIfksqaLMaCsARLxXvVqRVjUTCyCKvTR3kv2A+jFjxCiMwFT2Yl0Dwsumx3PUrG
OW3mRZzDSnk2A1eegsyEH8TEcHM50j+nHltxCRlGt5oRSU0MGKwVIT2FIYNrVFD8
1t+aU8NeoZe5SyCccmUkU9XLun254TsQjyEe+rPNAhg5ZIPXe7J836Pj1TA7zrq3
sZqRUxJswFwudYkFxHBFpU0gXWmTPuECztfkxQ2TmoQiEIIOWU7oybRLFxNhwmPB
mwIVX5mzB+JkebU142OB68mBq8I43+6JrDnBGEVgPxkTu9cUWesPvYe7yqE9yL8I
4AkkwN4EQ6wZY24kjLbY3TD57T08dbGrS00ChJUPL3Z+KUqKKF+xEYxtZ2qgTlU9
Cv6IXzzgSkdLy2eZdx1mpT0XO0MXLDvndclfjtYMuU6l6lx4aXtnI0V6L5ljd+5E
lc7qELKWlA8mcgN0b6DrzMFz+yBppevAArEUsxAaKTcjzXBewECfwa+4BCi2rWPF
fs77AZNtAqbRmGgO76ChdAbTUqAakefyUeNf1ROEXLdwsiowJ2GYFVMci1Xgm2m2
e6XqrsyhHmgoIplcrQDzi2IwRQJmexpgZ36DnFTsIRqtebzyj/ivY07sNtLFdssZ
o/9r+rFEi0GtRBT62rzm/Ee1V3nkvS13A4GgUre0TmksrQ9RY362CTYOT/jqeaXB
zkQ+KkdNGNkqrOXh+5BNoM5Q3F1XEGzJtYOPgFbLAJTavESHKM6zplWGm6tuIK2l
DRD3FCyaTCzK+aqIPs3XhEO/HG46teiGuRjkI+I/DqXUSmqm/lx6sWxdxNAOHaba
IOAQ3pgXmVv1LphppEfDHTbt9Q7ekVS1ZXQZ9nVN3MW/6fr61Pr6LJGVfOPwN2Hl
GMzzeA0Kd+y4wATLsKjWNAOWQ2pcAIVu4xJnRr2dt+PqotJAOwIAW+Q+AQssxgR8
mscnmuvLmbPV5EP72yqrFghR/UFTzvszVNelQ12G9GEKSVWnbIkvIIMhzeBMQnTx
9g3gKtGeTV4Pq8A2ItVhi0TDGgUgRCyMl1NrVHJBgK9RPjrz20mH1vaPzfZDs+yC
JVdT84a7wn2+yEL75TLc/+848MClvgAXzHxOdldXXNEHMR5KI6Fail5oGBGp/J7t
H4LxR0BV3AI8jMpzUNeieZ60LdIZvqPs9JMJw2sdeTFsSjRI/CpxdfaCqT5mfO3D
82/392ut63v7cgVHRMqM5PxKl2V0WbNqxkE4N4c6EdBRqad800gctrFhwMtczZk0
9e+0amiofVmbO5p6QtHyQFEYiz+nOKHnmNwyDSCRMT8YrtrBr1DPLiGibBT9ZqnR
kBSAwj4UGSXqdlrsHgpxEsBaz+1bScjPKaUsf7qv7y0dWICn7g/4sFk9/SoC+gVK
dFt1UcH6MuEKZrN7UxYiRR4QKb0g6eZELc8DVe27mUf2YzGNr/R76EX7Q6eZ3TNu
k6IshKjaZZbyCZOq1Rzbw70IGEaA+1S+2h4Z67uH8uM8bmbzVS50qmwlq10vLN5Y
sp8lMRewurLkwFVfIhC7PGSQl5G+8FUQdN9VM+AL6DJ4vCry0VfRiPKlBufhDSio
IIfiG4aAdL5ilVjb92Uy42fwkXmod5czfL+H1FpiixW3Oo4loBzlCJOQYZuIU9L1
mqUaT6LyHfnU00MJxPcUXmOVJtCK6aRHgiQH2d3eYyeMsh+9sx1BKfxt0AQOfLip
Ae9G1ltnUOisETizCRC4NvaK+asD/sSc+WfZvclL/qmnX9TAhvMVm2UzMJpNNsZT
sgA1sqzFvpeW59PLgDIKP2gBPzO48azQJtjwEVohHt7UQC/FYEvHpXEjUHnAtgMu
U+505Jf+wKIWGjeCUVwr+hUc6Ez5OMqg4x4vZ0grexPGG3fDMIYkCrlyAoPQ7GES
qQmijOMfaM1Bdc6Bl+cThNTGDYpJjSa0/jm3tSs4c2jaC/YHKFgFXih3SX8ndT8T
5XpTXlckbbuHur5LyM9/Sqe0kn4qxN2YG9mrxrnOoaGpfRk0rrwjlDFx3cJrf+m1
aNh3DWgptMmGRqks5OqMU0DbuPG6+7GB6BOxGQJxDoiI0JekPwlzjyqUC5nsFODC
qsFGhdnOJv95+owZk1ZDW1/cxayl0lkadOmc4IBNu3N6oebd2L6gEMxAnKEaaInx
BfhjjguZLa0DnbabHzmjlfWD+mBs1wlWNJsp+0mJxHsmfVecIYI2pqgYyiddQ3Ph
GOMJRep7k/e9hhLFOh37h5V1lvhWKJ9d6uubPVB8mAlol+t8L18gXYlzsnfpDley
0v524VS8PN53pogRaIGQct8vP2GAl+5o8P79Rwt+C5hoByvg84UkER2/wy7zcIJq
N5ozTVxIOJpY7re9vCsjBZaVzZQhRe1m1vmVwEaXBtpSNq4muBnZ5cCCKsKHdCcf
GtBX/sdDy+szNKPGuRqdlUblCA1DtcVyslJTdWgCnBUdV7i1kvIyQTkkCyoS2Wzv
mC4YXCkO8a36AWhgenjESx57GvBP/+zdxUq/z4HcwW4f/clF9G2ZCtdKN9PpznED
N5MuG4STeJJUrHN8FKJyuoP+69pYJqSOESgRPHyDALrRBt23Rx/bmDqMU8ySjZWY
a/CKENR48ROsvFO82QtRC9gkDSWwVQE5vjLI49ZnJE4rgn4NuPEbzn3fUy0vwU66
sDwXu1kgdtmYOBG//QR/BJ88H17a3KVlhStFvwxP5sbtgAfMaQnzhKOQl5i68Crn
bqGIgtoyjQEWfiv9Xpp7J+Hg+DXZaCqi3d2K/h0Hu5TkOMXU7vi82rWnKbV3F4Fz
Oh2+EVFAny/SfTW9znhy+ETqSzWE4Km+0WqdgnFWeIs+pDCPTCRLO4pD+AmUlKA+
WGRIY5m8ke/uCYpDijhIMiuwuhn9ZHSUDay6jt+ISC4qiFdegEEHfTsYt5kPJhe0
EYBMhqMSCMFTgLnEp4CcoxcoMyOvWHFYl2bxyQRuFbeb2XQI0AUd+IIxWjYDEEP9
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
JvWf6sMOJOuNLuYAHOtKQB8HVfwC84u2RIPRNg9kijVW5Kw6wsIEN/+C+wEFk+Iw
jUhW2Rx1j76hbe2i+KzXpFa+1WP5a4vnNI7m/PLquQUDyEPt7LuNb9B6QebIyzZ7
hvI0oLn5N+I5TMrJOaNFCmT13pDilrcYEaUZdAmeyr+fpIfvAWcobNCIhwJMRhgi
74+yBiNM6F51OUgT2W9aWA4pb77RPJzJkpY1qB0tZoopuTTBVuJGg6DOp7YvWC3l
Yd4T2sAilJpBv2PcIMSaUMXvUiFrumzw1wh6T2dm0O8lGAjxzYWgRzPlIGd+W36M
8AmJemn0j0hYOBI2GlkNIw==
//pragma protect end_key_block
//pragma protect digest_block
pXIrEo7Kq/P53Er6kcBbP9bqenw=
//pragma protect end_digest_block
//pragma protect data_block
qlEG8JKxiRGPthhlXYqkIB+IyXVD64Lu4BPRUHqLhAxi40PdatxtB81B8loNo/+E
jb3jaqksiHYPg+YZZjtk4NeGpmOq7+slq6MVJk34ddd52SJ7bMVDleoJcprQ26ut
CEav7nO7vk2ui2iRdX/RtyC3ItSROHnfPLve/sSMj+T3oKlgB9fcsREDHEjrw/om
N34tX2gRsx2luqG4v0WDHOrt/xSqluDNqLqo+/mUK7hNbUp+RNWx7zp09O7BkhHp
K0Ht6TWlS6J0e5IopKYKjuPjfhtGy9Dgm1+qLWw3QdisbLVghnNuUaJ2GyPjV1sG
5tGsuwuoZEdot0lruin8ZttNYsJ5CRyht728AIixTVxxDa6TQN4cR+C1aAmJAUhn
Z1cboeoNXfdwccP3Bk1ffOPy442Cj3tHJzziAlzyE9l0BAuvdCTLNvVW6AdoQItU
tNK7XG4sd+nvlAKWPkFUvr7Yn4BAUgrYbw9IdJTdSSZsdXIx/gTEGykt8kqFPFa8
4YY/EwI1vswKiCYkahhx5hiKdPGjpo+mbPRHkMOFvrOzs3yc8M/uxF2HNsgaWp3m
Mw0HLIuuH+Wh6HHdmf7ryy0GOjKXBshkLSubBMTbxES2/53GIoJNJZm8ngzj6DMC
eP2oBssW88T8+Y6rigYQtukIFtfUUEdxxKpY3z9I/wNOIG3mC+u4pQIZbSwNPpb+
xRnL61Op6lw9VVdPXawNpUyHDwrdhB0zzBpSqxUR5hgwN+YUy/8oQ+EodtpansDP
LzEB1JMWrG1eGE0348PrsVY0EiPB07eaLfClCpNovBWFI6FAooJ9PzIez3ll/9pI
/eYe46a7m6q6YXeUyYM3p0ueaFmytsMTQsSUYOoJiUIYKt8o59oglq/ZFrkbDL1v
VIxXoBCJokPTQBkFtHpjYxcIZ22++7q8QBAq0AuXULUw2AXb3uYRy2cvXwXvmAeB
uEd78cjSUwhH/Z2eltwyRIN/a/+1Hlh5JIJG7sWcYrTveDzXOvRJixOyuheoTthX
w9VCq9E6Eal0ybPbEA/1DGmrkIokrEj0DKDsXu21oaPGYOCZz++SRyj21IbGQb8l
rH37Sb8ikESWJK3agpmsGhM60sLpvYmhXUYmDe7nvSiL/AeFwRFsXQyOC9vMNqMY
uzIvNvV2zA0NyCWdSQx3KIi2SL7BwjljAAjYBH1T8vOnLxsB9N4r2soWhdvQQyzG
IDGSP8X0+t/nM+LhoQXsGgQAvciJcRYy+vkSp6yPZ1OAHtsgTRIbxa/xy/3172it
t1W74Olmqk2Vm1xrsRulynrjEmOjASTT3MomTDwoKU2t3BJ5Qv5mk0DM/IRxi3SH
dEliCUP8dRovgxlrVh+skDHCefY728oH1u9Xu1bTsHiFBvFlTSQKNaskUfAlqlx/
bNIMqKRcjyTOA4rH+/qfeCqHK0r+NmTM20ka5Ubez+hsI2KsnIpCKf/QsEKgOTgk
b9H/VSO8iJpWjrZIb9g5CaQ3fCpGjx2WXxR7MSBOd9cWWXa6vFHqi30556s6BYeF
67K+/cIPpaUPxAYbpoD2iaJknvv7du3/UMb51g3WnD29b8Ea2bWqsPVMe8IkQtgC
rtYqSYf+JSXY5CsNyZE0Co6Tdj4pSNJiYDEOV/tSr6GmlxHCNYJcsbnkxdhxNtGp
WqxfSxDM+CQ9RGOnfMWTS0bKAF6ZdQguSVZuryyy/SEI7UzCBJbK3Q6xJ1IKih9+
WfwVR5QkhDtm6ADTAbz4hAH9GdM0jA6ZW5eII8lgDGdJrNW69q3ujzCZFKJQMZGj
YTkoNUL/+nMM4/HZcETplW3n3lUAsGKGX6vNwjZdQ7i9wfnh5WQB0lD85e/HCP88
Zu2+WbJL8sTqJrgjnadhn5hG1mkd5LlNMXUsoTJ4hNjsiqc+iQ2JB2HRgctKLo+G
7MT2KoLD3pMVLWwdTFZdx31X8ADd/honPXQS5wEhEJDX1hSOgYdEIL6/19S3mN89
MTLBsPN25IILN4L3FxHmSPdd3caxscdNqqYHIERad4Sk9KFViFnOb4dgPa7bFQhW
i/fnhSyR2+nVmcWEWaxNCYINSadxSPF51FnAvSYNtyttqJrnks6o8IR3K8kPlnKo
qzZhLG7vDD3O8AwyE3EUusjN/Gf7Ka9KzMWJCxLbFux3pamkrVRw1o7wdMcCCXJE
1z6habjIcwHhhCB3WVvRXFAen0H47B+y/DCZz4N9MovTatwKgDHfnnlxqvJvYPk+
ru+VcOxAwoeDqWUNsQBd9M+QL8FIjx7xz9qrGfNQ0oPoJI1uVkTUmwE6jKdq9ayE
US71pJjb1B8tyTqDbboi4ETuIEnKKQZ7+xTsIZI2iQUuguBnG0a47XWeVWZKiDiC
7cP1zTMmLMHXJ2tgkgloo8goQVRMgA/4GGcRpSeOONHgzgP+TyJt4HIP2VoaC/Sb
2aJ7i7/ba362f3f6mbCJuOu7REo0YegIKdPMRxYcGc9U9wpnpOhLycH00eL3LmyC
2oWVeTTc9B0V0+XiV9hIy6f9BOmTUujwmzfoL+OIwoN1QpNN72F5m1I7eHX9c9WT
fg9eLJfnelCQgOGuLzDCcUQ5XJjsAcjAp52SgSkkkjJbbIbEfKRrE7KjC9z3q/DL
TXKp49uVp9sLNGRQt3jkoGEkH60MTMNSEbV1EJhPU4cawkYaQIh2jl/D/4dP8vz0
zAJQ7MNdJuiNjT2mf36lOn96k4GcQWMar3QSly9CTFZ74rXR0w3PTJGetJHY/c8W
L8vm/JdmtbdQoLN3ID/xrGYQB8U1IKufJt/1RlcfVL1OUL9nYQf2LoyI9Lqu4xJU
24tBd3We/rxkGtHsIkY3x0ipCb9SsauUWjyvRyPq6n0JglYli43QnBfx0CG3hOZ8
mXKRZkrdD1xmMrfcQ4fl0mxx2yn1ZMUyU4mPtbA+V5rNC9mwJypXaGd7jA3swXcH
Cx8lWwEk1k65PwmJNHZMRoRPqRS2YWR6EPm7Y7DKZkuYMDPmYJuJCFSNrp+C7beY
iKgJdvJwmabOuO14Xpq/VoNln5ZFYXZhPLlVE2V7HqjaWoPJ93Q9sFOJNguRXH4u
xfnNnDGgnonu5GrPZiARb1Jcp7pw8JT5P67jePMUM1hCZ9QGyYwJewxDsT2MmOXB
YeyBXYrgwdI8sle1I4HyyaanIUtPpFEwbQWZlkqy7IMzVpZGxKyT3yvP3xp5KxsN
nFyGA4J9AYzeaZ6QiK5b1vQoktpJIItRRkIz7FwtKuY1IV3tcBmZZBOI4Vj/GVYh
kGWvDWa9pyutJTqZuNC40Ded+Zhzl3uixWauu2yPIfDKOurNVPmNkSMicCjINFWP
xcTMnx+Y6GFeidi+A5BHzYSlpT2a0N3aopocOXBQFaMbVvrhagp7/SazTpNxZlTO
gv8j8LpASjCLUr24mANb2jD1vfLY5qyXcx6h/6Rue0iwd/m3rfJdIelmTYYUrS+0
YsfKH2aVJ8tiLwSpBX+89crHO0+blLrIaRfhfQEl0YNudn0E93MDc6DtiHnIYUgQ
gvwdw+3HZrVyXpG+CwuyyZ+O3mgchkwmggCXkvsDgaYuuhlRkL0ND04a6bC/d6K3
jWhFIPbe3uXM+B0ic/38qxVKaeQ4TgKTUJfIQ9M7FWWvZ8XA6Rm+uPjD9HtMAl+B
ISvXsHMpRXcP00lEpgXEPugjopDZ9X1xMG57mJELkwaNcED6jFmH5sxUiBBrKqA3
PKeRSS5011KH7TSqhaCa2W4Tl0cyjQs4yhNaGj7X43Yn7+RZ8a6diNB50FgO+Qnm
F7YpuN1lQN6Z3Y7O7PhKPaYo/u5TbDEzBXuMz6nbrPPSi5jQToBTIZNNqviarrIO
b4FncoVV84lkNNWRsqOoJj8e7ZKKS5NTdPSEN8mwmyyKWRUnia/QxS/d2oMRdSeC
xAaJu563WjM1pTTcO8WStGxqdoV2qVqzaF5IuvZcjOXyLCFrZCRiK0jLKWPv5pDW
tFU4CPi67sfykKjI1qtBnFVBAToNnjmph+FlF9plJgvcTzXixTl20+jHoqYbGcya
IxWdNSghslkhu4UENq8Rze40k/i4eQsf0k0f/Eu6k2/9TyzqlQCFhmxc8FSrpCby
f4nNa7QNPV9HJDy847aRRJE/2PYp3MgX+gLnKgZmtjgfc/icdwUjIY//4eGTgn6c
caUzMnOONgUBjJB+Jwjb7P9VpX1WLF+9LRb+e4lasn6v+Oln4xe7JGxnEpUIsOjr
CrcMgW2g0VwrVceoAJSkJajIv+KrkOk4pIHmk133+0zwXOziOkXKLOU8OoIsqZD5
ikh+6EpLVEPb4yy/Eo1X4wc9DM8kBw5lEwd4DSn0YhALKNLli29YIL02+i4OvBPw
QIzEzDavvkXwySEG7w7AEaLb8/N2rm/mqveVmuRpF/TX6rSyU8RKBPUHZurfQco/
mg8yRk5yZTIXiBAUD+v1aQ0LhNZbAoR+rcYVA2LdPGrLi19JumtTffXG5d7ckKdG
J4KQcUmPgFgaUI1PoMM+jb0dy7N96634UUTmIbeWQNRi42KdgK5FFnN+kahrMOXN
3zWBuhgnooiA52Lxg8xWiGpB9Be9tp1f0LcH8ynHjdmXdqd3uIvA1qgChhTHmuaj
pewoCr7RV2AUwD8rTToPbiCaCM+FvzkiXBsY7jvFGNuhHXreTF/q6U8kaZnKw0gP
X+1TPRj307PB3Uw10YjmiddUKqBGDFKlPANfVei73K/vj1BnKT22eTAMV80NPh8U
+GJ9+UIF1D2zWZoFMsnKvXN0aeDzIimaMyQoB2T6XC3MqUxXUB8QcrsfObryd/jt
AE4H0IFgKoz5LpfBbqZr00LEmQBFN/F8ZgOo503vp4vqwRNGCmfFDMGZRexvJtDQ
/TZav55O5mtBixfDpmYkWw18oNbhGpge2rx3SeX+PX6BMU38kUHXINMNjQZX0pAJ
LodRij19T8uKeIh0Wa7Y6k2zk2BbnppGvM0SFHBHNHE1GcoJSf4LUU9zBveh6I4E
xuOuhW+c4hdGOgmuQgJyW4kYo/j9kYlANNJ/zVxGxIKzsiYBqAzngQdbsAYYunUN
Yb9fob6pI1yjuXR2OaCaXCN3agmcK0Un0WSWsKkGgkr3ZE096O5YtVypCS12OLa1
1pBfe00LViQC9XRapS4TSe70oKX/HFYAPZr10VebtX0ghberbDl+9hja1KJpFM1z
8tmhmjmOXdAkfUO3w/gyTbDC720NmLkyoTwYnMhKPy0mldytj5ZYgI85lyUWMwMs
AjZD2+5wlOcRvY5pS+oryLuVqrAin7l15ebuuBxryddBeKiGofukJsNYmwtVxCy/
RYNisMoAPPbTawwp4Gc5ZUjNBUe/MpfKI5if1zdJjHRos9AEsra4lB8JekthX5RY
V+VQcG5kaAZp1mjWvkMDU0mlMGC5zlzR7/wEc0RZh2J1xj5YnHT/Tk9o6OW7eZir
Vq+zJYwPpSfEtVTkry3J/SfmYQAnqMrnHm+aSdhoG0Z2cqYgtnF05tr82CSoMOap
jVuM5TUrGMKvv7ZOnI3uEPqsJwAjgDzrm9hadxLnfnGKFBAB3Gn54MNfvhyvSd6K
g5zCKGL07lsLINMdUTfHecp/syYyeiLKxIkKZa5uGfKtLqWs2OV7HIC+WgGKOvee
dY1Vd2w91jH+W6sGV2ONWSewyerVoguR4XqLRoT0/sdK5a+DXewwd6t2Cu9nmSwu
DFkJJBx1j/1K2hNVMv3XgF3PGHuegXu1BjzcyYlSgwwbEr8vmDbu8vXXg5kWlKBH
WL4Keahz2Kb9Q+3zk98MYou/fiUcnjHwee4HtKKlsD4UhCyZ90Mf92l1qZ/PQanz
LnCT5ci7dcU/gUQRdt3QjA==
//pragma protect end_data_block
//pragma protect digest_block
+Kbz5Lp3idneL/Flth3+ubZz15g=
//pragma protect end_digest_block
//pragma protect end_protected

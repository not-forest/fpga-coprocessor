// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
vSQSbVP/AqzFxY+4ITbiHCZ7eItX+l1a5llKntzjh3oRkrMwZGk/lhTGruTkBZwmZF/aw5hTwpot
b/v5H1+8BsOIhsUfMhXbMjCiLaVu4kgzcwV5bzI7Wwjt+eEvYPBTzOSKjSsGIMA7yhWNOdWz4LKA
kOLVmRdkjwgvJK02Zth2unbrstQTsftlYTIOeLmuWu+ufULCmbam/u3l1F80QfKrvfGYw3d+dINn
x9Ztw4qE2EpgC97lhBTDH8FVWvqGPApvV0Ix970w+9DBQ/WWm7RgiNPrYEBBP19bqPPgpRxWafAK
QtWVh22lJseO0u4bNgWn3jVpyoh5zVZzSOmruw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 15456)
b3sF3n/9wEn0jHuDSipqOefs/8FqqIhMbJ7AAiO7IRITYzdM5CpBpjL3iX6OoGgcriLaVAOkMxV7
5L8dRI0sPCkNlwPMfbT6oq90bBcf3O6IQ9NWA45boL2DV6NXu7x0Ca5stmL/iRCy5N40PLq/8tUV
XDPrOk6iPCBec5rFpdIVKT77FBkDJWzxEuSPvTm6KVAZD6uqFvAexWYDTlnxEJ/9bGLVlVhsO3yn
KPbrTqOYrsIFQs7ld+XjkHNFvq5w3/JReUIZqXH1rUzgun+JG7tQG93HlR2KP3/C+HiRiiDFUkkK
K3N5tFucC0B0NrVSfhlkJh6zGyW9s64Lk91m/9xluWTfbSOEQI6ahYTAfquRWfYE4c4OIODK9W8P
6Xd3fzpJ/7BMRqjyuid3ApFlhExLy/1lM8fR12ZFLYLEhOlzs/+YBdAwh1O9m+x+8juXUMcuCu/5
XtDkX5z9oeC49LzIoP0HuHKAq7oM03+4cTsoi5ivzvt2xQDuVRxQQ7jpYpvYxixhaXBRhxIsYzpi
NtVimm50p9D/lR/GuFyDo2tly58Wv1lnLHza4Ctv3RNBTr9gMeHesaB21xdD3z3FIn/W6OM9/QqR
fbTOh7HGcRxYY4eBQFW2aXOST2ClQMU0Icx3R50Ps7b9iGJYoGSFO1DJ6hMql3yVnAJWD2+D2+OM
19bkJkB7++Q317xSqQ5SjGxvWlUQZ1jRfLZHljw4/f6qN6m790F4/z4wb7JbTXMm3Xxf+mclHdZB
B9SxQyUVvKdIWHyEnSETaLLY1m0ecse4vh+GlNT+9NalxQ9CJImHP5VK1ZSgnwNjaKWXJYDveHqK
z1LZd1vqHz4q5qhuammugrX5Nqk2LhfG1d2Jw7t8Ayq4wSrfsCayKAOQNbAXEiw1Lr8zKcQ1P9zL
BazW8lCmH3NyTF9gh4B0m4Fm0D3/ZA78kSAEzqQREoQuVIoja8izPA1CAuHzf8t88k3jEl6vVM/w
riae6z+XWh3snJKzmPzmLHA0jF+0i0BM7ifRFYtXseNPUFgFwN5S4OEudHGqEFWeHes7ifZtFb3q
v802mGswDga3fXKmIdH0dkvIV77ziuZTLXW5m3YmYeJ9fLfnbII/JQTTdVBHOwok8jEGtpJhjCrg
zzWHT6+8CCKlGQgI5OQXY1C3SvTd9Vh/KaBJ+vnlZzQv2QvxzVh8Z6vR1+yO7+9v7B2nOOmyHsj8
Uddaksik6HFSsp3HjC9TCsDGtyZf8g4F4I2JbGdJi325qvAhq/W8E+fcoASu0CQaDsINSR9czkAu
kFXmMmT3dvE+H0JfiFDF6dqRajgY2j3ItsU1vPCgXJyO9hYEP4aQdNSuxgoydEV7ymiTAF7mbRGz
UcG/El1ugrIa8cnPseSIjnElEFK7RG1CFycE/slu8UITS82j4e9BBlex15R5AxBNzlWJ/AEXZvHq
YNqH61ECaLnc6MLoBmAFlEve9ep6Bwc+n/GCaNc2taQByUStZPJxuU5ga+3kK1ccDFfb4p+j04hj
yPPtaCekbA/osjhdAHPh7kZHHvbVayIbglibhNvLk0sUji4fdu5CnVLPF8GxbADaeWLhEwGrPMWC
fZZvo8vBkhvqqZHMZLBkBk6WD85yDfv1wPdLwoLx4ca8XtchL3hM4MiopRcU8/a+NP31lW4L64O6
lM5vTPPEc4WUGqu8wuOh4PfFDaJtMhlYQI1B7AMrN9UWWHIL3XCwjXWlb1wn+4rAUw9XkdfVo34z
8UBOCjHQmssrdjNzJfvNxnDju3UA4aOfR2uk59udyI/3eooGVfcMgzEHE5ivq/ELockPfyJDBbYg
vuvWogUa7bY5Pf+O6/UpsZoJwagyHtAT2gnu/ah8t3DefRO4Q5yFvefj6sit9KP3xD3+dpsOVBWA
bg6EksuizKO+uhdiRxMz4aygdmdIaBKRO0ABv62XTX5R6xYdrylfKg8S5qPHPOXROlztn3Lvahzu
P0fdHatg7/PYpeW26MxKvkSmUcr1QgYhvmb6uy9J4UA4sieX8DGC6WyRffiRC5gus6MUWHxJ97+Y
C3j6LS3pyw2NDoUxRwHxkR5POPE2caFGzNg1tgRMmCPgCRNLaDuf4MwgfOrU6hoPpkV1wO5uXg2p
vTK7Bv42S1dxRx+gJpqYvouQtKio3XKup9Y0BHHMxc2ZGPmEPN7XJ2UwdYeZRFNbjB4RR8fKY8lx
7GHvcaalKBGQ8PcBq86vFgENmQCmHajykel77lQ8BsvGRFukmgejxrRaGN3NQQDjxOEh4xiPSrrh
ki7lF/dhi9DVj3uz8XY99BK0qBKPWyICP0HP1fuMbtiwBroX0PZeMGbPReYm+oCl6Of7HHi6UmeH
Ol31nk/hkQ2daZL/D96rY1jCwrIKB3LOWU4mGeOW5pvfN7XhNK6gazEJDpIbtTnxLXX6fy6+Auad
Z59Oio0MviUtIcFkYQdoXPlHeXAbAVXze+ORTB2Ae2Y4rWwPcUy5F7U4h+S/uFzBqLMI+Jl4zQ5/
ubF8opUfvQeNVjAbiq9aSY6TU0NsGBvLtjPSNkkIdBub7mc5zA8NNl4IR4emhLYME2w68YG16mlo
Vh4aXoQ1KjUS63zpUJHkHy9sULVAZkezV+e0CBTiZzVq948otZ3F+0BKvePQCTbQHbZpUVyiVT/E
Hs/vrvXMZXLXWLobRao2X6KiTw/YVSFe0mjpWVl6am6Nya9832tKy760CqeJqHUUQwmJVI/lWAwn
whMA5dKB1QlV1shlyu/ajsxdJoS3wgUAGBZxX3vteBwjSmvp8Ex3QSvQwcXrk+ETGfxeneuBNqw2
DzdIvgzNZvvWUZkK1zgKgaAZux8G8chMNjFCtkrb9TStiihery1VEvNcaYbOLLzbJR/ig7hryEUi
RwT5NzuDG6anX/+d1e/L0zicTeb0tryf/BZTXrz8gOTH+AVNrSZOn042KdO8YPuMaFSKdD98phHW
/BWiq2EIj5Nfi0f7oLvz6x6jH2wu6ie9c8au1lIgDd9qnbao4EYXD11Twg4a8ly++JnGzAqe9/1W
ugZzxQhaeONvZwz/Jyg5EGElZZKbBrQvyIlD6vhrw/F4C+q+E20UA8qfVIX+icj/Lrge7a3Hru0+
gmmHO6vs1aRcr5V7IAmmE0pP6eL16YRA/0UXwmswJ7eBvXuJY8azbilsIml4JQ11EBECtBOJnzGD
bcKk/mxV8QJUBRhNqeYhW5tYxJ7FM/n7iicRLggSjAAWGvQLXBCuDiPdeChjRnuYepBD2pMaVIxT
oywYMdUZydPvZdGhiuJccawnWmHHJD0YEZ4PDAuoUnzURXdYM1TKQXvGiXihRDtx7cwfv73stjp9
IShTbajdpKKjljvXjvASpaL95XfkUnRR8FMmUkkOJmwUQxwpaPh+lLGuJcA8NVqvIWa077TARdh7
J0LGuYdcAUBnYTBiM3iQx/O9T0qyxUfAWZ55TxpJLm47O01UoYbdvAVQ26XxAggsK+v9CaU/iyNi
sqmBFIc4o/aTt0O9C+roQIZw5Kws+2QIc99h47uja/DFIks7q2sNYH3WPM3q6WzNkcj5T5yNTcPM
S5kceEkbqiY/flto12e9n4t5kx9rO/W4rN/owaKzUWVNOD9Y7qPEIXM6r808XzAWTfUJB2+iWFtQ
RD7bXcEPGeU3UW1EWSscUXsMbXkCYY0HKf6lVKsagCLQw7nbz6OKI6E6tj4zZdOq/ymMXQbZcFvN
lK5Owi6tQmZ/rBWEvDvLDTqm4rfsyktp/73ioTQMTXCEoRs2YPFzWkNFWJyVUgtthCWmyGmpu7qe
HKDAV09zXIbIyCLQKWKQmBhlM7OoLbl7LDtXyQiyvgi9ANwS6EbKMiCwg8T2ysS1OE++2GdAweD8
oFFpz4XGTudAFbpYGfHBkIzjsXhSbmUW1v234rolMCy3ML5iV7avdNvCQQ4/Xf45XLcbNGG3vKpB
WhG6hiua0ORuFMv5BHvBSYZkF9d51S0ppq2wb2Ggb3NSIz50iV+jLJYyLP1aorrq366NniK6/ERd
uYVPdfZPsGzmJFZTktZm/aHbN7g2vMqDJ8yfS0ds/6ebi/IMUw6vlqqOlKyP4qGwtZ2JAhRqsKwt
62rBvRCdCAs72hQxj23yBA8eS9/+bX/wij9ZbNDgPL4iUg3+nVoajGmINZ1+nA1klDwlkoT0cATF
K24k9+VkxkG6AypQ3bj5CsV8AVt2fo5PNBogoFw4UrcMA2nNmelRZ39N89jMUhVUdxHHf++UXF3S
kRtO+OG151XLMQ0u8jLfdA/Q7L4zLnqoFXVC2hdhgzASPrPiFJDz4BSvgPyCwufFbrHtxKmRUis6
+TzH+MF7BGUssNn8vFtSeJA0A4oyffuPxhD0DRkgvrJA6E/RkrQdEqipdMo3RIlMbOsoabgkzG27
NgJyyeB1Q+3kgky3+gxKqC4+vV3jXWIqR5NTUM3gyaq7YUGQbRfmwLl7kKbg5cClL3sYksVh3/9J
uZnUpss38LQh5uU9kRqBqDh/44QkFrt6hmaBSZU+RNDfVK9PpULgYF+3C3z+VcTv4DKlc5Tj3PVs
uodge/8ril3BMXRzCctVjUHA+R6GrJEaKcrhWP9a0w2tQsw7oBssplICUCslcFEv4fHtuOQ1/7oR
MP+yS6rrUlMYlY9vlyuivi72VmIFU6FKNN4r3562NtkOlrUw0KmseYoDPDCALtZMcXKIvVDNKRM0
u2NP2ZnLpY4dtCY7KaRCy5wbq6So2UE5aJ+W4lyZ/jpk1BU7mokUo0q6vvYwsUsflzuOt7B0oRhC
i4KWY1uUcdqltAk7wFSwz99vpV9wafrcttZc/4cwnZpf4E/tbwixMXCWvPRiSpCQy/DDa6TWwWTw
0NeD2MYr3j2BNkpDxjnBLrz9tLkW2rVJYk00T5wk93V2r2zrR6y1DnheUBbEx+mVitZEb0sRr5zF
hqS6Cdf9eq69kiWaZsYPHLKquLpxxuc1xH4kARArESH3pEZ1XCUd6IDZOgo71yILpeoSzNT7A7se
lIrrd0FNvp5/OMWTZLoj3KVIzHvft2GpLXq9Kda8QUipf3fu0XHQ0K9uvncSIZRflFMCI0JdMT4/
vsANHNhmpbA5kOaGYyi6qCyEvCjDFOZX/PHwIh8wrxu7HtYlNU/sFOxOpRE8yfvXcEYhrj7JbdhQ
zekUjAr9TDDZqROkjgTMlEV5xVXcN8EuAubG2ie5WLeOwvUQFjo9xC9++XdRNkp13bq/J9vgM7OT
GgWz4amzNKCgaVxYRjDNtnyMFT2qkFWelYDtGqLrWCZD+WnQxPrENb+dHFgc48z823e/PCQWAvE7
+if2yNELbLSmPQ4h+MursC3udCeZzujURgd9iTBxDOHBrB6s07NGUDZDHev8eDNwsEKV4WSaZaLY
R+/VNWFfPCiMgUI947HEDtyBSh5J6OgiRTq5TKlPsNIBuB4kQfIoPi53ffmOTnHKp4zPZuliMCTH
P4AlxLemXW7vUsLH0c2s8iu1b/4ofjqpSTHfuqE79NPXBS++jJpguNpokO3QkOK9hmhV2Oc9x3v1
vsiWyOfBJ/jpB1nJCvAeLqzRw3E9ARolNCyMIVdoQCyr+ZpKTqwLM4gPM8P66gSNjRTZh/HZsSPC
Dv75Vuxq7b2+BC98xpE+BNcuQ7u0QtDmoXv0hZC72HjL+kjcDWkN1dR+HxS2C54icB+vHsH9z14n
qXeiPVgluXxjc/jc4ar03WCsyJpc69/gVmg8ci8EN9txATrGNn0P6KFkSr00j/hpONQWG+53QqpG
R2wCg/njIKDVxu+0Pg4A6/UHPNHoQdwMfcyQpckxfZr5B322/TXDshAM9h1ouETj/xDEWhmkCrnp
A7mHETTjMwM3n1TdDa4P1BlmG2zxb+CSpTb6iVV0VWSwrml+j5MvxbLA3q2XPxDMryVD1B1Bf4ZL
VoPKQb3DOlVUG8bhNBeCadYWWQpzlXxw7an0NC7FoU4HiFekFKBDkPHmZ9Pelw7CjwO8SZ92d1oO
lUuu/rYzrLngO+vVX5ozNAqcbp1loluxbfPbC+RYG2uawK2amIdaOix9b4SsRvqlVYONGwfD0TV4
p7DWFo2EkR06FEHzoduxoRSi4hQeLmIjdPxnsw1Vmo/GIbSQQ6K3wnVMgkBH7WSbHb3Pb3Fyf8Do
EHCVOi/LYgYORz7iXgLmGbYvy3IoZdw6ocVJz1CC2IyLUwFkyE//4bBy8tqEw4TjGnIDSM1/jaJr
zMSkhZAMPB/A2gOX0IB3XJCgjuaNss0UEfAyzCTD+Z6YodJK4uvQCpgT9pnDCbfw+V4F29fiDxHq
C+8C//e1ptUAQEwW7ki7nNoUruZz3jY+PyDz4O+eAOOqNUxNWMYxy9XGHIXpzHjtsov9UEUjJYPN
DBiLgbsYXiruv5LcBHewxUhNSvndVFMIvJ5uC/991+ccuMSHuON0LO9xOczXbc1G8IcLUMHACnFx
tXaAPoKdzSjDTXCVgb+NFrBsvbcN6yT1NC88Jcw/ybAgAnEyBYvWvBJtbGUodY6uFc/cRooViESZ
CuvyA9Lbb3/TIyZ0+wdB6nK7NJpy761dpu9e2y0JLtmIRrtlnkLWWV6RgAtkLU+XAFndNBvTwsnP
BwDwdWIvml8bRlNbNOFHOlXxKZAhz1571VjzBwpfpuuQFTfc8Ki5AHgv6HHfTmlOHOKVzUUT/oK1
54FdqhsFh+7zZfGQjuSNC2dIsEnauD+tjY4hut21Gt3BwINi5JyF5Ur8UFcwTBWm/4To/l0ZN3rH
FKwzTH17wWCRw47eAH63CbOfFS8/Z6MOZOw9Z0zjuf695wLjRlIdg9v5QCMM4knUJo+0TVCNDELv
U2pV7MsPvLw6Ggm8jLvOvHgnKIHgTP5+NZ6Lg6kuHjYtcqaRDsV0k7AcDD+PQRxBPxmFErgHBZSl
aE4AhiOBLlhW54+iqmTZToYP80cWSB2rDvxAdBzPpaq0xzZhmJxJcnfclaaVdJBg2IX0ZsVlQZ37
GjwUyoA2Gd6xHw4PBQZvs1bcTBB5UCGWqr2HeAc0/NNEJGvOjQweskNErYm2J2IIOLuvSFTdzfqo
5WqfOzS4Ox02tfENS0pSDqQPgaFSAbjCuZaYCDnMU+Hx5a9TZR7NJjfeJit5SpMhsrx3EzOgSrDj
lGkBTxD+K/zIryA0PtTycSUrR6PmRIau5MxOkCyCZy5dakVgmo/rPPDxuYBmYSK7pQNgfrp6DJ9O
L9rZaO8voXsh6cXUyClvpTJMG14pindDlh4Ntc0X79T72r6aL/Pf6xzRBeRpUV2UwPBllZGgrbYb
Xe1mECyoNj5XtSa8SHhMAHfZGvQYRRz11tg9uKPAeyvob+T0FJGD/AsEcGWscGO/1wimOWJdpXB5
0sirVnHjmitUCm+e5Mm77W6LI7pFsYHzkhrO/i/+L0rlzQpVwjy18bQNQZV9tUfgHlJJu5hoMg50
21vidW7HQ2u+PVsXu2HGJ9Ko9nnhREEYDmCWdaw3NdFredJcm8Cvc/uJYOt/u+3UECOq97WBZ6CK
nrBtNPhC0yqtWy13fH3Bza1PpGFWuBbTHSGJCtkc2Qv4Ly4FfF1sYCy9L1QKNiUV6OW6WEdHmQ6y
FBxl9vZwZ/5YlynSaLFtFPC+zwFNKKaAgT912Uqz3zT0dpCXpwbEYzyr4uID217eD+bhEfJgkxHO
5bsZjL7CP4bZ6du5kdlrUuRBOOrPPeFmIt/csfZuU/tYix6ECR0wvHtnBI0zOCRO166cXQdCqYnD
qSwVbcNYBIt+U62q3bcl4B/lq1boC6Lgww/ET7mZq4nhPoh3qweTRyxYcATqOsGuFZK0bKJ+fBtX
aH/1f97rahLsUs619OzkXMtlcDja6xRBCvb0Hc+OUlLbvTUzYv3crj+4lUd0vR72cDdPXSxUDsns
YND6SmKd80KAAZN/Z8Ppp3AfytLkiQ3YNrK1Hqego1rpDuF1UDjjrGgO5NKDBG+Ywubd6qdphe1K
BQptXlQyCKdZcHPMg5+6RqWAow/I+yDWETEnKODP/mNEMhXx4UaIDF12kAne5L9F8E3466hTaIAL
0QgHw73hi+4o2Z5A9xoCw9MLR2WxFQQH8Bn4R6XoBIGiu/hTMh+d+Dhe3KJDyMKdCrPgAMp9R57C
xrPlJG3igMnYhSt0eENklGQIYlkGFJbv13Qg5jKXQi9g4sD0ccs5NSHvelxdty3UA7HguIdwfcDy
cibXqv2NgXFvA5rN4f0uLGlu2uvT6ob/qoI5jaPeVbyvRh7V3H5Ga7JuEnytKdJEP7sOXx3R6anq
EtxirFepo5YeFEZiDYn/iD41aBXES2bcnpvT/2pHV1e79t6PnYPdVu6jTwru1PXYbecO767+b2xh
yMhTEoyI+Gnhl9GOEeCVzr2fWSYsaIU06Yq9jYy7XGOj0vNBCLGPYKfpVvH50th9NVG+n8uLt9Eq
SxuBxrSXahnA4XJB7BXVnXnLKcM8AXTrovrfgxFYaiMoCs6nis5GSg7Gdiuu+hzFS3fk9uLrAQpR
q5LCCv8UBEKmJ3hK/7REZ5jJ90w74bAq6J3nRLKdY5uhW2vaDDiJmjjCUHYDk/MM+RizvhgO4VNi
XI9eoQAXbQaotlFspvsEcOf0kMpl/wWJ/+HQFn5XKNSql5hxSCwsUG/uIaa75Y4nKaqZJVz5Pcjm
dN/P9gXEXs3M4MZRoN1Ht/KgOspKvzgrc7eM/JCBcw0AWBe6f9E40iSyC7RwuokX/Oi7wU5avcOh
NnMMX6PqCXHp6C9kz3/bB4qhL6fik93wDyzGoPa2wXTjd55EKFND8UDgmC+0rMy3CF3i/mzniXes
6hho/7m5ZbfANKZ2Wz4lYX0AUdO7zSpeJfbkbSIUtV4YyBoOAjQH9F/Zo1wsc8gjJWPi5SzCePqs
7Wh88xVwjLnmpjAs+LZuDmg2qxcKtlbq6gaS+j2354Ab0U5pRi+GKhfcMMn4ITz6QWRZ1hTwJR3y
8OouD8Szq/8TS657/SXEnwBOEw96Pim1zhYXqT0E6SPzzdAXDlvyiIo9rVvCd6ku5nhn/1I2nM4y
+jXSijiMO9q4x6cqfYX0nOgUFY/2tFtkmB9VBu9t7yE+jb7pQ9csAmOArtbHSQd0pZlPQ0RosbCy
NjvsGwxAZK+REfBorsxbhKQrJIbpTAyTmK9myNKQE3jD0H+MSxqj92osMjgU21qtVLrzAKAw7AZ8
v99hz7HTm1Sdr6wWvrPOzkYITeRIAciG8CYFYcE75KCSmWBo8Noij99uJIlPNo9KbO3r/xNYbrhH
kmWNIujn1eg9lb7fYcOzjDptlbusO0JlTSER3Y6+Y3I5YYZKx69KI0G2nYg5ltHqRr/jb7L3MRdh
Q9EO05DwobxxqIEZIRIMSNYA/kiwfJSF0TOUpmo5HZn6Rv9/kO6m1avU4tGpBWKxnkjzHqcdYmds
AflZwOCw9V+WblO6F+GSt1LKTOuWWTs9JfydAncYc0wrIXEBvb6mUmPz3j5fCnsks+WI5ehBU8oJ
kNlbJJuudHnoEFurBCVrMdF0sWKRAzKlaMgazEEsNOwTPUNiXGp39Qp3q/JXroNyquZiDcSE0gi0
m/xtkYpwJPqwmJE0QfklQArRKlM7Vsw35H19sJa6nD5nNjrfN519b6XbG6v8Uy1VIzGwG6VxhtA1
QhHQ6uhPtm0WVmdry8VLPuESoLTa1FDsrUr42pcitNeTnfCRx0YM9txOVabX9ztnua+u+NcJrSOo
XwzOSocc40VUzYx/zr2uCbI6o3r7FB0NRae1Ja24VZM9Msx1rGPJExXsMr+0NlKknGriBopcMOuU
3TmpA7WT3UwkBSvzq5LtsB93UtBgg22AEqNHEGY3GptEfYPHOaKgVFL0w5/JlPCmHBH2VXLGZUy3
ihg7lGGxysOSkrKtaINccaZq/Vvtq0JAc5K6WZRVpH3jIPfs8DSyDI/rW2L0XH14e/MzCgiUGh2K
Vqihm12qBcFwQDpn7Ksz8f3wiaPGXbC9cqRg+yn/GiNEUpdlFZnskOxtYpFSsWzqoiSgzUfWN3On
cj7xi1ni4DMYa+9NzgNdbjFhkPoG7ExV4l0pwXDbbBxMNcMQSt6M943vX2c40tafTrupU9WsZg1z
wifsLNhfd3PBX/0uT6Kypb6ArhbgAm7Wd2TQAo7J2QLBQc+VcnCDvbx219bk7kqdke5nNgVaUgmC
hGzq3Ek6MSGlPM5wUf5YP+7b2h+aDOOuFo6fwbzAYxpH/2sKBddpeAPbcc17GtiGZDX6JcsmOCEe
4cqY5RQYhGrJSC0wIupPUzbha67uPQDhNCwDqOHqcPe5RVH/E6QBtuT51EaCqTpmhNZrN0t+mzCh
pWnBkOKGz/bMQa1EscRUzt/AYqTGVujL51dT6sKipw3HT8GCw1r7QjpptLpDRurO+UxG9WOim+iq
hK3FC86aPpFaYYPrYvUeJT1GeBZl8fLO29gUUAB2OsWWkI6H4qG1RIeqGZiqSvR+tfelo/UlsAbT
8lXRa3UYgxKkHA5BWAu0AECoOrjv/X5ILBHaCuZZp6Tg+LOLnD4D5NaZLG+6k7KTkO48ATVVp06R
LJ7CEbuAwbjFpPaYtPJa5rK5lC6l7woXAjmdOs+alYcEW0lvcxSzVbb1G1t64kRZk9Ocfofder73
NyJS8WKo5vFCxJPgmwKGFL6HLO+kO95UHclWB8LLj2ShOejvLMYN9lLHb9QozcyjPmpLYRjdQyQH
RVJcXNoQjhVvUUmA6+iwq3nB9z27A1eDY97UHHwEeGx0R5Kt+YLNZFTQ87Cd3C8p9FFjfOnH8Zgm
4Lm6L6EbXgTDvK8JNUIqIPOuxngpKujAAtO9tCaL9/kVHMyqmQSJgFpbrXWAld+nIQgbMKHbNtrq
41Ylli76GTu+l0B5ybADmCi/cgVSdGqDs5jDqqOdwShDlz5oHhOxlHPHdwXoM27qBYFbXatg21Op
r0hFKLTWYyBGdrs5Xu8FFla18zg2iYlhDf1OoPQ6zBA/RVi2ag0CfIZ2dLWsYa8hMYBgl8wLi8I0
RmDHbIqDhCz7+YQn9yW0uQFBCLMLhsZjob9S34OXdoS1x9zYmBmfwB8+Xi0jzjuVltsxGMkudOIQ
IfnuCaMyqKC2JxisQfWjkepR5oHS4L6Vkxg6Q1NL2IsclaIoPnZhULVeVxmXG1xxF6B2x3lpi0Vk
PQLhAmWc03Q+95X7fp5bU5/O2DFl6/C2U4LtZqFLpt74UTIDCBCi9zYYnqFTUn/3R13bR987HdCp
ATODYdaz1bqc7agadKuLU4/FXG6pG/2XhFUqU5IS7OjlxMLciRsHHsJt5wRSjTcddyAVONN7hnJb
kWjxCJKAv3Wee3OtPMWnOYa+99YtvjX968jjNbJjsx23lD6a1FJoduar7FbWIrPw8fqxOnA90GDT
YEujgkBE5VddX4sBdGJKQ+qx0xyrjY/V97UgUYbc2quRkiL9qbrB5Lzl4aSPidWFsBcWxNFj+ZGQ
O6uTYq3G8Q3KrpvI+v+t7d1OpFq0jh3eOEvrT6+oKydaQEfwAhZpBoFcvxDJc7ye+2izpyeV/cLu
tdx0H/KIsCShFLcADUEZNvhTwj4h2FZQbotN/RiooyOV1SrQRylOx29jOeTV3f5xn94cCWLfKQoK
QDxRh53aKKyA2egskQRsYEuPXKEyZbzDUP/Ud3sT9HVYt1LNtbGS/hQbazWFJniT1n83k+XCtnSh
eozkUt2Ya6JIIMIJu1ZboCC6JKPPGHXVpz7o5ItFa18TVfaaIC5SMEQMlebBc63O7ZTQpf6/lOE1
OH0Bbo0eIjuV6u9sAM0Qptz12YdPsNCCxK1NpRphXWssAuUxAIlec42fkgF384tBTYyE1CEYV3vR
ot71Bv2LiJI8qHbotjH08+U+6os+renQw3t3z+uCBaJgIWsGFCYEuHPn/ri1NzXPKiilgVUwoj/a
rzGKWKRWwjncCIaHxXNldrkoxdZtKzu3ROM+ByHccwM54qmrA2vrVt1RaUkBFCPGnbRuAglESmRY
Z3KwWCOuIEELkxszYy3FQK/eKhcEBa4y5x+DY3ogkGfiqKf7RPjydHCqUtHGlpLoQznNTTlhrd5+
wDGYLTrNTvzICpHmj949C5sCav9LaXRXRG0nUg9M3w0QJtm00LjX7ekLzNtc/F2U1cnMYb6at/xa
3Q8Jk9RpANTd4bAvDa52OC6ECFBCy29XqccEsaN2F1VAOA2KRLnF8qRoL01mjfXA9je40f5NQDA7
icCmkP97ZPWaTqLO5hVG42dn9AlaxiVcbIaJrtEnDyFnHaJPkSCopdjXto8b19YHGYlZl5xOBnYD
SHwLH7aa2b967a2j4QCwRSrMDkdYTu2t7AAGSrm06jV7wSW8+3aic1lgRhBV8CfUb/4qnlkehPwp
gGl9Ts631AlnsCn9FKlQhCrDDbwooNoit9+XpU/101btiVa8b3tqm37D2ruf/NqZb4xs/riTZefg
Wvxy66SGN2dwStUJ4LELQBeJMdmJ8R2yzYPvppaZ9Kcf1GJ89n5sFVtD5ts1h+0ZEzlLHs6M3L3v
/nFopzN+yBjZwOwiYLH96JezWXBC8e6zYyFmwaAuJ6vRmfnfYf0AShobZKh+VFMBvjzbbBfJxTK8
wIIuLqNr3p1KpZ465h22znPbRhUHO2VxvvGz8j4KNTFdxX2/84qt/8x6WvPw4MJ3W0Q50hf+d9YU
AiYNQPt42Xbwspcm0W3aHhwVCXVQPcDaGmqD61RI9QjcsolsvUlhTAPdbCttdow2oVK8KqdfPJ+h
oIcMDKkg+Ch14sKmsjIGEtD+Rc8rw2Ip+yaPyxGbykGVNtTk6OJ1ujg6vsDipq0VIFtsT2Wghh/Y
AmmQZRQYKvm+izmVKBM6LWE3/xNTkBqJqF/N7wR+mM2DxRU3B/cQekiwicoHg4gVwdv9RVwt59Lm
3Aw9IL/yVtd63CY7SVb4IJywd7VNNTqtMSGfqDdla9klR48R+x1Sk6dsQdPstCa3K0ikWS649KQk
d12PHStV2j+HvWiW5HRWKLomaUUOCPQF0oSAT3xM+iwG/Yjl6MxmLrRaWl+8tSMRC31MrBakxcfs
Q27GmpsCtrxuldnuXSHrGRidPCzU+mqguS5UJpALYH0yEYhCaAIcMMG0aqHhva0HP/+OzEDpiKcL
aIRxBcxThmMPYzbkisI/wiWi9sf6WlqK+WH9AMg/pI0KcntUfoboSon/OwI3hUlZLSABWYmtWfgk
kHcE7yq4sXrq91AptUzZrx//ArZyZbCqqMccGvA3iSJjVNMlGa5NeoTAIq2a2sw+VMiMlfLyU8vC
5i4CZTVh+3HOCSsMgJJS74T3YRVgM2BtgLIfjPrE7N7PHuaNuginQkvNEyUwsThrixyZ5XnhoaMc
B8Zai7v+R5vTz603mQpKGSzguvPLomi6UKmHwccV0u81b8t42DMSPaQMeqTTCc14vEeKkQrWTwUP
Z+Jqh8ebW50i0X1ck6jEl/vjNaFYqmgVPsFrgsqQV3U94Fw/6k2FHha8+hqKF+pRrrbS4652/b6P
mKjJOsBCMVA7z6Q1i20Akdwn50z1NcHQ/9F+sOH4Cm7NDnaDPvAD7k6kZ6EY6ThpJXF6+ciJAQ1N
oARcE8n/yEYDVKjtEouhNvIf/4Atko75SKOEpgOSbgWC5fBGHRrzA2eCUE18vG0CQyP84cAbs0Mo
G3p40nRu5+DYo4SEe/TBCqO9GEsK+VuoP7mASvOmwsCwwGjycFjoroVo5kqZREg47rvc8oBQ00gb
319MKEGK7EwJPFwz5K5YWtDcAfsd3DjUyO2WBQtzICreBIKzSAdZg84YzBsLf4WaOsizUCU8CZdI
6kmPH2bCkjlRmB9CcRizGFF9VWZJSgVP943djqrDFjkmisqcuRYTJfGNFVHIx3r/KZ5MPlCzCBXK
nUaaFtTaF1cpcEQXfPUn75dm4I0Zn71Tsj3o8t9hL5mQuFlEuUV8DwcYx1iJRgnBbpEqsMO+B3qt
+ScI2BQoIutbk0osizVavyR06+NRv0AmYIUmOImZ4mS3Al2vpy8Y//3x3C6rjFaMHUlzL+CmJeGK
lWfU2enSih94kgNyj1AvxFe9PSRdp/jRpFk3r23r68CeNli3Jf95//WATerIqb5ZOPdGrt6MU6c4
A7hihHGZ1h/H7XBMBIXTbI9Hs/rGmQK1XO6efzIbkDFw12EhzWdZQ+2i+ef2o4MDAY3LwoaV5tfg
+frqLi4x31l0bhXVV32R+WosteigfWprtVrhYhcRhf3G3nrsDPpsmlpXwkJq+Tz/l/VDqKA1103q
d+FY3GuYuRdeeu9syoutjhasfZv/Mmfz/uyjEqKqqjSPUlir73ZzGZKbjxZa53L2S43oWxGnN3tm
ohnBj8sWIFTS0/mSwWFJRana5vqUIqJtMpfv2XC0jAVOaRGXbgBedvvNsMESASeTrqh9dRfgJ/Hk
oZ54kZMwJqClg8acexIC1cN2rvI7zU5xFgbUMPfuObpT46ufR08V9s8AL4b9tUfq4ZgHgYaQ2DN8
6DMvlIGCZkWfPUgO3mu+uU+s+wdqGscCO2yciZ4K8WE589zpftg9T7Lnqgp1b8pRm4gPUGEPgKSK
chTwbVWjI1JjzmxeapJ+hjOLLTnzm1tEP0WqSAnzekpZ40/Dki7TjLjHQJ26e2FPjCIFrjvsqJ/O
1pamuCV+rjkUrF5LZDbQA9MwEQ/4dL3vGl8f/f19CJMBF4gvgUyln+vML2YAJNIk1sbQRIj8dJS1
CqQ4KTR8SPnvFFb4GvJI0tSkKKDYArRfS1xTv6zHLCYgbppHO3Xgqnx1YcYAKYdEA6zzMaI5ZRGI
wjfKHZli4FE5kZC8wARbzBWw5jqxuykHJ6S+SF9XxPYzJRY1vufN1gE4mXOcOz/aTng01T+iw+9T
7nW8ftLrc4T5xCe54ObH8wXJlQ0dekpVNOBD3QYKSdBYsrFipc50NMSevQ/z870+iSmyE42tXYrQ
jWmKq5T0HFyii67wzHxazJw2hhd1tERDKncEYNW0f9u4uku5h9R0c1regAW4g97uDnToYZq61Awp
Z5pPSbxAmphKrTEGITh8K/Z0qMTobyTPwXqJXRbA+nKh7sCUVqujfeDnVWmowdCvLgmDITLua6/s
bMxoO8otffJ1ueZ/nkpaJiUcKPKglTGaoKDOhHa6XIqU8iB8nFrXyuCBRWujwcvfbBphUdEMSvgM
sxnR14B4Q6lHY9u/L+p/xz5ZjVI7x8j3exDDE1Ib5VkW1LVld3vo37ft0/l8z3SHjsFH0FdfUUkh
K9zC1iJj0aDHsbfdBGsUp3Nch4Tn04Lc9rWXB4WZjAeHsReR2ntwHDWEVqnjLh3LjsGJiBmC1jRu
urcqlkIEQ50vnYAYN5J/dB+jj8DqcoNgG4dAHJdMsDiZWhbXjXlF8HKqEFCT35HCq+UWujy9buIz
nQzLYzE2BnaEhA3vmaYcHx5KDgwWvV5hLix2vbfsf4WuGRmedakhWllQeEKPGYzEX9NSrCKC6pNl
upZUxB0EKQPNXPqTjVhe/AKN7GdyTFEQy+NxU/w7PalL3GFz7xyMHl0zjMWxEKcn4aekLN1yLU7k
TNU1tAV05sa7zjTkUCRIBcPVH/lnqw7dCObxID/NpC/5LiwlzhZ0duu8J/MD0Arz9vBqWsJXovBX
pEEEUtJhM93TOpVWTSP4Y4YXXbbJu19/coi1SnU/UwCeBXj384R8/D+XgD8pReVvbd8dv6wLxB5h
IBC8IkS3Mzp7Gmv4HCrRm0IDZrK+sxT/sCo6olJ5MU2f79miQRGtObUPnwIaZcb4xm9G5mmKZOL+
j5GAHS48oRo+F8GIj3+v9pg3P/64RDgtwrKoFeNY1D6UzOJKQd1OBifbtHVgtyGvy+O/NG67Ce4C
/Nw4pivB5RPl9Dy2JethzqPCeBKnsmw97N2V6qXnZ2eOK6nJGf1m6ZIzihfxKyYV13rIGp/boq4N
mnMBRGlvd0szksuFch5p1uZNucwSUfl8dWSme6o9EHIU37uVr15rx8guyUbWMkUStePG27o3J1Di
CIEO+FGDWFZtwcBw1fERstmsefwta+MPMkrwb0OX2i8keeRTipfcXO0WoELXKSY49RdM24R40M7I
wEhFltXVoWsrL3/0X0k+8ICvgRts/ujfezwxj55fbbMG52ynP1ek6Tx4chclNsxAwSIJmdeDoyf8
GxtXOd3eJWRyfKe6XSm+mFuxhlcjbHB+Ozb5VxA+VNB0iWlwJ3XBQlhORnnEIoG3/KaZv2REjx+s
bofNdFsMkqUnEWx+QGFlSpvNSaFEFmhmFEagpszbd1jFnlqtBDNY1S5VYItN+gD/8zDADpIleDOl
fY+64aZloe5snurGzi6K3RJb3SEIorV5eisD6cyLRsNfWkNxGkF+vDIIGvkSXqJTctyVV+rRNVrp
QaIq4lgfsDYt/kuGLPqjjzmrUp3dz1KTxuszq2mcNNnP+rB4IBW/CskXd9Tdn91lADyDJhHg9bMB
BjHQtr6zba2QoEpknyRBvXEdBOQDAbnvsaUA5vtusqHicGkhNzbj3i7EFa4peYFmvaaktmphH6V8
N3T0L6IH0bMLFVga7vGC5dAPFCc2kOpdoL0FZd+HwLcpQoI38K8GR9EfpVxXN1iEEp1tYx9eqDnj
aQBnQkGIc7gcvo0FQeNSgZs4oCK+vgt+8pzSHxohuIm55rPbxaYQgeJUfZbtKkmwT0zdsWQ3Wa/j
7n5enKu2hnykBCNyVhKUIA7nMNd550Ew/9QriVa8zxbo5VV684IwS3GEm+zhyaWyFbAYMsCEMQ9w
2/gxFaQjIDu2rFwzvX7Gw777XgiL3evAVTqF6TBfCLTrXhMsYR+HxSaN80ywTIq5x9sPDIlQocYH
jwGp39Byq0vPhxCx423tH3nfOnb4d6L0NYRYoJ7e2feI34wWJIj30P1T5Ae1I7VrT54lxAtQH7kq
O60q348ZxRbB32N0R2V2trluuRqK/UgSbechynJXQBi07EyMQRs+d4Rh0TLB7GcB0PbrY38jfkJw
VOfXhVlZgpTwdF0soKK0ngd5UXwDmrLhxhuXIqQgGScirCHpbhbZMvqouY/XbB2TnGXG1CpuaYeh
v7u7pgg45SDBOgWtiU9j4Q8gyNYjI7LdyUrKkhAOhlv5wKDzSEQZXyJkraGq1b+2UmMjaOWtPwAX
Spy5pDQXDPlfrpYTY+cop4iA4XkWowe7WS56OqJjSwgdxa8Nv6YMRozLuytewCx3HmwFHF33hPCY
+VTs2uameFRzD10C6B25x/ZH5+4VBMJG3/FTMyCyijsWTnLLTSDadysc0Mj1Mn3lrbW/bRBz+qlJ
KwWX/WbbrNqiwe/MXRf2NkWnkkXNZXuGouuZYk3fw27zF9vqsMmKF0Lx9R9uaner2n67JyQa7bLH
yZvANNkY5s1VQxk6TJWT5rVnZdOQnvbt2CkyrwyreTYtqSN0YcUHa/WtpqJ9IIEOscqiqtIIWolz
kAW2l8G5H90C6bLLO2GwVXpGhx2kl/vJrHSMixRMxO7JKIfTqAG8eVe7heO50nepztm8m0PANbJU
YXhAk6D7o7opx67ioDU4K8eSURvt7d/E2/pdEMjq4gtfSe01ejfePD0moLCoRlKJRckl0YMy1X2Y
5nXzRkaed1+ZH0y6Out377eXp/xD22pOi6Ja0egwuSm7pWBeas1lhxHZAqjPMg34aSN+mH5NfTv6
4ch/6DOsUhOzHKXuvUT5QzeJj3fc804+kmQ2npBsomJ0XOmG5qYHJIC64Flrp2vsqwwM/wWRhvv4
BMD6d1RMdCk2OPlfHPmM6MUU3YAKDliCQAlD6geUGAWZjlMjGaAdxxo1fSDWiJSOcfjdY3r+8zj0
c5mG/MGstmYXRDGpKjXVSBPWC/y1HcBBmNTBip6VO1aPlAOUWARHIocxAErOGrfd2ODPulnEQEWd
HLzKSZISmGDkV3jTMVF+SlreiCAVDOnQNhhdwF2AxoXVOZxGKLY4xYTRXQdpzv4y7UDxuvbU9K+O
XDp61hcCe1a8O/jQI81/E3zEpdVmUmg2SW8cepCi/CoSRHO+ZJNAWJ81mv55StORudPeeP3frIJO
RgujxCmegmqxASnth/1cg+ZXO9ftaCSepcCvfw/7/dihoQ27zaM6TYlYTTVIFF8I3k1vCrGFBGdG
36OnX26bSOVMtNvHx9DInj3g+TRd26R6wsji3AF+dl44/k0I8ouuI33myZRdAaUb76okzWDfIJTH
LuG9l74jZnI98PTGWVEPYUUXjfSHACcVQjrVFAWVV+hEAA5R+shau6uDAYxVez/QH81yL2kydPty
pd9X/2DSBoCzDyIAS1Z9sbPziZy3wzySUba3QW7+eEQeHX8AuhhkJNv1CEhM73lRijHPplCxg0ng
SZpggC2XLu/ThKhH1SpZmen8pOnx4swwnbsCo7KPXUSD3s/q/e2L2/HQrayWxOU0tFxFajYs2REp
Ov78ei8J2xLXhkOOGVWzFYFzVGIAvjlbnZjiolwzFXTsGDuwxnkQuaUyHq2dkmKbYRQUStqL2XTQ
UIF1MnHBp/u2JcXCQe1xEa4smCNpCxNgudSNooor1ktRV5u2C6+W2MnrXWQMVQqmKBgVC/byfAJE
zOAb7VxUNQGSvZOGdvX26JHbqIPF72aC2/cPSqGHCdBpkVV0o3uHdyhJwaE4z+MGfPKZh8AyynPG
Q+G24vU+3qEfnL9ul2tu8k1J5J/cs2cwjK7JMoLQHeEpqn/LqGbxSkL8Uu07gdAxZJCIlcKm0zRw
hoC5fxL4aI0mgo8dOVxr6m7mzT5QbdRVCkp2V/F8ILVccKbnq+qg0ug7+XBkIzDcTAHsYnX8w/Ai
YOqNXdTirAHc8gCcsjBeXOBdWLlYhQuLPWe4JAafGJk1tdaBD1Z8z3AqlLX6vdmPNlygM7OEifku
YzWQbLTMtr96PCwRUNtXbCc9BYsRswn/tbbz7kyU68pv5HhoKTYOkUDlOqq7l0r9HcG8dPkpx4sj
Lo8QfrNtaSntmtOprI6PVQHy7DpyK7/AWa/4IjB1LgDM0P0HGrfn/yxyW3t98Ww1D7OaFbP9DA0u
TLB9EhH1PnbS1I8WE9fKz5FrJVdy42ZuK72cfXiMUyinrFrthEo5Vz07XxhZ8VXKIEfkTnViXV1F
YO5fSsf4/dgZ7xAOWZjX/+btDRHIvNhtdALXHrDLnOXoeIk7ZEgzbxQELotSdqFBFhhaDv0LvLb2
3mPrnDB9xeoR9vueY6FM/KnhqqCwdn71E34Uuw/W2bEQi2D0GohTdXod0qJmKpwUEMK6DkyP9+sV
jXiX/6vztdjxbEjd1dNgGV9hhA8BL1vZVlxtP+iPUqWlBojpc5Jrycw8zRSWNImveduGE3aSc1B/
MazfLu/6jFCzTlI80b/pLbc/8JOUbWe26gfM8nxSMCa0Ybdp7DOeGBmoTfLnqkCIW1xtmVsei7A+
ANldwpotUruEsVKh7qX5A3yUEUpnNZeiUDyplW6oHIdi6+Vu6KfeqlfLMxOpr6cILLZyxGvM9Z0T
gKKO7mJ9ZRKiK/njhIFGSU/aWv8hPOjml2EY7osZZaTtiC5pbCKUy3eb+sC9raTL+/6I6rL9gxgy
ubRR+GaG+fkBqmGXcwVIhfdpzRyKcsd8EPZbnoMJdaHabV1dRImDNCruaMJKQaBY/097Ky4M5Bpz
ghZbBTI+EgKcayb5hnpkJndinMkfNcRIJPrjT/8+9dB/ISsnubXRtsN0gocyGhXjzqxRTtCVChPo
DHnoo11X2YelHWMw3sDcnmRRLVLL2C0HQZdWES3rdA4HZqXFQO+DulvR0u3WBN+yclmKiAta7NHD
Ps5CzNC1RklaRkO/xFiY4suwPm8/wm7IxkiJ1nwdjq0C83+Cmw361uLTRWR7N6IFRsNmG5QeXqgR
5qZGgFkdafax+W9dlkVqNqi1OL3PDMtn7zn2z4hhSfetGRej63eSbxrJSc1M5gcV1E4Htu8JLOzK
xUu5Vu/RvOBo9zuhr6+l/dYgxSAv5gwOpiNm9gwlvWhau6mmgo7fURqP6kci1zSixDbPJNK5CnK2
jXmeIhRnyi0GzRUndxWoE8pLfVCq3ryhsyLLolhw8z7KNgk9sUmvB27nwF5RQCQ8T3zcTVdrjeZr
0lpKTYLtSohHf5BSYzjszwiOgUGbTX4I6DS3x24nKNs+A3dkvTkaPfAUirBvGHjglpobHT5cOJDd
VvPK3uf4d2vTi8RXFgIRwzk9o4k3nThZmZnFGQlHc163l9mWNLjTbN/2RJMXWtdHSqcv+NVB2l5a
RTxLSUfj5p7nQ+S10b1rebEZUi2168fW6eog6FNp1QXQMxK9VfoPqlGm2E0p4edlBuSE7Kt9kkUa
Y0RNrQ03xM6DAKpIe1w43F56WMjAMSh8/cNaeyPXeAUL9CD2DYKBH85CGcuIC8r8+mSqNRquevXL
YnPIPQbxQtsfTZ64+3/k1JQWgqQO53/WPijaEWNmY742KUmpBUVwCXQjzK/m+s7zDGfWVy6K41kx
E6SaZd+fpioew9+PmNMJ9EltI0Kiuf9RlOi/ypnCBhXp5IfAX8nOHgHWlCLBq6wlUXsNZ4vuoiBn
f4oO/TfjbWwv
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
1EWL3ypEWepxMikvQjh6Ia3l0atyduuWJNnFu/LsX5omaQpBl+hmDCxCjJZZ9kw/
sexUAFT6ZajGeZIZ5+OL4CmCphnyfRwqZEzxFqyeiTN8+kxBtMajwe7bhikzVIe3
31UnsV80HXNRAFYKHrYjN/soY3/uePpaxd+l8qY4cIo=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 10784 )
`pragma protect data_block
JnG7BNc6A1b931nbCoXmmD4f17A0g13EMR2rFcc/iQxe84XITu2fRN8g6XDzAsja
Q6J4DAo9MAW7WAZ13xYPSdNL/XMRFvckKzwMvcW7Wyc0IuvcSCgCTzEFBWO+W4D5
yl41/ftWHb3TssL1fK5TcgwqNYppGep6FfzNAF5vTJSpn+CtUvetwn9y5+JwVGbK
UAvOYkejKi41Nf076nIF+fv90Tn0NtPfQMaEY7VFAbmUYalMDue8aL4pkk79Uwme
viWMtx0y7uDja8vaUNUWk1IqOBs4zMvUEQE6RbuaWy9syBme1xMv52pyRDOjERPT
R4y+5NlZYVQugPz5aj1sS96V/7zq3OYHssb6FxNhPVRC2oeW7YVcynl5l4PNtkqX
/s1xC81yiYtd6l8V/oD5wMVdKwv7a41q0xeJ0FvfZ18KEIHo8BHYhSTQbKvRphOr
WiWy9D3Z/wWTYYyhJrax5Pehpm1IPQ3d3x7Al+IGH9qLgRmNU6L6MTVetVF6gx+0
twJ3hCBAnB5SL10cEPot/1Ya84NFwM3ib+DU2+5L3aQR8efo0yX7vaEHKv8YZ2z7
3dwWYd08XEcLNERMiySfsrXnlLUofkfPRCaXaPBSZ/X0dCLw4pSgSOh2BktWJpBb
7bniYY1OFKZ531LX90DNS0By6SOtLGFKYi/sfleByMsyjQNWzmStVt4EQSzt9dzG
0GQLa7Cp4BhUfYHx/YyQiY90AxzQ+RnVX92NEWq9iMYcnDXSdhTls1N7KLGz2b9j
quW+emh+w5z8nELe18aqMIogRsOhPZKprr7ss/LJKFE7DW+1S4cK5p2/bW9CnblD
lC7m0wPG3nFg1NCg+pk7c8icMQPOyMrrq8b/pnPckw7cLAnwNXYmxq9KMNObX1RA
tthiDp8tgi8bNfFx4OrW6p32PJPtDq4JJGhbmEWJyopM9V1mxa9WhgmhIcGc/h7u
B+lZd+FegsFPJeWQ1CtWnU26szZVwYXTHs4CG3mvFZzvjrGark8SB9Db1MogSYoL
S6DSDfxqqh6aJMNR4aGoun0Ssm57027DFBtZs0/h+kwX7xxdNbV+1DpbYKEs3Oi+
mVEj+YknVX6k5bU4QZC2Eg0F0WWkrnIXdvlPAHdULn1Nij/XX2OkMmJEQHwfK182
ZE5iK6amBqWuxUdwho6emCIvp5UOQ4Gv5V6UqU92BOaRrmTRT6j1jjAE+H5LXNHc
88kbQn78J2qb74vwZjtZfTyMzDhgs6DQeEzUACrKHtrbt3/9W+oS3ClR9Avp5DFv
oH/Za4zZ2sPiDDi35lV3O814iYT8APwuvjUPbBDvryXofd6sphGdjIVHUBPr8t7h
EgCUB1RGfQGr4r9qde9UlUFtaZiEVfDQtTl+EIIWlts1ZiJMAgxtKvJk1sclcau0
riibo/bCLlsnm8mFtQCJk17x6jPzhLDZawRGyxTHKtcqjGSRk2c0pwTzNyMjatw5
Y9VPZagtloeggK1p6hsYhH8RNv0iyoZnKvI29NOa0JxECShp3+2zGLDSYQr5AXCx
uL7vBdtHdaDY3vVdqryXUw8r8tMpFKYFaeVa/w6CQGqg3F67i03131cy+CWzG2hA
LSP+QQoFOnQ/5kKw6GjjRUyQ2a6b2hJD5Zb41nvrZ+R70jWW2or+tfR5rL3sqk67
Jgm/H8mm01gNp4c5DvEw62QW1NZHZZWkgD6pSrhqbRuTLDuwMx+Sydbfa2ko49s4
01M+SGF9iLkCtB6xd9agHmVVOnhTp9c1gymwXYVZ/7N2Mnn4gVKKSLpILlm+Wvgq
MYYAy2qHTS15KRMiOD94od2URBqZW3Jg7lnw6B/g9ReiAmM2HuFOBJSJq8/Lbf15
dbgxs0K+7TRyky3jwjDprZBl2NhIHno1oY1lwBxVOd2nr14/oQ7unjHvNu4LSR4R
TLhNiObgTkubqydKo6NTaJrx1Mp9coL+JEkO3O8t/z4UZQGLlgQTkhFWyKotgsDM
j2CDG7dGzPoMjB6YLRx+/gwJn0REVEuzIgPO25m9BGPbUpGfZ4iQSKHyTJgy9U7U
ots3u+vrI1E0IZtWgBsw4GvCHnQefxzpGyVGNwf64doY/ISU3f6F0oW0mecpUfvl
8o73rS98zsslCEavVRjKU+8oiU3b13uRMe2AYBXyCiUUCWplI635w1mrePTuKQ41
03WG9oEstavkMjv0xOeva1Y8CYYD2LpOPr3Z0xXsvFDL4XEl+sB/S9MONXqa3KoM
EXvnUM5AlgpbqnVh23jmTw0q9CyeSmBKN8rMbnu1YEhU099E0u1xZ4yk0JhuWpVt
du74VTJll3uFCamiVT0Z+xjrF2OZhnlTD8/TPS8tZVdSy0yozLyxeYYua9GJrk9R
+jhFXUIQF9mlsHiFtJuTAibUBrdrLwfazphli8Fs+fqu4UWVuIOeG5NlRLmfreBY
kLbBt5w74GvuBVEiWmgOleijJpyM2ooy2lprCBQ7Fq7BpFVvt6jg6W5+KLWW29Bb
Jya/4H/r2rRgg7u79jQsmx3XfU5Z/Bz7HV5rQI2it0g6NCEX+UuTZw51+KZNTLBB
Yl0nudsLtyxR83PUMSqIRZpkY6ouAjBU2HFkZH5DwUTjbqlD5+p6Orhdim8UMHdb
Kpm3uHXEayvCQnamb4jRG/RfYbK//6FmJESQgM7RDMonDWTrt4s+aTUVgdDzZwUW
cHz6SOgZWTxuPuc7oQCujyLyf4OLjgFr7KrBswtrzlLwWPSzBc6JfBzBLv8ySqO+
V2a8FpUXljBZI1raihkoWfGZaKnl0McRxvz9zElVQW/uUz1+FWP/Io1blHtsGN75
0MFhFUdq4KcLlN9yltJJKjVmWO2+yKss10i1frCEdCnjsya+gYEG80n3Ca/WnIII
yx4oiLYvGB8SEHCR+7BuoDjXbQeREYhy5LzI7OqzqtwY8J6AmVSelIxRaPXN+ca1
zqiuig28vObWkY47ecHk+Y+RHXhSu9GCYvDznXY2Y41a+KhYntVXX49wNH7+Ptxo
7WqwVI7tVE5EEF0N05dacKLL05j44OQXkrG65CVeMdjrw/FHvzUDxsUiCV8whD1g
aqbftBScfxvJqa+V8UXAKGhrf7XXLWE8mQvQotN4YWiUvPps+RUtxet4BTUM0rdr
zaYY7wLtqYGsc+Zhzlzydx9+mAWy1w5zUhenz46zbd4uOZz4tjggavbQPTVDdtkL
UqkhJztuFgulHrRTPJ+TBYf5H8feGGYiwbcHgBsXXhPFZJvvaaiFf4KjRLkOmFiN
YTN/jSU8lxkRXIgt+hhEXjG5vERej0uEuWv9VzJvxa349SrjwuxPNRBjz9tjpWEQ
o/uUXkhs3KvOAq2tJB70OIKmQDbR1/MOsun9BkaZqmt87JzATdzy7nBIGmEIkjpo
IdHLis93ogXu5comjqPyT/QMxxW/W6slKGcnC/8tIT7DNGEi31DCw0mQE7svtyQA
5gxJrBzo5e5NXEqD1panMdIUnoqZvh4dBvG0OQMFOFWQkr25ejhulKbAF3nWxB7i
xNX0bfxYsQXr1q4LUjAo6zR7cpa/JxgMQkT9G5M1FinqmM9SQtELVtDfrw+XYMgx
5v0n/3Nw6dr0xMjr5TPw2FmjZTaP5EQ5NGdMgsKwy3GdHKVFlBGPYhKi/AuuZ0bb
USujp07A37bkGQbMzsd8zHgq7d2IivAXxryIczNca6YO/9RYi8kq7dlmEs5K13T0
QAQ3Jada1iNCC/RcJJIUiTMuPrqHeSuONsTKdnP8A3HMdumZuGYWRQjyUkefuYgg
FNHlgpl+CrbJeRyGYWk37hDVG+yu/njN8sxPsX8YGvKtP2noMdzndJhB+8Ty9V7F
wdC9ZFJ7+xuEx38hH7rXUvfKDEHRXlYTIno1Xa07JrWtxQCN8PUgcFcCXAP0VHvy
DLRaGk1XRcVR2TIedoqwdL51wROaEKH0xwvLdZ6cehjZsd4/FpNJzb7tIer7UQuu
UMhHTTLWYMoNU4FKBJ9lrf0xYZHIxLWCM0LTXYx+RRpYFJpRY49kUcvgwDAOfdob
Y2GSgA9/9rJs0MVOcuRkQPlSuLjI2Ix9yjSv7kCAXmXc+S/F8qQ1HN/SssDrlsDv
HmgyQa7vAYy8lZ0VQEZz1KyUOPg/cQvjQaZPqc8tkHutAif0jS+6qGctxXpfhmja
8ejzdV1rF/b5yKQ50TatkuvRiVhkFeUtciuRMU3uS7w37lolpLs+ZsNAiftuxino
PBO1G2X8JG1iQulGH3iHoswfb9yD+9igAk+6NdpFDddLbL6aKgo4mES2YEOIr+ih
3Ej4jTy5iyTmYOx3fM1vEZOLCR9ECq6gND6FYZeMkzksfF2ZOc0WJKmQ7JbCOVVN
C8Q3cWN1Yr7qY3L3mqNlTbsva+3IGNUkrBlZJW7gD0wrpJo3AIUS9GDtcCzgjK9O
vzZxreI7MvATRkDfSSG9Zt5PnyNkW5HZcr+ZgxH2uX5PO7TWhM7o4BZUv7CTm7ep
l45EN+nXN2hw3EmjminDm8aScXxVmxVfPnr6bHntRYHpzjDyHfa8I7zXaCRHR/9H
aDR2e9D0G8I+fZfBw4Y0xPUIQaLKfdT8kaI2Vh7f/2BSNoN+DzK8GKFQdZUCPfMw
jKb8UvSJkVjIBuCuZp5pAcY0joJt6Io46Xf6MdIc0SKC8VCWHlCeWJwlmOekLkcr
OVIXFrFdKM3qkmynxF7/1jebirpRBPqq+Y5S5vaDZ1AcWScdNgxplr7gWVvRtTRU
H0PZ+N6RE5ur1QqOCAQbeGD2idF4B5GMrlCbP6wgi4a2PBDqXGVWLg3HdtARqxuJ
E2zmR/vRvGnAe8RjjlKRM30rbYma7NndlI6oqid+pF0O745n/t2gEgD/rrPFvddu
wJLemmZLGQz2DgTd1RYN/6dUyj8o0BG6D6n2mP8adakr1JBx8yJvDr7BPoeoBik9
giYkLjn7Rt2fjkg+07uE96KnNIr104J+TeTh8nwGeICtA634g2PvU8kKpnptOTC7
IVryUNurDsw7T5Zs5sjdqH/WeHAMRFfaurpNqsQj+WUmYw21izsgiN1absy9BkWV
BJRNpAJp5MlB7yAxOO9eiTNRVjWtLH9GgalT1/7xp2F9Yc5H3LtTNiy2H3IFV0LO
eHVT6sRM/un1e28gSoqTzsy3IgZDQwVVCUqfVoBxc0PPv7/pb2c7bPjvDnJ/HAeN
s0HX7mAOmnDN/dcFpeDHihGyAqFvfwOYyjauMXkOtKIXRZkpn17nQmkn3xz9Q4fz
rJ8wzUqnDfglqivsAHZqvnsGBqLx4Ewg093PUq/ZWGGeJtFH/gGGwJIunCrYTdV+
3pRtcvNGpvnNxMYGJ+/AHBScCvOMCFrC1892WuhkHnuVY4uXuBrHw41eC4iR++YM
E1A/XF4rxVbrf1/3nNZGZ7Zz7mf8n12Xi1Hp5pbhVhRTRa8dgGXY31uvDcxcdadi
5VJ9LKxn3NwOe7szgGm7qxbYkY/qhU4V7QLWj9JXYXriDmoknA1HS7EmBfxaQI0d
MRZF80IUMURaT5DjvzyQx4aI9jOoHbeEa/qoUfgUZCik4Vst79iIx7IQQXjE/Wbi
9TClhFqT2fU4fN7DyRgvq8Njs7/gb5NEpGY4p/0FGoetUbQIWzEqfftPZempnxC4
xPLtLpJHlm7McjB3Nl7yMl3eTPVNINHqxrnc0Sw1/U+yTB9M/u3I0iJ8rk69eYMw
nFGjVYaZho/rpgJKtGUAUgkn7JW6sA6fLXoXW0QIEvJDtOd2fFXfDyzKT6xVEa1k
LUiwMl+GP2x40Wl8nVzn2HlUve7HaIl2fwt44nl/23G6PUBIEI8yqAKtH/Mb/2Gs
W4w/21SYa/ct4YpMLzpn6il2LM8s8h6bgt1PJlgB82ahxgL71/5W1N+Tj/1yCu07
Y8oMjlLH7yOod9Z54AmK29jgBk3EF6sV6bTM8b8VZ52FPX6Ma2tqqrzg32GTdqtA
1kvx5D0uziuWhS0By+CDkjdSeFJUiGJTtlquuMBA3mPA8cBiA9Agw+ifTudd+sUr
gQhVb4tR5qIOpVATR0oP1kLuW99tgyEnrOpR833NUz3DEhQYTLHcX6mSBg7TnuOn
cbzqwJsf85O2844EzOmbVVEB4ihdurjuRKMZsD0qP3MVjg4WPdZgnn4i0yqCL4N5
WuUF9L2Q7yDUPrmk74nJSvD5JIGwEVwSVHgRD0Z8PkEzbF+JGzdmpE+JB+NWsY7F
A/2vNYND+2BPGmGBH1/+b7mjiMOznSSZyM+41EIvxkGEpY2ofaJ4A5rMAjJC/vE5
e72ygD/6a60u8KFTNZRuMKIihinjZAJ8Eao9jBtWwa+f/w2Xng2+ZO1Z0MO7u54o
LmsddkYpdBErc/Lt1TiB8BM3+jB7G9oppu+zsaNbWufJV2U/RN3y+e9067S19drE
Cq89zftwH8JKc9nHa8zzgEq7w4A5hwRYdBtEC8IMpVDIG05wdl3CNFU448bSyARO
FEPne1ExgVXK/zIrNVrhN0CIyZiF3zCk/8bBSA77fBCp5gx5ScXiXKHvz8xddu+v
dMc6r4PvI7uZLaHVzMyrI1mMR7NIq9STpaZw9VAGoJ7i1aG5eecS6rV148HbWKBA
EwwMGYLHEgEyyca51fi8FT5PUTwjgbLRuRgC43HfPkKy/abYxMyQ5aCUS22GVb46
3IAfPdZaGGdSjBe3zE7du0IGwxCd1p9HXlxQo3MNm3GxXuHe89UKzWjnRex1OTc7
dQO5MMcOjNuYx1Zw6cWD7vGW+9sgYIMEqoxa3MYFHR71kq/YhsT8xGzP5GT/n/tM
FJPX1fTIAuPLybsjIM8c3WHM0pf4MjIWuE6zxPZLfGMSaYG59/yhXocHYBvZ9+6W
Ef0UM2KfEUsMlav9COSUC5+tTzsOUXo5UgNnhckYEqhZWZn95p3DgOxNlrGyyGVP
ZU0RhpRsytLewUONBtXoRDCJlyUeughqhcBX2zjz4zLj1M02PHwePdRop+2iBxbH
WgD55zt5ZQWuGABQEYVjM3gDuC+YU9b3ckC5B1yFM04s9EfrSWAW6KKDq0fnE8JP
MP1iyzKi95i/Hj8A0DL7U6cQyAC2WcLtSDajirgz9cbMLp/AFr5ySHPZK8ggsKD7
6K38hwjAv7yRZrSjSrQFwS2d+Xp56jVm+xtv4Tv/lcJ/qVnQiYIPDnQZhRV57z19
mSLPOZiN9VHd/0AVdl+stBrPJCASOLai0Q8U+dbbFV1llcVN8hKYfsqdW/YmnZzX
kcWNaZmBJpES5bHPW4TtZKcGlqPevun4ls4LZF0Sk/cfLxmRAv0VVnHDNSGst/yw
0FhGi8WQ9go5K5VgeEQLwtq1See5fiO6oMTB0Tk8pPFJvmcKZairIim2b54ejnFo
wsEXR8Yu7lHkrjZCb0b3K5eYU5crYnL+Kl0p72BYfNXvTseqeOLTW1Fb9IEuMqjE
tTDFhQ0O8bI26imB4thm4qUVDvQg3Ye/PO4hspjVP9E8rP6VzGOvu8OOIxkbwgAV
sj9q3rOU285rIlgZd8F16ICLMNvpBnKw6ahDwJJLtGR0HEvgpDmt39S10NacQ8J7
Vac8TqwT7aAH3/yLkXhpsruotP09kTYf0/rvztsQDzIARBkqn9Llt7I2o0HW+TpF
GlRnrYF6KnmrJVUlL0fpQ+iWEkgyFH3/Imb/gD34ue06sNQdhDJ6D4/F40VugIpN
FO5SqfBml/svNHztbkOqJRPMHJhjasCD7ZWVfMTkp4az+MBTxcYJ1q3dmatjyTkB
+ZlWDqtu/oxAgYkmTDGIsVX/pOW/PHrYbDacDUuym396fCLp+vcCKgGDqsGEgPLJ
twAblyP7bi5JNHm2gQwIfMO28/t47Q8MZxQ5MlQJRm1aTw9Qy3UeWKKssaIrI8wu
8XX3+OYpFj+F+SYx34vQtiMJhFBXX/zwLNn0NSfuc3WDRjB/uPabFnl/OMKpDBNf
7rUdvp9RAAdWnSrl4Gc5SnV5d7DWnjceacrYh/XJP1eKzE1UqXkGY9MjzAupPDh+
M8E61l8vNGUaEzet5TFkRCaz7tWi+mrTMrmaQDY2JNHzQAONRyucANeB7Wa0YWtB
GnjBegf9jA9wa2RM3V3RiamXMpoot3gegR5ekOja2lR0NRNGGN0rn5vKz0MDg80J
aTfiTK0l2f3jxi2pandfoLX1/KnCAfACaB1BVgfTNOPDXOimHzFpuN5xtsoHfKqc
t2/ARbO6lwmZqHy+kcqKe0k1dKbcX5m5gh473+OlRe2ztvucTbHXezI1COA8osW1
D3UiLFZ6GQSSFeiKbgAM704i5nIDHLHUN6OYwkTgmSzqYEUO7F764J8rO3BDNslM
Exi2N7inTZ8zpOaqZPIdkmL3B5XVO1M60NyWFvOu6pJM14v2apMGw1sQWu+5BJs9
IfLoWetagsXmCnLyR0MLvI2JH+cahl+GXyLJJgcEb4MktY0v34P2XqJOmvSeUDnH
0zicKGd4T/X0kTm7PgeJ8lD2KjcteGUKJprdK4UZPmzH6lCMMwdh6VD47MczsLx8
NgKOzTZLkJvXZTibe3UxgcNL+Lz2uYohNu3BI31NZdtKKhajYZeItoicqUB0R04Y
ZufX8t1hIvbADpAdRXwy0qfj/piigNujD8Cs6wknX5fImnH8x5Bpt+A367jhCdaJ
Vld6fFJoQCGcQRbHEevqhllNzlaUj5A1U9CTWZ/0K5CY2hYL3uE7WJ1ex0KvzAD3
2ffdCUOMRHWylS4dVJc24BN704URR1zGpdZSb112nVSY8f6xZpXEvqhdLeDylI7A
yxgBGGSLKKCfQnAgDjV4wUth5oovWkqkidb4y8CsC+wAexlKrZTkPdE5a1Tr+UqF
Al/mWWkqnh4+29EVIOykyHSBcsLa+tvE05AtYwKw6Uk7ARUSi/elOEH6uQakORVZ
mveV7S2X4mHXtVCLdT9rXARGxRhseiRAiEADMOtCPwIlI9U97pazNU2pvJ0iluMl
ho+koEDuSryVfKXNJfZOX3n3qBJzmXZBJ+EIZoSSdO7rmSiDq1BI0uQ8TG15cEmQ
fcw8BzkDZ/dcjq93NymBgQhlhznDx391rTk0RY3ZCpW2KH8CNigL72SwkB5Ylnst
B4R+/HOM3oqZ+94EcGfcuPhqd+95UieXtOLXzqsmN66nLCje6adQh/WHC4mpfjvH
L7otck+SK4dS+fGzSNr485az2T6ICqpZCgWO+OQWE4jVC+kuJnxTXKRNUCnn/Ldr
lLflkH0oLU7mVlKAB2IYBrVzRD3xe/KoLp/uwIm4O5dFKpDbGWzZs2nbr0wyRHeh
WL9gjW79K/Q59ticiM+Ca2ufiXoBwhhT9GvzXpSBdM76juKM1e0ipJ3Xkg8eH8UB
J4OdXxLwRzzwQOB36OI8pN4RwE2CBygU0M+MiFAaSCgsQSf6Qn+oiFGWjQV1dieu
Hh3ctUcZ40oMXxwqphOKbKZIxYMxAZgaAkXlK7lIR2nOIdeP3uuSxYuNRubORfvb
uzI5JAAWWxQqVLZVwy3QEuKWPYsSJNQwYzchuzcQ8W4Be1e8F8HCJZ+921eZOGiB
Ri+zOKEAOdPZ9i2ctpqUu2DKckKaR91AIQv/eaEmLj+NRAijGbTThneIWAN6t2d0
FfBvXPg8E/FOGSz+pERcaIfKLleOEW/8euDakmI/V+M31jYn6ED3D4+QQfxBF+qe
XL36sojAHYs94sb2CaiXE3rBI4oLAeAAEKxm4EfUpyKm2fKmFAqF5JWWxs6vpesg
9wlG1PsHHHCjxqnTVfaA8ZwQiDe2ZRlYG46bPUclKed2HIGR+ahoxNY8zXmsVWe8
B66kjQ0b+eDbDP42fvZ0cs0C9B0UyJwZaXxloIGGfBlRFpn3mtGQsjrpXUWTenRR
rnyY6hHfzy6t/T3KQlPY/cCz8fitFS46+TZPJI3Qp6nSE/Dn7XAOeMQYneflzVnQ
vXjI2DdT2k7aNSRzfokAo18KwovDzSTfCSmzm5DCkl5kdqCSaPiGwfvgtr3cDApD
IiCJ5DhEU46CdQoXdwZF9VGiegmdhWYFg3/0Ccj9Zu5J5eiCYDuZy5EZEYrvcgmm
tR0IesJG9PfErXy5E47g5CJd4fQjL6kdYm6fwl1BX1OforOCSouM9hFXqE9+Y6Uw
O9jqQr0XBSk68GrpxwQqrMDzU+bC/CNhb2D1v1CutbpDvVgFBvV4XsuWxCzvWatT
Z43W4UyE0kxvxK4GKZc/vea510FqfwxiIeEFZqXXVvXJO70km632j1BEnBXGMhrU
SPVgGknUu0gxMkvgvvrNHKY81bxPgiNLxnFHTHVakLUHUfjoES88/RyHZAqa818d
YqwCfImC29oJBuCUe7KDgeUDijfc2NhIZQzKdyp36wsMRg7KThYBsGRIEPECHAgb
pSIZxjIDmzMxsXPqLo33KXDgyHlHxX8Xbn6p5EGXZzyXzRV2LFDV3GZGvz3ow7QH
bC54eiYarShLurYPMrNqguJXWljVmsOtfRrWYcrtg1Fjmr5BGDrWmTlb+G31B02l
RZOvLGVbszeDHzLjVVy43xCosd0To8wKKakC5Lx8R/MBZHvWy0/vAilK3Y5DlmB0
VdfFF3ArSlcRobPg5oTo3zQuDWfjYKJRWDi54jk4nkgRadDMZebRqGGpfhfVqiNt
VN6n+Wy8NFV/xIDJXg17AoqoJNPBP+JTiLcVV5J3wXHdF0sB7AcYA1X9pDsQbZoJ
XqBoBwRD0DGIyOIEute0qN28vy0tU3Eef+47Kv/VgwUTS7eVIzkCoQPTPkd855xi
B/Io8xYfi4UB6uEtWyTDjJwC6Rwg5LDjCjrrSK5L+LvTRKF+WI6przSu65SVb7k6
n9XxEj5bw1HvJp9QtLOayMl544+HT2zUTHIrey5z8G+urDyeJxTwFJA/4zgPb4pt
pNYIdD8gJ+NrmLHutZS3CxQVnhj4UQCuokFaTeH0BE4VhKlKrVEZfihvXbYYdBRu
SYaSAn3lUUDQ+jvBXcp/nb30OMFTQLIH05CqX5DnMHV8J6uzN8BLkogadCqD9Cxj
8tHw5Se/JLf6tooX/bNZdSq7k1ZyE+598B9O89SdZmj8lzcWT0eab1q/KUkzYGzV
TKST0lWILl/UX+mK7MhikEpK2NkkTcR0Ma4XjY1vQGrfirGSIVfFLJzzGqHzPHFm
qonEmgBAP/AYltDmrMKluaoXmQgb6GRkeXCCO1s7NBJxUCY+ABlyYw2AmMqFcGmu
fcGLIx9jGG9B/upQ1ZUEa0ZDSFLwSowCZPyEDBdCBqTvooJ7bxIN8QnqeFCcPgYS
iwjCS6FMj6ZrOvGQhuSUjRw5gg4b3cc47opn13HKTkE9d0eNIa1rhi+jT+OVE0d3
9wMfqkQLstgusZot1zcIdiJ+0i5ZrduOtgTUjzPXMq/KABrc1gfLsDRXufNXvKJg
k1WTHNACJodHQ6+luZk0ebBWH2Aa6qc8Az5j/tt1UE+H00+GTTkPOG2Y+75TXWfS
PQUKPQ/OL3zgov+qjZjkyupW/jArfYG27ZHpVXtsfjk6aJ0e8GVMo7lUuW3CX+DG
XI0Z2tncmFRtaerVinJyolqJivAlKIeVcq/voY430QD0xfp1N1WPc8xYqml3CppV
iwB/xXTAhntQMs4O9oJtLkqpWQ47Fai4WJsc90k5uakW3AeaKclU0gDjQcUPNNFj
xtA0Pr1MfimcWkkHkOld6hbjGYNe9RFwc5d0PZJV3/Fg8yWmzPbAQPt6EmwQiAlK
dT6uY/hEttBVIRI54adBZ/YA5nDJdKRu9zKHkPGpkmE89ItEKrBA0j+STYjVTUH1
t8aumoQRAIbasba0ulMn9C+5kQcq6LIM691wrouHHtTlGULm3z/jHzxpirrpqdlt
EQvyQZyPJxB1QG+SGmJJrc2eKoaLZvMIuomPKEr3UXD7mdVAqP7JO31YUeOwnxo5
p/AdyVdWLkItqK0x30Cd00fTjxhx8As5fsMXmQbFynQL56srePg/wzoyVShKGBn8
tXXgRMq3vlnTC/tbez6d7udim3vGL5NG8uPgLdQjIklSz/PXrUrljPVAuAJqC/bG
DPpNVObbvUeSVoV9CSEn4+NxFQ++CnovmYfNxGybo9SUs/eaWyckAojIIbYZui/d
NN5WVLJt01o2LlxHA7WxK9pqMB3UTMvW87suKYiLMRG/JHcDsqEwlfmzTjMY96n0
CT2hRKHqitWVPffNxVDSvk0ONNQcjgnh0j51BxbCYQEsyxWgVXm1RrjFOG09eW3r
yTAbRytIlFmy4T1OinpR3N1MCerlPKWXfDmjqsI5I3zcD8IUkEjrYhbbPcyfhLtt
QfF2HfaGMKwxiB9Bxl8E+joN/llxgAk1NwaWHH7hwORMQ+SU6+Fj6iNRn+xbyPfu
wuLbaIrCPSpwlWfehhdYc7/zDgarUECAhzztjk2bRjMdIw0Bk2OjPkoBeguYkyeF
3gHv229Jfm39mCxNG8ACrmrBt9EX/Oh38UEurq92Ha9nTCN2pqzCe7hB9DHJfNzD
eVWAmq4mGHX8IJm7n+89vG+tUjIFxlzB7P9b2f5T0FLYXfoMSgrhlnDs8dv5/HA0
dPvV/OdPAzWlX7Lq3aVJWtHOHCA35YhIMvuR6DOFgmtLyWKh85938bsbfI3j24tk
8G4qq46NZANARPmHeQuBuaca2XcshA5MuIlfis2+kk4TieAC1a6Yp9QY7OnUYl5g
YEGArTpKjC7AQK8vbOCAC+s/tflZ3lRcYXG8stLIkTea8S3eLEyPKhrZVRPjEgDn
ombcjco7L6nWji1JxnA+Xdw42993pwH82sMPhN0RswOktCbyHkD8b1II1uuwO3Y7
rrb9pIeKE00rcJ4ILehaIANKBop/o4INOuPb31on5/G9LenSLSoNDvxTZmCtNlcr
CTBUN0SUwA0l0aZhZBNrG6EIumEwdWSznv3V8T4K7HTBl+AyE6+XLn3w9sZXTe3E
p3opzyZU6SkcurF+h+dmjOvWGLRpRWWts/2RnkrR6q1XIQFQav2qJvvnHpJkNwId
nGXDP+gTwPSPWatxdvuz8jQuPi+IK5dxybNzHaEQXNcD8pVPumk393xcTiAg9vW5
Un8szNd9M3SX4JzSlBIjz0YWSLX4OQVmaCo9zsc4RVmq/PNGSH6ywgOWHDI8ByNL
iX+iBWAhaD2QzRUXhoRagXO9ZybC8ufpV52xuNLoVgjLDxsG8WZQFI0E93hOpVYP
lM8TQXDwuW9B+6qDaFyCwXLJJueW9jey+moXwuHcrdcv54AdFwNyIttil6gC2sSm
JIJjxtnGSnGEkBHiz4nMnhdJehgB4liFgvzVOgnyN4wImn4agZygD5Y1B7DUhqsT
lzpVDD52A7Lb8ky/JCjiimYRHBI0elGkwTbOr6v0RCBKnarJK4BSfUVfsXF28ohL
Oc5/cYc991GEJyNbNcfaa1wPaajdxRH6mTMkBCuNCpVsXML/2Ao+xttt/IO5SND9
9AXL2YstPgLIffdSPku8+YjxwyKGhuwxNAkjzn9Y1yRVj+7HbaqJ7TUM5qooG5DC
U93upLiSzA+4JRZnkkQ6vggaI9NQkHmOfwRKvO+feFFq+EwdsVMFzZQXDMlU22Hx
N1M03lUQiCj+T/jMWD14/5en5DqNSBEAXYlbH0mXzwm/6nd46kfad8DEDmXxu7Kl
RZ28BSNQUvn//Dl5/Npr7r205s3AttHcaufoWn08pVqhlV/FJSnqtXkoCzQnDXf3
2rgjZNFgEzKRBWcg4IV5+VmQsSKuM4W9AgbT5MUAOhVYqUKFvda0IRit/tOVIaLb
AuHahC8X79/sh202I0wpZH/sf+VQF8IQALF6VJioFxT+AnjKM+Uvwg8kEmmahu7s
fK6im2v3hFqSXziF6DrTOjBgBzcI30rbmNAslcjfgoNTCENpfsh67X7QKe8001yU
+N/yA7cX/J4vhqPrc7cGZ7LzHl4Nk9wK4WFaXI736qPF231BVEHK7mDwUnz83w/Z
f9TpPYqxem/fNjXSsYsWFtP0LZ0szKu//aiUGwI12s0Rapr6A2Geu6/ZXVcVXsJy
VtvyUzmClIbtvwEONytd1yvly5Qwc6YMF3lLRX8rdMAZINc/9n0EX1IIBXBtwXNe
gsBs0W6GDZ5e4QL3PFUU8Qmmv8eo6VVovj8LbnixULf9tUSG/iZkFV7AIxnPaAEe
R4QL28Fvtmxjv8geoPtZ5B4GUhOXXoLzNrpwCG9PKrxh8sIRajxu5b2X6w8H4ACT
ueVPZ0rmtH3kaIa1u5IG4o/wPf8vVj22XsdiurEYTCUKWRGQ+AbyUHSD4io/UfPh
EsvSQZgbe6LOtkHGAYxwsICRWRJqFjzCEy731ibpoCfsGv0wBTFmGlrERpGrAf/W
cZyaEknKMgloR+7ZSVMr97+C598XuUJ5T7Y4UHJkI7M=

`pragma protect end_protected

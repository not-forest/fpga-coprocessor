// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
Nc9G9vqz+p/4MZ5n4KePn+adkHevvmx4v5+JHgic0GrLQ8ynHTztQVvoQWbyF5Hn
Ml/2RiA5MJAJWXPLMTzrv39Ni0hN0jmZS3obhetn95KlsvYfyAz3mSqA30Dq/PTB
n95FZAJUA1k17/aCT5jRtf4w0dvpGcfB6/T3pkLMjTnmNUHsyma+Q4CxmGfJUPuL
qeDrEE2SmQuwnTjSpSoDUd4PDxW/3GoN9Upil1NN0JSGBtvsce2S2ZmEngVsq7Z8
o0Mw82nu3SPauWrsT8Oqq+yt2sF21XTwmeLJvkEQyAauMCp/bGBxrRHAwGA8krZ3
C9Zh89TlHyRV47pUSxxmkQ==
//pragma protect end_key_block
//pragma protect digest_block
4bBLNlnGMQwtU+aMruPI4Id+qQM=
//pragma protect end_digest_block
//pragma protect data_block
iAx7HKvoKj1lPoSdxdSWekV4cdBLXyw7lBhJ/5CY/7GoB0VW94F05OEFo/4hFBfN
46IUqE15fjyF+hqelAn6Isd9XuA4Gh4iL3dMeIgvocGWsfnwAnoDHTuNmw2Adexw
ROxyBKrQSZsjff4tB1keFYEKrLk0g8n0Rl332L/dpH4rp99sqDGNuAPDcihccIdP
+XTEOjY5IVvosS46YRHgn9yATXNmOQovSj5NSwl3I+Bo1HjapHTsJAft3MET1Gfc
rth7c9CpT1qCfH7vL+3y64s5d8maZCmaIyBztVsFX48jdyoayuPhc2c6fy+cllXl
R5VVY+pOvMpyftHGo2KxVse9aLbhScYpqsp2z6LDmDd780zJ2pZmLnoIxw0L3+j7
FS5UN09K6C7+ZZqtcS8LNAmpLuKrNaRIKQIo+XZP3oJTUJktSyor14IYdrU8VXtC
Pi1WKgLWJMBE1p3qGt+mTbOEoD+EFkyu5thZyhxgxekZmcNWxE2p6r6gS33zVJQM
awdOwxt6SzRP+q8791BGjUH8P+yRQNi4/T5dPpqnB34w3okAj4KwBugH61wW+9XC
UFcaVChGHrxfQVscPKw2lGgwiqwz3Xt3iAikoLtd3tjLQ89I8J3BAIsKtf9AliMl
1aMbp+ettqAT7k+cepncKlf9q6E2H3zXPHCy3cE2ynex5Z/04DgutICsjm8AoxrC
ugUZU74yBU6nJTuxlrp4Kxy/g5C4ZF4aHlSY3q/CLhjK+P8GesqvLqoQWh0rpMkx
RzjTfCz3D4ZKfl+LfV2xGFvSe2vPF6sVH7bkEJmxApQTo5z4d2oVhKIDYlcBpTDA
jx1P8o7/X7VpYheJ12Ds569gSTO0YfOIFkuVcUCxOqM96EtfqjCO3ScYpi89cw5q
QtFnzRfvaOZ5aYCKVLZzfCcYEYeaTJh9tIXgcvpkpGpHMbx7EnNOvMOttY8zuWwU
BNRb+y85GSt4OAY9WZW1bqjzmFBIIGBeobKsdZFODW0l6gGAZYSAoljJAoFuNZsu
25UhmZSsizk1k+GKYHB2pyi3WPxZaX5NZjE1Q1yXBW3XSj7/gHsujpZvvawaduYp
nTnO5yhkHC2v5+3RLcpKivofMDEpjGdNAk9eET6nx6sJjwFcpke13TsI6cEDwM9F
+FSSGcmBRtO+vBTzN0gveXZF156qcEkjSNHIksy09qrNSui9VU0TFwiV3ywDy61X
KHFyDbxs0MGa38+6KSvEzNv4b55m+ozSAfpZY2tXGT3hAQ2ReQ6eRzVmpnfcf8d3
i3plSaMzhvEyfX2vIRf+4nfvbPxtxqoqyHrWa6jxPxg53FGwwGRF+Gr1w0mNzD+r
VBaano7UBpafd2yJt4i7M6YFUk57ts7yFtss9ooz0mjIXaES4UBeXPrz99MZ9dch
w0iO1XnBrn0BVOFvQ+PeLqu9EN50ifZ0CH84dkixtct6jDXy+NIwSgnOTEMmDX9c
uutWph+yJaNAPEwDXfaKgpi931RyqKqkvHAtGNb6ECRcGj21qUW7pxaDIni948j7
se6TnrXffsReEEgxTeSUDqGyZZRWJMUwfmc5Cpu/yySa5bjLgG7NzJKx+DfPtVD7
hhVMqfjO02ypei/OYhp72o8qkMoZfQKkCGT+A8ecsrWXu2ga5U/dMMnq4umYK5f2
TPOvzDIGRhCyfIAsimxTd2jKjlttoehg1OKrxT+/3rlCTXddrsnYnlSvIN2J+bti
tJo0zmzPR2xRGEV4j5Lvi7F3i1Im4TW9zpRcLWtL+halT9rEqs3pNHjVwnK+G9mZ
+FHtd2jyTxxFZ/PvHyBGHSYU1hoyq0uUyfQRbUshWmgIFHLBpeBBMkwcFIXX2G0j
Ax/0W78zmZN6xQAltSebGfBwBmkJP/4Jyn0203fj3a99az7/a3nxM6NqY56dND72
zSLxsq5rvNxq6sW6wtBU6+0ZpyzkH31T14S7KTBjawukqgsG9h0nnAUGTxy6P3mj
RE7LieE1wVsMkeI42QuEUG/zFOptjfzYQsBou7xk96M1fr+Xt2GAfqlsy5roMF4C
qZgRbh0Ha1Ze1EEqKXynPGXmJo6MxgFki46vZOXq4HrsuyGcGz0s8YBuueKRQIqO
yk/ZQHdjKO9fDJVEA+X4+xxW63qvIueTdRoKF5pXtk4cp78xYQtatI67vIc1kqrc
ReQhcW55/GzPsO6bEJZ1OAW9k/2OqSmxJQwzlMNd2zwvPyavJDHbqc1BYXdeHB1c
IkX1rj4hmJCUOJeruYiSPpbzR5uaJko76D0XDPhejnmceeRO6IyCfEx2pwJPHqVK
3gXHTVqOoU73Ck9GNNmnJu6PE6kuVSDqchotQIi6VCYouvaj6Z6Jm723VQhF3K2V
uSeulX1kSR6Dr4ZpkCyLs9mAM0xVozEPmXZcyeT5tRC0GANv/hZr9fIsPkTt9cuC
ebdVuFS+PNJntyKi6UqarCNUZpiKxO8kSEjk3Ehp9E1T38lLUKLBfF8XydO2mc83
KQdbTtJzPYiSZCkvw/JuJttdEwtZH6gm4bK6ykBdklbSX0VTWmg5OlR4uNvrtetH
ulzIZcUf0m/Kwe8FzO7TKXlZD8Oej3N40IIKSddCrU9mpMPzS3U2cvMXjzjCFW4B
Fnq9172XgzA2+gnBBtmodrB7/PWIVqPSTHNZhRnkASG/8mxFE14nJSfBl6nSODT5
TexN2bW2d+9LB+pSmjValWZXSfiwdmFknEib5eH1WHjoDH+D5QgjGpIlbWC/5KMt
syj1TwzI8JfxDzbgv2jN82u2rf6ssTAcZlBthxk/Mrg/fPNptdBKPh9jxmf4PTGH
pO7dQT3pFhmzfcxMIbPcjppRSIyjAMqjb1J0nAcySqlx6iNOZvy9n3walOldA264
Pt6tq1/RI6bMLBT3JsOTSq4JWMdzOO0YFJva3mUuaSGywJi6kAHjsq0y9vUVbK7S
7onADfQNX4tmLpOyMoFP8IyyO6nL2yzbNud20ZQei4QfMGOmO7+PMMorYjrTvjCR
rPc4TwVRj1mTYAoOLi3wUkiWglja8UzHoB20UgowsyobqKZRG1M7z/NRXlGLwRJG
TQLPKLCpa6/1lUqt6uimqibK2s8d+Wrv1J84Cqiq4LFn35xeuXfsaYdy1+qhsSOT
Wxvn4vo9677mKoZfo79iAiB6Wg3uqAXNdHlm0kBRWDEFaXM1WD0GFISMcKFFosVE
z0xYwnyiOL1gt3MVVLBRZ/QJQ/GHo3byGsntglDM7W466UsWUd+ZoX0w6hMlIxG1
Ft2eWGznenhqII180Epc165TzBQeIF6D403WdBvFNdmkIqM8g91y6heC+YHjKp+5
vdLNhIcdjoBG7FrecH5FHHGibIz0k94oBwYFWP4ClTgXBQLSiK0bP5bPrAmvblWa
kWKDf7dvIhqgpnZnr9G/6wX/ErXePYo3wMRvi6v/87LzYvy6BD2fIeLIvWkXvi0R
3QUOa/SrkcEOwOc4nCTugROO57jsWvahvEdFy4j2o4XHKCPlAiXFqb3Ga0GUJzsk
9VE6569H+xOstBghqmepppH5nbYFXAqG4xcbhhhqIld4lnnIuAEtcgCOkR1ZF3O4
S83Yx4DUwKSccLDM4E7zDnurROYqJi2CjFqamsr8eucOyuoOj8Hvm8ROFRxYMmfh
585+9jrE6sVWP25noS0dd+vo54dUxUbYP79ecxHVFV77AvHfwWsObd9f+V26Umpt
OsR/pZdQzTWf6LohgtgahCREFZeUP5aInGIMN0IxiqZwdwBfi6WrIJnvhZqtgIiO
bCWZPx6eGjz9l9DSGc2WhqPr8PK/1vcZzhuubYA0odPv9s8jQ2d+mia98H5wrkko
VotYEhkJurKnD7MHdIXjrFUMlQW9ZHLN3ZsWxx87cadikq7V4g+h6RJTeZxKxw4C
kaVrW5OM/XIz1tzcqvRDBBvGd5mUUjVnKnSCCQPPIhLtS0GNs27PgPKWvFaxSj1m
8E3WcUQvjquoA2Skj+MItgajw4q/qqrCsr9fdXO8sDSa6qrMe7FJTjKHGXCQBYQ/
TJsvLFyi74Di/2Y3AUDAVt50/Ra+/5wjUAEWjVO2rwTphbXKL+cP1eTcX1A144GY
KKvvzMZFwMTeR188mJlbeDJxHd+SjkXLVPsC02ql0WQpuflDxhSxZrXAtPs2O7y9
jb2TbHSXKP5nH17jrZMt9OyLs8egOqyeuWt8YJ9IQKL9QPyT9bD90zYynKJjxtGs
ZT+WHyivatLwO0UJpach/HIuMYKkXlxmC0jjYAyriVJ6r/oeNux3iPRYdKArfX/X
DUeEPF7sx85KPRDvElDimcDSes5IHvI7DES4P3x/ywsEAbam44FydFkCo5Tgbxis
FHtn0Dphgu7iNGAFxL9N4Fur73kE+B31F4/aUCf5F113GnY/lUPosrc6GHK3p7lK
ogvOetgSpHE54NmSlV/wxwgskGKIzViHyqT4K7eaSoNZd8fN6c1BNs7MTOqtIZyT
/BaiaSKdtIhY9LcO5TJhLEJorSHOBnSDiIujW9GzJwH36AbvSq70z9YeJLdw+mcH
7pOReXeGopQXmogfxaDCyvrjLCN4/i2gX83lGLQUIM21TwCoPEcFua1AihalFEye
yYiyC6Xh59W7wm9ncbCWZOwLXGW3gHJFOo2oHej7ZYTEY3vxJyzZxIitBaxrXuvk
syCrnUS4yeCehHc7GJJQefCNf4cfKzq+LAYsO05/t5lzHGqSXtpchpeb/EtrIlpd
JY7QWSajMyPeGVGeES9ChLZtFK8MA/569lm+uKrliFB2np+QA7k21xOb9ynbgy8S
zY1HVl+54XkavoRNZTgmDnFJEdbPcrv6C9naQ+YNQ+5zhXuaS9DUa29EtIN7ZGVy
PfJj1oFa3YLlnp/VIFxQuTwOKZSEEYGIODd4nAdI4jJf2bDtKZCzL/2tUtaPGg2Q
P/SPUvs12iubbkX2vXQqX4VDP/8iSUctMVjvWu1M5BkHRaZI1lgyTjiRlDf+hHrW
Yg5tvB4XMuK/loFFKwz7ml2HPXtKooqNvAA1qKwoqDNbcDVyHLucp8NX/cR+3aXT
sZpxE350m30KRyrFUR0zOi1/wC+M+S3HOJwJfwHJRxIvPniLn/5v8hzoiOqm4RXi
3PylrA8l6QtkkMsRRTjZtl+TwHzPNztdG4NMnfTPExkOFl3NhaW3IRHnS+HrqnfG
FhJvbog/A9CQWzcLNK67RYXKafbvVleoVFlqa+Y3D6rmx1JZqMnvvUJ/ChHnqRzv
ILGbRigz6vBUqrljd3kdKoVigpCuadaB5/7C0OhADasVmiyi2Jkl9ksHHY2N2CBt
0xPIGnc9gjtrQERlan6rAB0+37nqkwc+0TZKXreHHENuI5E9K60Bi1oJvvZA6UKx
/zIN4yUxGsZp9K1Y/9IeejPOgQkt/y33uv4qTAJfrYRmrleHeZUOgXy48rQ/bn3O
hHFDdsNN0YjJGWtpbowHygkHsrYD0e+4vnRC+dDO6POa7d/fWxpXLTcoz9P5Nasc
nI6AAnqbGqmVDejMg5jF8d7YUwYAYx1ZcTADuBP5N6GIy4Ce/SpUgwDlqa2SAW+S
H+iGsXGIcetYPPiT9xRcOz9RbhifRIalkkaIH/bAlzsKx/HTkXOJeSQ64F1JM8Tq
4VdsHiRBbPpNlFFu/QWiLKtoE4Glq1OG59ORWZgWOsh79VAw+u9KdRu2sVW3aOMR
fOGRhSMsH2VkcgivBSoW8hG440aGFjwLAUmAxWp213XZc91SPFxvurbIpFPX2s5w
wZVL/jJGN7KVTQnCPYS19M125Jo+9qHk4DvQaK4VVIAT2xIT3eIkzPPNdJGgUHI3
yK2C6wuHrAQmVRCJPbw2SDx735xC7RKpxzOYgymGP54kbY95N3k0GjzvBZmANdlB
3sefVXU0Whsy2e1oGtzVma4bUGqafc6TBW/oDr6KNbQCa9LuWS4VlX/6jiRUCWSR
LLiyNU/iJO/spW5fTR09kY2C34hAuvD+pVV40YIJCweZbfYq4ylxIR2ZIpWYLfwO
1/KbErRDZn8zvq0Ay5ri4sbOYXl1N6xPv5iV0nTrF34+yQVXXBQNDOQCq6S3T6cp
8kJxOfjai92DENcUiRZiXf5tv9/ibEcHfy5xjSu51uZIVIE/dq+hHdP8gv+afbUe
FVsiyRoyiV6nhGbmiiDObakjw8MLKs0O3G4g/rnjkr+QozRFNx1suh3aVtFkwYA7
a1CsS1LF105Jop0xRUaphF9ktDhycndymEz2NeWx12e54P92yQTWN3LzsldO1ruO
u2M12m/SVuw1L+A/qKkStoW9NYxNJchPca2gMVc64AcAhvpLAIzwfRQfMuR48BEj
MnzXKdc6utcs8Ewk49we/RpCzMJdGVyNBAn/OEyVIuc0A8vv8AOfh7Fd7UdDhHQS
R/9ba1PrJ1dAw6fbjrjvfZofQqezSyhVaa6z8ADacSypGBtPdy8uHMg5/0sjgmkh
WOMZUoV9MmP4gp0J4QLKnR3llSWuyhH6VSEKUhKE5/Cbr2ExGmqlcSm4T1ziLNGZ
1m1WoP4X5sdLisBWgZrd5JyZmWpkvT8frBvHvh/+4tpC9IqNbHNDCMEJGZaQiFek
RVikRXgcAYYbcs/XYvbIvue0bbmaNrJVrscMjpGd/4DJj6cygjyXHC5LiyQ9Bd9c
0Sor94fb+fgapvOajVqDYwmTk492gw9K/UWkoFjdgKpeqd+wtb0KQ6rUZVcKX0EB
UOTuHjqHtr7MyRJ9UsTPH3GYx5NJGJYZsZtZBs7V7eUvmANVCEDRkU2MJv7nhmqR
EcrGNN7eLZcIDUYzBYrvlsdPSZPx59E/XepiYsumOjqDRaJilSTxFl9YjucX5sTk
rmoIT+oTLLN/OgxeAYH+slc3pZa7a6LxxMds6eHd5WV1q/TyghZsVqfoRzRXps/m
XcwIwAoRpg/A76Fi3dma4p6jnppF+lR0bxKHuNghbVFfsBxhwSF/YShrUmUr2DG5
0Luk3Y/PcBICx+iqWhrM+tj84Sspf+zxIlyqtqo39OZChDeOd+pijInasyJvHrzx
iVPK1QtC1vCBjDc5EefkumyIv29kw/aYQpbyhcUYhRyFVNal2upa/eEFq04pyxMG
r20o3tY/h1N6FM108+at2Rd9sO1Cxo2dulzXsGFjaX+MqFwCo8uLMYAfntKRUgky
JQjT8fXoSMIdQTABwk1+MjkRgXD8pWSPaoXzTDNfzWPQ86B0g1G/kVwOgSFMH87E
3soLIsxbdxWIvk0oBUFD0WsLXBW0o/T+cZ7+yx16gtc0KuXijW7gpwG+FRCnFKv0
Ov0NQAYK21OEp8SbUfrpv10BZrjQHR8lOruOaH853MNqSIrz1tPO2BUd/uRqzpWl
JYuG6upgYkI7WsRzHDVTBr7RYNLHdYSTtNaWMEpOki1xrKX55TXOHifA/ZNPkba3
wfEjhEE7Z2ds5uAdl2THRg6/kjYNGAOuR8jf5IThy/8XqzKGEhTzvP73WTVPbGIv
WN3dtQ1mivT+T9jvfUNMw9HtL7ornAMkF3zWfI0EG1QbwRNOToh2flL4nFbMsqij
F8sSosxUPHhwnPzqmIiSmnrprDegw+y+8eQFOH51ncNmSyvgfhjVOPEoNIwn6hWQ
StnTXBOfmKjdrpxInwNiYG/ryOxKSOwZp/mkvcZs56XJ+xm9uiC4D31DyOKENBwr
vJ4FnYhJr/yda59CCN+vDdcgMxxByKxvLgDgaPOQPERaAVnkdWtE8UfJUO371RKJ
+wnxuFP0IHp/zQlXnm5EDOQX62zi/Sd21ioXgbOoHS3YeJm2ATYhqnXqnhHWJvk3
ePLmQ3bFYLDIpsJKx/bnwf9MnzWLHjOMJD6XEKXCXmcUx9BDan6ZRE+BZrMi5diY
xY3KJNRsroVrA8WXcxJsvQO7G+21j+Y+aFVvpu9rzN1osS5tp9xmOuAUCFWhWmNI
SPC/FvDNvSjvFfSZckVD8xsLtPb4mvnDLpPtMD4UeTe1rYijKsrPeJno19z5e/AK
eDoSh1E9iTGQMM67GI/93dDxDAox0wPSl6cXVGDQthHBAhSIYrk4Yb9I89Eq1MxQ
9bshmxysJTuYkvm1QZNzUNYwdzvif4hR00oyoJLlT3B8DHmLZf1J4B84G5Y+zlq4
bHFPq8Apf70DcuirxyT9Gn1MyJIgMWtfuGdSxJrX5OgKdby3/9EBkO1C6Z6nxmMJ
t6LvjIf1RueqFW/x078+yBPcbORyW74B/gmBfPIU2Ke67obPZrOatcEVY2kt+O/x
Xx5zyJKttjgM6nxuKGC54gtxoacGBP+GeW3KvwgAt+PfxJ9FmU88V9yeotskEci/
VN3dUcLwlZxlQF6HGuX26DySPzOhsRyuIhqyJByMynpcgZ1jHQmmzhAZrt62xzvU
m30Jonu9wkPPi+Ka4Tzkg82nxDrEKIVz56XWxDQ/oJkyEVUMQvKHQ1mpmII6QjfH
Xss36pm2dFJhmQw0NNYEzg7Xs1asUJMIFpU+hQLxYzkw+H+HdgHHfj99hp6nSsKA
Z4LahXy1bPSAeoxQV4zIMp44wPhbeQLAmNI2oisFT6ZT484qh671ojsX1C9jG03D
PXjY37M3M6feXhVAeMx/Keg6a3hi0BFRJDnGuTgB2ovAxC0QkiB2Y0TdlN5RYLnF
f+HBK064sm8au6KiC47GEo9lukUOjEvBd0iOblFqRhVrNbznNq7+hMhWUf7cQUbE
iSmGy2gWCCfP1jtRzITHDAdsMxYdCN0M/vOgBShDUXTJmKpUejrFCzjJLk3ml15p
WyeIWzkRNV2ErDB1a/NYZ850iXNJwwSl+8s7gqTHxNRrLcLWa3TNCzNfiNdVUDRw
lV2a3+/6NFvffCWnfK57SN1tNutRrxQmpUWIExdZCd2ZZ9DUm6QvCmlzXx3e7H4p
LNgMg+w0wlFXYIGKl1bLKKGWpu/NagDhehfhVFLUFRbnpa3UyHMy25gDWJVR7b9U
jm1RudyxF9xSLOlB6aFQoz8H3l4pkCV6Z5VtDiht6piQdJwR0hlpipiLc3hj4Jgy
dhmK8XsfeUnMypXGjL8rud8T5OogeTAP2st8mtyYChN2QdrqH85S8KbHb9+G+jlA
L9b6FLnpzAfsDR5t/+E6hYc4J3f7fNjz06ytq5W92fblCyWd8WF4EfRnaMsgHKJl
3KkZ7PwpHBgz34h2jBpDNT9RfCK4lOdVqBbadKGdYQJgX5nCr6JQFVAnFRI8qfG8
0DmtdCuD0t1h1ihttkdqX2rXoY7fA/XBBxYdI8IvX6WhIeYY++OChwEBBD7AtOg0
r5OdqsOAMA5S8eYo5kL0T/CPRJvoGO1FzsVa/plOXG8TJvLp1oM4eq6Do/Goo+Ju
e1hORbddnkwZwtJP5X/POlDozXwC1xSnOLasYEVKJc+pZNo1JB3rKVdSsedu1swZ
HLdmYSEaqecp5uxRV/qGdNR94pXbXGSMmobBbtQUi4dBWsKktJ7IPux2HlVYZr4V
iCVOYnMem1hFn04uFQ1Q+1OpevlZuJy/9JGwwGhEW52qRq2PYXn3H21aR9WuuqRh
asBHHgtPCKTwpFVQZOw7lapONfpsSE7EsheejIfZsPTrCkXjOtcDqO/VDzVmEz2h
KfZkUpaBZxZm3fYykAq7IOch0fFFCnNwxmDkcUpnJQj+g160W2fT+Ib1jqPmW8/t
Ds3uTsNT7dbhQCnj3Fq61S1oUd8gDjSrpZREQ6+xD5XGXjDtKMCdEcJCqilSnDkd
R3zGRAgdYihNi9vwlhZM8Zb76JaCWAu18888+3SPWcy8j3zmGjqanhXysNj51jAQ
NAR1xka4EkC6WezlmLhXI4HR1Nu6u1LoPwyZsfvWZaRz6a2zOUPgSj8UkYFr/jx5
0JVtG/RjOprCXP6k/7+WR+Fc1t5DK4DsCauGghNBkJnUjscGVIORjzrd+iOCYTBp
RElVb5Z0cYhhYFQDGiyvtHAgXZv1mGMCvHitJY/hW+DzphGViUNWc1dabAtN0wk9
NuD2B+oEUFOfcZFAQTXP8QMk7xJdLtkn9LCE0QyyiLWrpGvx0qYawQAYd6K/wZXc
lctMHtpSxzjaxPncFmNF0nYzZJk0msq8HnrGFYfUdFDvkJq72jtt3QQYh/0QkwTx
TfqlpTYywrH458sUdllkCQqOE+qHbEmjvnvNL8/CFKpBiBFNDvFiOMsphiIsg37p
fwDK7sIq0M6B2UK6Qs8F3wPDYyhjfdBQP9HUuni0SfZFdpEpSjAmWHwbgZg2pK7u
cl9ZfR0xqa6/tP3NmJICXe3txD1gK0JxURC0CQuc9WYoIdtHPGR6fHT7cWchm8Rt
PVEa8RRpsET4JzF9ULQ/yxwWATXRnCyRlxsrKemhfhnes21RpXV9ayVb9iD9Uv/y
sYk0PW7jMRn+29KgO1McZiP+evFpyv8ytcg++OlzRXLMF2j3YmUMqaF+pl6H+LNx
h3GiTvMKdOrQ07I2NJfJEA9fa324lFagzcsP741hq9AukZO4TOKcnbtrllteoojz
VbcVm1+IZ/g4Ogdyge+U6d3krJz9p07Xsp5xQJvpN00h2N1DtbpaJWrJxVq0Ibcc
qyv7NSpJgCg15LoiyMMvfnclHAZ8nrvUYs+JiTNt7Co01GpYiZ3pWQhQmPUTXI8P
yYtN8L32+YR9kydWuT4+iTp36dkO2KCv8xCHF2VsGH9LrAFOZnqT3L5AKQfnzSC7
/XrZ1vXHSCOQn8JbA0DTwwTpbDjTsbtul/gEm3OzmEYQMc0o5569wEMTrn0WEP7M
8y8rHCUu1Jo07Jl+RL9ZkCqFQ2Stpca7MeDyXDu2k9B2oE8A5aDEnZBwOdGJljtx
Xnxa2MbuuD5RN/wIO4Gtznxnhp+aiFFVlJIvYKxrLm5ck1BBWywQTbqDtbCyelUn
K+boM7AQFb9FkEB8X/Ldt5XqzZ7slU4Gl1SZ7rnXjUEXRuI2VPJhn1sZojNnZaed
9RUD8W0JrgCJVk06MwhyTbDoJ/inhhEb1C/lcUsfAXtB90vsrsSKYr6/q/LKxi/G
DOEq3lf8BAVWgU9sNxXi95rus8PdzTRaM6Qn9zt2KZzgsZUSzx0xFwIN0SWaCvKp
csf+CUQNPCmkI7nuq3pH2QwOzsdOanJ6bhLQUeOpc2wNUWONoXJMI3dL3s2fUCQa
1Ueu47u/nG04EY/UVhtvm2gQErp9evUUHQuAxm0hmuwF/nYmysGucTBzUfZ71CmZ
Gs1jvsERHXJ4M38eoKyjneq0A3bX/cN07p0iFXwwT6FnsOtbbzYcK2Y9eh9+3Ges
iJxi5c3JO7afUwzn5u+B/Hr0PwY5ywPaShv6rCLOw6fe2VibxvLMSbsEiATnwPFC
SOglF8Ljrx2+Y80YuX6rdq/puQrOoyUICalxbscnDsKH84wna7fy3ECTfCTWB6/R
uw0s9zG7365DEn06AGj90IZEtGuJzY/HJFLBG7P96tHYUdtb7G1JoANUYQQ4V1RL
F9CZ35sy3AKj0hajg3HfxVFbfED8giod4KgxBJjQzYYI/LMw5LuhP8v9CVipmRY0
Ek2zMFz50CNlDTWpnYpbDsA2Jw4u5TIFA1jJAQhRH520r/KEcOG//mWEZgcejO9G
CZ20GYOq+7rw4WxzXq/S9aX3kAG8HHqxPgRe+Ojg8KwVm5qeccS9egi8JPnYjKUc
mHVt5uu1zZWkiF3DDkHYacWCWpkbd7u+qgN7jHHa6FlCDUCdvKgPZ+KFTCcipg/b
IzH9JlxC+89TmsC16dtrXdA/SWTa/xS74/krCyOi49JBQaDVjLbxgORYeJTEAnBZ
DxR/BU9rez5mR6aU5ybT3w1G1uh4nSvHNtqUkVAF1kvJF0tDStBCn/N+VQgXD+3m
tm2v1658HdeFlX1rgf08I6fyutYOhC3Dz1sda9Tx6yre8QB1apqmSAuYn6huIeWY
QzRokEL1SwHD2FKyoUw7bE4TUH8T8LxICix4ob4zzmtvdiNKi5sQeZG5HdkEEczj
CVcfgD8GF2i4tySvg4hISTNI5jWHule3ybV3efzAlRpd1GUMfSZLugcYJbGDUGsU
2TIhEfnO+/n2Y7rMi4e/EcRBdqM+j9U0dp03e14g40MJOnMqGHxOWCw/MEUO6kab
JZ3SEvaMdBHspE6p+OtYthOaQn/EPg62SvT+km/xIYGlzR3mOQ35mvd04M4UrM87
ZSwQWLrhTmYYe6GPXw00QK6PsNJmEQLMA90JAxXiR90B7JY3lu89h0AIC7MLuh7m
xq9BMGVJqeXgbycznV6k7K1btqEqY7swmAnsF/LzxnPfIdgC4MlFOJEFZHik59FC
8Pe55igD+wzEiBP8VwQigl0Lr0Q+PHD6Ke5fmmPE0yZhksw1GoUTjih4bs3HvpKZ
2jixkCRdGYE1ykaPAUGKLXqHsTEejYBE7feE/VcspUufI3V+knLXNmSUYCjN4rWO
My7Kvz9pIJWd5QDNJGXJ/zXRQ6P69ar07M1FyM9QZdm7ED2tgcAAsw73/IR10tSZ
gYpuiI0G5+DK/DbwUKFNpzsuu4XWkYAAM1nPQVfGbSQQWJvrQrUlvz3jT/rpepLp
pGd5xxFpw2JSE9Z3eqhcVvcfkkTC9p7R642ztqJZ2Jp+GqCiFQkmUay3HXXktf6+
Di0IwJAZ1bu+adJgCOiJDiFJXB5piBScITqiyBaSMqcq+bGdge594bM0DvgnZij+
d+0ZAbMftSXHmmT7TEzadWkKpULZo0CJE3aXL+bMeRMgR7oojsYZJaISn4pz2wjk
g+8LubWaaZu1zttDhmvodisOWxe8X3cXyIaAIG5LCbpVn718XOI/RzUs85C3AorV
UIS/syZE0aP4PdF+Yi6uI7fOsfgVLyyt+0lPfIXYM9GCQCns4xiNPvA6/Mn4rYYj
uRVS72RnRgm2qOWye/IOjMaIgNd8+w3NqdyPO4zsIOPE8DVEZ1zYrl2tvlvXZT0G
A+jNq12AzxwHqW61jG62g+prBr55vJ2O8RjQzi2M0a+WeEjk/xKpa/9rQoWwCvXo
rL9BS3Ko3R9e8MOXgy57aVsiL9L0K+35Yp/XfBzdrxcHNmydGfiMEVgZV6Bevalq
C4bAArceNuyKkftJqVZiXbHz6mT4JsyO/K4x8z+N43jYMljk/GitZnaMnDnjZP6d
HS+SOPbK7nDHw5WMCiUeNW0KtEz+aoUNMORC35oLNwQlNgtloqWUNVnkBbdH+DFU
S1s+BmU51YKkJ49jBgV1TfCf9F1A5g8lKbIc/tRZERM3UEQY8TfreQniCPe821qw
/sBoLS/GSurhG6k5VRc1sFoyzOsHA2v1f9ZS9KBN+c1jM6d0W9E9N+s71TqztmhN
7TqbK+cbE36+nW0IZiTJ/S1ij394r+xMJO7+dHm1XTJgAS2LvbzP93nQbWvWXP03
bX8TmriLg5MbLb37FBrsVnP25LVxl5uy97wBFZtDN7cp+CldSnVGIpjyV2Ig8VFB
sXR0VA8s3d1BumJcXbaZRrCBKLMrpQErQ7d3PMjqqntBQX+F5KG6fKv0E4Th1Dpd
pdBUwkXp/7oqZbfzbozMDsT3Rhvx24/foZ6NGzQWvWzODbK1xEjCTQxE6qwuerSa
mQ2muiVNnfHPXQJhMYcyuPbVSpOMa8wm13uxEXKHpHFNpcZ+fk5oGkxLX4GCAPrh
gVJgE6MdjMwg8/4gkc+OVFioHuh7QnUoN4NlQX2gQNwxXtxUDKfvUrnQTaWgW0Xv
xB5S5wfo7GR6roqZctSTy5k9UPLFne9Ip5v4xzKUTZmPh6UfnRQosOTAjhJnsbij
OQlxDrcipVarfR9wpf322kKs9Yf+aedtFyrErT6bMkptoyN9FKR2L4aeW9c8Tmd4
zPq2OUzkGGIQV5JXMzbTYnYiIZeejPnVePmD5+A957IIIvpaKUb7c5O+U3O+VmYv
pF1HyuPhMe+lQYLXKnil54oMr4uojDToeBRGBGT4pNYOMNY4T8goombDuecK9kv3
aQC0df1ily488ZVm7ibw/wvrD5TjinJMpTLrMTMJtQikEDgOEBwHj/ONoXrvXJCj
YWmZ2yxFpl8K/atDG/gRt0TDWyrJElzBTRqAaxN8+d2ThpEmSfISl75q1JWnwgYt
u/IFWkogDI01pk7TtceZMk2o9Lgec7vZ1CDRGZW/kL/T8mrdE7WuzbcEMkuTJto2
u+GvbbB6VceykignSYiDjVq/5oEeSh/KW0/W39/7NIOi1zMNWwpYrofbD9AHAh6m
zZIa45Fs9CTF2Uk6FjbMIydoh5TucCqAtyYAIsRQqsXrN0DP9q/yNmSvzx35ym6j
+WJCUudnMxWLTYVfsqBI7xforfQoEDLfMVN/TGyN7DpmcHCZJKN9qonO8XpD9N7O
Wh5O9lgcYd6raeXReUSEMaH1lDvBaeam4cSPXaBlMR+OLzH6vAPslilUsMR/tNuI
J4ErBIUBc+x9kzNjjJkf9LsEJwEpbQ3hrFbFBYSpFd2iWR/IbS2OiyCUxIMa2QoX
cFJZnfUaoD0XmV1qtMQaNpiAFbIZkRp6nG6Uvibiawg9Psqqv6UV7LceJAtKn0te
g61tLopyazZtpftc3f3qtif6SBA2kNANQXIzGWvmxKMYS4omrF20ulKW0DerdzDV
dHyCJKgz0ag0XfIE/jAXHzeeNMcYSDjrOeDj5hNuK8sAT5QtHtGqsNMVQ15wGLy2
IWu0DQh6e9yVfvpabcs5FKVLJrZ9mxqOfATDqT4ajk5gEKItqPYgxgRgW5ZsVxz/
ySNfYKT1IDBRzMozhdhpor95EZ8bKvIWBMChMB6A7F5J3zYUsh+Z1bCMv3DYx3xE
7PDIV4rBjNdIj/E5FH7utAXO0+821v5mFbgm49+FMtociS56+J8NpZH1JeecC1dx
C5YdUY1O20UBjmVe0YqUPpHp3k7mkfpqVunuNf7AQlRVuKIrObvhaiRwpSJu2OL+
8W0W5YOgow/4wGL7gyYt2vpafils9Brs0ym5W9qbUdCflQk+HOrRXR2xzRd8syxp
HWqmqs9HwlkHwL7QIEIh+he2APl4kXapN4H2Qw6Or4ybzYLovlTL5OHevOiBhSQv
fIVrWkTJ+o8hFYgs8Y585I/46F+S9u1G5n4sbyboyrzqsH4T1v6ujBjdLMzp7Sc2
tyOqlZyvpCRymamkDkK7Efd8VAQwdgYE0m/bfC3Zl1qblD+ZlE55FgGYCb6RxYrV
MkLerdiRNV05FQAB8fZd1EvnUfUU2ADlFsVtvPGQpTELnat7efl72KzOuBQdnPas
tRLK/u8W2RNi//GxVtMBLjixxLVSzikjkylCVpusyl27GuQLK1X+oyxDY/G8OCHU
oYMyj6Z/bKYDcfYIg/zYystebI64JwzTg/4n0q5jEJ69jUsJkFwQFM100tMv6JXg
/uKQf9Spyxii8neqb36azTW4vgmG2yMDrLMnoY9wbhDafDrdDJ+vuEs1WyfF8Vmh
iEHErhHvPrPnKNbk4Iqqbp//sla41KF8nB63q3bi92Qng1kFAqOe2GDpBVcQGSKA
aesXUwZLdwuXg4HfWL0VFFFc6fxCXXCb45p7yaw/Ryavk8KJhfdd4DzK+a2uZdh5
Af1+egtAloHzK5dMFMBkofRxoVE4LrY+Nh6YHBZdIpmsY4e/Gz2qn+Zg+db0xBEK
8LahxlSdQU13wcIoj3bFBZQLiIXhnQI9uOduwR5QGbakrGVwPxSPlM57wPN24wP3
rjX64besuSsUhpHn7k1oX8KakIqOLaO+icuoFTZU7XLIxodrXI/b8paSJhx5rlXk
K4376zdFr711j7BzG5Fd5nHVJ8/WmYK6T2NxQq3pfMkhcPbuWSd/PlABHHSYFTPm
/ylxHf9S7xVV0cLjw3Se5PJbrgcR3YOF/ONshKcwkOuWZfIt1c2+SFj1j7WSaqLF
03wYPU56koIt/dad92eaB9FY26YI9erRS+DETpIsFpO0A70z3YPe6RAewCEdGYyo
wrio8y1BiHoc10I8y0gTiTNEsIARhnrPD1TlD7Gy2Qy1zG8wONmkQbgoB1Jjiyzd
Kw3yrBE0V+FBAOIMF5Zf5ivi8qGu+QD+dpbQryaxwIOdBtun9A740meTxG7GAVZB
+RxcpNiHrHZIl+VIYpn4raNb9zqoVIyC+/SJqEurHgOahLNRzMM/HMfTmVsURto3
jTTBDa2S8lY1zyaogOMuVd837Pv8SlpEXNGiuPUiXruYz2h9HSHQdajQk8xyOVbH
6fWlLq3D1HiFawf4+2w8fNm8hPgk9UhXPpaFKIegc+GhpsAoZtDXbtT3QyPMVlbc
gmzjyagOyVq6QIasnum5rSy4SO8q7MdjeJbwMtCnWnzuXv4A0u1iJnDhtvNkNU5q
pvTbbNsqBXmQkjn+t+acD36q7DQqUho6rhtXQR6kADw=
//pragma protect end_data_block
//pragma protect digest_block
QgSWINyP/qYcB8/+fQI3EwdRsuQ=
//pragma protect end_digest_block
//pragma protect end_protected

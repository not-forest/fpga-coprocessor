// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
c4Hma0rUTLAqkLB7XjTMVeL2nK67maOwSpUzLLoztIDbd+d/P2599e+ANwaRekTfmBeegxGUEzPb
NfAnbafO7aBJ3+ycTYDzcaZLP//fC/Tp429/YHtY0c+sbiKxQSycHtBE5At8TpYaLfWMkGL/CVpV
ZT1/iaXdI/XIOQt781SolEqH5YHUvFJ4+C7dBePfl8GVTZcZltFxQ9M51pFtduk2suYaZRmOhc5j
qZq093RGVFKknaCUO3Kn0w5NbotEJhehub9etIsPxDFrMFkY3EUg4tyK2sUPGs2OY4xqK34PtlFu
+46uGTIoxdjsk88j4nLv0WIaMLYo7VtvXMRK+A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 31296)
D2DzGtruq4sbb9ApKsd52y+FA0Y6kdeNQ0h22abo79gQj58eQuLpCyC3a/6w22TNEZV9RXYR4OTv
wwoogvIpmf+S3knCqB9xXc7kZK5yvpnlqckG7/UO/DZ/0qhZAXV1EWxoFk9fDQ7uC0zEhZQ6iEx5
B5nQgEHGLWm1HozCe1tq6CNpCDaFqiYcv9y80j1eUQ1OVSVBnsPoqZljzhYwfetQJIQYFQbQSVCi
weVROTDrF0bk+EyB9t4eaXkBIHva/svwN/QJAVxC4k5aGbDcltBHEviE+OpFDTj46R4q+umI+ndP
VKG3zAvZudk3E9ZyDfrFW10i9Y2KozyNva4XU5iB1eXWN8X2w/JBEnEB3Tdm4zDf73wfitK3nHpl
bKNDw102SUDF1GijpyvxVJtOKKyTlPCFnaFVQkVJyYwb/MTOi9MsNYo7Z6tLObl5xANxX2mY16jA
K/fBd63xPcW6O5fbI5YM7a5dM6nSItq2z0DV1xWfjQh7eJcVgRQhP189jJ94cKdszbxHbTWveUVr
K2hH0MZZ7/YQYgFYR786cj3dEd5DwjCZW0TYGfYBBUqy9K2Q8SwAQvH/65IKhfLKnYbW8bHHomJ+
OoepgP1nQZi0o7pqfoxOcCOAOME2bI6xn3PHO+TTKEw7HtZp6sPgWDq/DWMTQbhj234GBtGa+Xq4
7zVKqP8pBhbA2PIqkQkkRcAccktboBRo0oqIsl2gcclCD+c8/dRnBSc05gRQSx1Iu0if6phyFImV
PkPA5R3LOK+5cxlCw2M+FQsNYvLXw3RQgVeGAjcnLd/c/NLZ39beQDchBnQ7FcbxgeOItctk6Dke
GJaHZ52WgV1GpuBmMaVOJPFgRuS8+7E5fDk1hmqsatfdqXNzKNGtJF99C2s2QC9xlgUfix9bPM6n
MxR88OpAwPdys6u95cwQ2Rp4mgr/XItf6GvF90cOGUhgErDy2QoS/rRTgVmMTmxiOKCp9mco1GU4
5+g+WrmznUUAd68ptIox0LT4aaK744bfmqnlUnFk5+ZAfn3VYTN4CIy8CnkPqCRDqHSEl0mFHsrN
zzhfDwsT7rsLlqqLqZTaQb+VuCYfKXMxcCwANCEJ8y486BH96kSdQkOkGzAq+tVmIdxdtn9xl3FV
wTIUX3H/Als4H0zrxVLG251YqQ985m2Xwrasf9b72cMqfwU3PsBbgmCWeyTAZpYNzUPMJV2WO1Hr
OJcR1X+y3yVHSBMeq752wcW8LEKiYEMjXdDcKT8/tL2brbACsUjBWYKB/kTMwXjpG2VmJ7eLqG47
lQM8mKiM4CKS/QSY/UR0GsrTRuE/xQ6f2Z/CBnlnhTiDbhEj+x2u6u8qVJWTS5F8tC+YmXs8yBS3
0lgbAbgy9G7tqnECno7l91bKJxRHic9cDxUmNk6Awb0VZG5n0yOIdtmzVwYQZtQSSuaMSFJe+An1
MI5UCpRzpb6b1+APrzesFyeFDRweIfzIegCs0YJbAfInzXkPFsCQaBUrZUl4WEe3MMqlP7LMKcD6
pdt/lm0uoukDXE/9FEj3mu+XPzSIcVBoYpAR+T0y05l6C3bPiS1i3wAxhw51I31s0uIS+M1XxCb2
E4RemVpSc5RgJlBzZrkMeoPnK00qQpyy6sRy8ZRTDNj/Bv9C0ex7iHIOklKObAL+fpYNubWQNP5K
UODV/8FV7fFWZQmeTWQz8wF4uRHJO3WwuiF5zbcTbxaIR+OfCrWDYAEeKHL8u4yoaDdTkS3vSjQ5
cgQ+OXlsUXOmf1aeN0J877O4TmvsoThoDDMUJ98R1/LXYEFTexfBkZ8IYUEwlQ6dTrAlOkt5ZsJL
eepFgU+8NqR/4PLFcaIDKBrZpoc9qE3VyMD+5nZfbjFTaZ2WgULARuoDDtf9e0gIYyHutSf4fgoH
1vVHZi0MJQ0WvPEM9IcyYk5CPCFCTX1oKAfJnWgiFYyKcrW/yf7xAUDNdLD5GtkJUwVb3cV1ufKl
iQ32IQCzl95hs5AOmKnrfAo1mouvjWImT4Rqd2A1t7yaAfGUQr8RyUSVhHec268YsIHcnHCgBlKJ
TLsQ6EMkDRPjEQtxCLc0X9n/nd09rnHZtJqHJzHfX4E/cbgpYXXvdGgtW9HuO4sJtSHBHZAXEuT4
JRMi177iUGIVPP22hc11v2YrfQX/OtBV/fDiaAQDoNI++kuUk67IdJKNutoiGPDlHNZ5PN1lGDeA
XN9HvrUIy/7XLLD0UjKOXGwB4BCw0SGAHDr2E32op+VNpeuYDvHurWOpioiS6Na1QT64uex+JJHY
tSrs8baPwCk2g4ryDyZ+kuC03uOClAQqGdik7klCVCWrmrSWl9rL/qfpAMeqdUfcivARs4BSrQ3h
y2SehwaXSFBfDKo8q4xuBWdQRBeZiPCbEExUAukzGuTgYiDTaVd0hHkD24CWK0sFZ+lD/1tOMtfU
/MIGB++BYH8RhBlBwZG6B9FT7VQO+3T0KCasd+y3aPFn+4Yb8SMtmKQnY9PeXqeltlonGjdZC9nZ
6vcjLmBv2NHwdqLoUSsCKXsrVEAnGHVRpn7cWaydFrj0OUfKE3cu3qdoatEjlnmX96ar+3No59ez
I+nG4cIHyxrvSpZ6ZYBGKiPVCJoTlCNWmDFj8DWJxsMy9rHavqbQZtT0vHZC07x19W8NS0HilXxn
lMa9S1ThpTTMDC3kM8pIcWDn//8GurHgR9uCH2l+N7Ok0qZ2iRezqTVm+DLAnXQxPCEX+ukLlOA0
QKFU8zLDutbN/U+mlB0cpu0C5KJDNd0Ol0Dws0aDOgHDObKcP9wk8jQuEUjg4EdPZJVb3C7MjfCa
lDoQCRh0VBAzuQiMEI/OKdnQAytDVzcZt2Owr6rOVAxDFHe0+tYC/y2I2QLnNX1wP19oED3l/AFt
l4Y0jnb5oWju47VJ9Qp3kzYUH0CX5AB/gB0MUrw7O/tfBQcsRS13HG/x2udrFVr3BLNFL1cGCuSJ
neb11cXIwDwiJzzPrEVxNL/QTYPUb8c/B/6ViJ/d9dYFfLAqmrmbm38NmZBLKY6ky4f/MM+lpuYG
8mKgstQm9OCY3Py3CkrVPZdFWtvPN54YmXPjpONqC6SGN12E+mZgLISNVrF8KxWuW8G9LtHLFkor
PJwkoDPf+JGhvSKjPTRCQOw8SMS+6huHF8X5MK6Ih9aywuBKq7o2qVW+109YtxaAj/a/c3BC7QeB
cspQIZlDmDMwQ6qS7ZsxeDcSwp4z1rDXlrVtL9nfzXLeuyeEvwE19YnFSsAI0ZOqIvRRhC7NYEXW
kfj84pSE08arWg7RGZUBFgfZ16wE7n2Zbn1D6NxUK4n6vPs5vBrZX0PAd4hdAM8gHGeoIpFpPlT5
9K1VSfRrVk5M88IBdvpuiTUz5zhRhPCS8tfaW7wp3DD1/ZuaZ+S7neeBYT+wdxRV6XJrTMEoPiFH
WZIeL3BH/75i7f+UPNpPLV8Y2YXYgo03ttIMLr02a2I5pj4YN3zz7y2vlFFvnFY1M7hr9pxtNpS5
yPto78at0ojXprAdPyEB7IDycRv1vqd1DPG08Mw4KRSBBgzXuk66e/bYrFEFIS9YcWO5K6egug1y
pNWIdC9UiaQGG0StrKEMGJ8vIU8PWt/EnsjtJCKUW5cJHVb2Up8qCLeO6I+Nb4X7IB2F+oawrB7D
tZP77f0nJ2Em3BNOwt3kJOoKVEKPDpVtTxVgRoQcWdeIT501DyugNSVgJnk5QcuYxrZnQpfsxarc
Gf2vWtOmrxyssoWdB2kUfwwi1mvZ7keKRkSaamLrVyMmzdw9ubrCSkEbSV3bE2VDqKDWgpMYmAXG
BFu+rJhdgnlZB26V7x1gK1APmEnhdHLoS04izhhs6iZM6hOJiVehKVW4AI1zuivYNXnYvZwAyJBA
ODmNTSwsfpz4QM3j8wy74tRCRFnnxKvwjKr1Mq20P3RApGWLE1eTx8UlXUmv8PvFsc92YViWnL2X
6hZpEazPhhi2qO6tfnVlQq9oHhkX+FSpH6Msq2ydTHCALhr2DUFVjCMoJft5I+nBs98cKAdg56zG
ITX0tIB3gOrJWui6J6P331WpGkACcJmAGwvfIyOxgi+RxX+dzEZ2ZJ9gn2EmJxDBFg/d9amDTUy3
/lFlJouGthvpTZN/YY2kDL0WnCrWbjojIKyG2FgppZShz6BR0+/20h/Od+QG4n9e/DhR8k2onLkf
I2c44+U3j/Vr6F/BPW2hj3pwMV41p0SI4UITOVEZ8tLUoADX1oL6XJDs+MnmctxSN6n0VJ78NhVf
kgCzOnf52YO2eBKM/hLc1Tf7lCe02SqQEG7RIzoNE7e8w2vHJ80/IjtcwTEfXMGnjrjpVz4+Dxew
i3oy5OmSxCZcIEKfrNTguHAFpb6B7r1RLCZ3my9OvdUh/hYKQc9CphtzGrLL6bwalWwXNA97HHlg
Qt2EY80144iIF0wU1gfBx6wuiuuNXIpeeugODbZiGdWErKvakxKMONLYbe/6uooT5Opv8HV/CK8+
cQ3J/SatKwti9mkrBOcYxlQJPDdvd4/KZMxdpPZbgNRmSj/cntE8MbocBcbeA0tntVH7qO+o2fC0
rnZg3vgrAeUr6m7KRttm8bEA4qj72WBq/vtAiFt+HrJu+V8oMTEmatlecAv9mWb7y/ZBOZ1o9BWj
ig/RB/u1uhPLfGYT2HrjluqIt/bndX1y3zpzJNUKGDMCmQ0XIL73v91V/sltA+0mldfz9eFY4Nmu
nqoGrv51d5CkpKlKSrNbmzCWVTLODoIcUJTlorurmd6R+oBy5FaXUUOJZmZGOacJwfzO/in1QZgv
YD6KbRT84KSt05nDtdD4e8w+DsARt30r0CEtQ8eIgVS8WV/XNpL1kPy18Ufzfmu9s1doRZ7J+WGL
6X+At4jnuof7Mm5seB9OjmHI615ttr9URaMoHkUZ6GhZBEE6wuRety29wv56ccbQKo1QVAeZzI4Y
VVde9GKcC/cuAosxMHMrxh8wXyQ/TWdibdEyDWuHsm0gdNVd2vL0RggqB+T2xQVpgXCyha1jBmhm
Rqzi7TsE44s9x6hb3xLUd9OX6RHwPabxPLqEcAqjYMJJTOP7Env+nDonaH2L335zb8WvTBBkhsu/
vC/uogxnjh+5Bby8XAZ2nSSp7CQF5G+kHBA/F5W7oPKd++xYDm1aDPTr6JGtEnbPFnfXPCMR55UR
XN++zNOkPYh39p/QVAJwrGk4KXccpLPAvJIjui6AgvLUGH2RvrwWBCrujFVgnCiHOj4mqmcd6+3B
W2AfHVQ8SwzMkpTG6bgympWsy3Ah/G1YsxTmpDR7nfV8oNkYg6xnYn1TvFbNhRurCOhPjWfeuDDr
XqzVqC6JTUStZ4jaR1E1LFYY5j5HymQmhlpl+BuzVnJDReFPrZl+upfYSqD/SADW+Y1V7B3swiFa
ytlLGDe7PWTmV7Vi56C9drNdFG+Sjlf6AXn/1LTUki4ng0/2B9Zi9NvHBHxNVOpEQs1IXRzr9aJI
2utXOh6ypQDfxk5Bklhw/1Dbq750OBKLQ4tcifOM+pspdAyeZnrDstCgnkNUSk/C357/Z+68ADOH
1CQpOP8rKZnGAeidRYyIP2jkCBrR3M8z2pyRUrQ+sbAvt0OW54RufAG50RgUjW3kNfdtbKz+lyao
tzJ4YjOUrWYZ14kfnqXZKyJMr66Ef+TSkW6VKfK14ebbxZJB9clqaR04/1sDTlgTVxdR1iYFctB8
/eZXMfDEVbOgX+ElGiGL3j9degVQGiy3AkbSytF2UixUlUz3EhpLz6h9uTBfrrx4DDmA2Rc4VFDD
vBZWNt9l4upMhdvr4cILNjYyAGUceuR67TDxOootGBeNnErYI8VzbNk43Cdo+s20hhqgDiVyBlah
m+pqPtRixdOqPgmQZAXPCLKPNvqzHcRkljE1/1ZfPqtHUvIGRCKxsNEUGA7F23cIw4mCWRjfOEBY
IeLAMYRMWIJyuu2AUQnF8uYXZsGtRiT7uGod5VIE1OFMFeMHrl/qzN7zyZttzfDdIZjiRGNpyldP
kXB+nagAkgULCPiAjfbJNsUMtFfplkgVDqrPnxkWS/MhEQsmRkOqJbP0GRhfgi7VUsnrNstwAtLt
bbSR5IcZrLIrrYANY1NS7J/h/xB+xEPSTgRb6U3hEv/8N5OevViFjxmcJD7ubxDX/GB8EYtNrrHd
XC7ywb6cpPjM3s0sS8u6P7/LRuUlVUT7WffV3mYpabFeSia+RvBngy/tJLYzDxe1xe2I+gvbpf59
lZ1j54BeffWPHjy1NZUvXZTpQjCNBvCcZ/fOi2HEAJeeYx/xcMTwGFRzuosMF5fjBlOjKjNFo6Th
FHH1X9KmbwD235gRsKqr2/eeGzCJ52vxhYMW2k5ucAhHY5EdvvyiD3DkfX54cRGfFNkr/Ai7mJbk
3fd0oKmxzOnlfLZzMCr6QAsLEkmME2kuQuYaaGsS2bheeN3nXWgeC2P8jybUy9oXxDhddB8rKPvD
/hS02Tus8YtVAZhseBR53+HsJvbRdgHEX2LYjct064ltHWHDvn5VOVx7iznTT2Q5y0R7zFzEhVcG
Y9xK9kQMnQhN0vu50hQ1Pz3ufPvJuTfR3RNwvA4nAnqCOXqxEMU9UFcumm6jQErxZpKBv4MkhqVL
UEOOwK5dxs/s2bPdClQo3HAdUqcQvmfbBO9e0d9AB2/O8VN9SAt0ucx1JTCpaYYx7A+MAf/MyGcA
6rnnkxoqlzofm0cX7RL1j9+6MTspYkuDXoOejoJRHLY0ImDuAFPmjjgsB09R0Kg12lTauYjC2HGi
Leb3wsZUd3v2dmwxbq53nf+03bwgmRmCIWCgeHeqb6BLO0VQO3/fNECuWDP78vxpcF7077lldikd
IBS0U7tOIZuFJZ2cgygWGmM2dsvi6T813IzTzhvCd+HEeSC+48xf1w4esS8EKlMDL4bceQ2oXaRP
8J24wmaeet7uy23InMdFZv5CYy4zmwcG7HnOzoLaXGF2ewNJPAbsZjnZFt6tp6MREibxwOVt7Kil
rB2dS9jldZUch5SjS5CzF8nLzcLdabhR8q7OJnCKIx4F6zPefhLoSWTZpxVYNeQoKn6JRTxpYd7y
C8fySJ9ohrSOAfZXcDSDBrXEa1O98cC1suGsWZuvfYoAp6EV70WjUimwu0N7aR50ZkvRfI2gIl4Y
8VUNFyfJCtXuzNQTutTYliN3S+f6xuTBPyXhND0pIAV0hNcKpaKOh0T/VMPXV/bC61ZCXN7QGUxZ
ZwzwsBx0rmQdnfCDY7/sfSCaRjMde5wDj2k1exKPRME6AMmz2Wv22QTDr4OYYN1dQGQxb3ZcqxRk
cd3sP5h4JgkIKIUE+LYcOuSlIralaTMfdsK0aDn2kE4L480AqxzQ6v7RxM4sb6vwUOWZdvuzvdE0
uky9ZwrS/7XTYNZB2iM6gqCKPG1a9MQ7LDGyZTdvsllvp3ryWTBPbvIRBOtHISDz0gVN0NtPbvOn
JdOmQ5h5qE9VmP7BK9pobF6NbOLw6OI3j1oCCyHvpNzVHWH063EjOUVnTs+0D40C+R7rZvfjiZG7
ljDar4xO5uARNtgz973e94TSZJag30xEyVpHpkj4IjdhxnnEC147l5F6GRWmlyaOf8mM92yPP6c/
49v2JGkApOM9WaW8K1Mx2QAyk5QeYVtzKqJTaNN2BG4Ek7o2wmwagyPtP/lNERLvJxYPJNZ1f/lG
dFXOG2pbpQZw3Zv8hHwJ9JFhDe2UOZjC60nwVQHGaUt2CJIxY8V1Vl5OgqA0moouOy7JvVia0aSA
LDs1hEjS1YFd53S2x/AiZXQ3ZSHm/sIZE80xHRI6NZXYruKfyTclozwYyEAJ/AwbMMBNXpzRqerR
2UyvNCB2zaWAPAv/kC4mKqKd7fQ1Fvvz6N64wGyvONvAdTvnXhaoXuLUWaMItV1/eyoClzCcyMxL
xu05ZuNPBYvs+IUZScxZz/kPFM4RQJfyS76oBImlEN4gvpOoPvsmtrLIirB8Qo6Nr02NSx+j9zy8
ODKDa3TRuddozBJAwtXLZkisvxCniGIrRi3cD79x43LUKtKndb/tdOTTnIfsv1iNggjYsGI3mTDN
nJWFdqRheFty7eYkd8gFnKZ2lNiMwoRzettcl0FgrViqBWK4vmAaoKu1kaa9l8dqV90kayH/FD8J
r9puStT7X36FD19IfqmWD4JOiSe6BhMcGUyyrEqovCBIIQmKr2Mzh/+HaDQ8Tgv9kBktnDxFSflx
wnhflmY9Ujhwb1i7TLiNiBR/llFA2RVHXun+gDDqsk4EOBW3+H/u19cjdLon02i9l05+vhjoMhsH
P4NhKe+C0+IWU0x9k7Il+wjV8KPiGeUJh9DJB80IsqPmzjCY83J/TPvUHO7srekGZmvi9uYfRg2v
hDGIgx6tVQIiU5Eg5RFW5Zhx3kjEEDmp5VpZ1ZMIbuxNarl7jAJkHlG55htyqxkTIajRr+1QFBl1
K28rXdiLl1WKPwOs5SC5vTL05175CMJpDBaMcanKgxBKB0XlMkXOlPdRNZUbqnJj35wy1f+JKGsi
XTPhqG6KWzXb0rABeO3P7K//az+Nn5g1fDQFA2wDNtklaVvekXK282ZH5deP+q4cC7RMl9HMLgJH
LS0v3bWnd4qqKPKoUX+izUkX8mjqWIx8PFR7HZGWpuVPayebs769l64mox3WoGRDbxdCz5zdb75U
j6ByYnvRY3PXbm3JorhqJZ6pC93bd9w7oh3YqhBXyH8Nqf6SnNpSeAivg5rFdPq+k8sngzYh2JN9
Se53n6XqIn7FkMEr+WWv42JabsbfXtPcGjLroGR0eabfzvPmA9dtAFlb6pkdGGXl3P/BZwcGYj6f
e1GAdPu8qfWoVG/lXAwc9iYx1dMVKaGXvqHww6uufGDjTTgXToBcWHx0eY1WDX9Zf+NxJbaSI5L2
Qr6fkJ4bIx26Q/Vqjlue61rWBdoA8C2KJcS0Ond6Gs0asHwRyPJVvoHWPBKp6lha0khLci8zjLTH
2tLHMzPPen6QYpsC8kBk5fgC9DxVuHJKzjIoQyMv0X/NQDAPmvZjXd1TNdt44D2EOlFedcXkGNMB
wAVcFsDKaK7AVW3JULR9aYqWTOLeuqM75yMSqzuNNGHkzO3R2Pc+QNN5heiHJVk17YRBK7IBPtI2
H+RL9AyhcHMmCcdMuCRQ2gSC2J5IrsJRJVcEWkgOICf05vgMwWrr4vk1vCGlMq+FJAUxC1t+KREE
XIt3eA6F99EjNJB6E+aOMhiJZeOMWVZKbV2lMgl+fZ4lRmLwpbvxm7cE0MQdLJXvgT+GWj9JJdhg
TP31UTa1IDpkf8g2BcAWEteqfvm38etc4cQ5OHLiGDNmbIseZHKq4BQ4zEhI1+XlYd8jE9GjhyBc
L/wI0IsyRRt8hSkaAXPQwzRb6UaMywraOanNhn5A/joKRylhtTaY2wy+ucGsRhnV0CoVf0D7THSd
zRqjaJin3ZRQtKqRctVtyfHYxrJ1143tnDyafsgwWE5ndTTrEAtBEYYKPSUNHiNJvYw/hE4T9dYM
L9+Y4FW12CzFs9uvMGprQgxWTT2P0o9hJO+18fezXZ4Jq7eIOTE874+Isx/aTET+C3KnVSttuYfc
4dBd+mIqTbCh9QUXhOoB72lPVtkQJj0G2TkZi3zBjCD1NhBVsVp+v0jx+/gMWtqp2+P59bhPU7Ln
khH9W+KcyHLJOaFwSBaMUJ22g+73ZMsATXOTtsjbiH/CHevXVH2m47Z6crvk9h3gLFsH5kQCcD1x
8ZEqqeNMIZaM7dSgsmkP2jS76344HYLm+k0S1ly58tHzpmiVjRx0zJXBgNe/yzzd5OmWcJtfvWBP
PnlZ5ai3dtX67OjQ/RXJFDPD9PZmsLbI5Vz2Aw4ODzb2Y7EUOmJtpwPRSMKLOczQ7k/99t+vBOvC
Xl+xsERPdOdsKjL6nnGGiQ75acoRQCpobxuYUVzIfgZF6H02j1L1e6eeU9buQ/i2HhUGkZ09HdLm
hCgr9L9nvbYH7rvmw6ekjRZA8M8NSa0YCOW+AopKJ+d/BBPG5DyAznHStvb/f0Q2gQi4oV5AwAkD
ZCoH0xMdvQctW80jm4MoglIQGH2ZaGIXSR3R1qG0HHzgPrGjIJjLQdg2kF+/sl8DiBc9jIY4KCFI
o1XJJKTEitIZtN/2YM8jR/RaI4xtX1LF4plT2kAIoN8SrKO6Yh+FbWnEv609l9HJ42Vpz/jqQ1Mp
RUTDbfhHrMCXoejlAiokc/Ysic6sSLiEPAUkOFNPMtPs2nd44V1kKs6sSClBYMbieOndAnnIwyXO
B71Ga3cIERl4KvnLTBYB0QC90waLFh1Rn2yPyGPtu7D8zZMu410JaIChjEyj8wpWz1vp9BwQk7fK
ctzj8HZ8LuOQkc6G0CcIWii/6Vvi4B50zEyhOcDmLAjVxf+GAfQrL+BVdJ024DGeaWlkRAaEJE6D
XtQq/F3dKYUXfdS1Bv7mVI6FjTbwdurkGhHcoaaG34jfNwpU885mB5wXIxcEGsWwxUQu01DMO0B5
5ZqdO6nKza8Lq2TOOIj8G81LkrY1ZRkS8zJ3vLWJvK9BL86Bl04MRac3fe3/zXiFKXbL15RDVlkG
PJePoL80Yj4dRUhXF+FmCjp1bL1k2S2dIXQaXcB0smsocB1nmISKHW/MJa521Bw3YP/2NjyeCgir
ItMJXR6cbOYVTBBZo/pfdZW/gP1nsH49QTCp/If0exXk53/0bzqwGumMe/Tvp4WcV6szzp8b2DzF
EoZhGeLPm/zsZrrFgjdsHF6ySRFSXlCQq7keXcET0ETnIkIRT8RyYitWLRGLUoi3Vwq6wAb8aZZn
loa4wzC8c+xbuv7TKreMKDVl9TubfwXRyLGVS5qNSoG37V4IlD17ksMnK2GliQB9qQeFUH+06VJ1
AAxZkdDrcQlHcJdT2vriUhS2evNRM9Xt6HkpBLCVpGcyKUGPUv8FRqc9VfZvmjbGPQmFenLmqTz2
a1tl8YzRPw8oHrhzMERw8KkDu3FF2zaGxgoG9XsIKzkmdYR9/Hhs8wJfneizJ2rDReBps+5fj8F+
zDP0u5FXebuw/KG00Qy6mX+eHo7HSqteVNFzXwwnoj54fOjndxqn3JYXHXlwJ0xwlDIAW5uloyxe
Jh0JTGiu67UEYRh2Fw4Hcos0Cj+p12bZ4lGf8yazesKjthLq9yYYz+tDP4Fdf2J5TsHbTTOuMpjr
m5W7dKlTLHthSHbQjMAXk0dvnoxkPs/TtCdHLctfeUmTJ8efVwwjyV+4t1MpIedU3I/jM46mEZrs
ZvYBvwV8X/Cp1g/10p/uCFZ1nSHJQQgEHAHDn/DDeRhaw962hkb+d1vw0CsrLgaFJ+KTLpuXr3xL
zxNk5NqLNEg2IyRndHIjWIxRr5gO2rr4/9a+KCgAFEEsHVY+UWohKYPxpRikd3RhHwKvM+k4W+6j
HNFA9x5e79qUY1LoOs0q099LIyMCX/Yy4xyeNvTOCQ1uuHVi6BiT73JStIt5XU+8R+wmD9rExWfh
P8c81/agQICN307f5vDNurDTOpSV1nrS9svZnpRfYo+dCXuk2eczfW2YZ3XTqBfl5Xyuq9xuTNC7
ndZcjus4BEqGua5QRft+enAxwqSO0IxnCrG/XztAKMhWds4/63WZWEE7LbgQ821MLpKLAvskCvN/
iPAuZQZhBoLwBXmI1sZmaF48yibp/lLnPVixU7EtgJdEa8hvqs16oUFtztKuscXgkFNtaHeZz7VE
uFPaaZvD0cipgGvW8aiYZHvbFvwIGkn7YjTUeIrjNAb5u2mIwUnktYj1MyNCUCxCtCmlHZbFn/Yq
6v1v9ZTeJj0O0ro6OsEdk0PnLQUnol2apN12a9Ukz4csTj/gc6Bs+n2oE80bZBgwlRNxILN1Yegu
i+hdHRhailVgRcgf7ov8esKCxAYnrPQgFZWBEG6zNb9GuA4wMqgRV9MuvSfV2VQeFeBk19Px1bFB
mW2exCsB0NhbEJYdifaXTaE0ioDeFf41o8JicYi/X3RJcNsndnWrC7c9kwXF6zb2mk67sN+dwl8o
UQkvWDXaSY/+tIop9+l4su++KIWSdGRXz/+Di4nLNk7dPXLv5q26Rx0+rAk6S29lFpaCO+OCNljv
xRfnF6gDwKvz849ikK/fPCW/jzXGLB2H/JPOXCG2P+hhdXEgHixotKAk8jxassA7j7rmRTMe3Y6P
WJ2UoauxHflCksD7q4cAdRepl94c95FojtopDwSaQQ8Xu1T4K/aWYsm7i00IND0PRgMokOhiup0Y
bylVc1OkV0W14S0Tq6+M4arMoNNO7kdeWUM8JOBgn91ljlWcj51np2CJrLmrZwOlIhJHJokfaF+X
c81PWUM5UyxOq20OrJNf8tRx9hvCEmHIUmR5DT7DNG/JRBQ3+UmTtWgXmlYI82imca9Kr4FlTwcm
faMohwp43ZhNCTPtQuLdEU8o1ADsr4uFFkmX40vbZrhhojInSYGsAo+ZYddBHy4djlA+3IBRXuSi
bRmBPWb/8xz8weZH/ITZZYL3s58I2fQ4UYsF6OC4+y/PfSoC0KYVcpWGsKg87w+9fMAVri5psUBj
KpRqZLvTeT+945+LidVLdLA0jrsPnPUyNeD6R+CimkDQo2khE6hFibSLS5Ljfot9jo/+TcTnxErA
PnDbD/Hn2MIwkF5kWQtDoPq0fe5dtYk8No4SQ+NpFIxA4F6dAmYWFMU7kmbyZFmw5Tk+kWHv6ZJN
/gyupkqUKWEESfIJaHBDUQpT0b0REPTeFbUeFmjbq5vmi8T2rZCTT80t/6XlGxrsqSjYCdwhIbGl
Si+GRVY9HOvgPvXC6d0RW7Ql/yfRc2oAZFsOwR7lZIkIAHY/e9mmFTzl5IfPiKZTdOPw6xLqp0Uq
anD+zEVPjS3BZ2UpY5kOMCftAWWN71M+v6aYqLuXnYm3E6ue9pFSlzY9CRe50Y5J7+GNGOSA+8xZ
58umdHO4zzlNWy+uapl7Om6hN9x0h16hkC6UtD6aITeVpfrToAOlMCL9brjRNyvdbC0vxtf4zL3+
9686mHDU9cDP/pOJaSsnEmeGTTFbHlcNYU3mFe40agzYR2A/lVHe2sWNeko/UEx5z/Cf6CHuzpYd
LCBpLwe00mkS+T/6dnPUYRJuZ50ashWHh61AE77LMKNR2wjexcIMfouUCEfp9eBWvaRrrtu/2F+s
JmOuSd1rh8hzbdPqkC3/pkC0pe4oOyTgh+E+aqSLzGsebqwcp9HAt/xgyIQzJsLlaSHaV/dq1gpw
zwo373UUsnF2m1NMK/3fyTzfq0TiWOS+bJXozoeanXaWq9OSOCjExhN8PhWF0jlvZQZg97kD7Joj
hA6WVJJKE66cf5aQLOCOQpAnUfITV/JI07NpNHDVJqUOJ0VNa1CQv0z3+kwZaLLMR3hbvmasLURY
uQ96zVFVQDjwtCbHBDYTupgV6imPoJGCi6cyzWT8utLgK0XB5IDvKY//OrbDPuXIHJT29NMOe/2b
f48cxYqlsQUpAAnrrv3SItA4QsdZ0QiyT65DWrhtwplizIudCmWsW8l9Owp90f42UXa+vxhje4Dv
xewNjD21icoC3Y9ey1e5aE+Ne2rfS599AiT0yxDxJOMfza9MLIYW/a6Af38oXQg4xKRW5g904Ob/
oLee2wfOnmyGX6WzT5CJNVrDgnWyvgcQGOx3NOEWzp8MdvTzggXiRUSyBMCr7R2cJ74dDMJghq/N
/VF8NgpA5JvMy9UJq7fhVUUs4TizoEO7sTTN1/blE44wIHgthPzGGD83K4dALpzzVCKhALiQ18tb
4d4EeF0NNCLaiMyBj97r8yGCiQhUBW3hDdwDQ0rwg2aONHnPzOd5sAhFCEIhoVIXNC0zVKyLb7uu
kE9YIjbZ+zjPAvH0Tqzx6O2GedlWLFXZwvNuMR+peSV+W1dyr5pcv7tFTb/HmRoNTFYLKw8Xb2R+
VibS34KBUVkY0kI1mVn+IzqFBEnDfI2GBFUru+r4fDzK6XMn7TWSq+nHKYGUH/zT/UUx8sZvMyHv
Npjl9xtnSUHKkurkR+82IAfaxgmbn3fgS9Gibb8fN6hZr1Xt78psLjTdLkfhmhc/LUaerJSKDGGZ
C5+ms2xp4aotks/X4M9aTABjLgPG3Xkl6CdWeRIWNw/00/6zOzDfM2iqTGC4Ni6XEpWilW6W4O48
YR+JVPI3nlyWpV5m5+dqPtqsADm5HFjUdh8nWk/k5DF6/Li55RlmgviZN/mv1KpOo1tYvkwy1655
jMfd66G4S4ph+g9lu9Mq+igOgS77M9mU2QumF340y0M5YzKXsSmY4mFjIe+ImjVEzqzrIGPIJLtr
G/Wz2xyXon78gIHfMXI67iOcZmwLUpFGzboCDV6n/DTMzSdh3iiAMCZh57iQ5lNAKYzTYUsZBkNi
btL8lpmSXv6oBP4ucTZN1BLxzrSLHnOl8TkzkltVDve8rSoTU2zSXWba5ULdfGY/ISV+MIdCIIUJ
AYoWKqN8VkwSz+MdicUFowE53+seRKMNGV0Os0PeyxPydOP3MSZ8oyMkBa/WyWzdsb8E8lyoXjMe
3CfwXnN4QI/TcdsUtNQbADIUJyf3OOUn9/hRG8CF6bzdHJnHJIlOhLvESKIIy9R7I3658oo6+Wwp
DGn70GYck8OZl+hh94mgOssMaHFBbRB/grAaIsDSaLX1o/79oy0ORsrbcAQhWPhBB/Rg68zTnkW9
iL/gF31Upbcj+rbG/lWcPGae6RvkZozdQsov3IsOUu5K8FqWN/qmUAo/h0P2fxs2b3ejRfGnUrnI
AiDT8LpTeQ9QpQcs4Ic2QbcxceJ1K9WK/iS4VMtMTTJFb+W+RjzU/l93MEVjNmRU2ApoXi5ISDdt
m7cUcNR5VY5uvmwMfsmx/Pc/qiywRl7peO3oK7SVeFBhvXWxpGdl/bOcvu7cTDVhgs6R4KqiP+qK
NUTHjIW/qFnFUUPTLwACSyHjQ/28wyQn5r58gX1z41zcdO4F8KYDCe3Gk35Rq30x90cQbgitZ4wv
pX4MkX04FfMCRx8ilu/JWFIVyIYFg7trDl3Vc3vDxp22CI/P9YT2o9aUhlHGGZNlwsNjfikskzEr
JfMO8xYMZ4A7cvMAibI/5aMVqvdH0Bp7+K6VQRVyQ9ld1PHloIMkTdSY1X3yRBc6A++m/4tr1Wdq
sBNiOju7mNAU0+zB8DPGzKURpxIwiw0pk5iKJOJ4d85NcxBccjT3venRWv26xt/VmVady+0sYh9M
6XyAtKKyKGeShYZ/AojgT0j7aCOr0Xb/0iHOFG/wSc9ORMJeqkRn7YkN5EcXt5ZJLPh/5/vD7zqR
j1pUOfIY4k6E4f2yJaMmNlk1VLOjeDaps98nGoLVvfTMsxb153QeTq7aw7EkRIyAZEhUjYEh5bFq
M6XRiCQzaFoEe/fiv48DhwsDlJ/KjMh1AQzv85tFPCM8dR1sVx5bH9zt6JEV+KTkNWIK7RAiWXhG
zGn6/VZxsgIeA3AALHT1QgxzZqb71uBLUH+dU+451v0+ottEOitn/Szb7cfbuHejavOcBRQR+vzH
7LsdeLdyAN88OJXOp9vEgpvqNU6nd0lzbILZm+YU4IXbnOHvHUp4+kC3vCH+sdH5GLjEj3Ucf1+m
1bM9iNYL2keIXhPPPLqv3tvMq2Td876AHeUgovXe3EY0KHD4blVSZmRqDAiYx3Rn5kyo4TbzdU2e
UilZmABxIqd1kP/B5mH2qXDxIVJzyx7Va88O5kuXDj53TGtUEut//f1XNMoWAdQ8iCbCY5Dx2OGb
Z7k8PT8eTZSvXjFuowIE6nUALaNG43J5ClT6kIJL2yw/abNblUfX7+O5UbAsbn6Oomgz9NbFQLNt
7BU9gAHZdC2vP85+OzMhbqI+smBi2mkvl+cSWMvabi+X85xhnuWf7ld2qH9uB+4bluxh7kf3r+uV
XuNlHOBDUmpLioMkXpqZxpIvlObdqiTvkfaY8ryubTo2aq55h+5apr/wZ8waIggP4Dn4YyK3Ectl
ScEInH7rcMXX5FMb0mH9qRQGHnh/hMyd8p3rKSjUW4Do1JJf8C5llGyR6zrSj2Mx/YMBib4CCJdk
pStUF118W2u+3mJGGSM9L+dh0ViT56HRTl813zQ3kxUKxprYEeES2EBcek0TlzQtAoQfXrQ9Jxyn
8S3cuksfk8baODRoFf31INSw1P3VR1ROe26M4tqP2OYube1FanWP8I0EzJsTWZ7aqkQw/xrUWTKB
zXod5q43NM+YnGnoLzTa8zfheQMgO5Tm2aSaiF9D0KfRzgsB4MSTIYNIJMF7jSeyvHnU0KOlPaPx
taH5ulhp4nGqNnC092jgNYOvUp2BcGg3b+M6HU/+6MAuiyqOYnaUVtMieWf1Boet4Hnnlz+Hu9s+
9EmAYYMjHPaqcXfpPCJPqd658Mhry/sC+ofB2D60YlwWbrE0bGjuF16jCBo3HfGVTLzYAVutTCz2
qonzAaYhHbdkmJ2fKFP8RE+zqsfFibl8wlCTktFNRSCOqjmspZ3jxqNBKDwd6MQlfPRDSmtUVuUy
UuUF0FRRHtMoVPRciI/qJtOWkcXHv1asWFS5BBGtjXlkNGcEqxKVPosXy3LBiuJgEn8oiqktkCsO
oNv1LyiBAS9T7mLG3nr/hFgEmx3gSh6bczLCUgQiy32vBDJsuD6IwAwgsBVFnXa2Amj1J9rfeF8x
kwBCx3Ma9JuyvOC2+IuH7XnsWooNIFulUixrLiZ3APc/8ci85jG6e8N/6qch3SLU3gQ2kLmZt+/v
6l3VlORqC56rX+zaWgurMk8aDTsbKj+i/JAZB3Hq2oYOwxIcwl7/BCDICA98XvNyBNqQ2vUiLZKQ
jESIJiiTU3OF7w57S0sXLZXQNHbeOrFOIIyj2LcmuqopduSWneVxnGcMVxpR0RYVsdjq/wN0csb4
5qeQzS6F6/genXwTfPJmrhvqM+zYHm9mH0LLs+AV1DWt/XMSxV3rQzAURsUPQJjUFHdhNPiNbEpW
7PvHDIbMhMwAcw0SXx6Lr9CFihitPRWunriszcw/3wHaXKK9OJOsaBRgaga7iZRG2CKL05bUuH2Q
qNwk3JAwixajbYKMnD0kmhQEY6OW9RMNz950UQIQOKoBkjxhvI0ZvF7GLHZfgyobFCqCuHLps9tD
PlUndouvswK3FwO3yhq722h7FgeCkbJwGgby6F/BPlYXrogtB4iKtL2YfNsmmUvwlkiDlxHV13mA
fRxRNdbflN8cZqZY580T+eLPg4zYCK9/G/gq6RXQOTO4z9zyrATXxAiyelbOHBq84gXz9WeeR9n4
oGk3NVjTz1h+Zs44DeFjFdE8FfjtXTmNSph4BWOXfZtkS9tzq9BfXD85NI29ZGk9VKLP2hWF0ABx
FbyMFppq1uQ3DtewhBi7hf3EphfVC+tR/8jxP3yVFVidgEH7C/g6mJF+hnMqjzIDOecqjZkSC3Kb
P36pgQUlnQS9TUBGR/em9xJzga8ilCTCSCPO40kbEO6LMvKnv1065w4WwCXu0rWFnnJL5K36zdTY
OtlkfgeldTtRYsDDlRCJGA6o0fO5efg7Hxzh8r/jq75gZC4CYE7V8riP1QwcEWdFoTziWZXg4mR1
TA34/I7HPNi+/ON/P5sNhlJZ7vYmiiTI6o5vu4GMOl0W7DGhUpCdV4wn7USov0nb5oGRx4ZfeKH9
zpLHpiNuSADlDTyFIwWDb7mEOvDXRhBljO/L3/IfOx6MJze+3G4ticNEq06qL/Z6Lpso69AkJlZF
9LZT61J6+9x2Xem+ybhxmJlryz6j0SYW5p1j0whlLwW8Ri/X2Xjpd2ZVnLzHZHaSarzl1VUX9gsB
7QIPKz+UQp/3g7Z6WkFJlx92NEeBC7pej7RUE40ZckWn6R0n0LNn9tu3MjbbLUf0Vf4nSOZ5kehW
N/YUVPltCNNrIilUqU2a68nG/lSYLawjX/W39Zis3d9eaPFHJgUdHNgGk0hV30kJkH8TzU7GTOoT
cXkyT0/UoCQPX1Vmst79Q18K0TqKkLCL79fhk+8c9WwM4S6S3cGpdqMFx1emWk2o9yBesyC7Tj5l
msU2Xu2lJ5m2YhidVEMnw99e1ZJWTQUGRv8UTgNvDjJBZMNZJp6vjVjywyvtHvP6D2ZO6svfF04I
Kg9gn0DtVGkPDWriflhaO8arJleF+4K37EieWXBzUEWFR4MkCD1a+CGRRJkiU8D17qWZeA0u/M9J
wVfDWPEcAUhg9zN97ukns98XXWmc5FjjIGAIoW+vhEpuSK+TglvMZKUxuezsIU06a4JUEWwihryW
GnyCoVDe8jKJYrNYsIR7Zwb7SRIRBmzFvMrl0UJMZKc8nqLhpA81fakg8OD2k04Nu+ZcVUAyio+x
rAj7HwSHkjB1hDgTvXAp+I6ZbDX/Tswq7BQvvvSCaogifkjJlPnq/M1GR83vHTWejHHD38WiM4L8
P8hs9ixuT1HdtS/7Gje6Q3OLoLymXUVC8kanoJ5pqn3KbgRXCi8UXa2U7mRISKgNEWlWby2MrfNu
Kv7K9RXkopsl9LA+yDwwOYZ+7Ziml1iWbOZI5ZFlNltJQxzs1D8Xma2u4YoDtM+x+s64zj60LyBh
Zz4e/0AkGZycsFZs4cP3ecgvPvzE8ikoDGKmzx/k4gohVvxQrr0bs4mwfaWwmenqw5jfanZozcLe
yetUFy6/LqZEEqBn8J+IPNRjcAomh90SSrBUV8nJKepNw1aSA0fTQP2gcxQD85FRWdPUg+avU79B
k6ejxTkKiJT80sPQ8ER3G418XonaucCHVOoUJAALVp1kXIib6Kwa1W0Wyk2MNvc5UbAPG0hi6Dmr
4gRI+itlW1YGBOeveBxXlnwt7BPSZuShnasM2jWnUpjgUGk3P6kxfQjNkn25Wuaeh0wtxCjQ8o6Y
6TFIx87+JC+F0jnY4Tp7/yehsXat9QQ3NUHufXJY02Dz7flxVBIB6G/+fk7ni+qiS2d1RhvjMMOw
VJDKo5nNROEpcpk3eMXXwcbwnv2rbuB6DiRIIZXBXdETxdG/DzshFpchXS6oF/dk3WJt1c3sfbNA
NCO2BnUh/ut1vQX/VvP+g2O6Op7s3Ty/oyNnjXoZvAndXhfHzVrrxkxK95Gpu4zPfRQ+BI13scoP
NfnXiQxWViobVVCjt4FK7okmEz6cBI+FwI3Pqe5WxMIXzAeSvHwzW9LiM939o4jXUFFZmudEecwg
P2TmP73hCjqEr1wCiJ23Xtl5aZ1+RJvDqL8Dd2NIiv6sSXS6EuxRyXCi4JR2+mgBlzKZ9jrEnw68
JXXKCLJCPfFUP/BxpRrhsI/+poJxh6XNg2coZj5HYTxq/z8Hom9iyHvQB5/2LJn6fIIrEo74gGN9
SPZI8dcqyMWt34pRHJ5ZMijx/sHO4JCEp/zcfyP5nFqOtaZUO3nKIKsoPiJMIwW4EBZqIq3S/AoD
oMCp6HB2ri3LqI/vWw75VbvE+EZAcyBd6OgcmuXtG6PyQl15Ot8LyUBJskSSiVw0hMzYKD04H7sS
i1quAUkiPSOZUxuv43plHDK5DMY4dQYWSmb4kSDvp25rqCRY3jb5dBWL2rqL7Y9ep3zRrv+7qRg3
lwPedjYVeA2G9ERZtmQt+WgJxTa+7EsUBAtexY6Wkr6nKfZvfsAG+3wwU5eJxrD/ggzC7wqjpDLS
hpjabTt+in2FydMqBagrOkfO5JtyqeObTKDC7cAFXQCE2CLoHeEkffb0lSxrRQxtazkdwl6j6etd
VY+xRgNsYyurPhonOMPgKd9GDRGzSFjbUObTAYHnxojc6wQsa5nc6rUYzXZSOCkyeXbmU4sGlgGN
JTBdk80XkdULKLn9JxdkOvfK5q3ux63UE9rMJa/Tnpt2ku89rFYyHelN7YFokFpwzScSyQylBg/e
8nzYhJP62CU0ARkjNSADHRTdA/jarhLE9Gntf9LFpcooUj7plqmeYkP+FxC4ZW0trMrxl561ee6C
OnJBmVX3xBiik7aNWJl2VCdpsSWCf+S+URL5Ia7agNp/IpK9l7HpBYpch9FTIrUQc1HJa3bhu8CW
EJHvSVdvqPr9lbrbPK3PO5Jld4nzfTWMlr5AEYUbZTWB1B2+5vNyOL+LVi8xe/OwOSiTgJHphaQ1
AsfJUtxzlKecm10zeLA0Q0UVdBuh9zh23/oHra7XT968F58LG0mPbt7HsJx70UIMaCeAKOU/EVSB
Yo3rWmWn7ND1P/5nDaj5TwvZDTLL4cl1/OHY/DtkZ3ZoaRFlsOdJDELtELNeolmnCfaLl4XVnehL
Y2dz4A2I3SK3YhjL4EslDbIO4M36a5J9QlkWhQ/0TCJKJGdZ8M36AagGlMT3A5EHemEnOCVjKXC5
jUZHryslziZoaeNetwTJtBPJa24MWdyEhkD9HmzjjotcVdHbXUgDvPhoXkJQQA+jHS3LenqWR6ES
skVgRQj5werwuqBDfRIB5UwSC5YzOkAfutYWJVw1FVOJX/xGfrb6y/7lEETHYirYaW37132KRYXR
/Sxvw8R5+juwvrHghu9DUtIFgR7VRjum3Bqy1uys0ITtcphBYmi6QyN3tLvNwLmVLN/KSQHz4cXO
Bus9uDdzLKN5LqImuthU99jV557I1gqOlVU+qhcCZtNOspijJPYZPsLKx++PpgcjrPQFOok+nOXI
6zAU2+FfRKgaeJYuvtxbr7mLzqyJcuI0jXyVhsXgHiOMszQBVHJ3H5Fe2jllTo194Ae7De7IZe5s
jQnoltkO12WvIaN/VrgW/IsfkDaFXDdBJ3U55R1eiBqyWBPPLU37LOxAq30lYDdIqu0bBYGST7Jl
LPs9EVNYqHAhgPlpILEGmPNVgvsBqbVROtDMeLnr8GWDH5urDG6tyyKzKPnDVVfAOCng46/zIC5v
9wFePtdbVdTFSwXTf8jHSM7wPh5kCF0f5WKLifRcRJH9oZXkWML+0wSZJh7/8SzS43zwWf56Q1Zj
cGCmzJWFDlP0kQ8Iyo0YHMRA5r82piaXJM5HGJk0V5eKU/XX7pbNHJm45oNwkZ7SrUrPjvN5J818
K9zOyYSsxqfj5PHyYRJJpARBcWrVTH5rFlbut2Vwbaj2pQ/Im7ZnpaURBTucMgSPcq6zUlOJhd5/
vmUmkA8AkG+HhgMiNGkYryNAvh6rtpsm0uNo8U6LlQCJqMvuc9LBlCcodMBzAAX1UhdFZ8g+8QqZ
PVs8SubBR+j58ELbfEkC8WWLuALzCWZ69K37EHkG3lGb9DOd7a/CV2pglPeK1vEGZMABDzbbUo8s
8NED8Z0VC9j9uRn7q0AAiRorJsXqchdOpAZZhtIqlmxQDuceF8KKMgUuT/BDa8IghmbVXkNkQiIc
pMozLmMgmZN4Rrartg4ajQshvHp7Z0vMweTXmeLjY3EHmyepxctOIGGEg5BqODkgLLQC6GxjnjQd
/tS3b/4KGqmUrzGz31U4OsgrfP2R+o64dokDcYtVvvk1t6dXWwivNskJkaCGZa1bS2xnzkBSGbE4
Yv7e1Pmklda3HAj4LB4Npi7LzCRBdw+E8QnAForqGoZMKsyq2YnPUIJ0L7k7R8Pl2cU1zmVNx/xs
YaQgJl+ihgplq53o6UFNiEr0SboZnlTxKMdG8OX3k+nC8gLjn1h6Cw3bar/Fc3V5vaSwswZ0c0mL
tsvkzleM6e9xMEtvoYnmDU4Up1qU4uyeCR1uOpHgRzctkTYlGhvVSBqSAXJfA4Sg09RRKSpkDYvR
qd+b2GVTyzJc+MIoo8tF1wzOv2ok4xviqNS+qwxQ3Nh7Gks27kIT2nW8b3gDf0S7aZVBXTQ5Rw0s
N3KwY8Yl/vhiQko2X4Za37nUnqRqFALAqC2vQuAbCSXtQiyvdpgY/0tdLHo4uAUMqBU8asjciwVq
LDuwnnfynyXuDCMH0IiveeSJkcZHk+4hIhfC6PwCxacNta9Iuia+LonIo1Qi2duzz2LQI0dU6QSB
zVDmf2VCjBkFOOvvhf5huoNGOrOeeq+l2BOFXTHv23P20hVVPZ45KrVm6LAwQDy6D6JbfpRbUWS7
wyVY3hIK6ZpEjWANgOGiVtY48OGlxbIJAMyKCubyxPLRqMfKFquau/yIUVMOVbmTMSNE+/907+td
5do5muDI7LpihOqPm38+vgXqiIOH7YBVsP+g+oGGIX45N5lNVXB0iEFDB2N0lYv4FuoxtxQD3pJ6
mxBvU1gJSTrGj/p0hn0oakpWC3s11WXaptIPP16WdQVU8vy5/c6CqZJzQjioN3F6lD1yTDcS2zeT
Xds5P3vBvXK4HsRQAE3gUakseE4EXgHTUfXgqB6ZzXO0LG9rbL5wGNnhclhHV1TLS1GBcX1YRz3t
46HngLBJzsfYFxzdc/MCHdJf4QyVSMgzFVtAonWxHRQZNKf612tXkJg3ZsfQLYTse7uhE4y49DIi
qoKQpnvO823DWOsZaq1mGw6rqjTLjfscDyCBb3RdYl+mve7yJK2l05CBBjjrpTs/Flthwsb/L3yo
syeEsOoG4Q1vZxtU4IYRc79YJ8mPYPDF8fS0rp/u64q5LAGhsN8/3GYO9RXIIRi6kkQnbYEY61VS
ofUcxvWRM9dUwnO/MuHPqnBanEfiA1TJw3Khf0JIRER8eZ+g6Ko7xApx3VcUOURSamBu2CiYBI9A
0JqCgFCBnIQ1dMyxmYRjmHgQN1YrygHfVdx2nn3QDXzj0G20hL3uMV4nGSNsFIN2Juxf7g+6Fjm2
BMgmF8FlwyzLhs5ZANMiK+CQPCH9GkNJRBPT9FOZnBTSOoTU7TCY/61ug/U4s6EwtC2IQPkWEUDZ
fhRgYmvOgyNvr1MgXtkIo1+nUK2fbS0H5hHr6L7Ae0sIweDKHoXD+kvdGbM3RkASXUsDYhR9hhh8
geaUod4WxK2LaqCNyZXN8CQ45izfPXJM3EV04fc29maOF3WZycj2fjrvGJXDHr1lq+bXiUn2L/GC
6eNJqYVC+UrFX3pzYePKRhfoXnrtFz6vGNcm/pE7RgjxUF5bbaDmmROG/fM3/eKJjnocwl5IVoLV
jAijYnAYejE38u/szNdfVaOvYzATzZHgqlPCe6It+4fEHZbR5BiR7MrfkMqIuceSIXq1YRT8kfZn
X2QnDsLthyhkBwtBVH2ayOB4bTsCR4qrPlS+gAmIHtblJRmYiF3FMSFKKO73hq2ZLIO8CHbf1yF7
1y8JU4mgozOuVz/jz3QxU5HqVoJPVOqcoCt3XpDa2cFOtbs/QtfF9Oyw+VS3g4abFQdxjv64HViB
+urlszAqfABGnyK4k17xtf+JEd3NSxtCF2LVFf6UScT0lafXY7k3BvB+vLo4buqknTioiYP/TxNh
Mqc6ylbg85lu5cJTv9exS6eTLe/kLnY2V/r4hNGx0uYgTyLM64QrWcu73nJxYbwfqMU+QWZaQTmo
GWM9Pes0uGrn710BTtk3splr4dhigjCn4Fze0955NABSpFNrRG0l4fH47ObEUuipAAAi9WJTRm4l
7Nfz1pmhMl5JNskNJd2X5N/6gKj/kUxDFn3EfsEU3mp0AczidY4OKGgfL82afkx25JCnSTC4eRCi
Xu6gXgYoC9mL18wKL/d3imf39arF10Z9ZZlxdIgYYEk/fU9B1YTDAwaQjMfvABTYDLTuyQh7/u6E
J/MGL+cKLyxtl0vgpQMBfu8BjvfdehslOZdU3dA3PBc6bJ0Iy5AkF+koKdJkD3NNQPijW4TN9cx1
4Cii9AOhOMiI7CV1gJR1YYNf48Kdpj7Fbw3IJUVzwPRUGRo/8wFTSGG8kSxK7gjVbuQS9gFiY07F
xxCh+rPTEx1OuIgMMozeo6r72IgtEp6D5Wfy5HvbcLwXH3mGtWT7yWEgjr+V27uySCmDN0mehiNe
pkrhVXVNGbhHL3uC5luHzSGtBUWCrLJYp7+e2H6ZMNjitqPafYFQLHtmAmRqcC53deWp+RTW5A0N
y5B4Y+rpFqr41idEVMbSVvAneQTkR4/12C3q574Mq7xQOYHm2GRiqD3nnI2BkzEwwAqS0ikIOqCQ
3HK3alelyHVd1LwKFPKXtizb0t5FYQ8Zhpcr547SzTH3u7O56rAvqqa2nqG4/LZlNYtinXdn5uNP
xnyaIJA/pQodbIu0De/xbgbgtIJnjz/njvabg0EJy3sI9PbcMUqF1thY+okSYekI3Fm0tjpz5ezy
cWG5NK8akT+7hJuROSizkzjwKjULS9fubdzmNuI76ZvuxkAenY7xflbuSYprGbC/Jl+F8tbZLBCH
nxZ9VJ87AxDlEWrqvUZtkZYiiT/M1vzT0f6AjosOyr0oTui6TWhsGH7fWHjQEXIfZGii1f74dLB/
Gsk+KI4KV8/PIFHvsEqheydIXNSQ7vA3m+msddkCoGd3Grr6NZf14+MwLiPKBIf+1oSjAOvVAidR
0TQNyKV2DFdtfxJ48BTtYpSs60ONozNGlat75DSCyGNn5Wc3aVpO2uZtfDIzFSvghQRPHRlDWX+h
dsLcpWied20QjrElk011KmvgDQCckipzO3C44YHfwyiz79WFN2ys8WZm3CsoGag521RIkhni4I27
gf++a1NRMCVinoqfHKq0zch2HopiSmJOAAcxEqShvUr4xEnggxHDdZqeX1G3oAcKsjEKyWVQKFCg
uFnMbp5oKCWgAMab9PcNfFbi2PJAXxy2dNGWq+wWTVVG1+kZE1YmHgtTvAK7djUER7cH/icSdEbp
/hJSlUQIt/OiPGLPo+VbP+EHgCY2uiF6XuEuWMshwX8G2mZf+vseul7ZNp+oEe18PruVDb5JedlZ
CvL+j48ZzxHYCrbyMjMVsxYnRR+LrDzGsMBYAo8zk28bnucJjQasWCNZ4o0qYqDD5oaAlmGHafc9
Bw0Tmx4DtNDXMvtVieCfO1vRFqH8HGZkxBHAefRLUk+JdVHiE0Zv5RgSb3wOY829q8qkjT8mrb7z
jUhFfl9ZgvzVNW6jnHd9PNGQYuapUMcpYk/3WPXvte/W6G8gqsHe2uYSlu7T74v/EvZY2vgcDBS0
SiIc0IW5gDlXoqj/8xiPDfb/U4J9Bo/7b0N54QRgK2DR/aQHLThSTKme1psOl4PW1FhriM9uPP6C
gYNeG3XqiWUj0foCOe0KV/kcpajDiPaMvIQ4exDZ3hbIdE8Rk7kbWEaqavHjkDYZYZkoR+3tdxfB
eUpGtXwxZSoESBJsN741eHIoOlFqzjNGlYRpanBtV0hqgDwcRBFuhuzyQSIcTKqZ9Nnjpiw8h/6h
kx8p5ZbxhCrBuuxdxSzwRv+KHzIEIfkzc/E1kt6TxHVjewGGRk+OxNWdvpBNMAW1jdhfHDFai8BW
4q4yzMAOKXtWPZdVTtQMeKQ35N+7DRDcilTxcc6XyyaFF1zLczPxahybrZdXb+j24Bd9CzFKySsH
m8UKKLDK+54M4PqyUMh4HC+dxbWZLCptSakhrNEFlEiAM63LPiwhk3cXdxh4U1y6gzybnNVkQvO0
Fxza8HXCn+xE8nVRsOnYNcuJqDgi84gG1+GzXrtCD/GmlIXyyzbnocgQzlW8Cqec9pPBwvBp4S8T
bsiIOMoTW4RPBOW7SJ6lRYfQXGPPtVkR4sBwCod0L6VKPR2BEzfRMjuacX+afqPx3w2UTArLyOG6
CtISYfzDoJW7c/5+SOIXJfFPLxp5QBeZX5OHtfzjP6N11EBJ/PiB9ylulDwwlmHzQKGHTa5V7sWb
pEg2DC52i3Oe+BXrafZEXvBbVhProhi9XIn+fYK1FwDqvfnjZX60D4zxyl8/cyAuFRsvBTNhTbI9
FWyFtStHxBjNv/yNmfYw7LHeuimmzPDWmu0JFHwEpsKPy7u3r0yfXH9tgpYLrV7/v1OFtCtdHoh6
wMZ84VZVu+B1U+OJSr8c9qt9a33ADHJE3gzYE3uQOh0NphTeF8T+AFYU3C6SXgt0NqHro9+tI6Dj
2qF2OJPBBhMye7h2XZ+qcMfzTDvED1vzx9cHI9TPxl4YZa99gEpw6eKMYwiWYb/puliA5IoaxG3R
d7Icoh5kyU6eNir0kerUI5jW6r7CUsVfTwDY+SVymJ927ZzPJl+4IfMzJrdprL7s5fO5g/En86B2
qy0Jv8+7U5YIShTclInBIEEaaETI69t3b+AOZ3hFEbDR/wqiJEvzzbEw8cTduPZ84lr0JMhDjAP+
wiDs/N9yV8V80LqNY+TqytyWpH+UFWga+4W6xdvJAqnLBJp8Fc4EP0ZBsLCi3uPFfvl0K5zQq5FY
H2ykX74ZlYMMiGM8g5RXUfmzftb/yoLMOAj6l7RsHxeQJrwRMl70u6qiUZdtmxrNL5uMU6H0lZTc
Jt096VrVp9HnCD3zMnxZCTqw1nv+8zsYIbfgPTEHngsyStSdU4rRg9PJaO3FjzsmCaZYulLNWbBD
CS+JxITa2Whc3bGvwS1fKcQwRBkYKKBC5L8gjIgawYMX4qZWPlNT7inZuAbCdoMSlssNyevox8TO
Gvgl0wdiCXhMW6lugAfRpnpsA1wlO2alZNRvhHHAXZz5a3rSSZtKLdHaEjcc2QNb0v/ikJMwFqCN
efCUZLuBBEA0+pRFXrEt2nD0DM+357rirNnhtG3m+umaBVREZlRAJ4RWQzdk9qCKkl9V5RWwfDIl
EYs4n2rSisfye7h0qIeVKyx4s8wq24h+BtkEaG9rpL1amFpHtpUZ6Q3Rwqmghm2T7NeIzSDufKOt
XLTlcwxy0OwmuK8clqt/k8Vv+Sx5A7opJ/R5hHV32nDN5OC3qHXQ5SaKNje1rowrT65kcDiDVd/2
hO6HI8JiJq8YDJhdh6/0lxBbkyyr1rf0s8GUKONg9XoWUwPvyXseUDfSt4l1VNXCcavxteQ7jNhU
Y/hzkXuW3KmpEPwH1shwTi5R/B1SvNI5QsXS5Hpx8h6msxbIgAESoMM7rPMxdVFehklrYZkkKGmv
ZIUc3tKQ3G+bEMgkQmpls1iv5zvi/IfyCHIXlbMYh6R5k6ZO1mZzIrX489J4DeAFlttOoB3pm+Ft
JYWJWMxSKsXjfk8cg2jvaFuETn1K33Yl90R2gMXhklPpnp0NkAOlL2MrdhpqVmRWS7ZUcz6uuuZv
LikDpUFPbNpxC0/O8Q/9RLyPTo6zFKVutHqh4bvFHdR1eOsOAFWbH3Lk58cu1V9RsiDW1xuFnk/R
9FDYpSwVtc3bHB15W6JE7nqAB25plJ/uMzq7fK73PHTpMT1RfOqW1ttL0/O2PQGmenQK2iBJ1vI5
QzAmAhI7H/PybMFu7iklCFm3xeiWPBm0nAPVMPCu16Hkk4TNUwkVRb/Pe9ACIfgBh79Yal8SCrah
UVA5eQKXH/lG2dA1iHVhoA2kUT7mvAj6/G7B9hazJAZgQWVn2d65GtGTpdq0GP5/btfWwyVT7JQH
dg7FrpUbTK33pU2knHAqN3ZWbBsUhxT3VSnxdVYBRSEKBUhXV/Chj1FuaQ6hIgtBVanIk6QUDd34
95/OL3NRKJkMRrSbxOD9+S8ttcZ/Lpiafy+bDEd/W3DGDOlusvzr0BcM5YtmpsvyciIFiIAFjj9I
T+usKycl/MJnl5yg9cr8OvckTUu923m41KCdeQZOwtjIpU/tL0UHVtBcHk9MmI4V/V5uJHiHIaON
/v3577S7KZ6Wc3/kmTj7Rhw5x6DBMYHzLTBcZbA7GnJa29XdheI5k74rhncZNSbArIOHYko5GH10
pvwsM0rUJwQ4XECagzpkBKlMVglwZAR1u9LCyg4f5+rUoP/y2E5p+mdd6OHbh+T/KgM7FInID4MJ
ijpAeZMRFs8fH3v0hSCRZRqan+b9gEkhwjSWom5HB1bItHx1qt4gLurWJQ3sFfxoC5w9SAuigCOX
LXEKpT1lU+EJ3aKbZiXdAf5Kj/Yf+D2sZ2qcxoOcP1NaakpRijdbKKvRiCeBmebwYWrbNB7aiGpO
tzHsTRxD5rBPWgwV27OuI3iwaaNRg4oD1ySkgI7jGlZPF3dcGav0AVbG+MFQS82E7oz1A00rw5yz
RYIFfOgcVBbmdPVzPNEMMz6SIk6Fi9L9/4BgVD4Fp30g6JZvabIO5dNX2sGsonsqVx0oorhz8JRD
QC/SYK4oed1RTlwmXlWQUgkbmh1PIgpgoUJes4X1U3hUMYLjIOOMCkrh3NNYUEXrMVkV/6l0U5Ug
447UJezK2rxlmcFHzI8iv921FHCh8L8StHjize3xV8uwfh75sW7QMhRRxjXZpKxCsc8CaUshPHU5
DvzM6Xtzf/5nsuzUOfXojEkLZiyHgbtSih2KfsW0cfbEEY+LlXzk4xwiW+zM70u8329MlBlGI45K
bexEXItEM1O0+4DDaMz/2ChZAZz8Zn6Nfea8v6xZYGq9ji+kqiRISDYDoBJFRzscoJxC+T5YB2vY
hTl6pCFdgu3k6GFeK/Korkg3X8yOHOGIhAEisSJtfb5pQxLIvq/PdgZ3eGCJL9p5zbjPj4Kwrdsp
IxXCCYiiQSTJJ4q2Ljt7HeuyWG3In5Jw4Ght6mVxilc5/9rS0OQGL7YL8IP1JplonD5G76krvSth
aJ3dsZdMkDiw55JjwoU+WtRqF2cNNRiiOo4BQGXXC75VGo3I0pTNMFhsHadfZHMs4nHSXYPw6bm7
RcGo800Y7veRo3/VgKIV7nOdOeKTTN3PBVuqH8RPZtbVfNYWtVqEm24srROW5fV6KCmBf5CZwq3K
gX8RuWkcSUpW1I9raJJFNas65eevzIQUHDIgP8TL9oGsIKW3Qc4i+5KUvB/mqR2SeW0sQ4MCsXtR
yGr8p8ogNJHGSsdiYJia3DJoNwGXHPmuyaLcWnRrS1f2lCymtwKwrKheG3uaAZgjqUNZ6AJXL5B0
MbiZ/MO5+cCkuYn0gSA8xGbUiFfd+1ncT0t6DSExKP8WsWT4KJNCLZoKRXKuG2xiTkBRe7REdx6K
RX+2VzjFi30NiQGQ/sBlGXqHveXQ0EkGvZJCZnJfR1tCBZXZE5KN7WFw3qc8BIxC1ogGjmD3uQRK
6KaJ/BjsueYvWg2G/gVVwWsePIUqU0NHzSW+qu6QXLTiJSdEMFray0tvzQ3gU6VdKNUKTZ4SDWmd
adqZxXAC19QaCkP6yNaPE4ZfcN44WpJYYDJFeQkKl2qXkEuAZwy1pTJQ3WTnWLKpc8g8XSvXo7EB
UKvzH0+LRyQ6NN5vxjiGKSMRniwREOM9X433zaxgAwGwDVWMC2s4M0/Ag2R0gswLevdOK5tTWKaR
QGwb+IC055pG4AjtcEmkYSeh2TBEi2GUnWE7a0uBFpnfDDe96PXXpvsJqBhXnhmxAMT9lNLTIxIB
z262PH7m8pESqF86DK+vuKUG/LomshwAP/9ro9sdDz/h0KhZb0iMtDdN3jmnnef+H+OfelD9XCGp
T3V8uTGWlbPreQlnI00YYQd+ppWoeD9OKThK6gfq7dQrsfPzIYxie6NqyX5nrCFQhkLobiB+403j
VNhpvN9tysMzBmaGatVLBH1H3zvAna8WsChHtYAx7LvpZHN9cUb+RKAJNoliF9nH8ogmrFv7E0cL
kIyTlJ5vuwkpAeedRRVkUrKpOqM/qqVIPAYqN2PDcDKv719JhdlIAZTbWAKDQ3l1J1505l/A+Y0h
LRgGwAcXYz7s4SbG6oNyeB0Pt6qKABeIAY2OYpHeRI8GBsHVgBtmCPYvEjjpoueI05sobgsWS4AP
QBTSFtarQd5utihaZ8YqrAJr0kLlGD11sesL3yKVgwoON/MbA15hKutYkVQdPBO1MhwIdR2IgYda
mAz/2BtE5sMkVXcF138KYuHlbFsYWiHTxItbrE2EKWjh94gto8Gb82XM6S1ws1052cN7ynVvruvl
waL/UydgjBTxVP28uMnEcQEfhsvYu1DxXtg2f4KDL93s1ZQdDMJNojIZhTdP7AQNzIfsWWCA9YO0
ohxCIpVMJp5yPznOOWGpPjQg8uG9No/KeX1MAVasWd/l6UUukZlxXL4qfzSvovcRi4ZqROthmsKT
2TyMzfbftNqriL4nDT7O/x4o9OvB0zcxWvkIEdjamgk9t/VvgiXfs5c1GanH9yE6lnh5pRJR7mkg
COr85PGTdI+9q7tr9gaMwz6wVjZPdvHFzia6Fzd/78LU4LJs9dR1EJAoSjHsSfzKRqUkeaNnriOu
RG3jJJiiVx2AdrhQ8k7bmZpUhcJZL3ifQHw2MIwXs4LxiecfGftocTcL7JlxGuEqkmLOdGidlMee
2cqpN1famjRnZsVNbOJmv30jBTCbhbKQxOt94MJLdaNdlSWsm7duTXqQu3hbUQcTn1YUz7izxW7g
j/6g0vO+qOmv27iItljbDl4tUVPfcAKWlqTbuR1YF/7fDzWiPrAvMuRs4nJt6LWCPinK7xykgk9E
AHX/9Fnl425+Pn6g3Y4HtscnPZ+DWSN0GKmmShFtIbdQSoZJoPmp57KESzGe7uVSmjfrcj5vwdYM
NtIX1jxnmxR6+c7FHsK7fii7cVCethAt1uqq0d8o2vXAAJzw4GpsPAWXmjmiEMWlZs/L5YO0li+N
KKEj74AG/nFhsXxDhB4BkfOQT7SJV+54qOew536iivkLRDakEZw9tuSxfUa0NW2jvl0O9nCHZz7G
Du9ou51bE/VEmZAJcrjBVjMGtM0s0C2cUXcMJln9bdxEsRPqhj+TFeLl5cqf1J663c8w7fxsWCq8
yPtzphX/nJCFHC8Srd52/4DlMWgbiRKCDTAS74w8Hb6LaCfpJYolvvLvvGQdWbc4lVdyPPMTqRy6
qyKzIog3M/gjNClYAmcIb54L2r9ilScaVlwOxuY0vqKvsZg1+qN57wcP6EjVXFgILbSgAXwIauFS
G8Pa3YULNWkpa6ifxT7hgxt/AgSEoeHRjiCvqrpC7fGrA5aM3RgH9KQAZ9vI1fSpXcsfOgUk3Ib9
j0RszRXAuFc1lPzLLtXM1YxDNjaw/IVYe1kQD1DvtWWGFBK5xv5xVCH9LSxrllMELIJLPf8UahAF
jUuPESiVNzezV9wJ5dqsIjyUKfpK6aK1ZDWSK98tPPnvYmV2dJAzY2hblJaJ2B5T3zc/rozjRo/+
4H5p7AaQ+PI4qPqOToznfY6HK6/hShsdfFg8fSVfNcJWm8P+laFv7MZeQhqJNTfM9aBG1ICT/1gN
nwP52PJWYrRwtZsUOj/Tk9cTvnNQtFk85CZ6iDANq5+T03YYhcE+0CxFiLRrtsJ1Wm85c2WqGnaG
kS+3lksnuwdKINNBfz/BeJTz+xdFnubofpF2w6faeXuVzCeddhcgkDNgDllSOMYt6bl4Hq522yMK
tmZK+po4TKnkPtz2S3aVV0JemQGeTtnjmQgZCakEhwGBq+8X0bdnn9PWAIMy98aWZeZVlERjIuCb
0CREqiP+IsGuoQKHqh+ccAbEt2LuL2xpDKLmDRtYM94+1ffU5Hmzbz+W7Pq04B5gr4xrG1yEgphZ
ppFVGnEJlcmNJpDW1Id6QwpnHjSab/UxQejUOFrTvs0bprbt36AiCI4L7VBYjy3fG0kKSYTt6tbU
cj3wRJgh5IfB9hQoy9mcWr3BJw77o1w+vqeO7Eqa7IlDMe0GeUyUlyzoBkwJ4cvcfcWRsLCTNIPi
HjIekMsg37SjZ9RjATiv+36G5GOgx8WHgWgaasRGjOY5uqEtQkon4qJxU+b8tFMrpXCZm3FhhWNT
ZE1Dc8jQRlmn7EteIw9VmzkZRdH2VpJAPe/1qvaV6Tn8KYmpaEpGCw3QZjSg0uqVUideEgnyXIEb
+HEbt1XTiqMC1HXjRplnvp8PmxL9WO44nZz1gTyOUXbFJLF34ZfovtLYwa+QzP0lVkpk+2hfEMb5
WMQ3oYoc3E/woCif/M7xOw4CP970Awq9DD92q+kqnHynRm06z+SV+0ZYV2v85fFTx+5Y//C/EgfT
da8VOz5aaPKnV6sgcD/mNcjLs5TOVe/LhFYYTOceuJZjvO8BC5H7cnAPDS2pnYY5lvKFozLYFG+F
lj2GwIb+nFt2ufReGFVmhRlBylltMOzJaG7xLr8CGx1oanweLi57tlqtU0CYskv3lMe1zsNhcP7r
weupB1R85Grv8t4avbXgUKKh8ASQHp2ViVRw7O5TYf87wRJgMzdQ/T6ctY5Hfdj7s11cQANl3uRg
BTi/tdbqbU9OHu0Al2srnjDxxmacebiHat/h1rHU55XbjSZrHq9TvG47NdqS9NVp+vZ81JnErzTf
P8h5fmtDROuqjH8FvJSW1RkhaU5DXqYTfIgry0D0gx6o6yeJpQoiQPf6sWc3YxeNxTvoa1XEqMfE
4AKy7C6biwhGFB6ux4M/BDMnBdVMazu+Mo2csdbNr7aI/fHsE3GiBQc7amWdKsUFq8Q3U8Wb256e
NFnaHTdTL7XEZH/7D5HUCwr29ILU6QBFWUGCuzuNJYR+sJDL28kJSFS1yZi/T3cAYei43MZocqJE
zQpCZiTZBOg6HwJwh5i2zLvHBSGYtXmT5yEmDHTsRfE97HjyGzddUg+6Fd8shlGcDJJ1PNYQZCRH
oiMT72+ICJm0xueMVQD3QeKWUDIAYJj72XS6pcPztAIn/C/o+w0RXocHFaxLpk2p1VKyMCEfAhKI
LxmQmnKFxtpeIqazaUB91mXzbEv6iy46OWKs7HZ4jQ42U9Cx4Yl4zOh/ET+tHetAboj3GnS81for
7pGZrMDq97Y+9Rc0APJ6/C7lZiKyrHwf24uPkUa9HWr1AtslcRIWBHYfICRNutCyhUR+smdN9FHg
b3WGjMFVjnllfMJ6yXxwzSHU13Rmd5PGkCjqzRcAGeQyaCV6ZjDRB0ek3sAIRmjSJ3R/vc2/+AHd
eWZt5vrb6iKA7/JlvtlccIzP+1woURwtR46TxNNcLf+MppFjrmjPAHIFh9dbpPuad0g9P0DXpKjy
XPvu1NSG0S+SrLTWRswK0ucVAlOOHS/zyHofr9D/iMCmKzL/FC8+26S7S3nnHPwBEDr74XyKvrAD
1Jd2a5BRFAFd5ZeUrpIwc7S6AuPolVTpnGqenXpa5s942qYE/ChXBxno9MPaIbnu+HgwUEqPKpiD
+LmR3ezYXcDk4q46uXH0NXds0udAwpv+l6ylfRxWTqWX1cQv4RQrn2CQCpM3tXORViQmfN4lu9dk
urrDXCENNQ6bYxchL/qHku++GpJM/xASvOqfKO6ng3peQDqG8FrkdxofJlJZXcVvv3K1rocvP1w3
3wLJKKfx0vGvjcmdq+l35ikEZ7/x9r/EPAEYIckUiaUXaZJX68eGZT2smtiLIDBt7dTZRbGKH5HB
wuZhO5OfukeZz8MFftnL5jowYimymS1ycsU9uAZFw3G332AZA3URVE9ngIfoqUtdVA9jp+ub95km
eMzyL8V8OJQYOiUMP7+bp0A4FH19D/eJrigDNOHZuULzluMes/YXNE6v+1HISZRv7aTfy0FKanvq
0vFyq+LBkQvRxqZR7FMOmn/YnpYuRK4QzZ7HGMc0XfaakPXBkG2xrGDox9DlnEaoq3Un2cOPQ1YF
Q9+j5GAJnZYkcxFffm3ccuy3tJ5kse3jgJ6n+mjvN8t6BaDQMdjf74+ptIH5GRGGukJKGTLZad8p
v1vhj+dNK5WvzrzJdhdJAuW8OBbimbHGQ0u3iV+niHkEPgpEu5dPyuApB9RnjJlAedI1OP9xeZKv
V0fzi60qRgLG33EhS+33IydEXpBlbU5blEmvx4oU0xmg2uc0YFuIJqj51pePtp1q6XWHqQdlUNrE
sN3kTHVFUFZyua/Z4aWmBEayFTudMMzeHvTrpbuxFvylyBNxSvTBvXJNAQZyclMXTFnjKizKuiQU
qbPr+SDn1iMqLl88orAvvjLQv5/bwSFPo5Fy+4aAoTLpiPuDlTdQalX2/9J6iqU44Q2FarjbH5tK
q8yB8itCakuHmxjMu0xlubEMG8MVRn409xYtZLwYrEuABD5+2V2L5sH1dekI5S8dxMODCZnCuaLL
Ql/JXbL577SXMq7mz60mH+rZ/UgZV/k1C1QzG9IN6jW96+o/1krZC+UJZ6usJanAMK9v9BlBa2G1
FHwZWd3xW7xZ2UZtVU4EQtAOUIaOtzmH34svLlk1cjRh+HUNTFfd1xdh0U80g5MDeStVKU+RLFnd
vq4j0pmc6HetNeU8c7vDqSj81ceRDOeVbS7d1lNj0Nj1fSoCh1t4rvgE3oU4yoEqRDH/RifQ5IyT
fVSmdRa/vWDcuyqAmQfT4llLNWWJy5mi1SnXRS7qz/l/BjKu02QgYqa2MhtfSmeZRaTta09ruJUP
gZ+YuP8ZFXRyz7hvexz150yvE7dSZC3SLikidsj6nlv0Y5HjYn3yjUIqxKeLnQpTVwFbTd/yii3Z
F3f4LBe2flRtQHttIfjigZuY22jGikWAinTZVEVc1bJ1FoCL309zgmsQtIUFd+RdSH/RiNrnSIrP
8LcGKPWLzBf7vbBqmZ2y2vtloQe/sdNQDU5CUCeTaJfKSgQNs4jXGdaG9G8Jvf+feWQqspYRFtPY
R6j6SfEJaeLmXFZAhnK6SAearNZ05WBYw1U3isxgpB+1ECqCgJGgAoGq6Y3xi7czpOXYYXPtPngw
kfdW/sGLB5dA0KZ71M0kHT3N/SEtwb4wy4JDwxfJLN6nhtPjZagKq+FpA4Fl9Iyp9Mw9OEkE7DgT
2RvYmeziG4uM1YWCo5i1FoSqNCfggCueWLZ7RX8n8GkV8Bw2DUGQ1AUW9pn5xQK1WtEpA5b9ebC2
CscIaw7qNNsv0NWzi1Frd/xw2OlyXlse27UtV/CO8SMaDkF+ILrrhGVyadYHkKujzMRFVMDagDI8
tWO83pAwLPfssSmvgH7Oc1pZRjJPQRbR6xvpDH6VfjFgjAKDL9QaZXRcl9aAxYFjDVYBi3KvikUz
CelTwPgCud62SHk5mN40pLOtT32JQB+BNpmuBuMlUUaOYKCIGlekCZ18UUEhxyKVI6bd1RsAoklC
jLrFXsd2fMLWwuSD7MnWTbmupHNAih3k3HqTIYVoZH7qSSsRLrRr8i1f78zJB+Llg8soNs57Z6wf
/wjlq6532z4E2k9JE2ffZLc7DDIwy2w2DxB35+rsnzw0prcXdWdQGFEYXkXlM49Z1aMebM1zHcWV
w/5P9NJPDslCRcDwjM4yqwziIQLVGluiU0JIl6jJ+lc4lPBIE1TmbzekTfp1dbL1o5Un9fwIis82
npaAtzaDv4ECp+867uyjrV9PjedxYB2pYTOI1jFnez9DmfTFDtlTiOrWbBhrQr0qc/pDHBrokvqU
72KvjwTv5PyGo6nHYot+jKeQEzQkyIhvf79dPTnM2RvXXk8LdTo3ktb2cABh1bMoIwjHxolYWg6Z
J1HCOY4B6PzogmqHMQJToBn7EL9enZldLw1bBb+rihXDJ08jWFM0iohSo9dEZchZN1UCInBq1tMd
5p2Di0FO4xJS+oiPqLzNn0MoAs0OJrugMwOXhtOKEQiFt7Qjs1vs9fCcgcjI/rn4/6hYCdbvi84X
3ak4gSqyLUuiilBY3VP2BSpPYgSNa/4Ff2rS37wqIxCAlANqw44CdSwbyJzWQFnnvo+9ADymMVJD
vP2Pg9M6k9b1DSvXGlIOOkzenCGdd7Dt2D7RINmSwijBbhXydYDhAfSZBZYHFJGyqu2isc+O4DlT
IIBhRig/Wlua8jAtaqDy8NJi3Ia2PeTwtdu7nFBdby8p5J8ohZpK7ceK5mulxxG571lmkBUtW7Lu
OlaMI7yuwQ1/2THZwj23lU1bUYCkQMr/do7QnYlOMLnJKRBP32TkfTpunThcwq6EkZghJUqWDgXF
0By9zqs+ytM6/aL+KUfsTrVuSTilt+D6W03ulcEAIuucjPDO+2BvGzjEVHxX90pVSZMooDFV6F5u
jchlyM+KrRn3cgamdn1ZFmJzXmhTgX9ZrO8voZ4tah+/Heo2G5TQvihVv+buiVrIDjd1O9Dn3Znu
Dsd87ISqJCfbEXlRJJuzhg8q4tC0NlKbHEShXisfD/bf343QQB9dJuuquvcWWpNTBZvYolzdLCaV
WSovK23w9HCEQmvgSp22bLQ7TESytDMZZnPsl0RjQB1RZc2MEGpjsOpwTjbllb2cNDLh1kVeUAJ5
D/kXy0hXIp4QkYWIjcvDk39e/ogPhiKPQvFko4KF+GtCeOWFzlvd6D/kGkOi/l803KOl0wwL6H5Y
qkal6QyJYB32Oql/pHM88x+PDPt33T4RhKB3W/pJLa+bWlZcjPmWpJZOz6TPsh73r7KkPfLq9v6b
YZTp2jacnmteRmffFKjTQQPAOdJAXL6c0nZ8mq58axfmEcxgHDcwUXXQSxDqhSUZZ0FKOJuwI5nP
E5uK72JyxYZaSuOHT+HAIxvG4qmApkJ8EkViJWStOEZKz//rAgWwCQlTq+QVyh/05enCj45fsCdr
Y4jw4kJq2rH+FhviijfHv0muLDl5gzZn9+JF7SC1ZRN1kR2R0FHZoNA+j8qZ7fv49DeAnw5kLZmy
8IEdA8npx4rFqggrlUcZWdYwvhsMMn35rENPsHEO1g9d7cJYfUs4JUnfwyhff+wCGigHHmhik9ET
hd0JYgAyCmY8Tr0sX0snn83BELZkH+iYDNQImzHjhVyJrO/vJmQv5hdEise5Q8bvACKpuSnzQZUy
4gQy/zNUreQNdMjJf5XJGNY7eMk0gCb6XwhY0wDxgnDyQgsMlZvDT1Ulg8yDejCbidZhWs/gDy+S
TUKql7UxNjCLvMz+5yCd5zsT7ymTHgjpz14+ZqhqsnvTMKl9tz7pVjT3hqNz/16J50TNYAhbClpA
YeO0Rd96gBElMAvj04ExyA+9bJq1sRx55i3u0FEFaJQBMYf11kXetnE1bIRTpYt+UFKuFGYzPE3/
Yl6CekGos3cbAeDxHQxS2wZ6Wh8hyVOSoCsumpQ6l0/0oSVp9bc3C0loIFWyod6IaGlCud3/4smj
qCYe5WwSlgE0z0yRRPOcKQDrT/tUfvQpE1XfYj2K7HGHxS/umsOgNmQl1DD8KXHRmWZwpYW3Hsl9
15vrkpa0aeuBe8iYRGQR/FnrJbFYwZVF4/vlwOFasT+N9+Pa4SieXu6Ai+8u1iJcdUHFFfjJelnN
7RvCLA2IDeDT6hgd+2nmFyIs7bFD1JGJ7M3VmarSsiLqFtz0zbM9oCcX8bIEQf97hQ7iI3mvmgoL
YXrb0IiZzUhDAD+1HtiUPkusBbDGnS22+hiuIi0N8K3R3/bNUcj6/lMSintd1WdLkqLMZRLaQvca
2lAzgOvKo7bZtxtkKPELoywRi7MFcmrkfKX8C5vj2sHhE53asn7HGMMAX30rUODnw16LvZwpmFwD
Wu80OJvpOOZYsZ00HXuCO1VSiRxv8PIjfVmEXePACOHkXyP1UmF4Yi8E8fg5v1E33sIZCqHs0z6j
wGup2Remgdm5xugxXUCBqtjcAE4+zB0z2SS3Wcreu4VkRftwoM/wpGsoNaXrrWiEO4ThGPntGq1U
BHiNzXmzaPQ2rrH5hzmFswpQYXtHxn+tG2dmKtIDAanEx431shSVWG6oztp8+FVN8QUIo4tBy40w
q44qkLrSqP90PpK740/4EkGaBWux+wCDutSUcG+tNnLWZd7in9Sa3o+xdUFB2HZjp8qY+T1ic2ih
39xAONNSZL48OFhYZl4i6lD1Svre+pSIzTkDGzY2wXsRLICD/P4S85ZupxX1cAT5p8RRYOhKIWdW
00TyZjfTKG68l2Zjl797sR9ayLDrY4Q2q3RZx2uaR+e8xYiLjqjlM5dLXUAZxmh+EkZUrejccVAy
3RWhgEkLpYc+i6IEoqroXgicirAyBlnfbyd8q6//XO7novHQAvw4rDjDqgT3HtI61XvYT2YjZS09
oyvxAtJLUk29lRE6ZwwWW7j2w16+gNIFVuw2dZi587gFRjBBQjRUezxjiU7OpWh9kGIH/evMbPqS
QwLdDs1WK39CcB54r8aUNWduX2Y81hxUDyWRxVpXa43pJNqnCk6iUuzW6LwLX8Gx/JYGk4D/37ua
pXHZEg/kwWLKUVlwET6Aafbn8/amhKVrAtig/4oAx5CzjrSG5ICN/0nukUsVQGvTMuFghN1XkxGq
hR1m4bZybQcpFgVVA/pgVQvjZN7P944/npP2l5VJQxfCaprr/NWRKMy71S99Yvn8W0Igkz39tmmP
jdmJBuqJpNEU267mEXMEPvpPky91iTICd8szoqa0ojBgyIQhl/NEO41zHd9e2SDEbtZELGAZLZKQ
FPN4Ne/U7sYYYFYqyI8NzQf86zUcY8wxjMPjn13q0T3g9NM1Cnm1mQwz6uKOn+b0oNasowV1De0P
6F2FJb6tx0KRqhWGlQuKIk2PtgPUpsJkxo57eCCLKJwW1AjE4qGSg9giXvVQdrV41w1lbVhJ17r4
U+hiiRwfR0Sxe5W/lqMg444S08VTmaY2oh1WVu7WLyYbxjzlfDSP016blhZ4lducfzyXuYsprH1k
azJfXgCpgR6j0N9/BpStHA8PA820y7zCtobvwsHF1taswUBDrxu4+PKQga5rCeGxr/0tfoSy2cRD
XvFdpQkLEtnx+bGnOSa+SbwhtP3RfheE472EyxFck+/ApsWREJlY+ZpHbLOd3JJrtc/CJZrCnOX8
Cq9EXh0F4Zf1zlthUa+RLhqAHRsSAv6QQBrMrYf3RPjBbNdOsdZqpBadobMCCLCeWOoNPpQ430DY
BJn0qIvyE6A7onIN2vEFVhQ4ohQ/io3hMKlUci4TvpmrG8da/HTZANrtHYI1QwNziXHIbuDI2aSK
DtMr0P8SfMIfvIOs5t5O9R5rLU5+mc1bz3UuepqLxj9FbkfQ6e6gtD4Dh+DP45QV1hfrk/7EygKm
2ZOTUf3Zq23/d+yyENyllwZUIYK3AzVqkltBLc6EiYLArx9uKPPBYITgM4yGOHsAT9wCL9dJ7Zqw
JOVazeYxbiHLtPk46h61LdiHX+dj4J6Q86aHen9yF7lv3vCaksDvd7BEITvEijhO2q7iNqP09Z08
qOimTNgQhZjFuwlsYYZ2xLuRcM673xsEx/tnBDiLSxWhQRoeXRc/vnXo630fEtPR0qOAciKpJliH
Iutr3qEhwSQMe5KfixLFEIzbPS76zR4gYnnEAt0x4bZfWCfg/J1zoPAz/ddOQ/4HEnG7LTf5kUAG
5aV5nAiFvwjwvPlG0G/+DFGuDoFLFfRpGUEG+0HIEymPpv7h+tQlw2KW1YQJ9Hyo2xJ686L0TyXl
F7aNPc2TinnMKAsLvTwdIWmP5PPiIGNf4jqDT5dX/TNuvNxiiVnOVuSaW5DDp3LwBeEfCYLiHN4/
yUujLJ7pCeH4cKp5LvqQeNSARqyRMS6AnhXAjqf16Ef9/8782teBRsNFwuKS/9q/D0qAqh6Cqi/I
JNe+I3cs4IIl9BcP1XdK3fylnrQmXpGg9v5Rm2/vNpjvSYX7zEAv7xnePVWVjUZMoRs/zVsg9pTH
iXF4AU+9pOlCndUHGJKlrxWPlfYL3Ov97F4NHH75yYqpl2Rox7g+9zvZz58CMrzsLH2OwsTc6MOl
Tc+BgwKXKpwdINaf983piTkEbxVRaZTNfkYbW8mq37yFauKOpVDJrdBdfNRNcbVCHj4jJN6JKANu
d5FyuTI8ouOhk7dBu6Wr50ABneJ+gP1fiLzKHybGaozQ32RCIL9uIZwU1p8Mg5lJ7ucPgMOk3Tvt
Ya13uDTpPRjQEqU6Uf5zwJcckUFvRZuj1aCuoaGO4Y9ezUW8sF7+Ojlk0xtrI5kW6clNRMqn/WIW
ovlPEInh2ZhAdxO0LwB/0bJ8rcMksXb3998aGKqiwS+xsJU2a88v667onKKmnA9pmoa1CnydO8Ct
mJ4l3I79mivpXxqcpln0cBPt4cjnR+BsMOwF1XGWXmjQqNj1k7qE4dENB1OT80yKGR33w1iZ6E9O
hW+aoNse9yrkpIHDav/hTruj8q5GAZQWr8LycDAmjCjfQ35J45x+Kw0e9uDlZ5Ya9pulbfXcbc31
JodzqJ1tL8SDuWiSg+vpnE7WEpQWehdEYv4Emf3UmL5lRzNRZEd68CzSfIO89P7k3T4AxNZApnsq
qG/8YcmQaSss+wTJr/wymtiM24tk71tdZdeaOsGaUANOqxzLzY7Gpwhh3ZDDbbyuyx8bzkwFxMlu
kBLsh60XRBcM5J7BLGTFIaJeMnsP07WuS/o164K693dd27sfw0hYo/UwwJ5rrWJbQK+kaXipWJ33
98iq+Z0K0dsqanmMTdEIkg34u1rPIoDDPMisoV6GXZ5Q+SaSkXosd7+QTcLo8763o/u8StjfW9yM
wKFjXSGA1nL7A+g4ZLKNg7B7YKzEGqAMUJEOAihl1L20Ucwxh+PhRW22fed0+UJzJ4g/rXw8E2Ik
k4ArE3vKKgNEbBzGTg8FnmAJsnL9JnJ8a4LqEfFInBv2hRP4nDpY4IQKS1vg9FCyKhFI6t+aHuia
5GPCWUkAskUrhtOQUVUF/6awTDPV9vehnddGrJgGXJ6/9aK/Qc8KlRAbVa3aw+mUEbKqYRUggk2x
XmyFw0dIvbFcsno6m3VV2l6YM9OKwtLuQmtDqS4dIvV4U8GWqs446BhMKdy/reRAjobm7Yqx0XGh
8gHEpcJK8Ipsj062oPjgauwDQOlKpIu0WoVqiqobfTO3qmIg93t+CEDrLKNz/FXYMC1jSIiytJu+
4qjXrvZrU6Rk8iz9CGr6UbJzLKuRN+lITFli37W0bGLdM+3t2kt1CoXq2XVwmUAZvE9v8ZuohJIX
bQJ1zZ0mZ1JVXDNcJ1pZeSbvCPGz3wyDtp/dzQ8Y0OdGCvYYx4x+/JBC8UIjbsWvBrPGhCOdPeue
m5KROo9RpKLj7fS1HfooLiy0yiFz7Njroz3J3YX1aQJkeCOvCix/d1ATCBKb4DPCUwAAIpqxUEX3
Q1K4+LiojK6m/KNKi0ZvjaWGRfZHV8d+ZeEfUPr1BU27e88WopWhiz93Dv7ddmuuHmgQAafsKxVa
UBUhJBt8KEjN+U9z4nPmRln+adB8CxGdDgPh973BhwGUyKPkvj+UqAQRY1ZKiBnTCTw+WkVvoU1t
cRD05FsCkA8s8CbCYCJ3U7G45fJaBWDXLRoI0SPUxlo8t1+qmvf16l9n/nq+n0JgL1sYOtmolaJG
hlQQnh63nG0ejgHukMzYTx8CBX64++YiZ/dRWYzttPAWRtoLtE8pWSt/8tmx1V/NK0Wwnyszuq+E
cmDZ00VS471Vs2m4HUDZBmcwlB+CCU4kpDAqiK38Z0xyQ5Vl1zrABC9N7MMkVKyD9zeCNjIhgAM0
IkSTA5c6KgJQOj2LPuLQ0z5IX/dHE+XudXm4RIhXLUb0YgBw+3xXOF5ulkI5JOn0KwD65R7Ob6OK
C5RoC7TtfbGeQHtTHpZnVseM0il6L9X1EQMQ9ob0f7X+H9Fpt3q8JpkFdLGgSfzFVchRCIVD85Rb
+SyaZPvoO3YTfi9WfrY9Q5bN8g3ihP1/nKrvwwBcXQ9dj7n0M2wwNfWHVUnwlRtROu49tLG0AjYi
oT9MsQP9rCXYWWNwukHRY3/vaATJzVjKO4XvIdatgcMTquWWdyBZO94NG9IH056Ge72bbr0Pj4uy
gWLgu6hcDhazAgSWQrfi/FI6q5U08Se0sRjvpV4NdgIxdxPnHib7+mXiZbFQ8zWLKSpskdRjtGcl
dTL5YiuicpSdLHmnChZu6RXrxtompsZUjhKs/Drso5RE6d7m5HfHNqR25WEPjQa8pJdbchYfJNnQ
KuUono14S1R43ZOjHPlHuN6XcRDbih6RtTIlagOl8xudjf2C2Vxpki7ZgQsiJa4GCkeRqboYh6e8
syRFHMPLfFAtjwo+/mOfladH7H4HzJaqdgeusODhBdwv5ab/maGGW86AkRu/Y11YqP3YGJd5YBcT
pYlG
`pragma protect end_protected

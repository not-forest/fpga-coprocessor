// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
OzhAk2RLwffQAsgHyqU4/09oSEjZ0nmFEwFZXniWtigqkDdOTckCUoeLhvMKOErL
waOu//2eyPhqNa6HdrXBG3jI5l6IKM5JxHvDbZVi0bni1abL34/WU9W7yDSDAx1Q
p27Vd+LU7CpwOZBrxxL7UOzTcnDDkgBeZzTPo2uHtVrDmOoA5dVhdBbcZ/5F06ZL
En1iCiQAliYUo3jnlxel6SwQp+Gfu5vwO4sPr5S2gcBpyF1Bxhh/ndjjJVw7M8FS
XwRO79K9Yj0qLUlzyu9POZaDvt/bsCeEHNscvgmWiJu5z18NHE3SmAzVogr6eDGe
sxGtBbCO8qeu67TH9xSgtQ==
//pragma protect end_key_block
//pragma protect digest_block
jn2FYV5gTqA+e0IqOpwlTQP4Ry4=
//pragma protect end_digest_block
//pragma protect data_block
pHF9uapO5BBOSjcRC9GRUyPXOD/GmAaJFurZgZ6eoKNHZxo57gFH80xycjdFLnJL
temTl4T/iFL9TT8XkCaSVWE/jJjEj5y8WqAIg30ATIwlzIuZFd8j+THmTuIAmyDR
lFrXHsTvcUoXqfBu93X6X+cExdNu3CmrCBX8jqKClUN8BKy3eDlmPodUMC6NlcqD
Ubo9JN/o0FVbMcR5dDr4hoGbL9fjnA0bbz82vR/kwtWEu2jGRWEDChpIDUx1L3xe
AebAmKZuVduBntfGtPz2AROXmH5rcLO9T2zTd+LPaTSfqdd87kg8L+1pT1iAoRlA
IfgPJMcSvRvco5bU4djuG40Ziz7s5xsPuQ9sFcb2iwh6MqVLV1pCbEPjYG8uUi2b
NCHTCkmxc0NLamMTkLMWoohUvbqs1KN0KZbw/hi7fUU6gj32FdaqDsts2qUScOpl
fhUQQ1TZLuLSev+VTbWN02UB/z3mR9CKCLMqFMkXa8mmRNbtoSh+J03bRKYTNHLv
xU7idKc9SR9fRpJ2yOwqxqHoylMSIgIZTV+whPnjLr1C95KAor0cAtW0ZnbZC/2M
YyN98NbSpQEiNHK7KFJyqBUmLF5SpYxDLvHG3/ZSMD/A3JvCgxDnHVO9VGl2Fpk2
US9dWOuLKTEvGdj6UKGHYEdvFIVRn5NybNTgPw+qi4b8HkKg/2szxB1uyXWLnYEf
05qMHHQpqvHM3hk9+r7aPQXXRCPD33tqJ0ABhdOn61zzMA4mfwx96wzJpY6CPETI
9o3M8pTLsQR0af92+ScT2TxAG8mCEaqHxRaqZ2x+nzib7os8aFH3Y9dTqdRq2XBj
Bf4DdKbt3LXU0RgI6pNGzDksXbHZFN1J70W6pmeErrEuSlgMrc4UJZUfba456Fg0
nEvkDZsD6V8vuEetlsbPQZPuq+3C7Vu+WtL1c3kgEzntS0y4ly+mz8bN72moy7QC
17kivbFkfIc9tWFrpse7NlhxidJ1P1fwBx9sCv4WGfDUOltlUoIhwokRhqGbDPjN
o8nFmRZYl2UA28EPe8yF9wVDWVxtM/Je38rSupkpyEvcOiQM7s66JzGKMZt2xZ2T
VSaNrQM5EwL7tTm+uNF2fTVI+NyvlCZyk+v6u59epOT3LmHOYIh/XNKK/miuVbtk
w3ow7q4l9TEpZHi2jPzMFvkBufei6Lem5hU7bkY65hjwOJM5mWrVFvdujGcwmFp0
nErZcD2g6YWlpavJAJUV6/IFwSxvxuH9PtUo87IWCJOe1eWqtC1kaiG/yVb5tkNF
YxQmrwB7xvTgZhtsjXuapFPawoA8g1mZXGtmRTc9g7UDZJHD4i/Cdq2NvbEsRppP
VAbAweQGUknB+Qr3K1rm6TEOa2xZSAZCZr1Bsk2VwnIW5jGvKTbbMJYZtSzWSbjv
QGudKNZ1b1npAIZ+9Fh/x0vCX28bMI2y2iQCshWaM7diL9pjGa1r7Pq/3RJYQ8j4
XlPIhYQBsVIiF75rI7pXlhYkycvheONWnzkPxP18ckaARJ6k0WKFcvd9NK3AaPAc
w4NlKziQmxMUhKW4snep9Pf65rj6G89L+cxpNc1U21iHsyjLamaBhNWbsN3yWcUe
4VRCALqCGuS/2UjCr5rHxvHCd11afEqXeee4Fcvi2Xtxp8RYmGJnCxjdcjb3pSIX
a3z3y2yudL7a80Op1DCYT8vzVBzQ50cNOx3BhGq9Vm0K9S/0/NaL/z9xC9LHhecE
NgOp+HfcZhBE18nubLUZcBDQqj0dJ905q1hpoEmbhB4rIo0jS/O8+bNKH6n/Jiye
BNW0n5CBHER3lAXI+VBQKD6jLgauH0o+lGNeKQW80C5MmtAfwgG5akfjbAx1Bez8
3UuI2cSubHRwx37gUp4nF6gsVO/HeTACzO9prSici/EURpMZSLCh1VRj1X9Mi9mv
e8LSQE6LU0+n+SAlWuGNI11B7NU5++y870ljlqGH0s9V++a+/Hzu5ZfiTiTvc8I8
RXKF19bpN7VYNnPwDIoDoiqSY+FtBu4g0JZ5zPDIWWx8uIrNWD890XhprV6LtmlG
L/kYy6Bp6VAdW3QObpwR3ZBhX9Jw1JfKWX1DG48bFsmKKcmSRErYx4x6iqbimv/N
3e8bOp+bJF4CmXjkSXdgd6XdQlPKXqLz19ri9MpdHZObxD1TI+srmU2CWNu1TNYf
3hfdbSKts54uci7XOla1LX6XSu1hYH1WGk8b7Rtvg2yt8VJgJ5ggV1ajUMUM4eVs
6f7vkZr1oYxewrHg/VctN+0lsHB12cCnTlLfIR2ssBh1IDm6j+VN1xgR0DjjxsEh
hsa7bW+5lK8LW5SNKcOpYgaqf3eGSYWvnYXqHS/BvSfed32+kkEA1c+RwVAb2ewq
a5Di+77CKW2n01eeo9ntCIcoRMc1Jt+RpcC0WzMQMVxp2z5xPsxGWCy79cRvKxap
1l80UR6YFVHGSz08Q9QVj2je9izHSmZcgoRXtQqkim/N2SJdHhuHA3TvhDOFIbf6
VqP1hec3TMFSCkRkILarkW6pBrM9IRSPc/mDg6ETEEtYACfQDGWmEIMM4T2/Pakv
Sof9UOsbPnU4JjXkXbBWmxjPnPmoL4PFdmBPGRqGxqzgIh3ur35Sx0yAZanpAr74
IxQeBH/wd8gAGSRKR0wdgvRKWrYXNGeZmfLnGqNaeRaPcEeK599MOVz1ZywJUzfw
5F+BPfyPMCIjx6LyQL6HQeV4oSUCJwg28wNfoarLO6Vsu7sdRFgnWlEAJmThL+S6
8Af2KW1+SCK9Tl0X6j+SS4dlwtHGE/nQa9ZUB0D3TMTqwo9K8gexPC/oEcrL6M6L
HkwyisZWIMctiK5/6hecbc0FoSqytVFMkk+FeZ81stLUxTWEonvq/2cYqjGVGoKO
2brR8S/7kbr1QAFNIf0gdL2jUPZ2JdNjPeUYVN2gMH8d6RN2ovpPpufTz3Fduq/p
rP3t9QUt9XySwVg67isZsKavvfUU7HXX9/L+jrjRdIdC8zyBT54/s+HXSDvOCnbz
MGz79NYxW72cS01V5cFHtax94z2xHJjOPpTTu45szVz+gSkWBAxAhx3QWxKVZgwk
cSWaCGFdYCPiqgtNHYPblkHuNC4YI4DqHaB4q3dn0iWBvnHSbK0CB2GjU3M0fq6h
HLyyUiLdmPkFpinhJfEUawsxfomO9aEEme488EjXuFK7+mBGOHitSUQjVE6DbO+m
YeMUjaVjKd29rUUt3VgbSW6qmUzn+XRxeRYBwy7f4Ojzs9xhntro9+4P0GEZAACw
ByEN2y8EDC1uzghrZG0APSHBBxEZ0CvVNgu3tE4jA7bxIzJtS2QSn4QNDNxvK7ed
p+BurN+RfFJ3znW3mN4L+eRlASjgcXjFh7zCV1gjodr170jdg3u7dhW6Kt0WzF9i
DR4h8v4KdWl/E8UD+H7ISvkB4jSJSyBBVgCBkBl2iJ8KseA4S2CWv6E/e0gEqcdw
GZBHzU63XdjqVwEFurs58c4KR6o52c/DmUXUaJOuaQRc0noDIVnaBOklkPcSCVR5
PDwNxM1jlc/ot/sAVAX6PBV0n/M3WUHjhBXHLfm+RWVwwEhYh0gNQHExhjsFS9jG
oYXycBF0a9lGZN0evAUjBaR/7JntudkSASwY9K87zY8G+av976eot41Nz5tSiH5u
k0FactedyLUtcs2XbXctb+IidxmF4IpyzSk5LuOaQXtsTHaTmBouuTpSs1CUJTs9
S9icXYOGwoxOcAweQlOtT6UnaZZmnVWfJqpPKfX942xARHVHE3TdJWbVnIcf1rj3
BhyjqFEQ+mzs6Kt9wulzelQoZGCq0DpxMUye71/0+027qIETy34tpOlDUbxdjMdX
QWGukzyuC83CiLHROnt/SXQdZC5vavnWbKKv484urXsHTICqqTQu6CsRZBB2k2KC
ijK8F3LkgZznU7AzXI3RnEMb4qelX1AUZqTEIfp7JEkJmdrCI5/Dbrt6ZAWSlqrS
lGe4QJBM/l2boAZR0mj00Fs1xH2BXJ3Kz3XxogwttyKkP3Pc0dJfOeWNFQnmavnF
5b0znL2TFx68JwQq2bavwFvpJjIDZFNHVGgMv+3tcMUugSWxc8jVKak52yOkhl2Q
ujZrc80RmLHvOi3IdJPtmdfWVAV7x+j2Qky4m2cchufHWmKIgAfsm7tPrwW3lmW+
ylnqZO1u0hJRDNhjH5KjNJoAkjkEI8IlLjZGzu4Cad9viLFU02Fnpip/I0tMY60k
GGR3Q29Z3SLeLqeliHKPQKdY0AweuxcgLzKiNFO5CrAbi3R2xCwUhNWrgZjCIIKk
pis/FHDWb46qmk4ndW1LUgh3uTGTUz0AerzSQyO+xQ8Gi4UjOUys7X+zTJZ6+YwZ
tdE+5++z5oSLkVKeeeQ0wxfG5PWRdTPHY9cKyPf69AQLtXdSkd5jijz1Qt+U1xcv
GWPyLpiNT9h7KEshA6VCwZCq+lgFLA+p3EsntWU2FmIwvLX6miF9KYFnSyuCAGkk
JcM82ju7izyLRbyroKE5lEJDBIUB4TNyRxy7mRsSrgQDNXPtKiKWgqVlg2EJYdGv
qaEtJzVjbcef7sFMn8jPXnlY5uw7Krd+0+pw9X2CQeblHV9pSrvDzNrbg/5Be5fA
G6u88pW52go18s6HaaMmhu2OXkAS9Ux8EAOCzX/lSIxOmoQ1Zo2hviH7Sq1Yx5aO
yIbPniReNp1HrXd3Po7Ef52sV5w8FFYvwp9nNOBwegdG27BhGC9Fgg/kkzoyflRK
8RB9r/DGzwbmyNPJeuQ5uhqZUrbZzzqaNf7aMoQrbXNhdXc+xoeGZmH3gltJXxgC
pSoZ85hfKRFqU+KcpZ65kPvVQik1mn55ppa+gjcKwXnIhb+gFsD4gQg0kS00NkB2
pZI9GsCpN6U+UXAurE5/aekWJ+HNOBIL6SVZOHDcMTHNABO8I6tnKFWQQJ+Ehyjp
n5OJBDXCtP7AUxtHXsXx7xzR3JI+7DbqzvEzGISl7AngZ7OjZHKSIFuf95c9BqXO
gjbT6NvUOJe/VQCm8yfaXPzRnoxkrJxDdJ7WY0Gwa6pwATLq7Vr1T4Z0RzkqbBrn
6PMpNmfbqtbWX+FDi2o4dXR7aJEGoW//3R0yrHh2E2DVwGHLUlYlJkLZLfr4ZSiZ
/tLdfxzlMBzAo3RoU3WGsJfrMigIdiXC2LGBLh+vKofBiZrvgv9v+F9RhOChbWbQ
9xHR4d7DvjWGrI0JQxYTOjNn3IGQCNaSl6BHzdV1Du/OIIzC2t+g4vsJL7RIa2Ds
dTLDohY4+WkM2um/SHCgHKR8sOlot0WLIQQFWkt/RFnG18zRQU/5f/oaVkFVhKa2
4FXuJ/iJ1WKzrwNysWHd3cjR8TPZqb4/47ekA35smjZ48BtZiSLRjNYWigC1Jzjs
cx4Y4oixD5VMI4SK7G3Lzed5GhFk1N0Que8LBryKH++N71QUDRogNIJRbpqTOOK3
yTbCDKj5eE7/DZsnzYhnqJ6TvC2KZTQ/5+s//+DKgf2gmOdHfpUfZd4uoMCbg24o
bvmPi4rnADqqAluWsnWsHOy0RyB5lAjIx758TKPHGwKYV2Esfkh5cTVZzCdkejWi
hu7KqjtH8iQTPa4DL0aEGT1E1nwRIJsCHto8u1rMpuifZFbjh4LrvTiH5tEdaPIo
aUZRV6SQY9xxXYA8fM5DashBiKgqZJr19CYWCIbveQFEujyNLvUoy+MHGolpzCbx
dS7894lK0pgqcIKrZybp+xKB+82VxPLsn5nR0Tk9cH2PpATUF3DWTBzsNs8b7I4u
DFvVlYZ9M9gtpeMQ8QoN0zAdKGmyZOoTxVR7LlHwe9oj6hoyw3D3XGfwIvXMJh9Y
J/9fpy73iUdCWNdcyZZHe+EDehqESWRt6p0Z8a1cyvUANPQaeiV28iVnAHeXTrkQ
DUtxk89L7tRG0uzqRjyFCasr41qpo99qlQXYcE444h1xC1KylrDSlaF2IKl4R18z
r1/Ykye6tGxjP/e0ifnIYWKaTjvTq/UwN+b8bPqfCeuhnInqSA06AQCOz+5v/1nF
UdiCudGwGVeWSIEbBWzGyk3ekhDu32qLpQBX6l+mtFv6UKGEv4A6VBdI8PMG09a7
/Fw4XURJzgVcMHOg/a7lG4nAMIcySeylLj5IFX+4YG7gKvvfk4oK3dKnm+L4H86N
Jydep9zM69Xef5aPe5cMFzK/YuHAe3AsZOaVdQPrNZRz7sqtmafA+bpMLP7taoVJ
7onqo62fbpQj07UrpZdHYXw3I0besvSiTCfU6lwtTLQe+spqgNl+DaWVMNHGVdT+
KS9zsexlKjYntNMcvAqW2Ok34UUkqN1Ah28PUmNHaF/yBFu8/WEDbDpPM8gDSBMB
LV8jONUFaPq6J+Lh8X+qR4G67hzAtAEPDgZSqKG/1i+U8HZufJpYJ8ptM+JKw8u4
7ht9FZ+7BHHvOhSzDPsuXIO5YM6bKqb+QDv9VczvPxN2oDL7tDuHCB1QiXfjVjsD
jeytBBXa+ZZLCTgOqCcmlvIE1ATuNU2iGjfgfvYdZ66WMKV1Ea1M/Gk3zXhFEsdV
c87FE0QQ3stkmKc7CSoIhcw826ZaEv5ogYa+79Oxywf2yreXVn2mO65A5q/2PzHf
M4TAhMebZhLIzRpD08k64FEb3ZdcTdNWC0XE6izFsCRuHpUYingie3YaP1oZuweU
05j0pKvWC4qMOZJX+2I+TK1ahAvoDnu5UIyaoj0bVpEAtWlqKFuYFDgv1G50ae/3
CSDczEo2D56Yq23/W3jjJl7+Q8aXIGI8EU8VhSaTVBquTbnpN+Dac8sglRp8FZqR
lJXOkQS7XXquzqJdbDKpgw4ynGp3ve1QLPyhllxiZ69ufs08NW53Z82tYa3Dqd0A
Hhy4I0cBIrvXMwlQzHELz1QDNtexEIiCG3kVJi1BE3VteCX/3NTIQDp/yrOcSOi/
Oo3jq8WQh6XO6+OtWKo927ZbMycqLLoWgyWggalyLeGdkvO3+6wUHJxF+X2014Zm
T8qBOeU2yvAzKd64WSAVpqfTjp3WJwENFSSqId2VaeX+XUPDoDCzeDSjWoGOAWbY
Oso8NPcr4J+SBht9eJxJuHpTmaZITKrknaVPG/1VxGQkrkIwfA8lV/yAqcHN8Fla
gnQ9QMAVheTBrU0Hp5XRddnhDxzpF8lBQV5gOd1QftS/SFLkkS07Q8R/gko5loXa
nwcjSmBUYI0o3T95PjHDxHnXMrzbCaLhoQR0gdW3DpniHoiPOH3ghIQqt9v2eP7W
TOkAviP20of/V7MkLMxBGiBmnW5GQKH1q26hJNvplNgXmwFgS5wfLLfFnNAX1ood
ZxjWSsuXpIh8bxntkioUvOul+MnCIXWJ5RqPmzhUX9Y2x7xRso0wfMb9jFJb2RvZ
SPag8kQZeRW8iztcZlZH3Hx45MgXB/VnLOPpjMxZbQdvDvinc/GNG2Kss85Xd4pb
Fn6KvJPNJcP4+lsRdVciKtBhngpkLHViVl2XmcC9g7kGGJ6MM2M5rqYRBJBH5YlO
NOCWYE53jjjOXA2ceD8MekhdrlLJprdIo3etrIxBgPg+oRzzU9tF9cM0umw4FCaG
//pragma protect end_data_block
//pragma protect digest_block
PhaPwo7JFfim66uaYGKW09OlyxY=
//pragma protect end_digest_block
//pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
j7nB100y7p/UQ6q8Na82mei0qeKT0/AS6eOli3Y3/EN2UvS02Y2zo5t7fATPwVZi
u4Y+3H8QM8z5Uk45AfIdgcqta7win/yBz50NoTbBBKtzxtmSBjm4jFGSC0H0tfYL
u42cWBMoH34DgbmXBR/o9kJxG3HFet108ePnKS2T+ElOKIW7dmjrpUVoZoDzZ97S
dkjSnwty0sDl4bJIp1GiwaWcvReEXgTFenu2D0fQU1fZp9A9QD+Kyev2R3U38s9O
BtybWrR/LNmGODAUOytLp2A4zhyq3SMpp8wV5vY/N0aIv5AzD/1g+XazDyDCAUtu
1cbPw33wP1gIqcyrf9/NHQ==
//pragma protect end_key_block
//pragma protect digest_block
gFcUJW6yBMtfa72qONGD/+8Qhs0=
//pragma protect end_digest_block
//pragma protect data_block
WToMlZSacAZY4hQH1WWs8SOhzCLfoLvp5iRMuDA/TSHNhC9DyisIjk1c1NQP/G/Y
qtt0+2MILJ/la5yRF+tq18Y081gCKHPEIHHnnfcVyjSBnIOOamsaFY8EhezPXQ04
I1PueeWJ+2tv0npUHS7+nJP0UGju+kHdpTrGbU6XxRQyc8ua3M/xH/FWkmylm6/M
XyhdJyi7oSsEhyOtLE8y9jN413KiCCCrjGPMOTX+iCiZ8FVCoNJPie/4bCpoun9k
yz6b7eZUfatLc/V5eOGgiwgZ0b5ni/EQeb48IFpsqu/FH5fgdxzWBlibzOa4faus
BE2Td4z3YeZstxK9sgaQmg2KUqOxpTyfzySyUiIES0OevYuB/HZfHL1gHYyQiwyl
hxCSodY37Qjd0Z8pKh5LQ57m3hNZoRj8eVdJDDVP49D/Fip9gbwCkTm+0OCQhBUt
TgeUFJM/1DdWt4683ORXratW0ZxlSVsm67LoVBlglT6llTOkgej21vTbwooS3fCM
PGHgbo7JyDTZUNTu97il4pD0m3+m9KPQ1JuiJ7ewkQsLNX7z4pmpSw5p1+bLs9ZQ
zEL1CLlsISYZNxPeKYPsJWfF4nfpOC0VmiE+86vHOGT5LfX2yogOOpBurGpO29FM
owEXiiayr7O2Sz1RM1CAsxO55INyXw9NC7bgvUyAT+tudGK2BF14SaV6rn7Ndg7K
j6dpbZLQZMkOHXrKYLqykNEXP/h/EjQfTU3vIoY/SWxHajXAqDqg0LItTkl4V1nJ
AjeLwGoQnxck+JSncO+nAJmth6L1Se0qwoeTr7I9cRU0cognh/4muasEKB0V0pFE
HjPl/Q3NC1WMLHZ/x76YSuLtIyJ0Ur6yqIDRK0Mn9FQXyM8HN3rTENOQZN/cu7/M
YK4g/hefYRqbdbP7Fb3OpDQtNAYFVN3PIYeGdoDPmRzh7I6tkzARJitw7k//zrdq
vUhWoxEVebz5XjmIB6fAPtM8ijWQJc7YStJ17I2WldmR2IgY5Jk2f/n711Tbe++8
kzvEA82iyH6mnrMNiUCcR7zUujDwe9WZHmF3O5vdlIuschwV1oLk4JUroWW/l+q0
CXw1rjJBAZ3Vvc/D8MEHrvT/IwHpKDI2U7zpxgcOV6vmCvWOnwCOOO9MaFRKXr4m
fEiPDK0cT5uu2PlUBjx8ktWMSyD35fuU/WhjNq64B5eJZZwJzTKlZSPXSNy9dxof
3F9B8qwpooHtMUCkwKuyRb3SAuNvKz2XO/4kRALKvEmBctW83ub2HnfkAFwXMeQT
xOdNW+2cPry1jxRecyyXau+sskOpYuwu95rUsJyQVCsGHQdJytrJy5Px5MIYMcbj
plDL/i3OvJAQ3WGbH6j7121Zi9pPZ3yzAsBMAqm2jQsZPPrRsDCyPXgra0JdYBNF
MVA/TV4mSWBUMlGmfiEU9iQZtW5r0otkRUdBNdxlZYfndetnhBouGXOdVZo9b9XC
7nT9ZEFyFuUp5W+U4O45b8gZyqAVOZPMPlwrwZ5bwvHJGm5igmbf3wbZhlUZlCO2
rfgC/f5RqxSqUc9rRk58mi1527EKKgcC9YhC7NIksD/YU2GZS2FwaTh+Qef+g8E1
j2+xlYrAdxOqGGaAjO9uZ6Io0ie6ez9GoVGhjfhY+o3clgwx/MtplMOfaxNlCmdW
uvp50lqR+f30rZ2gGgrxp0h27oq23E1cbf/BJ3km+D2ltT8e09d5APq2vWfP3fwP
PXWdPOKNOp5YoxotEJI0Gfiudp0ZQ1mnerb7Abc1b/pV8P5CW34bF8JONUM3npsC
124xWKLLAam7ampigyopWXgSZnApb89l+cjH1gaiUYmov8tEl4e8JB29ftwz+/Gu
+6C4pvdPWHRKMa06KZWovEcLq4Dj9JfRWTpkQOt3DA46WJ9KN9o5XNo5htpbqh+b
XZCjJQG8O5Je3lWrio0Agqib5cwy8GfBdA4idr3Khm642ZX4n0QotJBj4Qc+110d
ponbYc/ZVTO9GDKJWbnt4pkylvrTxf/eveDIk/8VJr3+72HmeU3bpxOSttBhstvK
zuttO0ub5ZZz6VR+AKeVaKUKf5rPYaUsRH13Q4lSoAsMTso0AGSVbqaEzZYzAmC5
b4/4N+BjBNkcIhj7I5Aae9T/8zEqE4qgqK37HC2qTomE/pDhGkBX44Qh4cY/JQN5
sKvKb6AU1tigBFmbPPqKmHryEXBPixynidvmisfAKvQJySydmQUKkmqh8QxaODAu
PAOe9mVTxFytHDU+q8dhYeFq+gbO6i8FZdDOsT2je6gy2PRPDoXO1u7YKhMlxc6D
CStgabNDHCz1puyqWISQu5OZOk/o2v595nguqFpaB4fUJsfnZ9HjVrJs42Koo/SP
4pHkD/wx8spTLes61C8bZXOTAtE6DwLG+knNxzoMh17HY0PUJIZkA7QBmc/8kD0v
5KxaRfLQ4zZXP3NXrHKGhkonxdUfokK224Sikr+LXqnHPRIoF2E13mewHnU+uB4w
5kHVB0rW/P9V1UxUlvuOrTA/f9JU5RTBELEF9hcve/qOe6SwctpE74oHJY55ClGl
ZBq3aFX7BHIwB8vkOddkIX7b39zPZzN+LObE9Nl8Dt7wVyBVlt+ewTjvNI603cyu
O/4qeawHtN1epV8LgBMmsZt99QLqapTNFar4kkf3VbfwUiiKOVBdem2HNZXldY9v
a8QUk2waXz8zqALnQ0nk5mSGoxxPQwSiCbsvCW1awVAOC/+WD88z3UXLZqnehFG7
f/Xy31qi/bADUYBJYP5ESYmapaOqG75pn21JzLVJAwzfZ/znwt/4uO1S5LEi6XmD
L73OlB4eRmF38fJmzxMIxWqZRw2IwFsDT3VW64t7G6bJKH+aGaKNKdEZDCspIPPC
Pi4SEuUx9wy0xmrClj7kRcnG2zdDrQ6bupZgU7hjuBkVLSXRHUYJcsQByvPCNz04
WipH/NBYi78ibzXch1D1/duER3t4ckYi0O+S/RJOVi5FmsIyat0f3wGPqpJBftcH
CZnvlkDERl92EOgml5+bJViuUtOTiMnx5tO4nqct+YT4N2LotxQVcg09IjNRr5Sa
GvkOMeNz6SA2AMjZpXBdT6x5qmnggdwYbL4benq7UjdmlgYvnt4OTpW2UtFeOAD9
7eJFPpqXDbOplskPu2/ovkPL3MTSjH77FhKEXi1U1CEu8mLIs8me+9/37TwI3Z0P
GzmTAxoSfCLddfqF/2BMCHhxPJnQb1EGwp6fOr0pdYidFK9GGopiEMWk/QvuNx6k
l2vNSUxUt34KaxQjQyfqAldT4FXfgUY3hp7Z06ORrTDFxUP9Y9Wz+WJdlnQLPykX
EMidXN8X/SzrGGNdbx7Fs9KMEzzKIlK+81Apuo4Reur6UifkE4bRWAI1OWD6L30w
X19oTepGJ27iSIyKYg36jJ+ZMba7u6HxA54qrlD4e0XBStOF3paCXG5XTKPendsz
psquQOy30mcZDEdZmTe+1H5Th6kTcIcLd+vOiwayk1zYFJucanoeiU4s+Ec/gTkl
5wukDVrSUKgVnX2EZ9XLzmO3GGm5E6CLB2foOgNtlA9IeRCPtyvj5dnm2reiEr3N
fmijtw/XjgX4dcfQLy5k8VwAmWZWFv7GM7JAXFOp29GsogC/A2u0ivfTAzQGmk9D
+zTaB5lqtYcSlc5Sy1M8HG2nyIzm/2Ee/mt8KUF5omNgg/AJ9a2qcUZbjyk9Mff6
dXIWfx+PIGb85zXqk0/PHf/oyV0uf65znj9dr2nZ5qa3RZLYUzoZabL8V2dzpmhH
hTUGaT1D9O3twkvkXy4LRSGsbx+WPUJQcEFHqtrQV9oiFggGL63I64fiWIjjhzeR
U7f5yu0H/aKyIGxlriW+yXsQGoYyoK+AxgFHkU7JF03yYpTENkcZAtXbKCzn5uvA
g15gK5+Fq3Tm41DSzjmvFOKfTzmBajjHZ/+AJcVzv7wWi/qo+lRA/wvLc0EXYhJp
9Fpor3xA9bJJx3GJS0DO0z1IcwyUfh2foPTViSmD7JtoutoCTI0XOdoRSi2aE8ML
JId4OGL7DQDAnA8hlC/TshvVQN1/BTGGXblLVld4tK4oc/UCbH/GhaW1n2HLByRx
9ctBXUQRDLAAQ8UhMpPfCOBCq5F2NiE+sDingFtqJyWKGu7GWT0AQVpFJMzUd1n2
19NZgu1faBkfVLassGgLavIYFIiW73t8DdOz7Zmp9XXFRuqierP2TMoGDK75a2/F
R0oQR6LyULnkFAQ2lzJPtAsYf50RH080thXk5KZh5ibbq7AF2rcwqPyovn/E7ary
4G+9VDJ+dWYLM0XWFE6XxM9FqlbTkh2O5dd0JAVEVhziowtCnZzXKwk8c6XEPGyg
ByqUoJeihe0f9Cz3MN1gD5KzLROwWsJQVBbeEJhsKNa1uR1vp5Glo7f6bIFTwT3+
rt/i+T0LOS9NXlwHI6bgk30M2lMM1VM7X4306dXTWSeJMCfWbM3x+oQN99Z342Ep
m7DOiiJPoa2ubZHWBS9pPgtVUfB6ayT2pbgaNcB2fIzXHNveVIsFT+HBrsvKoCzS
eleFj5bfeDwvWTOoLta8a++HLT99/L5YOhRjaJhrH1RuDkRrCFty4JFsyPKYA+Fa
jriAQmTJbNQfFs7xefLBgF3a48/u59Ije56vusyCDdgyaHXiJVemZiPgrOa3AM+1
qeO4Ol0nZXoSwperWHolc6zH9lCQRXEPJIlNj7+wMv1YfMRtIW3uI9JQZiTrzqY4
NYK/0FStDnUbMfCi/6yKcPvPNuegqUi1aa6oJqyaT+xgylBiZj8CKVfOmFLHFozT
T3HNNjno21JZvxc49bUqGgZ70TvvZlqVhw0OcN03ab8gxMEGaAr/eQlMMuAoEdgu
nVVE8av4qumCrLAgstsS37qEz4kuLz4zQzzDJI+BXvAXjACmsfFasx4bImnKg/be
rnQvej6ZIIpkq5Ujpjya57LMZ3JE+aJzqFNVehD6GUYOt/ddUIk756ttclvSQYzS
2vikjC8lcUWp79qqLSUBXqZo41jtc/XB6JNh0OejOJINiBhbg4AO09B7T5K1j3Oy
iveFIfqnJUNie8fSgWaeSPDZ8wAZzxUfK6huVSzQgDHUGGTOh7vT5vzKCHc2PFSP
0Ge+x7GFPDtfpNmrpQ/56k5Z9Jjf1Rg1vf7xCcXws8yZhUsCVB8glEI/kam1anuo
3s/3TzioPh8H305iQWID2G7NirvWIo6SSBKdAeU7NmMUKScZNyKKmSsAzrgw1J7r
lBiCW90hiGMDv+082XnBLTzhtwgcd5c+VRWnU8CLgIMA3qBA3VIUjMzylog4Gghp
o0KurSrCHbrU5e7/6acgoZpbO3CT0HRoQKZ81QnbwKmhdikgglSCComa85DRiYX+
rWJow0XjpQwrAqyYHRgUPqBvKylsJ3ffEGpm3FH5dn0Vwz8W/STbEfh4tDUwVNI2
/VWq3qUIFnYx7BkcNfL/HcSY4bdO+L3dzyhy1u/MsaPJ+Mnh8QPHHkaKCUC4d3Oe
Mf9YyAOZMsrlo6rlxOdGHKIt9iGwfOXoj/Q4LVU4KCSxio5rq3mvyvSGW0pq41Az
suUqgAUKl0zJSAX6U9ah1QzZr/BijRQULVJydIYmfBAN0XllsjIJcm5rk734m3XW
Btd3ZTmSf173VwCQaEs9wHpLnVMifchshCjBvj52eOreUwBGSOs/9ovL+1F3Y4Cx
Pa/L7MGt9JKMqVBa7GfzITfUL9TCg+oCiZ7hF23mkHlQ/RyTWw5vSU3PPHaBOSMI
y/9JKqFkxig4mZeiNurcPgNMfsqYI6Q1Txvg5v2KYKQ3F+OUqHcVEwozZRKH1CGA
vLGNmr4PJRrV1Ol0yYfLReoLpGA/yJIvIM20QW/puEV+wN8BcXJIxCHQ+dkJHLaj
PJAcJKI22HeCCcgqXvFICCFOpYM3CqmwQVO5Nq7+t5xz8NEkNv+JL4uHWbKejtVd
AZHYfsAq7ACP/sgX4d62QGrvIARkBKjOONzULPZNATBDedX6n5NL3iHEmq9X8fh5
2PcP/3CaLF+nXLLN7/EtDnt+toNV1DRbhZfvfD8CiTtT2v2WGDs86WQt5ewOOcfM
MXxNW/aZrQ7OjCT4K2a3b7uCoKNUPNUaof5sl45wslu5JIbCF7WtO/d9ymGUiTh4
1GrnPFCdrMWpm1t5aqDHnwNx1FQ7v+Xgij5UEHGneEfq4cDxVtFPxzMqvpEVmnEO
E/QGHmzpI0lCcV3AqrAUBTH3ekuHaRxhEBna7oBi8pSn8Lc7xHvRZuM/LTPMwQYk
Zq1w9W04aCy46ByeoLrGTxPcZiEyxZxFFTikLjQvSze7rDYDeB6KqRMtu5eLpbDF
cJt/muNH1RS5XulDAG6/FmipbGVTunxIzLeXix6k+9sei0AVhk4XTSmMd/xr9Us7
nInAgwmFoiGcNqBbGl+K7Ea23J4fMZqMwv5vYcrqLMRUWfNNL7hjQW5j1LcY/X53
cB+t1en9Fe55yluIwlY956U5pX2OUcvRnbi6PGI8V+jRCFbLQOAE/ks9nGuDjPwV
x+EQ0zg3Eqj+OG41tBH0KdG8qVP4YsL8l5ibZQ89nmdb5ZvU34E2QBk8z3wsgjOH
hEhuKT4H5SvOfklJcIuxlJv31D+QPx59W26/oV+CLB6dtLVLNJmqSONp0xxgwZql
UJ8zr6QqJHB+6XHaDZv4sGz9ixDipcw5i5ttclzZL3VDIuUdixpIaeMmVOgygcVS
21JzWB+Nl+9Pi4D+kZsLZG4QmWyusSnHVcNYWp3qIbRvB5ERTLHRMwm87YePBcO3
/V4lSsZKbUOlh4K1JjgGld/RJK8PmH6E+n49MUQvBjUTuyTUGn4W+JchpvddOdem
XLmF+XIenEc9KsT21ge8Z76kaDI/sdBsfM2vhV120bzBGDXseu4jwSCkbfgamDvp
9AiGkwPd1LxNs2uqA2P6YRWCOMKAHb2N5FoWL8nSsWrIbKTbs4vlCiqTkGhgK5FX
pCMFRhKrspYGV2Exhr3WZORc8gaSC213HMMyeoqN4rRGbUaexZpy5usDXv3ZPIWF
IuLwBNkH4e4xXZv+T3u4DEfAgNJzPUBrGLl03X0NEgUem9RqXqjcbb+aGdbwZx4M
XOMdR5YKSJwYGEiHIhtWqxpmyx4eZyYN4Q+q3QwYIbT+jK1y5u6ENg57lN3Qs2D8
Tucn0q5u28VfTb2X6d6pw/RZ23/rU3ODITDs0M0bsdfTpcUciXXzZjGwcHXn24rN
hFKEYMcDuR3hVo+HkJI6twZTse2iQmClLi/hJLW6YGmG1HeTxROikFeq4P2XmDf6
lW3Wni9x5Q1CUF4pwRddBgClCSe+W4Gt42WKvuNNw0F5bsC9sJsIbxfiiAANMMiP
ptObAKTpJo2Ote0XXnLFJVazy0ubqLo0zLOwWC8/7abL3iUqZ3/SwggctZcRB4Ex
flkwq6mB//Sc4S3LRSTW78LwSfLOIz/SPfj1uGhx3wO7OeBvcCa733WDh7hmVSaO
9s53B4btO5gRs37w5qRotDrlNN1E2Fr9lfKJIxQ8kZMrT3RDd3Jbl5hzcFz1yoeA
SvpXUnjKs0tBKe1XENUt4Pm+qBEmWLV90LqgIujWYcGtG5vvqWZ/WDSqSgUoPYdU
xBq10dfKlBTKfETWlgf4F39X5Dg6/KZdHI1XFuGgVO0/WyUavL2icaLdCYbOlGhL
zdw+8mKHfO3eMHm5AwDy9fKQT5xU1yA10NzwiAN8VM+K1cPlqlZWguRbG424Sy9z
E8TNUKnLgoU3Y9UWj119afuFO3Z9DN1ITb4Sf0UgIOFPGQMfQnU7f78bYUwszWL4
QnUdkoiIilp4nIEyk8om2iMoyZ/JTrOhHkIfziAw1Kz5t/QxTxUhcrnOCsxtsTNX
ixQeHyRfgfjkPi4hdUn1oWfAcXVhoqY8zE7WC5is7dY6JPcI9OS6pPJIocx82Wfi
RGHashg8xcp2JwYVPEPvOlSwIrBGn8sxYPk42BPeNsfVQmXaYwGXQuDKO54sXc4w
66TuuugKWllmi0wSqQSxcjNqHvEPZtu6xexsDvRM9+MlQQ928cQn3TAMyua/L2hW
he9xqC0TngFQ4bMecsHVVHDlspUFdMr7R+ru1p/0MwWg+aNYSldyKjsUYj5rUEqR
XGI1ia31iDh7Ppi3FsIxV2H09/W+pHV2KgJtma+SD8oGBTrvYUpczTQpEvlPmCbo
ZPOoH9M3VAtMSSO0XnmE0FPLQsvauiy61o4nSr8UhrFrpwBb5oiSz1F3kb2E2El0
3r0cMguT11Up49Qw9TTptqeqd+Vygb3wrvB2Aa48cb3tr3zrIuUYxnDG160nyMKG
0aG08sprInvhGK9PNKsaLpPY52sbWfMhip/iAcpHtSS0zpARCqyQq/jUTcmCuiSI
2/u13MDFGXz1xN+ZVSFgGxphwvOLbCNQm7xkI9hnAnqtxM6cPNKzmaVhk4dwD9+F
jAi1trbsBxF2/z5nJ72plz0uX1j54EuOWsoj0uAC29j7//358rflofczy8kQ1iIl
boDFFRd0z7cM584K3AnsxMdG1fvQnYhSy8tfCQuSMhSEx8ofmL1teAJ75dWxyTKC
YQPrXR0NowH7ClgIRdxM62kr3Y3EWj8hF8F9EBSV+jgzPMxM0BnJpI98/7Rk2ywH
NLxPGlVoX0bFkmJt/rpQLMX+H1dWW3SAsyAMZC30J7L45CuwHLpgTRqzHRlyJJBx
wu828hT0Dhnsn9Xo2ajSIHg3YkoRy4Jl6g6s/JOO5YTZhQlkEnHHbgDEg1/kQVic
Nv153YtDhDur5/BOMIVBcJMC2o6j4NOw2P04YobGg1k08lsvVQFTViiZF5aIK/p2
n0Xa1KTNqlusn4bppRf/yL6cBJSu/RlhtOUejEpOYwkefYoFLJrYLSo0tkc/YNlA
7I3gw0FCTboSPyAWFlWnEw2FnXCE7DvVR/mbSw9czgmq82GQipmT9fSV+6ezwXHT
TpUUj4V4dwChSBjLKDMAb+gFKUMxpAtuhcVHYQb4cCzHUMItColX/9pDOeFYB3r+
v6kG+WK3YvBiC11N2JK0zczc7+7xVlTKs+npX/ixutm8MFkHzcvJZ7A1ltqNr2Kr
+h8PWMEdi7toHJtI6O5agZLglMIuET87jb4rn5EiRuOmZN8TwZLUkxqYFNBRcBIv
vmh905H1t8w2cqOqZoFcIyRtIBJyW5GsypgQdEERoPoPB6sxFVGIN9gV9dsruCw+
h29GN5/BDTfuBuhQ0YiLqd446yhx2gXwly1lu+RphOQiy0W+V2Ro+UYzD5FcYdiV
WPV1BfU0PSSpAe3Ha/te0Hwxd+3Z8C2frT3T/lJ1bQpcxaaxTGSa/1WI7R62YfN7
MYSG42bt2xrSEmEPSsftLGAkauz2GNvUtlLKV2JJPyWCeUewaqKmuvzy/VWWOoHO
CXyu1kYMIGqu5trU4MGABaPgzZgRRxOtVHaPCCn0NOFz6nrLLB8UnYXUxFl8dSC9
L2Nm71doI7Trd/8w3h6R3ExbRirSt5krggdx9nlzD//Bl2S7sVbelPlaGmy9X8Kd
PUJ0GUyQjaPUn90B2mq9yZvvaZzpzjwXxq0sySN4wXw0mchX0eD9wGRefyeeVGVZ
PxTVGSo73gGp7kar7QEif+yB2kPtBytHfBHW5riC5QCFT+KJ8I9SYmVBeV/QErZA
b6zfU7wr+xyZ3ZPp+DCvCei0UADqG2faqrhJqWwodWzKnTLT1WdoaXFLUqfiFlB5
geBunZxjRYHKug0XJ/lWmyDvI7nJpbKjQo7Rc3S+oHSRZc1iWO31p2yOn6xSED2a
OPm/4XOaFPwZnx9jc8niLtBFv/WmAwOAV4ruZdKUwTf3okvhwMvakEPox4MCtJE+
ppPCih0eG18i0vv48dxiPRC/m1gzlLdTbQwF4KRmTg1VKkSH8jBAy076PXLSIrir
AwwPuO7DsFovUqU5XlWDHb9ltv7ViuS1YvcFh74iA+wOJ87pPAF7RmWKGR2n053h
NVVlYzT8Ex5J7RFD8Npv2223XF4mwOvXTUHUVw7UwBEccHFOcLZhL8p0Ne0QSwol
fy+87xa17TYDy3zDRPr6jO9a/7VnaoFJ2qFzDTKqG/MNUOZsS9Dtg9T7JpkDgkCh
uqulIJYcAJnMgkZL5AyCj6Xpm+dkNMIs11YpPX/jGbk1jRnR08mvwzTd1GZDla22
yCFBaTWr0RUrqZuBm+KVmZmj7NIXVMxD+YBKKmQYw4ho/hnKroQjQixBYmYgtfP0
wRVsLoF6Ze74UYYliO7IdrqQ2H9Bc3FRgOsggcb4BmfA/0xVLVRFN+3fkVaOqr38
ZRHgQNFWGKUpg2dZ8LKUEUMYOpDumA/F93D5Dzt00jnPv6pct2KFt0JGWglFX8YO
GlELEe6PRuAjxCWVkH4QBPwx3tRhnrVyPiwLZHOe9OZigmhkr1GhRo3gLoQWqqEg
bPfgYLaPYwzU6i9znRT7oVAf3LEk7EOWkQ9w3QGf8q/nJ4PpcbcwTBC3M+ZQ6IyP
vl/Cns7dGhiIO/6poW+KpvtHI3hWbZJa9SEd41TbKHaai5CbLlB8eL5E6XVjI0xM
gcqXj1CH/pJjahJPwb8l+tdgc7XUEggxpdF2WERolS/xZ1Ov2NU5cptAT9U2kgo1
ealS64giEpvmlMvfArieLki5wrIpkLMMd2hGU0j4O948l9y1pLt+pUIObyk6MZ7T
umzqxxc7lbQVKg99pvEUTa56GBu0AhNZ5NAqrZ0+h9T/FwWaz6jlhqphI3euZOJk
x5utA5VI7pxvrA2Jyb0ErantVFrbbOMMnoTwP5O+PCtvrj581HfX8aiSSqeDx127
z5jG+HvJ/JNpIzuHmnAEuyzDWyTUwM6Tt8oPqF453EFFLJR+4YoNCCqbglPe1S99
2NBlazcLkUpQ74VlAjaPYT1CdDmdA3xwK9Fp3sAIPjnF+TynNP5Fel3LhQoJC/2F
0lmJn/9ggx//PuetYvV2xnkWgdU8mMuj9ccXwL3L8TzvrvtyZ3FKayKOYQLXFJlm
XBSjv34f5SkEGKYGKxAZZNSVminb9YifB9+PfcgnC8tlTVBZApZsHT72gVFG8+zI
A/F8VtBtOfG4RDR5Di7ykjhtRc5Se2f8CQTv7W3dPoIACgVIRrmQTF+JrGj+FfIn
XvhN1bkkn5MJHJF/YWUIwXNEaey/PRuOVIx4nSLz16TB5FGWAvLGwbUe2PkfcLwE
32bXAowM40OzY1fzuBT8o9WEaWPxS/nKiRro76UEsAdlC/8vj8/J0dLBuFWed3Ii
D7jaE6UM+p05+usJV1D08KoYfBXhgXrOoWzfmwLe+/DTF+WYU7IRHnZIxkNT5xAH
30lBjPRDeWLLfeJtds4myHZjCXSreo2eTALqygHJOKWzPdxgCralXlQ2ece4ot1W
LXJhZVPc+/zOrT2LezUy6uFmcyTM3uqmd/V1/DhW8i+JZC6142ZuFtLyyUm9SGrN
fYzJbgzSqpPXsN2xwEPfXcKW0NsDCqDcC+8uvMQNMshiymvqPFBcS6NUSOEcRDxO
BlWF/Bk6SKii9V8b6ZyAg6ET6CgbXBS9itIa/7mfk52ap3GjrUqVfmHp7A5+4h6W
45DshAHZp462BpWAq7ST9LnwqMHHaiwhfyqvuiTaQbtPnUtwpkUR3jOLpLoLq+Ac
Tl1vClMcBcPQjNYbstihC9UGsEn/Tls76ep7eaSNkcI4JT3fUbjAEYSAj3P6vnrH
J6wa2Wnsw1daZUXSK/cmjjKMdGJvg/7DKnFmTmwz01ox4JkVMiM60rlkgyPC2Lzg
wYRfPEqDC/gbVrBv6qDaM0huht7QzNkciQ1HNjQbh650U4hANxbLeSm6HAU9PDoL
NLUGJPM2FYw31TBQzfO3ZSiHf3kKjG5gBGTZXHWqeQv5tVdSgCoLzeuSISPwExV+
P/VrrmSatPAsqDYwNDfY7OR4JG1v5JvAaUWUsdc3NP1onUKHDV8i3ibgS5Muh9wM
zv/veymdRxLQit1GxHE9bJo9LdmOoE6kNKeauuMqW7yKKFaQYVA48E7PKLMXOMiL
C5dIBFuisdDv4+Mcf/HASgfPbkfby2uy59I8mt+t7WCB6o+kRaxXzpUAjwYEh/90
/jDSLjs5+ByW3mHU+MWxb2dOzN218mJ2Bi4PMt+yBt3rzdlI13Px1R0ZBxh7iPmH
A8kGZmYwdHV6lSpgUwDZ3qmpyfHv/+x/0YpWIJtH1zpx4nmZa7yJ47GTNLz7m0xe
M3Nt5YX2aN+196kKT0c6sDjfivyoPyMrJkKuuCHvTQQ+a7bOBAdyJpfnNb9FYgSz
uJS7O4mSN5tA5ESVmRwzvc0ZKOt5v41x5Q0P7J3T3hWCopBp+/ZZlkXDBA5f5k83
Q24AcyGAzi5YlMFZBdILqX40hThXspn7AeL0hm7YDiTb+ziHQQMgT3soFq1FRIHH
6gUJA1w6u1DKirPKnmLzHbitGZs6X/hwZkkS8BvGqYIDRK9QyRPWvwtkGtxOIhSJ
XHMSE192iB1eBJEj6XftDMMuTGqNMZjrw3Be7YT9h0JLvWadefYotmBnf8hNo/GB
+meocL89RrPLAZkt7alkHfRmDK2sDMGcXoJFFpKNqwx2QnC46RB59Wfsc84HBtll
Ca7chrhQg5yBORNlDra3QNyMg+twpVeJrbCr6/k7TvFVxV/diP2doY4bnXG2ug0v
5/zUe8ZXEOl9QQWf77Jxhle08lVD2GzLJ8TrB3/tDYoBR4Fn3vsik4N9LTtTt3we
YAimIx1Af1SQy4QvUnSPXNP+Ueitcay4YAbWYLlFwArEPqaHUGSalHr/1CtQEgwl
y43ulG3s3pmcE/nLeGhThzRYy26Byur81b2kh1bqZPfqMUwSQKkTVxc4OexYhuPb
Ktrx6DRFjivCLNXDrv4IKn+hwLWR+wTmBDKbr51mJSEaS4rbz0gMIxN0I2+u4zQV
wsOrV//Hv2niTCRwVLU1yCD3t+YglfNQdT/RAmRsIbiZMlomGPgzsNJNgk/KUv/0
nbmD9Dkar49l44kLBHRRWizH1TBHkk2d0FVB9Yb+mppyIiXPGozNuSyY5796bdbA
k9NZT+MNjqwsE5IyF70lrocgtKi8viHevBURkbBPjpmpkA/+jxWTdx+GVdggrAlQ
IH0m0jAFjpE3F/Q032uh/ZLjVviSgz90cXIfHgNQj4bA8OTIphx9cTmUtdx/DGRb
pkdtFbq/W0y1rCeqQAAK0gF66JximujPJXWLAgt2yjQZaEVUqGmDei7Z06HZt388
+qv9S4pY8YvhD++xBGtSoWBRzIE/UfkZKxzG7KUHbj6ABmorwTzus+dGUTyKlnDE
5Rkyl+LrtytvME9oDLtE/TCmEa6knI+/piwN9DnBehBKO6qWjpStuSptHm3xX/Nw
phxzrEiOHMjSjp7wBOfJI0BJO3Pk6vv7MM8qQfXqYgEyKJF8vLApRs4Rby1ziiuH
1y+AbL63Kkfv3O0+K4r8eXJTqmOr2uO8+jJvSHf7C+WJgGfsnkt+R4LaAB/+U0Ew
vzXcJkQwf6AUOMKpad2qGvi/F9dxD6g6n9fISszmds5+T8hwnSybnHX+AxecOYnz
c8gbieDdmmGPSU/0UH/ks32f8CU4TDGbj6LE9W8FfyUOYuDPs6rQ/eQWzCo4rti1
Gw8HaW6AS40B/K5sUM1lnpuw3L3VD5REXGKVmfq6yqUgc9/cGYekTumEiisKQSze
2+hAxKTBIcN3jmo+PjhHQhUn2Utl0vgTnYGKAX2KN9x9QNk1o2p+H2V3Q4fZ/vb+
8Gt5L0VK2GNVYgRnMcG73WZgGAcl0N6pviIoFySVXrTQw59LThaBoboBgrIqTjmf
PgROfFzmvb3T+BRXSmPRzqRYxdaC/HFk2Q/evfIYzsOco/BDUIi4t2I8jOT0Ybqs
OzXGmd6UKfU4tKUYNwxg6FSniawgzcoLIbqhgYFb4wRcmFrENbFW+7etiHJ/7q3V
rC6QVU0snkAb4385vZoUsgimS7icULs6yuGAvkRDBDKmC5KA6RIxqDcrK2PoZi1D
8/b2/9EgtD4cin55yUUK1wzS1wmImLsAA2Qw3+vvdFXR/jg7RYuowrHD1LaMf43j
yUfw99ea2uytxKbcgMJxKaS3IUkMOhoaV5P9Oil2MVwwz2DrR9w7DjActtCZoveb
qBBj69R7ioilR6EwZUBLS/YeC52tHjYaYFC4JXO8UbwN5R+YICQGD0WpTTa/Buo8
Nl4lRgOhFpPpD93LYvySDYgHhMDZCRk33mGIjWdketpyXNBhjLzZKKh3xwuKY/uj
+B6nY3NHSS5o823pTivEM3+w/lWJB53UIes74Q9lmIE1nAgKlcpoa+rdv6Y4aCkT
yZ2sPHHMHvnBiEQ+no1SiRE7BYLNK6o09219INhO4xjn6W54ww96fXt9iFRTu+he
Q/rpc/0dtS33Oek3OjZkwC8JP71HqLB66oUXY8O9gRzTLuXYKNTEuhZnd27ee7Yh
9IhRcMJ0BbfET1mJODvNRInX0VBOMVkvqWqgFwqcqqebmRZCpOFz6ZJU5B6oCfaV
u+fdZUi8QJSuiurFJldLWcJeTkPbFqVjVqxSfEnhgX60l4uEJbA0pjQZR9el0WHZ
ehvlpB+BOyB2WgI8Swxi2s2v8MjWUw54GYtHhHGuesfXy4HG0aGA8kIeGfizqK8R
e7bDRNsObVrrjzknUSszYsIUc9TZ0rn9Ytkhd+k1cgZN7vjXRo2eHebKciJx6jKs
TwBxJmq/UXbxRPGJ7v7T6gNzSCFoBI134yjpu4ZIuC3zBrqRmkwIACLwGBsRWR2k
AwiHf9HYcfQd8C/kaSMGuVQ1L60KtIUwdbFGv7Yc9bE9vYvkRW/cg5KOFB/TefN+
KLbHtcGxEVBQRQ/kglwKDU8VN7hGX0dVGUQ4F7qCCZpdUBs8MKIfdw+Cm7/cG2QA
KetWge2GT31oDWsu9ucRRC9fZ2Ml6h9gI33tfQxSz9EKXzR1JS7ONrGmSD6RF2I5
nShelGWfFajUZQPC7HT5J2GkSx2zBAHsD08LsRr/Mk+ej+Iex2hvz5yxcqY0dvmu
p66JCGKtNzSh76H1SxclhmcqCiO/qp8cJRLED64gpPslDoi0mJJPjdlvL/7h9jW5
oY2ry7DcBdfK/hjns1drOT5s8/lcXBar94uQQDKD1xpbP6Lp1AjzXQ4+O8bGZ9rh
wo3AO4YfTeSDzHFegS4h+8g6WQBxb53fGS8xICOojjhya2+VWstzcfurU9a5V3AN
9AS6B8lYJmESPVnD83elspqkulaBdpCWtG6ps4e2TdsfOtmpbBRlSxbw6EBHg8y7
VYEGSN+4Ep5BXFqK0lKNcFH3Cz+cb/pU6Sd5aDEB6bNgU5eQ1UyOyjaZEShangca
JvT4TGirga3rf0dhONZN9jYnc9AxKiqg8wYUHFyIDjC/9evD6DSTD277+UVpehjv
yGDb6r1LSMxq6pljsexcRPgqKk2zl5Q52W7hQ1fqMPZATtV4E7cgk9DscVwvt0e7
mBZahicnLji/IpnqL8B9uwm90lAnZary3PBAFnGl0xxRe+/nztcwih/Pab6avDuI
g1GMZfWElwGIKRki7/9Oi0GWAxE2t00zgo2r08yZGNA26sOG8RAAL+j7E2Ja4Xff
abbbk52luQkTtI+n66uFgdue43L1L+cP5+2oUpQtKNB6zEJkqsSSAd+bGECAPglp
MN4XJGMQA2kU4F7DX7EPVgDVn0IWbbrDG2pCVJ851lSBtB2qHjX1Qf/rQ+Yj89/V
7PbqlmWREDOXRU6NJp2F2N6EHlhSiV+VuO4vDgoDzNHvzJ55Jcy0jhPuUozBTTaj
SV0/VRYulNZkopF8BIw6NZQFwo2eIJNXGFKzeupNXZoOVEEdbKttARXqbTdOiQkv
wSYVgXdRFRm1nworX08JEX0/wSC1ssi/G5wNCa+QZXYCXClHTOzKyTc5XjFSy/6D
jJ7CG5B+NCcKCBcpC1fGKHGQ2GR0ilIhcsmDIcQ6We4WmEX9KYs23iuwSYSoi0AP
mmgA4ikPED3P94nPSaafGkyABw1svePdL4E6+sZTg/zeAKDrsWBab8PXj3CNm5Wc
3sMFfEZzDXvVPaZ6QYtmJ+90qmxS7btjEtjVXL5mZ5qKZOsi0T0wGWbMvN+jDc1d
qd0X1HLuBYwHyMwVucTIl3gUCYCQgIOYVW2CgR+KcZvD+JYApF2DohJzUo9gF1eT
WrJCeyRImtfvViq8Ge7pVJenj+l5bttmW+Gowl33++ScvQvyaxofBFuL/qGeuac/
rOWrAFufIVlehR0JfCvbOlaQqqaS+tPKnep9UmlM/D1eFkpCBbhHeh17+tFLTtXG
kH7Dk1umew8tEssfmiB6wupKykk6p4woxiJidICdx3Wxd5qBQlSt/nqD+X4wh2wj
dEsSUXyIzNpbIQ1SVO6flra0/y3IGWe0r7KM/GXWm9/mFnWFmlApsvStv0WthKcA
55S4wGoGn4807HOnaBpHRW6W+vlSNCszIrMI88DCMSRYHZuA3R3NScHdiDsNWNey
RvMMgsSqNRuI0vJ0FzVrok0KRzGfXhbdKlJoVrzc6PJkb6KS71NpABSVQ04046o8
iA+S1fv5uF1WFYYRE3XcnOysVXV/jYPF4nv9QGFPE7e646mBXzr9x/J+BIzK7+cL
fGduxCnuLLj638tRU+ZtZsIX6M38pgJNfBhoV6Y1SZStNmJTTgh0UDU/jvXmXPXh
S7jV0ZIPN6Cor8bXo6gHim1XMLAHEgzmsjxhccsANhHiB4CJyMUWhxysP/vNL5MD
5AeIoVvO/+eLSRvcF78DO9wpizMW5Hezm/T1AaSEoJtktRQNH1/FmT87ZFL7F5vo
VfFu8zoRymZAki+SuDYyYGOoa9jhaZ9VwVFxqB41+6Dz0UOeeqTMu7b7wtzQ+qsj
YgqTKQBdEVIqK5ZxBlhTvddTrF0tkki4WWHzds5W/dXG3tHBH64TvcYJ1bOG2ozh
/8zZZxyqppeNHjAIDYabZ3mTPjx2iKFuzeD2+KT+jZNvw+M3zESNbrHtFdTxMK7x
MNp78Vbj4PtpgHm+xBfjDcqzMkMS9Us/t1ghSXJ9/BwbGdjRECyvD+YkYaHAR9Wx
ta5wTBKP/QCiEq7B6ip9awhdIOIt4oN9JlX7YbRZFcjLn8yoQfket7j4LIlc8laz
s+lNJF6/bl93TOgFDIsCfmJEO3bpxuGc83Xf+DRFjRUF1UUq2MEu42yEZvTku86t
pQlDeYpRMi8vOYnpM77mCJ8j88jcyx6Dg/8OvWoO3mwljC/bZlzvQunOhShEWOR0
XeNHls28HtdzgYXrDTO5gtQ2j/Rwv1PCpEq5pYXaayjGuwgxw+NbetK1HkeZSCzR
1w/NFMbJTclW0c+fPkoq0ZiTNrLWakuZR38344d2NH69h9ZUuCmhB9edMtvc1P4B
NCEne7Wz11yWhbYyq2R37GBuL9XHVwtKB0VKA7eojEqkc0+0nfWMUbM6zS37Mnvr
+Oji/Wowx7nS3rxyH8viwiG0KDxt1ONZQSNg5/R563ouiVj9xWXL5osbAAk1/RmZ
928+MryAYj+rgnk5GOjfWeea7ETJFkbGM9ucZSzn39bswtoPRQSZMJc2Qflj+MMJ
Dtnlt80Iyy1bf5HwJvPcPkiauphm0B5YE+HXTs3sp6k/FvgxxTiy12HnzzLWoU7L
CnW4Op3QIe9lr0Vv1hs1ZQNG90PT/hrJgMVD+it3xKNY9uZWDO/9lLS0n5IfAxcS
B1GXt8Cqb+6W2spLOylyCLQCppfsJiz6n5dMPXzbNYroj9nicaVYL79Iaw9Ty/6o
F/cibx3B6ro+fLMUO4c/ub10SVtPMWj2wDKQ+ke/jI+jbQ07kKjDrDdOh9qEBjKW
IulOj2TUOQhBQ3A1V70aimTv9xyuKDa0ItS3bbs48lLc9YmEeETXymmTwY2vHd+Y
gLx1qo91wiLdCJHkKoceqVVBq5UyQXTRd5uAqHqEzwXneGJNB3+fPD/cT3SCcCsd
oqesHQ0mVnmam77B59unKsx4K6S3WKNQSui6gQmjWQDSdnkkxlj1ysEjnIKnxPiA
Yy43bI3QtF3tkHqkOpUttyf+UCmpls4biO7lk8ghOhmbowzynTb3DMpRPQHy89WJ
Csq6pbO3P1RWaL1Rx5Gajoy17/eA3NS74dpUD3u1ImOrBBZxP6qzpUQ5TdOVGd7i
n9eBchH9gks9dc5Udy+LOgWWzywZ86LMZ6NnNWZKQceaI0MFasJdtjfhipzkq/+Z
70sXKqdHGasyvGefMws5pba+P+/Kvg/vHUHmnF0EpwVKSZhUJwwRagHEnIf+lFq+
87UOmFskmqZ1EMH3RgkUMzZtiwmenrbboEWbHOnfwWP0G6I/TsGV/FU2ol74joSQ
lQkV0fDLibvTHGiP+6rJto4lQG1HVy8YgoRlb8quCap/Mfyc2KwOTY0YOkZUjPk1
otYIuUhp9sYTOhxFTcSkWJCTsLmg2skOpHPCWmsyV1DLSf6CXaeDWJIjbBWypSnT
4bXK+iRUfdIK0iZi6fY3sDTlYhCY5mbtxu6LllmWEM/0jIVuyT0QYe0VYhtlWBRr
oN3katixDOWf5if/rQ1l17CZW4YLZ4g1JuJn/c59GaPbz5r2ctPeehtVR14kUsty
6uLhqdMAe3OF08VbQG+IijpKbAiLqcIktbT5ZGHmkw02eG6Rh5+WwPLxVEgEG0mD
iCoWbQeWfbMdSM67KbagJvJ78Unq7U5RhlJsBtOZIOcg+hN9UpRH27yDf1Y3TaKv
//pragma protect end_data_block
//pragma protect digest_block
Md4uH9QnaLP4t44j3BMvykSs768=
//pragma protect end_digest_block
//pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
zSzha0vHurzb23IuT96njezAoM5t4HXutf+/Bj3oLkHS4bx6PF62azP8DGVaVhQt
ro1kjjmq+LI+Pg074bFi+Q0jelXBJ0JjdmJaj8TJE+wYWeMnA6oD9js8F2Veqg4D
JFX9W8ewLnGr2p+MeqIAn44DsciVx25G++jDC56c0yM=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 22096 )
`pragma protect data_block
1rZ+xA+QOaVtxKkckVvCkMxLdypDIejcEdhYi+J8GKWO/xXaGvgg9BT/5Rh7ukRw
cx3ZlDRF3BmBcJtL2u959OJi5tL5mFa2n6OGroUJEsm3gQkZO0wT2FNcDfpKq2rX
qNiuTqqdMxnycXgEPDxHqa4dsqCgJtx1zjccWZmBPLzZlv5H98W1T06wzu/bGmL2
m++WQrIFdJhhDXA/s6wofyYKqcn1+07WXLYraUUQWDVXwF0IEOKYSQyUg1yo3HqI
HrGDI4qyaWTQAgIlrynspqvrYwqF1VIfA0Z+cHrl9D/emlA4G0y6qWYGcYlRPe5f
mmwZ1kQtpVLhBFG6kUXa8kYEa47QXn5sEqKniG3LKKUUsw+wMNdHrBKJmebyfJWi
27800kapE7eaYqo9dtfraGB+tOQno2paKnlW8Ou03xOafrqrMGPJOZOgE7NmRj6l
r0QCvzhfDGJKSQF9PPY8CQz19RX+Lw/SF326z/yBOqTkYVevj4kIIrPttBF1hLN8
6n/6HZnmWB2oYE8xRS7w5kQFFFIWLEIHG+ATw1RFIPDoRqgWfyc+aWWtTsb1z4u/
3ldWICDVClwPj6x9e0NyAoGxkQGUBJzR2l6fclELzeCPnVj6PWfNiP/QgbMxkJ4B
/AXNFzSl6ZXqlbs2YTEZ0pWB/pY09tVrjLMXiJMr6cyhQs3hx8Of4CdprDHFD/eL
cIxFFVVPow7XbUc4sBWAX7kphZsiieLoAiu94hKkYUmJTmj9hhsDghrWqewKHTGx
d4fR0uHWGOW5mwn1M5hdQ1ngwiiccsQ/kE0Sl2ranvCRi87aVU6iSBv5a3EJwp7q
zDFR7gWmsXoE9i+UUuWU0ztzh+FokaJjnQasZ/2PPoq/J/bCMGQ1PQp+yiy2FiYJ
dnpwOdYvlxVDyjkTw3+la1P6jxRy+pgtfSw28/RA8ubiIQ0j4v4Eup5Szss3JYUb
eWpt6n6A67/ixPB0P7QT3i6GiR1a3Ik+ctoelOOSZoKwS34SHCg6C7uL75YoBMp2
3dSZ7zzdEEcwOCRkCZMuMYgF45TA20qE++c94wi65cPIsQ6F42GC1tsPFPVlBJCN
gIvJek6mzvHEs2v0TXY+b23aDB2Km5QTbZKzAALRlDzMCWTuO8AEVQP72k5pOtYJ
KKlV5QKPIL6p3sTk0hLaABSBI72ropQVfyehAUAvhcADJq0yRvVtHQhhuyFX1yhF
iUlwFC/s2tvSN7tPC1AnZB2yeU5Yi80nEdXf/x/DZ9IpTshg25s1wunw7l/rm/ym
5Rt+/g5IFZMYLPPEL39nQgOmdkRXdPNyXBbbF5hzP+LuvrFbijLHH17qC7VkSTbl
2YXdGIgvFOoMu5xts6hmPl/PTxN00TiAtvNyiSrU6WtvmcJONjPAxDL9N1i8/GjM
TJjtrxzt4Ev/C4xC1ii3odmsQeWMuYj+zh+eb40eXZqkDd6rOcVNwymiQkeT5/Jw
sYLJNOvsLwm8wBPyuCNfe2PhyY9nWEW3FxKLmszqy8vTdLmCpy+qbXtkSxS1wUkY
0b5zxq0UzcPU6Hf6Tym8FATutry1LJfWQMAwDHdvCF0GzpbD17wzV/f2ObjNL1Mv
nyYvr/ntDlFhupIn06bj6I1B7l35gZ8UN1yuqJpb1VQYi/jM+qNUOGDoOBPeJPGb
fRYGIi43cLW3Dejtg/mLwniBrTcIYU4Vdajgu3Rc4/8wzwkEr9GQjC/t6G1XkJLG
yP4TbRjPB53By4M7UWA8KzgeGxWUWdHJZgQJsTV8/ej63Ox9WZq31n8NuizBCgpc
dOFOjgk3/6pfHlH5IQwSnOeMafMgs2sCKDJkpSsOlA4uf/XXh3q9lVNLjtGI68gg
AhusudIlSN+rriyvaIEdU3fQtpdTV89nCRh8s03iIZikZXJ+FTeocmUJwUhYdz6s
xg/4YOIc1Nsct8RHK46Y87xqkN2al358CdJ3tHPhiuYdSSiT3rlVBWfQlr3/Kg4d
djqhs9TwSULZ6KvcWnws1f2nNpyg6f6wAZrjv3n+sLdKYoQBzy4NQAaqsuTWfbD0
9QqVhVWXQt3mbuC4n2O6Zb2D7H5wRM+bWuET/oSv7i2mAXvp6JH4IQl1WJeTGmp9
gu8ETkt8Ks+PSbo2q/lffqYgJx7qJtmnSf7BymUL3D4sVlD9wlVo6TIsBwBNAIoF
XH2lk8zMNu/Nd42A2dlXUqmbAgLH4ojjwlOVc8hWyvYCaoEcyVA2+U/WmebLz3Sw
FpP6QL7S8nwAMsqpWnfYe3G22FF37bPAf5oXH2OOLbGfBwULEIh7pwexyHQAKes3
sLTqyjFEYIazkaforeW1DY4p32IZgHHjIDK2YrSu1a0KGP/ppozrNAZ2AhHwmj/k
eSXgNkFlFs5tcjK4gRfwvNPDq+y7ly+FYACs92Sh+yD1b51KfhE9CjDfOv80pICZ
w5mLJ3kqg3HsBvcCeysWa7Zx0Cez4bSJQ8khT0/xhPE2Umfls2gtFXdkQpYQDpif
Lj6ziV8XcZCD31mwbG7yDKbbPAet7dRRCV+8ZsOvzWc9jbLI1//8Ltaip61gG6xd
Oe8R6/Rc8+kGRBiNmBKfPZCi91DO9pQMob847BbluXK/JPlxOpZ9+yOxb8zjdmZ3
jXBUBwS94LU2ccjsH1nvjqboiIfmWuxBSaJN7tdZmTB8K69gCAo5oIO1FIj92/0d
7vezHG8EhwHzNYA3RSYIy8zrO8hS9hl5nhBFG96pVHJ5cD1oxt5Fo8NG2AS2nSnn
xmw3me/yaYhES1jeo7+LpGzcyKWEn9wrThwkMMOzh7oraThALHX00P7fmJAVRe/y
vzyJkVwX0XPwlIiijoMItrRyF063b2uuNmVr625dm4NK1SFDW4qRgJnKKBKLZTVW
ghAAWYGOuLw2zKAjO/jjDWTRBuHvkmr+WRuXXMuWNXJ7FV7/2whblXklZvfeAd2F
gA9rNV2DWMWXSlUi3+yln0eedBdVqer4BupWXeRyP3Ryh0RRTAaCsimAbdLGd97L
aIPhCNCs1xNpTD7jVRzvOzkCGyaiT/wUWKlnX+AFjcp53xGzlyesA+3+S9r9wwDa
PZPJOGjEjFVaie2I27K2Tux2cS0WjU5y9mSla0valVmr6+0Ppg2bLFpSHFcGjeXq
PiUEcGZFSe4y+9VQG9qPBV4gMK03Pg06X8ZV/KQN2kYGl456+Xxb6xM8VOI430re
hUP6P6zyKerpI7RIox0fiseTRzkfu3GRTvAc6lrbQZthGV5E36cvJcOSNyDxFdvD
szln+2tbggRE506Vaki2ucKTQsFI1tuET3Q9ZlsBV5KzqO0YxYCNwhEhVxaFprh9
rFKnHIm5HZFCJUrA2WuNgNIIPsCsTPhscYivberaiLSLxPxcqibMHBEhNuraDHv8
KrECgWb1mK6j2B71ZMd11QOCJxVXDCU7CY4E/AuiS+XKFeiD+EWnHb1lx/Ui3S8x
8IEQBC+R5M6ayylm+eAsaswh/zos/agZmzY143SiaBzxipUD7lm+2syCkQtILvhU
L6ZEOY55WQ37IUO5PeS+/mbePc+YgFN/hmeNYTmW5ArFq7X8ABp761aPMJxbHjta
+sDqpL5v2QWRJUMuk2ebVnDY0EeDsFp2/EGCHU8g/PU45jtykJ6rt8361QF+9kG4
+4xbCBFGWlbogfNqlh+c0CW6dG/8/TYB2lGLeBcwRu4DnYs1XVJFXVDCwj3wVf13
Mw2ClsWEOidCasNsoyl6DYDt9mdOKYKbCnbsn80ElcS/rJHZ6IuiVdiZN65/4PVN
QjWn+F/N9EV9r37TQVjZquWnfQm8lPSL76Nz3Eu1GfvzMczuAMpgorANT1kjchE4
0t4JujN7n5zFnZf8hXJEvS7aWv24MFmrdutPAEDiul/wW2b2sMdsE9rMRHKnah0b
DsqdHV/Swa7Y6f9PmLBra8gFHndI25J14nwNlPmgPAyqACvpGfjafZKe2Dyr2kDN
8dZwV8d91Q8HxQdPQfSrJirSuLVh/vxmEG0wLZYe7epuNT15fN4eJqp5g0VO8KRi
BWZTog3AR14VjKjNg7iVffHSA0zPAfp5iTdU2tno0/3El9q4lU8LZwhUEPPg/DrB
ZlydPqg8O/vbh5fg4iFni8YKL3DVCqKy5ejIGTjCTcRQd0gD0rIw6kVen+/4YdF3
5q5rbRwgCpxMP0U4zAzcE7Y9AQO1lVtTv6UzFD5to/eMaDTD856srMxVVATXJoYL
5DVhbunJtdOgMjBwgn8rOZPrZVDFNOzlDr/6Jp0mikmcvL+SQy5JI+zo6kzkm7mc
3DQMHl7ruJqM28kaEs+DbLpIPT/kwHTJx1TkuPndZdLuG/g+Bl79oldZn+mr7her
f1zGocSn3/nvFh94ZmpiQ6GZwJO20RmDeYfctUDRaDZLdQQ5PZbNEi7d5VucFgtz
u5EWGoC4vKv9Y54F666jnlN01xwmG+fKW+iVmiLsSSEOdBjVx58EdSPrVYQoWshS
owg+jY4dl94fapuozSPLEWVLLQejWE2HKuGdkv8khrq7TbzhgrU1FEyujtB4907N
g0S1d9dfigQMxAmXyeuwsYr6DT+wz0r9jlBi7vk5iBO2mSL9+wk5IeV8BfewBEyk
4+6a+Fw7vGR+wxsazb57ujNHxknC5aK2zGbLC3QGeFTSumwIK3faTNUOZiBnTmYq
0z9/jvZvxnfV1gvRFyN63K3fnvkAdFe6S/nsut9QRfgzReLA1nFJ8l7T3c4nS79S
V9KBVKDCkG0LRoMHqdsMVMynhSJLT6MXRJferALWElrpvGTWaPkdi8U2mKc4Cx2I
+/N9KaXL7xubXSGfSOGCT0p61ar/9ufyCgeBP1OumkwrM0ivIyutalpY0mAmMDL2
UzvkaCo9p2OcPMOjl3By87J/NgVv8KwV3FkOqHh3hK6T4o4yp/EX1AevmP7lAx0e
ZxfA6h2axCdNEOGfWT6D+SvFiD+gY7mmpuQgXGM5KoSaTcKjXx4V7jdgfL77J/QC
ZeJT9Vxs5YC5Q1ctwB0SpwnnzrtT4VEdZUJ4WZ4AAu3EMbjGLWk/UhotdCzbx2/K
DYwbxcXE8O+ucAsMxxPUZwdIHN3Kj3C3p11kU3mlHAARHXTjcXaZKGQdntihVdFb
cD39n72/1PSXb3R078bEWPuuRIm6RVPd1aKxZQkiCOWBYaAmO4bVEisskjjO8icy
sPQXZVKU1wZDDoEh3hC9QrtjZTLCyJfaI23rSud+/fm+DeBCBST6pyqaw/8CBJCZ
nW8Y6TRrL3jNe9hlFMA7XEUZvdZf/UaaDEuy3KzxYphR286nUZXzAVTLjEnh3OdO
jQjNGXT28DzgncGKa4SFofrMHEHJdSyHe2m8XM7sRbkDPh3RrqQo6SqVdl01iAmH
RpGat178t8BSc2txRPtQLGB1D7Klc9GBQNfDpSWXp7xsO3XmD8BkStGOvZ7ET+7W
3dEBfwKdaRyx5ecYIIKalOkDeL/24RtNenVMGrHr1nGPSdtHe2+wKUAkAi7kzICr
SZBlvcGY+a/1VZTt+JJFqREgslpZwHOalu7z16s7SDiMlT5bcT2nbNZY1rsa6bJF
VuenJ/6rcffVAuU3t4AExJOJ+1hnhPDoLdDfJPvYsrQg2tsultzPwrfzzbxOptRq
YzPSw5x8rXJuI4ymgmsmcLd0uEEowhM4MEJz/G/yZNxp/N1Ys+qSAJRhz6xRtd4w
dhCq/Vnbb7wgjdDgLxpNlB7OGj216pwIORezJIZ/wd04PMI7fHLcRnrFMIx/S4dS
nq2cnr9KKxbgnh93uXctAvV2gmareh9LKWbhcNzdIWrdSwtJqdRRkiU4pBwz4eT5
3LkmiTQXQzjKZ6MRIyIJwKogxYGI2/xhUm8Kis1FPT7RtKguVKMc1GGCBBD7/wtO
c6r15ZBgh2gK640U6aAeMx7MtyWBaEaF127sMO4qZ7qjdks4bva6+fWnLCgH4Yxl
UaUZePx38Ba+nC9F21bCrfJTDGnjp7t7IFt9F/kEJ9Yj9V5psfNPQEXHXrZvlo9T
yDRUUQBINsU3TP8mF/xAaPJiPWhMv1esIHvpKChqeTQIrCUSHvxBKa6kfrpUHxqS
CedX3r40M/RcDx3HCZEw5+T4aJ/x2NlLA9QGqmyUK27nmhduvpmp85NcFMWLP4eF
DwHRErC7XhvSGESAlk+c0ASXFUqaHxmqFQxwIoSzpQHuSHMMhhct1OpGJFR1ZFYG
gosCfsKc17PEoEJYJyel61aTRnMa+ZqtAbEPxJ3+Y6iEmvMpwTfCgqve3Lhm/wZ2
ziqoSvNz4gQyzp8UxKvfpQ8aRGwlZ7wsr3I1mXZdskKWLWk5YM/RfSax9QNJlsm1
hn7y0qeCdaWgem/ELhb6KrNT6sBrfux5bdogBrDRioxAJUOP/EA/1BXAN4bZfPbv
SebIo1pW18IzgtT3g9FhzzzHb91EOU/Z0Mjj8J1sm2aeByw/SF/u7hQ/7VD6imP6
WwK0jy7oVLAX9qtWVO26mLoGlvQbJbk0oG7umuIoPUm43IPluHim5RBjJZtQ3MRv
zd+Xrs9JNfVQHCKwIyL0pKxMAkXzBATiWIIDNOT/H+zasfv8Cy0u4kG4Xe+OBq+I
giSkcateY2c7ES7cAlViZAN/TeHDMjjAgCUbfNhAql6WkVISh2X4VL9fp0ep3mSo
1I2lTXcXm2joEEgVtt7qaF+cdJJM54JpP3cPLr+X23Wf2my3idm7qHJNO8WpMxVk
4//plNbp1bxIAqnsac9Sjj+0RLJWcjlrw4G/lZuQcO9qBATqwdYBiAWRJI5vUWch
qjMiQ3CF3Z5722PtLd7Likk2q8o8BKr9OCKciBcL/gfYKAVWZJSsWU2siSXcA4VG
sHO1kp8yGjZ5+ReW4GOKND3n1itxcKtp4C6+BNpTNv452qPtEWu+qvE4Yc8m45j2
h3I5iamcXxG+0COruTxlE30z/6ekuBqYUa7EvmRoyJYXDJkkFKGcIPTLTdrtZAHC
npn6RXrwZbe6wMOYvrKrxKx/dqsvhYyJr6uVGJ8C6KMg+uVqW1NWaFyCqKJgydKp
GN1rpggE4OntSVn9swl/337NsQx0suiLiv3FR1uDLGqyJ80jcmLguT+/Mfo74uFl
5H0ojtTzq9UZJkLMpRfS/3DbHKXGvpifurIlNjoTObhXQLI7bBj8cBXLQsU0hiBu
Nq/fDFO+uviVcRKcv3ChdjggOKHSeBpn3quwVpQyxzqRen9rW8OTNQRmnnSxSgc3
pJBAVUA/GXDR87Ax9mQb/Z/jV3mHgBWHGyfjKyNOMfDENiV9Ktk2mkJLoz1aU2tP
yaLyjckMQTEmalJD7gLQrWMFnKJ+0s+Het1syB+gRypmtimMlYhTPtoi29RXukht
mnzFYW4StKCifTSLMScIb1M8I8GIEKr1YlTSiF/4Gl01t8vbtl+JBK0f28WyXO3E
ugPiyrIZ22aftLU555JPdiidqC/1ehDfK4siRrmiCC+86chxOF2/+j3rcH6XSo9o
1NHtYRnOYQQBcDPY6NXqOZ1kvbccyKYHoXtbYgiWVlQPGyQvr9SpQbQEsLfDYYD/
w4nf8aYJoenhwt+DbkqVM7gqXJ8tDUhOHSxSbzd8G6x05Ef9mTRKWHRuXr6U4Q4g
k1yI++HbLrytoStJAHkoiMFgZYZUKZH91vjKn/9URoIRTQmdKTz3kuquvIxvlL+x
3zlgSPulGpOlZ2F2wNaYABmGKafMeNsPi1m1uOeWHf6MKTJnETVv+QGrm6W8r9Xu
vrTQu4D9gEYUvPodrdfTDng+yqNLEzLdeLpTHSuNkC3LXdVJhHw3lqGC5G/hLBDN
8CXBVjnIzzvtwicGZh+EiEpXxnajXZmJHURAKdm1R+2LqDYFbKWj9R52RpiEdHPv
V3wuLPnu5fkZib6gnVcjtBGxb2LFdsDtNLmQr5x4DNRjhuTm8L5wMQOZVkALBFUa
9c5QXDT/YSr3QH28NcEU7QVnqCjouDViMEESZoKVOKgkPWTim4C018hW7bkyasPA
utIxQG79ckODUfG8EnIYmffcFrIq4wrGO9USwJQlcD6LTrnhV5IDEBvVFlgpSrpK
h08cfE7HWuPHcz7h2sf9dRvFHv0FZ4EERmmuF+GMisM8mhLq3J8/IgmZvPHgIAYe
P9mk36ziQm7KcK+vCF3IogrGU5QuzQbW8OepOJZdGxY7rDMvPbfGOU93WYFidKd3
6uwioQFCBQqkDddM1+LUK3gpIaHaUChYv/QP+EyxOF0BmvEVtTLEh12MaXeGOK4f
e5BucJIl2kxM601tQaCh/YCzjCJCALCceTRl4ZQOS2YSCkAzZ1zT3YO5kEKtCsCG
kPe9M2su7/iQfbz/uw+vTY+oCVzYXjMTp2UwvWeduHsufEX/A+xWiA6hfDFHRlfY
kVIY0LJH7Lh/zcz0qaSwY+bama6rtjVO1/xn13YxFZJjyEd5PY89KIrIwV1+KyKG
BQLB3z9z1K2CB9RvqLbZp6HsuBVvX96SMtH21nixcNSF3x2+Ba8dEBFJxW7cu7jz
MowYXWOPApfyjxoQU1UORpF8DrmM+PLKWpYUunQy8Haay9o4WNb6LQNu2itEfKiz
9V5kBI9cxwAyJ3D3HROzgaoPsMrJj5ocbE2OlF1y610wI4bZHksUbM9Me2tJmHWl
A4CnY/BD9FH2IB007jKpKi/jPzADXmzGsqtqyjZ93xyV2NeZ9p/RnzWTVHbK8KL9
dRgVc4eWgC2XawHsuTJdYZx4BGk7CZQ64j3LL3putAjdU2EXIQQ50N+oOvfsOwYV
SJoKYTJQ4BL2ppV4sowQGmofWNy+YnpQilbQdxxB6Xe1Wu08XyDgL/hWuXS7SSQV
7pkqWA4A7kLZHOPLaGhnhJsXVHtbLCby5iu2upBOGjpnPtTH7a9BHTWLlAS2AZre
Pv6xcjfZ6Yoe53ulTG9A7RdFz9si1qOvFloBhs9R4IjcaFi8orehkdiIxXoECYgX
AgeZ68RCPUZQcQQ40t6R8kCBMwW6IH4W8de/YxwYsY+25mQ37FHGCyj6yA5NGiIC
yuStLt9UipxhJ4PwVG6Px7GOu8dYF18gQtvZCZ5WYVwWAZ4kRwHIpd/y5SgD5VPq
FPuOKYHnLXTt2A00E2IdeMvHYTetR7gYUusVVGyoK/FaNiJHfk96lnk711ovjK72
OKl2DBcx+rdqvDIveT+2RqSiGk9eJYcCM+HlYHWleqy8p7DzhjPkXOcp9DNgGKEx
d83yoMfnChMd1rXMMp7ucvpiw+Te+CFdKLgj4e8ssWDltum6zJlsWpEUXUSBWABx
p02YVI/nb1ZwS0lOyiq0t/jxkb2hQmnO8WZpP+zhn4feBVa+Wnr+oBEFcq3YV9Pj
iU6eqzQ19qXTA1xh5Dyo6MSYYigI0YgnC76AMugLcgN2zUcVXaNYfNqcWgLbCnmv
pkYSH3CHd0/gs2kM2lxqr8qAz5IO9q+nikVF64Y2yI+N+Tf4dWLEKrQnVYVloo3w
6wHKKjqnRmjJRAYVM2doN1IIXulxsoZDVPLHK/9V7qBTX2uHvpjK/AEOs0atsR6I
zKYnM0RAnN8jGx0ra25TXVNQS8WYCGzPhLeVimdaEhb5akA5rHX/WzoC53ReLm81
Zo/DliCnKQJ9O2qpu3p1ZLvSO5gzLoYPWvIsJcW78Eh+FuIPGF+QVUBNRbzZF/XO
tz3xcpbMPG3KTyYdKqhTCbYyHEyXhNNgdYO6EdmE6KhQaDi7GnSdknoxmyFk21Uf
8zj9t5LtkoTAgXojCGylQNM1g9+wm3oQnBkCbUjHglPOmIUFoeSa9eLGonx3pU0q
mnt6vjdWwBZ0d37S+E7cSJjDgRn7Rbk0/TDbV5tBCFVnRf+DO8Om76YRjTqz24lt
dfddxJ1mNXVc4qI3EH7wwbJ/99RA/i0ziZuiPB0vw9bNDeYNEPE7QAhGk5xMX772
vtGcR4lc6ZiT6QQVDiWUc0z37ahMyiLX9Pgo8v/BmEv0gJ/7R0y0/Q/UPWvtG2TJ
zNtVPHd5RHweX9oik/goNnhEyLXuZDBscTM4tlNvKQq3zxScd0pAbDjsZeIo0Loe
DUzT97TB6uOEg6vrIS9Kkdss3FGDc4mFZ2khy3d+uR8jNiHKgQz5rUi7M08As35q
9bkyu129Y5fnqc/9oD0Xxb7j34zzhfUstjE3PY8bEeRXZjHLBRjn+/tsM6Tc3Qaa
M7dWVlEKYakFq75V90jV2Mr5UkBaSIH7RcOlGMCV6cKQnRaiJQIrsfskjLmbGBqY
u1lU3j7uopYhIYS26XOa8q5SIt4IMFAo0eReHyhwz89/JMff+hZMOJmaruPxVyan
aj2+qjaKtqV7BI+14I+VhwY/RIm2ue8dQlnaAXQ1ohe8SsZErhMX09IMvfttwvC7
VDJGKGJe6az9WQBYDMCk0+YtFkBYp2R3JhhE1EgzFWf1chaQglgvTChOnC0wUU5D
vzpHGyPetbNlwvgqw3tFxl4FGQHYBSRfIWdFIFxR0EBXAF+XrAvhIzH2iGQ+krJ9
jskuVDsYQ3hUlI0rEqng/IlFzF9oYzHJrDDolurgWASKJK955YiVO4GF1tOLs17n
s2y5YAzcheOaD0FKtZcaQyGa/nWrKgwqUAR6Pf6KSQC9HoRrycFskjuETjmFXH3D
zraNjOIUDVqFykGFQCA5IbMOYbunbhJdZXiagFDXFUItDOPjg2icYvF0XE6UiU7B
yLepDB4Y6/D9MO2hd8mT7r2raNFz/u9scvUXD4zdHlQrjXCi7q/VlP+jEVFg71AQ
G749AdMDei5LN8hzQ6LBNNBbh6kEnoLn8XX8qQYl8X0wox1/LmS1WpA4GR8TaWEZ
bgx+Ku5VH1TQxslMoSxB+8l0HgK7aw5mR6nmFjUU4whCGfKEEyXAkMdu4J1I4Wsm
jzo3/0Sf4LVudIILnahLajL+MqupB/m4O9zuPf0dQq3kQagFypAwSya0315nL8Pz
QtNrBEXRBAV/Se6ShVhI4rv0XHQfZghI+Pt2+mq8pK/2vUNMhWmcXDQykTBMRpqz
072NRX7e2+K9DWaRi5dJgnEAdDJ6dPrYfVSvTUhVdmOpK8qjEqB44Vdv+PXx22jj
9Xsc/lGcAUaxMC/fN2O/MD1bWMZnkXLzR3KJArPIj7tVlHP/D4YHG7MNe4334mNh
BUMOozhrzKB6unKMBFfKGvR7DZLkyq4PV592DTk9XmEdG2uvbYdNNFC5m5/tW70a
0A+Eyzv4pDDLhApqUbgKGUnUfpDE6jOjI3gUM4h9DsobiPEdvqQjMLlvf0Au+9+E
6lqnTxSiA9++NVJCRqKfqAiqBlPXvEVlixk2COlzDvDI2BuWaCFLkEkzaktEFs7l
oEizHEgqtLxZ/MXtDefQTcTK3zffDsW2hwUa2DxM7skkZpTBahvBPs+C/PvnGJJv
hu1ED173/d7TJwJHLe9r+kyI+ilgDeEO6OYz8WR3GNx1A/yjM/qWcNTs4S6SdIuU
yCLqz+L1PfsD2ACNxovaFXJr02vYfFgSPhycxu6ddZXQeka1lyqh1lZj9e+cm6un
ZyWXnuGeaRbjRArNf23/tin+05ePqld/WsgFOg96FuGqAS0Tl8rrjOTL+0v3yPOd
qxPSGXqzQl1iXmVh1Q4qtmguOd4liwvhp/mpSvecgXsgHdfCHLqbpUxuT5Nv3Ffg
a98wDJogWHfs6TJBweV+6+hXkLLf9WsL94NK82RlY0TYANMuKQ9aXSMJDAiZliVJ
JkZCZc9ejmaHZDNo0WfeENrwAEmreCnJo6sTqW2MnFDXVAXvwSzZ+v9xZwgH+03f
z60ECh1Kt5/5E9zUAqsQdcu+70euhVrT2Nqyv2y7pDtcuouUnCnSiaRkJZQjo6xD
9jh4kasC/oGr5h1HRIAbp3H1COXbvArzGz+AIfIP9zif4+I2HhvBqh+H9xgBz4jP
B/xzdsDL41qrcBB2Hl5TAcb/4ZUN5SlPus+JhTBwToakbWx+H6R9u+xNW+HCcHLy
o0rCH+90jgmmTuPPYzdChbv0xkn0/D5dad5UNBSKAELfL1M3dbs7mHhZawtG70i7
mmumbvc2UFaXRzS+80D9wtfKlOuH60vC7gl7jiotHCTCvc3rX1OSUcSRWC9BFqyX
vOO24DjstIMejDpqLUOOF7piGvTE9YFlCduhnsTmH8QKWtb3c87VUisU8ZS1FT5D
rQ0w20C4EAMTLuU06S6izL8B8d+GvZpNQRljyPai40ibantGseZPFS5q6eylQVQ+
gxHDFgstECyVMZLm/s5OCB4qm5CtjD7Df2KnzFkalSxq5HeQApmxNVJbpx4IhDZ/
hvWJXClSRs1WT7VE++AQCVCmSY4arQ3Y5VxrIXHKtbL1+VRI7OaycCXapyrlo3Wp
/xK1NR/y2+J14Bx1svfIz6yL4+G4OYfyY3h/OA/xwf/UhcHH5VwvPFi/dbkce9EO
0Z0iP3QmIfqq307a2mmBn1e2ZH/qi5e6EFcYpVcUntAkIYo9MeTRSKMeyRdMeEms
wO8CVSwYPmrPQEXfDBjiVcNRKcnFkpFn0S1p/96Eqrt3riwxL+aLRvBs3MyyqBf3
QwarBqbuFdcanGIqat0szMeb8+Q+gZZUJx6nIf461sGFkyIcWaJ8IlxSF/C8BEDF
So1vOLEn3GwgZVfKPmdNBsc9UKShKzGFMY8Kvbdc9nVtj2LRj/Bo336isxAJGF+T
iBRsTI2SbVa7LmeuErs0FVkp3i9OCNIP0Ip7C53dTL5m/20hoEAFTa963gI/TDqH
Z9ysG62P6jhToTxKOKvpRvv19tjONCNM7Jp9BnJrWE04bv32/vQWh3GOFlTuCfwq
yj6B2Xw8D4IAkmUSAH6hctVNtnovcRup1ZyJg4wQbqIeRfqMuxFaiH1650sX0cXX
Ty/HoYt7XFNfckvr5TsJ9YpDtzAFFpbNJyxf5AYCkJcoJRE9d0OWUbjNpBRBxVp9
AeE/BnwuXsmNj52kE5DNlhSsKYX+D+c/dKG62/xclc69EtlSH9H4pe/vPd0H+gMN
RG/ZsRm9q4HbxjdnMqvCsGS0LSuKgRf5R4M8AxOhBn3dBchYC/0CEKutTBgG8zdy
DYKW/rpOztBW2FeFOGkJWtNIfNWXKEE9sgpDdzUpmfoUywXUgonznn+HGY7Tk60m
ujhKTn8gAHA2jHkaqPdGlsV6wD5KpiC8MH1KNI2p+v9+uagAYCMTzBg/xs/GT0qX
cfCzKhmO3hboT3gVNRCykGsH1HK1njAI4+Bq4FBWgHNFEzzKLeFloL+Y88t3EaDi
q3S+uMOX+XyZCaHZvFRvLQmIngwibFS8XKSTPi9OShmEHKWaYmRfFRWHiUPE8+K4
RAXneM1TFIB9rMKmDP4NLRqDKAvu3Qi+ryUZbusu6F7PD3GDdw2aILxkXGS4Lnr1
SbfYVXySJthbL6QaHO8ESy5/fdRN8eNbZR4+cwj46T1SNTwd/dSpM1UpRxLuL4cD
xUc6Q86YR3dBHzmoGG1RM6VwSP07bXVoU1tyt9/7bfte1guVz6KPWToZ2advxL59
DkK86uJmd+ND+w1l7/luUQ3QmHr5oGjeeFm4Oz34C3a+Mpaxv5U613NXvJH/nszt
wSw7myowW/MORG2ZL/CbgDwFozgUzT5nRksiBDkCGIBQadiU3b6iA3TPBXD5TAzK
aCB/sZszvx/PaGAtR7WdNqE1i9uKszgL8SMuZqXYYGA7nbzKfs/WLeec/TXokJNf
ve9eCbLVfmgpHFp7inJca/zXFf78qrzd4WE8KSy/rflmfTX0HSTXgmiuFxYTPMNn
WwPHRNIQE5FiqJMMvvd5/WXtzgPlGIvEKeitvEUIkJmlmindWE7RwdL1ryk/TSt9
85kjZ6jVYA9vxm9Cea8wbNGeS4D3Y2ditL6H9IQE80GDdEuMNaIePIzXXKAihjD/
d5rIuWQehmIBptyDpPDeusokysvINTvad1Z588sjRlySxuvqDIM+JSPR8It8xj1g
yOGZAQtTJc3P3k5NPg/VH3MeEl1GeQ3YIolu7e+JsH2ZmvGuAo7ckr9yZmTaCZdV
fNiYXsTRLF/rGOSqjwqvT7PAElQEHitrx8GXKTcp8VNq9mOXHYkz9tpfdZH8M7RH
XhfBZAnoailOmCOgtx0Owz3cfWSAiypD3NyhM36kksbIbYYb2Py7F81HwnI2W3iJ
hMordA2Ex/qoqyJNcJfDXlV9xU/6nHD8JH4uUxcUWKGZrtxK4UX9giurl09polOB
X/QNLniIryc/4DPGEF0Uuvom/cqkrytFBDgkfAz/r0+bpSsAky0r57491ShpgidQ
GZHuyN0JIt1C6g+bgAXRnR0znF7/CmIndsaMEJVNSewJEFPq46Qq55WyduvP+jb9
fxKWRsSVs4n01eq8o8SDIdNSDEAJG7AYuOMlm3LO1GFKtC8cx0CoHom7vccfa01l
odDweHzZ43XRLzft8Lx9HM1qzAbilr9sKwL1H7k94PjP6DvwIDQac/c8o1aa+CqX
b3q8Fq7UceCEflba+OHAxt5a4zokkqyVwgVu/Yrgdi5U2Nnwtw4IgB/qM7EAJOs1
PY4yBgp6RYkeocWMpHbQmxMa9OIduhvn1wtsVEYuIQT/d2OhiCnalqli09FQwozi
IUhJADLpw8aH8gyWje/dNV3b+cli5H9A5GiR1rbhB9mT1MSk7eiH6DPOfAz13AlF
mK5O3ZLYx6uUr09XdryDz/y6KJOkk52VFCMy4G/lxMZ9CfDwxTD6XptAc4KFyUiq
ZkHRS7f2ShyVF+dds4Vu1DDG9ttas34K8F/f02ZnIOQDu8Z2XKcgB8vdVifIZdtn
WiYMff5fREJeMTRXMZ5sBtYS1DUNDWOJV7VCPldORnIuW5XVhbo83m4WO9y7ssMo
dSRry8J2g7AVDAb4jvz9ip0Kmx5GZhjsP7+Wc/jdWgeovThXl6hM2rbO8R97/t/k
GvWQ/qjRl/0UKhzPBbu9/SGBOV9UAAZQzRMPI2917fyDzQzBx9/w6lCRSFFVOofc
aUGuo/nCO3zF+ofXAa9tNENoNDKq5Ag2Mr3Am4yE+xKLKus/WMupqZUtmAMSkAG/
rFvKNE0XYkwoWi9HUnz8+zm2sy+I1ZNjKKjUXOmcZN1b/4cj2PHX5McuQFx13Wcf
dnfp4KV4/IfQaloW82ICs9nLfDmr8ZoV+eU65SY8yuXmfSy0mcnVHWFfDmyvs9yN
J7dVyp2k1UTezKlZG+mvczpSP/YYuBMpGCUrNOcvjEA0y2sSZ31AJ3lgIevFxOFm
zEY/3OYr6MYEnO8lj15WHAspx9HemlZRW2Am9K7LnCaF6KqaZSG9JPDqEqzY+p5O
5w58A5EGvZUQq1ZO+vL6jWdlGhxpWIHkxpqXd9hCQdYtiCZUohr8s5xchWRyKkOs
xNxmBAqlOG9/CRkUA/u8yRUd1uKfRT/p3vgG9NiOYaZHJIwohplTtMEr3v8qDkQS
ji5QA8hEAAtn1hM6u2JKTaKbG1bqWN4SLvJx1EjbSiGNy6g9Qb7NYCTNFnXIQlz/
eYAxjbDs1cdYNwhD1lICEB/PAqacEbfBS4OUscy4pXoz7GkV9c6WpfGRiN0fAk8P
Qpe5VTW4+VrtbtOy0MiR9BXxkXov5zN+cD6umGN3AydwNCDomUuVvv4/De7MIbuA
bfFMCLM8CKwDnN2a/v5ZchJ29VYn7XVYLo6ZAVMN72uom9TzSqPrSpCML+DVdO5v
VRSbpJLyTvVpEKotfUrnu2uC6HI3LGH3Qh+OdnS2VZAx0g72GB8GHmLCo6KFiaM+
lcQWQaJFJ4rT7MO0LlyDjVYrxQPLn/gaiAmdOPnHR3g6SkCeZ2AehRbcSzZEPNyu
hCEwx093k7wxAUHxz3oiN8IF8fVWk5Ah50xysjAT1IXxABG1eWCa2h5x1rrcUomM
yMKErXZ46Fk4C2hj/yiPPTR4JwanwFIPmFo+wDJHIyKvl+6Z8My244eVBhwdf1nd
R7nddDS2R/fplpvrliooBtTfEi0sdRkysMDxosdmdjcBPrmFV6tgKf36E3b7bSGE
6h6ofRBdwPxZRLlQpRDt55m6PEO19iY33CH4USpHpiq4f1DdLiLHTMOaZUqbbEwJ
YACZMibINIsFJ6Jlc2jHqnjOPf2heqrGRkEblREisoEdYYAWP4vTyJAAOksdPsXk
SCYXoKcntkuy8ShjY8ZmrROQUGcccvX/+kzCygVRyZ3A4qXHGToc/EsOeO7Mbsww
hmhg5LudXm7hmoU5nTIZBbbsHNKoZk/yCWZ3fUHaD9yGuqB+UzEajbaVAWuNKo1a
kGGlOCJ2rByqjYOkasfyA3bsgZpHWD4iQmxVeZV5eIe+tr2zff7JhZKHc8aywHC2
IeW0NYnnWbrQKOYtCxBGK5UvH3kcf1JXoVDEXWZZ+/0qjNHKCWAim76daU3yEJ0G
5wuIuS/5iIZcbLeCC43sbWzuaBgzQOCvx11Sp1BQTCpGK7P+7sIRncFFy1wT5y+T
hoP8pbT/y5baeZoUF8fxPc/G7/DFj950Kb4Cw+uV9NMgX2hCTPSlCv+8nnegkItF
UqbTultOyj6X7sQe/2eRk5fta2mWO60hbX86ORmxi8ql+p55vYxSx1WfEel7qUzx
1lJSZNRjrPYAjNlVeuNAnVai4l2o4cDCxxAiz5Ryg34E+tikqC114FFKiPQ7Ac0E
feopAqy9dtsnhZZR3AwxvJWi39+vucseAdOvnohi8VXR3pMnHwhYBS0kstbbiXn5
Z1ymDC8YTQePxlFz2MIJ+Irm3/VotkSTe8hoD8s2pcyn59GrQLguetSVlSzWYhuz
0r/zKs0ppA6rdVGwAyA1b44YJ5C99V2WeQXHJWVA+TL6Smwv0/Nj5CHe8GpWd22x
JqAnqFdLhYfwQGJrI1EpwFIegsDeV+umoP9plFyrzDSq9Y6DAkPOmaxSNQPlbMiE
GeN/66J0GkRmQ9uAny8fDOHz8SrkWaQ0/ssZWfdFetMY+jVYk0eNkD1pjMAmPXqx
mWxkAwcpmCVFC6bZdNxMrPbLUKIPp+mqQxIKyOOxnTxuUJK+KBdvddNjHGXvXZ+n
VyVvd6+jlmPrnL8sJjaMlzmYLt41om7j4lPDwvswjM6+Op7KJBqZAxR/K8JchhPh
TgcVtUxohiXIV2DYTDY4p/ADyqVB8kW30PtBBun92DKW2AskA/KCHGCbj5ugBv6+
mnUEM8Fod8fjTocCzdlSiJwL4TcpMcbEtuHxA3g6DfcTmytdYULqLLX0skB5KDnU
FuX7xoYSDCVldhn7UaParDQ9gt1Jkh9R18OcLtgCPe88igCsAVTX6a7LIaWnUqtD
cj13rs/hN/xGzLMRdZ2Y2istjs1IgZIkYi08HNcl8qmK9Rw4znLvSKGuy6aByvt2
8FQ2bpoL+aoSruY8gTZMvAmyNmadtPovKd2JX+JGF+V4KaAJDsqsNv5yIp0geMcG
+3EftnlbqGZx2rsH2rADeIrcC3yA8PGYLn6SHaWkxdlhRf+5LeDgt+LcEqKEheDO
KSplhCXUDx9SCA8Dnf7vx8LsqiTJofww9IlBalI0Ch3Ir/GZ1LVsJR3yDqmZQfHj
/WIGkM/9gaiGRFlHWues8zO+mId7M+x8VUNccOLrwrjjcVksAxnRSR5C1m0OnUak
4oj5TnvC7pNz7hGmW0rGgPUhaZocyrC2Jnc2Uc7kSbpxWju5EyMQlvybJMIiyhoW
l8WXgTAiR3c/zFMta5dtRlU/F+RIsuP/c8kxTHUdv6t5DXMkRgMFQnCt8mnLawSg
9y59P/CpuOKuCMb+KxaY8kfVRchh3+DEjM4dPXQFH3BQkxXghIPx9WuvdVOPGwBB
rSuBvF272Tc7G9FzPMLpUt6Nf8i7fEqKNs/8E/J+xQvlikuyp8G0QDBgMSpZXOoz
lU1gjVajj+nBLf9WYS/7HO9OlDBRg0v5xzf6voqdsGgO5/2Hd4V/uK5V7DNlUqYB
eXuBszOIBEBuExKvzpyXpuRQScDlyf3aXM+jrJ0IzugqA7ueAIKoRRB5nUltY1vG
qQbdfBupCWL20LDPx/EemkisDIkvZ32sscCTb85DZy9t1p56P4DGTW33+r89rpfl
U/ty0fY4CL9tBKNFBe+M7CuNie0bIlXUGfCqciDTdZE0j8E3QqI5BaAecHvtwwxA
uV6WkwW/hp27O31bMFF6SjmZ4LsIaOIniGLFTWbQa6jk/dpr76kQE7//VCcsrrR4
3qdrNtDqxXMiLF3gqxaThP8MYi/nMydK72RNneu1sYYO4Co/CudqmxK3l5m1WiMv
9gyHG0JMvAhHxIN0S8p8rjQE8cB3oXBImo2OxTUcqp4397pPaa4ctoodvPw4MCz6
m1TPBVjLnRk+0EjlLl6fUMyZYoY+8P6+vAyYJ6lyx6LDObWqi0Cl3+LRvwJAqezU
W8cva2do4ez26DQw70zgI67NqEC/ERWhAxDXlJR2fqUKVAqO9bZZQ6pDO+GkKSDa
pXjG9Coe6ASIWP3oOs16OyR2X4xjdzBzHUsS3MWflBQdOiYqB6A2s3GEDwnW5mv0
zxCW9mJ77l4/BlNeHGVrXTgsz9VExoeqZTcTfTj8SRKwo6FN1ZBj2InBG56TfQqV
zJhPDW7ORYtS3vP9ASmMDpO+rmeOKs/8v9WyaV5uCQfQHcIWePeQ0+VI25/6Mk2n
8ypy8l3uGqsvvTqyvzmJZ/nHY7UvIELMADDZg01JxuloR8urXjxzzK6Pm62zcJFl
7IZ1yi5Nn61+/eLsJ01SGNbnzxaHx1V3CGxZ01rlMGRDrNpJ6NesOkgypXXaiTTe
d7gS9vt7oEHCMMC8Rx9VgR5YY0CMM5Asp6mHb+/RGodjnw6qlnUKP1NYQF+3krl4
bTbilgxvUEkUWqn2ct3QmwpDq5P7SzbXQJpcZLYGoE0QwDdf+uTPsREeHfCSuQ34
B1rXkhdybM6D5T6dWSNP7nv/d8+IFCS2bPhe1QklO5hAEDhmRPmLyR+FqtQKJfPj
raPzkLK9U3mvijthrja+yAAt5uYYAh1XQ2F+79+1d4n7EvsquwrnSjSekRkQfr9H
pN6hNyJ4h2fchQHn4vQCzkhUpreKADkchv+jvVq6hy5wWXfZr4W5WAdSqAbOLDi2
1sObRwVfyxXeBbqB+0k8lZfUJA/V8PabkXnzUCNvBmhEamZq7EzY5XLoA5da2lhA
i7/1AEEl/jRd12ymLejUdrxHBIhBz2hEskuurslOSC38tiZYm61EOmkFvtBT/fbl
MNJ4aKQNhZg4ke0XGpiOPqjUgl0jOhj5PE+zRv4CizqBsG9P5zXc6uvSS6grNiM6
2c2Dsgvqv52z5sXwNLEGAQfOPcUl1Nu+/ZrdhNhGX/Gl1W9ZqBRRgcv8xDSx2b7t
ykrYN366nHCjMxf26NEg3nNzIQTDgF1HmHmV0CWHQdwtgm6EfMaPY2qXY7ONlWtJ
2cz8l/51yBPuLizYvKX8bMr8J4oP7T+Dpz3Iw7k0Hq8NeiT2GcAEcty6qw+vTUcq
04wcVZwNtAPyQRKaPAIKDfzEJdJwmZdpdX8vFeOCadVQxOXggsk2fA9D925Db2oF
xJIu6I6CW79ymFpO3JqEG3pB3lN7UyQiirzAWNWviPbl+BUJR6/ao8p3SqtGqc4t
Ony669nmVOOFciFC42bshLgLkOfRCSaZqLBRX0rcfEH8x4zYvtPvdE6XbRBjHJxo
iRdi5gxHSmg9XnjxFqxi5gTD2ttKYoPI/PsThyK9dvLR5M/6xNY5xGDnGK2mx/80
MGFDpJbRyZf3nZ0HTMBYZ6Db2bseyGN1xhjSjVR4Zc57kPck1RbLYQ3782ta3U8S
8uHf0ZeqQd7u8wnkib+maMlqo5Z2kjgigfyuwyyFho0ZuA/Lj1cZRjUpHM8Tin5t
FmKgf8EOLZBsL5HSbLnuehI53rOzCZvJo7pMpurjyd9xcUUXvpfhXSLuC/Kq2lsi
4pRHf7m3Ecvr5m6kH/sK5peO39bmqapI1l32SrxU2i6pa1fNPd/p8yTX8rKXK3wQ
1LN0I2iDsHbCg9Uh1RZsYRV/tbV29RkPG1AWBdSuaWl2pWNCl1Qjxr5lX0EIDJ7D
xkxDgYn5JY7R/rtdzfnP0L741iXMX5guIsuaAtcdgfMymbZ2hZXdP9dIOGC4ndFY
8NcJpXGDLqE5Au40/Z7NytEM87aq9S9iHrRxsL395oB4b/POgvvyg4TRWCG0/TAk
yLqi2B4iP40DwTIFRDvmSLX48NtKhCwL9YHkFF8OS+bkSpg79hHKkfNaXto3qB8D
ho9z/epkpPxtvBWT6eIYaPsL1LO1Kx/dTLmH+AyNp5VdmBY1MfQNA/lV5E6/BZ7g
966PVTFwFWW58jZyUv4NHcylnytt02iJvkyk/GCDC3NtnC7dqPvTebVVJgvEvp2v
rsCdTjQixfHXg10vzdPw8QpvGxj9JlkJwnVEsUCLcfY2n8QwkvvmfUuge4LWJfRT
XKrhyEwW9PpHA+4HmEMwMzIMviY5bkQp9pKOkh1aA6gHgDTRU30TzFGcCD0V2K8o
x5sO++TCjaBY069bCtbM9b3QkgTPdx3hOI0uO5F+HD8DsKcVWX1Qe9EFqXxgHXwy
NuHUFEk47lfow4e2pzIJs5HXNMRtzagLx3+rEHwRCTO1kIq+qNpKQK2TLenrdn8M
DNV89TpDGTn2+tqgDkAAOkMVOARoE8JK3uZz5aaCfYgXNkeCrb1Dyg6Su4cLOKWl
Jquh1lbM/2pbPwaWv1TzlJk9Uobc/I0YQqZZlO1PCXiGEp/wBE/Zkxk9Uf4iVCTG
UMlitgDvQfuFCPj4geyg2GMtHv/jkjx91CtH/LwUFAitwxDKV5FFLu7y+j+l77NY
0bwDN7nKTc9q8aPDcK+tJAQEFzArV/nT22QG1uM7j0RHdRm4jiQiOsn/FnlasPqN
TKu/PH2yIm4JDzEJoS0fMG93Ah1JQZRWVkdGbS+hYwaN4sAhp0fVgBrFx4vU61ol
WxXM6Ap+sEqpkPyjqmhXB5drX5YPYZk2BzGuEDTdAKLHkohV7y0FnqmkH8yWfqx3
CxZkSWqYQOx61EGi9TRYy4rJK6d/9jH5RT+0phE8S60kBr5IW+27Wo6c4uQpLu9m
YjSuMvJ/TA2MRIGwoPU42JJgjpFIFAcFrlaXFd4T6vWNfcsLBYB8LvqeJ9rhSwiH
TOMzOiauSMghVOsAwlLQHM9WF4+YnTesv57nuTBF8lbmZiA4kAo1crRJ95Mrrrm3
SLo+9HprbkcZVrF3W5qpM0LV1zDaWvBHpIMr436LOUm4Nj33XdDg7QFphpXSnpv0
cwwuA5PmIr4lccxD0exIHgzrOBvFd+Wp2az6+uMlfnj2eQRgN67B2feCxBZmlOct
UVK3qugvzcQD8545io9sKIJvAbJ3fLdPmjlYIPVJL044zX3ZewJLyHaHzG85WN7h
XjMRs260f/uf9JHw6WNHLPLudooqYIIt22hG+1oQD+4QxwmWboWovDYpCPEqx8Mi
u6Zb2sM7eaBCacMGNIIrr+T3i/IS13lUU7W6cGNvZMiPWUbDNXYuODQ2qU6Z/FK7
i2FvaItOmAzqgykc881W265pL4Uv4/qZxdT+47OOAJ036YNFM44k7LQ8YPoD1BQI
TYRyEWqfEeS1GsrQL5BscqMSHPCDECPndCPQTlxjv4bdzFVCpqAJUsQ2hJGJlnob
K84qvYXCnlHQsluySzT34ybHXCzVfoYo9EcFuIMuHz1DvtWk4NC8hz+b2B7lTb2W
AMaGwyiZbAq/ckXz2vmiSaFPBQiTjl50Q/dKnlEa+YPoAgrrZP2vGibg3xv7t6lN
Cah5KyVGfTZmyo9gcIvYfrhMdIG9PV8M8CKe+0G1MhgAeguIwAwqgWPcLrWE1JZ2
Td617O9dNZoewIU8vw1M4uf3xbOSVDNAVmyuSPtQuGaFJCNS/U48i6Udf4v02r29
KZkXioTZGw0oflIfymvmAMttjlYJjf85ZoNJxIksVdugXzzQlCZ/7v/ZheCJDaox
LF9LRw3024MpsAQ/famQyjeekByv7kSYCVD8rrmZbk3brs4ai9rHIoCesaqZHQoB
QKtHbd9/IiAheNJRDu0i2bh0zX6Cm60rKRK72wdc5H6qNLqSa4bps6FEWjVS0no8
LNGb0V+ozgBPpEl5QYBgM35vEDRmdKw05B5bgZ9LAcIY6hy71o+OkqeE3HzG1MgX
jJ8dxsZ6hk27sW++nyc4rA+ox9BCIL6jgSlFkk6irl94XQbEY5qcqMlwNOFEaa5g
r+c/0FfcBX2GjtVrG/NLQr6gLYLsrJUdInjM+IR17gN1qZ4VGCr2B5qNbB8tq629
8AMASGiLhZrxnso+0Tpr/VBo9PM29bIvGtpjHSWqA5nrH8mGf1DYo50I8ooGjwgL
u/CnHNj9w7B1EEw76e9kaXxjEV2QSC3aPiepxWvOHLwF9m4P+SKHHL2zGKF0tAN7
OZZYV8s2byptsVQr7lrsHdY6fNeKs2hWToaCftfuf4cgjAvNnHPf+Aj37096MHIN
ls+95bYYTz2/DM49TnCuXx4CkNtfbeckVH+dtLy+isrTxra69NjIBTpSqgIEEyir
sm7OBVi+dWPyFUPA/g9zMvv2PXQ6X20zcky/Q8sGx/eiF7fQkZQf8MnCMpkmaOdq
akij9OLlQvW2PWIU2Mqc31TkCVvCEyQkHws365eYQv0NmWnIh2VFPX7ZHG5vNGz0
VEtbkhq2QWnXOCIq1pV2L9iOOtV066KZQJdDcMSQ385p+7VsW3Kh+Oc208M51eSu
th2MoSILFQIVdaC0LLw6vAMx67Hna84A0bcOPzfPutU92LpGf34t42/sTKo+luEg
jKuLd0rz8zthzQTzSXDGT+GEXVhM50jPpqEVCQaz04bvTGHioRDo+vkvfpqt+U1F
iCkUgWB2PXc7GuJxlaMzPm8CTlDH3Yphn3uiygYykUCuxSfZ4OiAgriI0/BmTpO5
0WKeZ+Irmn4o6unH3QKE3vBDdHQOGj5tnuOPxrR/L1PcRP4TWZWPii6taYKJcU3Y
YFXmw52yN8diRqaAq80H69WBFXKP54uAVb18clRGgbx+3tfhNhR2ahj1hiOVz237
iTWAUEau+YpqUbmvkJq3JlCgMn8ejGvDnfEQ+vODbKIWkXys8IP39FH0dhXk9Jk0
oLK96LBPmdsaDEVrvRd65cz6bC8KbMF6+QvO1/Dg2sHvZL9SiAgNAT2d3nXDnk3r
6P5j5Fds6MfG/9axW8DQzUOSFJCwzryUFmvmjORYkdGFZ07wJrovYvWUOxnbYEtj
WKHRG9nRb/0GBdi3YZkNiE9A9If8Yed2/q2RP+wQhL8X1gQXYL3on3E3pbw0eBOS
NHkNn+K7Q0VeJgzKVh0Mtcob8YFhEr+ZOKObFXCzh3VuWOpyJhib5DX+owQjgTY/
ot4Ram31m3nPoAjNsuvwkWkwlE78M2VA/I/fC7JtFfb8Zj1FWaINFfiwg0itAPDh
v0fVj53ybKwDe16vReGnfejADp/xa7Y+O/4SpOrYGnXou04FhClah5X52BBb5/kA
K5q+wOUumpJyb85hJwW3TyQEMt02FUdjRdpQraJcJTIK4Bwi6pO9CATiTJdojVP7
by5ypOuq7eU24N1uShkEW8zah/ZzSbmZrdtDzAOpYP5PVqRHrjk9aNvmPM3nGwU3
qJhXwzpjv5qVLxhM35CktELns8zK3cYFJBCW5xSBilX87YTtWwI6MTlDqlZdoeog
M039LhExFn9SXS1dZfpPLSfvTDWtXlWJOzfPE3QJG93nZFmcUBggYPBmXOFYooUh
CQgdR/AUdre5lS+NvlXbTF42JipuWuzomvTJZ9yTtssHz7MQmfcCIbq7rSML9y+h
xYIbiNl6L0FZtBpYpmAHk24UAOJyxTyFAlAQ6rUXi1DRElcaUAlB7nMQMb+q/JFK
T5jdnd2hJVZL2nc3borB8A6hii0k66pvCtTrlsfkPmwqoyxWfvyjZiMFmu7LPlLA
cPZ3aJERpEEzhSVp1n6DbLkqIRuP/mDhBm5mJ3ri6lbtyTZ8x0VA2JxLfuhKGysN
qqdN5m97j8qltvYFf20H0KJl3uX4nHHkr8wt8RbBEFHuiM+W9XuhvmcrqWepA3MJ
/+W3pFIzd32nkYlYGlS7AT5OV3U/pcY1ub4vgD+rGak5Vo/Z1KraZktVfVIO4tds
niKRawsKgmyqhzCb/lKSmMVNxG2Da8JWUwVAM7/0PUUgyxGp0K0ebg49l8YuwQrh
iAz+ENGRKku+CzO9eyVPXDMyF9cLCivUwCHIeOyPfrDXC4MAC+sF99w/0hs1tU00
ngqaZZy5yodQoXIOr6RIiioqpP1G9NQ4IMUtFRAhc05w99JikaQE/rjqxXu38yFI
jimy3HSiokwH6NdAD/1yq8VLbc0g1APN/e+uG9QOwlABHkGe9Xy4QlAbDtTq8LT9
cJzGpf18P0g5qLxKXg/2blZZhaoDT5UPQo4wmUDTiEnsefujZExvUSim3pigZ6k9
lH3gXiXoaR4PV8U/Rfh3b1UVvKNcpP9Kh8Gkh4R2QNaDbGXImw9rP9zAt2ndrmX2
NZEK6+COrWBIZGBfhAJImzqLhywRYDsUBEt2NxF/+rmXaayyAQKQKk7NDV3PF3Bt
yUfZb7POa6DyF1JG/zPUjKOBKUu2shDAFFiz+GE2Vwl4MMq2/2PtOLgMtApfgVi6
GQTS+2OREpCicvlqyzEUoCKQ/FEWUIIxeb9FrZFgTWbnytz8+2adaD55pKIDzbJU
Xe3qvJ4iEqdMZTNZ8j+iW8MLDEdvOT4z/PJJlbeAaR87vZOHnX/vtNbD/ixR0EAG
QKbrI58sohoktku3i91/iN28InErQmp5s75rktNwvfwWp1oJIWFctZWHzUwiZPyu
5VweMo8Lf0KHtC99xKqCZJpU6/gMUMMCqGaTTMZuq9+l3ZMSyPSkgQwcVkfAhPPb
zOl2rnYvXhfVqXX96deIktjYMRYEKP3iGybGQ01pmSP9Lxwlfqsu8kV8FjCVqbZK
mD4/r0rtC84eFMeiyvU+xrg7gQ5iHL/BbJFDmX55fIaL5MlXS1S4WCrHAmUxI+eD
Lm+2YL8rvhJ1AEaQp+DllUfb5EkzVvG4bFSY3G2DJVO/aBuYh1+739zQOed9Wgar
0T94fbpavJOP/uH/6nu1FI7BttUYhM++ERIqZSDFGmnXh3UlBKzXM2ok8437qAPb
qZg61Je4lqfMP4yyEYbTfgc+ql8fDHBANJHQ4w1eAq9prRTkLJDoGX8lzuUxzWD7
R7xgcIbD8P52hc5N/ukwTPe5UDf/bE6g6cPQ6vGZwNFIz4F5x0gGUE4XzOaiulBV
8k5vzLBmYEYLKoUu26rBNPPh++EsYUKC/BRp5JDwXr9mZj3agOwiWUh5ONyVji/w
kZBQluKTApdbvPjkb0hHQm82sqt01T2DbjFQinicvzz/gtxCaCpfSYzC/2xesG7e
ZJNAdyX5EMi0X3Ch2N0/y0UchfwCY6fe05NtyyHt3BUY4QRQIBM4WKEaRWJI4h6p
qjGeIQkmhliSA82ufyXnvJhkE+aedDL0b+3Mcijdc4Z0sTiUyZcNNhFugl21xVCH
y6LW3QNjEOZtY3t//SE641SzsTuy/gdqc8B/15ZWrDHcDAoJCaMBU5L1gaPFJI7l
8WetlizRXA21sf9vPj6DdqKw+7l5YIxkDN60i2xqJ/qsJ4ivDPGB9CUTRGbF6fEm
mOlZMPucPbMOZsRr6T+G+52e39md6NDwAiD3pV5IBqif9kMFLzX6Y2pg3o5LDLWS
cVtZsKkw4P513j+3iDctpPKjuUPzT9L0AbJi6eY/BHTGAGiiUniNkV9yNhYQ0JZF
WBrmbmMfj3YRagDPNBsRTgHL3kJX4thfmePRfkc7oBGOmFCxCbXwlvoTPs2bYQqN
ONVNaoevtVB6E6RpFFplXbjdaGHB9rRQp2bwD9flqe28/jJuQWgeEbHLih/hV3lH
lJO6Fa1uXen4SjTGS158kbu3kAPT9KOqVpV+aSd0xAuNMiOcfNSlIQlFrVOdMRe8
Kf3H3YQCAElCWLtHvm/2Bv88Ns427TG0Ki/d4dL3UBL+L3UqtLbiiBTtYh2W3ean
QSrVnEaXTG5Kn3WmERw7AlWdUar7zYiFlgBqQGbcm4XvSSUuFwHJAbJLZOK6jesx
H0y1dSSoTxxI3yVFMH8G3udhkAdZ4HtvqRjKBtg/XumY4MiYgb/0/PUl+aKX5eNY
uYDrz1RWHQjGWYXMr9Vgk/jpK8WlJQ1hhqOSD78qoodeyd7LtAoEJI2R1d/Mblf0
BCIvBqbBwYcf1zDY5cd+0prCBO26VX0PUaeKU1hghjScDqxZGGLDaL3wj5PjTKkV
l6L2RITpggr+RxVPWJMUbxpErgmz2TQgCaNWm86kIjRjKIucnxfRZdh/MRpxkmrh
74oooOP6ivT6Y4IzGDxGXCqH9rRa69MP54He0w9VcSbT80bMpw4enpHCVExfTiAF
Yv/LZMhdK3vfOdY7TWZXYMY9+VdieiIelHItpgFwbBYqEKFtfx1woSGpvl2wrQ6E
YXVHTrqnc5IlecTf1dFhcz1zJusz2azyDCiQ4BobXDBoNEpzdwzaMRJrHYENKV7u
E/1sZ7xLnV7y7BA4v86HyzIV+c726bTh61HwrRlVTxvmyTJClV6o8b6YLWA9kDc4
f+Vs2mBz8h4cJvjILu4TdlzmGB3J7xh1yEeZEJjbnkUMdMH5XCv9FH7aSN6+LDNs
iTKKu1dKqev9qbiVoNsHySHEmT0LYQTNrJSNQJ2azHta5Dv2uSfOJvJz2+ySwH8T
Lzi75RU/hzzfXjmyIz24N7pXHs/pTd3Xe8JHE3x41G72Mv5QbsQqnwfmSNGBl/rk
lXw/qyoa6maDEdhCNmMxU5SlKJJiI1JSJfrXeCkV89e55sHvhg2lzlEpZADSSmHO
qqXcz+pQzjQPEwBFzIbINTOvz2wJwaHp+4ai5glV9Vulu0uPGPU2W748coF6ZMdT
fE3KSs1xXBZn48XFv7uCWwVTc+GPH2wucyLRP8cncdUsMe33aqs3sUyIQgaX8j3F
ZhVQ2JpHmJdXS8I6Urb7uMibgYoC+nWF+Mgh/nYl+WEjCPisoxUWo1SxJQswiI+c
P8LZrp8QCRNlkyO/nBSDft6ozcoGgpW8t87aTjz2deQAnJI9Z7L27xDYNCkdOyMH
cDD7PT5oud719Lx/+EYl8XMr3ld1hix4aZ00mVgBtgzYraJyMXlBRIckCanjZVjA
XKJBsGdkMn6jyxaH7xK1Ho8nxMyTNhgQHAwmQy7Msf+ENh4cOAuGwKdxi1lTUugj
mCSPxOg+PYQ/EYBTUe1yrWy7uPu6XLzhPsJszz6TwWZqwfEz21zPongcG4CXL8L+
c9A0RdjwfP4etUAnc08dNgpNkDAmM1TWyMFoxGwSIQDyxG478Ih49IFdlsvHqkNn
Jzp03ehG1OE4XsXzmjy97BI7fVK3fovM33L4rZLMbO/7SqwAQl+QqNlvpbmEQcl3
jHNmSdovu3jjYYrgSrbS1btehgKQCI1dBQFYxp1ln6xdM8BjC5mjbFza4FbusGlP
ZAyQcI3ATB1WzK6GEZ7Kmj3+2U6mCuP0yr9fQzczT7O1sxbCPWMN5Qq8lSM+p774
IEhxLU05jUKNve2K6azkyaAnQGtLw42Xn00hKh1++WjqMzQTnUmz4XlDdzqweeVY
EFCtaMBhK/mSCDu9Qv53Pbx5oX3EFlCqDEYvy9sKo3WtF0gJfKYaDtypt51Ou0JR
Cg5A2HS2ZsS6gwnOigPyKWA347AE9GqTA6ZtikdVtVFGgVhynL0ipJUfl0f766ov
qwXgBF8+Xlo0vSlspLbt1/buuoe2rryjUaVxMk+MgFSY3Sf8Dv2xS1lYVI3IAPk9
YpupWy+B58YmZO/5CaP8TVP2cfc5kNBbZeGJjsPnh4vjDEZpOktNknc5ft56Caz5
dlpxjdD4JTP3W7ad9ervPc7i1X3XbX2GPNeynR9HngBc+mYlQWL+YxTvyjpw1KW8
cufz5XUrKu8HXhS5O7pVlNasHjvWfidJwz7FP/w6Udc9ekUoxLVX2fZXhseQyWZC
bG0bZEN0MXVynHlrCkxN5sQ/fSYRb4W7L/VlHvCuXta6BjE+mB83ic03gplenlyL
Zr/nTPqGS3xP0ljfkgB9d9DsmgClkpqIdgbZ34r+ARS6FiL9t5XK1wn/RxOaLVQR
7qLmA61MD/3s47X1GDXv4dE5iuQwuY+VfHViE7Mb1Rjw84CM0Qi7T1k4c+dTMm/Q
jt+I9DuKJotJrXZXo5FDaGHkT1+rM+OVscERWP8kC7eXU1jZnM7AhYoeDBMpwaTA
LzKjbcjtpQOMfDl9pHeU/ZAixTst5VulNJM7SfFIsDuf/ZwWa29lPTlylH38TOcd
dpTPtY3cuqKCIDHWAtK7yYFPp3v5EzLaJo0JdXy/0I5mxd1tqqy/B7uLThplk/lm
EcxkfVQQdumbtzghnzkPelJ91RQOXNYtwjtaCHbU55UXdUVMLLzmBbyVXVZQn3dE
QNIxRs8zeyy0Ig/pKofK2zKLjoT5fA6qhGzrqiY53bbOrh9/aFOO2FUYyYNHA/Vv
mSnflJ4kmYMFjM3VGEO3JNKxjTIP5ZIxcjwO25TIAQXQbayKFbhHaBsZsDC1SIHz
TfsqVVaS2Ff+3tO0VlLLc72cGBfJxndrcwFJNJbO4z5bioyH0O3Z6UFzvEdRgA2P
12KOe8jol0a7FBA+o1F/GOcnHqKa5vWrlVquM1/jkZQqdv9JoXAt6QflFqzBn7Na
P4ryExI2xHbF8CiXt/XWxRmwjaPFHZKS7B4wa5Dq1qs9IFFPX39Qvr323AcxWeoX
zADH4YmimXlH53y1Wt81H5vgFVUlqe/bspTuVaD5jv37bl+Z/nFzvGRVPTMw0XIP
OhQNX+Ane37LVU8F9VnN7luoh6WvFbnTPROKDl290p1/TFW1BbGJS68C6DODn7Mp
VFK4w5rggMtnDDWn81txJmgOwICWE5SJzjwKhRpjFwbVrVkSdrfyNo7CY5UlIxcF
g7tm/PPXpNspqj39kX9jKM3yxqadSjC3Rh0YxhErAtPulI5zBlWw6AtBnYaEVY3i
rcoSMhg45aJKxMfM7gOtFBw2f6amD1SP3xrwGSX1mW933TvE4a19LBEMYiiCO8kL
WPCy/AufaukQo0S2wwLqoDjg3DNmbHQLd8djc9VOnzPNSM7Pizdl3zMriQmahcYa
DFCRtA8HJTgd/U0eeTesFkvnaMfBwND2J4wWunMScLR0NCe9K+36eQXzhu2FIBJC
MuWeXyYXOyfOA+yUCnJ5ERoDHdq5pfL6UxrXi9ujGEAsL1d3EXl40OxdHa6H0uFR
krpil7s903/rqscb/bM9uCrNg4cwXSMulgZMQscyBnAw5Mfr+Kg0wlOybASAjiiz
kuRE1zlaqGK2mWuphVSUu2lT5LpzwdHWzZof8Sppbr/UPH75+NIHqv2zg6OQdh5K
uEvNz8h1Q9dvISox2yD/3g==

`pragma protect end_protected

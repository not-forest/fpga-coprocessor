// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
A7RKd9j4Hbs0VaU0JJV3pieRuJvAm4ekPKV4f0vjitWtbnJO+RnuZaSdM98W2JPWdxRUaGtXFdcF
DVrUwYJXnOd5w6zBpqzgU4GwPr09ux3BC6c4APmlCmB2mA7XhkxGWUewSrK9zbT767OKKoHhouT1
FRvSeEkfmWfWu9X4Gvd1OTq6n1nGs1Sf/BHwkMBaKvAAcsHKQ1YKOoMM4c9n1eiELfjL2+Xwf66c
xtmgsWgj/CDgV5a0dUddn1F/U6eVwg4tcdq09d6TIDPUSzP4ZovrtocvlTIT21BeIUgbDO8xMp3B
om3eLJjfIz7Yr5gnOHFF+x5/RymKPh261ORrGQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 63152)
DocU5QCeh1RS92UNxPNz6Er2VBUzl8COy5tGGVg/woYCbbEElzfuoJBzRLWOwHW+Z0gEg5fY/gZf
hiUb89fKBZbVqmxoqRIJHYt8GOCj8FWKWm7gPn0SEeNtNN2QWU+MMNZREOFVSICrS87VKNTtKEcc
62kvSFLzaq339S/o/K+XeNOEFF+I3s4HWFzL3/VmbbEARxLup8KjLC6RLd1dswp4rIUm5BmKIxtU
SnlUqfxZcaiWMdqzac+wZuRxH1Z7J28peGgtYsetlQf+3qKbXz8l+LPfcZ9Ik2AcDWKdwRsUISOe
oF9utXjT4eLnMlHV/r7QkRTAHktuZOEchWqITPy3iyirwBuE9ZmGFbvRlQ06JmNWvHRLCvsQRQ8a
wsV739Yi+NEBQo6iYRaX7FtaYD8XJT7t8daHDM00TTUbDjETMFCybECG0MLnsH4PWu+TH31OA1A6
EXKP5z/7g/uqpgDwUjrXmGA6c0DmVe1ro8E5qNdqMr67DkmvsBwVdIjMgPT+X9emBrXdwulGgqxC
wVfQzGgHNXjJUh4mT1ahylY5pU0bUQPQf91PQBJWHr4vexc8FN94HLpTMvkayrcpMsG01+nkZlSY
v6f7p4umqptcl9eMlT147WbwthkGH0diZmmkUQC46lwKXd4ky65TKQ3wqzPHrjYDjDKlp78rXXEr
pUBAp2HQwtItVnPrfIRtbIOyJCayK+K8q6m5kPF11QU/67sSrccbPxj4LYINZf3N5aLE5Tz+a7To
fFJUXX9ni2VAc9GPYakQ6rarItzoWs84VH0JPxsjoGKHLjWTOlsH8MOJ7qEIPjM8wIWiLMqqrpC0
mJpvNgSy0Y/JaaUSbhmXDVz1GpIB0GZ+HKQLZtLVThfW10Z7F6aYQIdoabuiV9YtNOOEXoNnvH8D
ibYSLH28f9Y2Csuzff5ZZoIj4urDU9lHHhEqQsjhKuCvcW8hDbIbsSnPg3i5i59BmN9ull/Vsk44
b7HcWm+MmOsNIwgYAqLxcO3IuJxDtw+Ol1K73UDgN3VBYjBo4bBh3SDj+46VtMRGDluMj0IC3ia4
ZNuJ8N8APMydLVpahily3vIODGNjb3qwXCsqeoymQs9KQRnxTPHxhKkkdtiBkHU99V4YBt1n7+3A
05qz/OjS3M7K3PSDmptQCBX/+Rwigur3x168RZgLgYkpOe5dMop1dw6b+Px744+spIdHpY2fquhj
KdU+jweAlS+xGTZ3V28lLxbvrpzG7+sfocpjjDswMAVYcGZuWlEbkn5X/dMKM8PD7FmXVc9jz+LJ
Cw9d4M/R6uR5vAX9+wFjIF/jmO+lE2vZtwkF9iP20d1QmCxvnh6J1JUmW9F093699ZNe+pzTHpq+
0C+ozQ4Hz5IJdecSMddOHyQl+LMNwLEJfDSydixRfvtnGnI3G30irSc9qB50ShijuRtYTQTlBL6I
R5qHnpduFRB5JOYNZjB4nUKJ7Qjc1nZIOk0HnTFPJYzkO0JP07M6gCj8CUiZktpa8GlwhgeqSm2B
DmtAH0uJD9L0moDAmKkcUt1wd/izbarTsOHN20aj6WanskrcXlB+VI3k+bcq2rbjBULH0ftEVLGJ
oZoKFpWeDgauIldSXlwHHNF+QGKaNTJFZ2WpABXWVpbr1fgaOPgt28oZRZCWq+wYCNVcnpxRXppK
SmKJjKUz4zXZ9gLu6bWBamXXQelQUq6JIr8qfFjoO/IQ21kIdlTNJX+2/Cvg1o3QvYIRWagQSOYP
IB2DuyFqkvmKkBck7Lnt8z4r3PnDzp62o48i4ZOqXA7fP/AKWRfTKjIaUReK84Ys0aDkEGtPFATB
GaK/EnYUhb+sbHkGrvZI9zElln4xymIk14rtMLLNT0Fst0ZsDNAJrRiBfFKfC33rAWDSRp4sEfC6
neYBBTjhZDVeGZCsjNFLyG/2wHUlu6Lam4Ike8mBFSUNgv6r/zmO/Qm4g7cfx02Z/MlZNx5l4ZEk
niUq4i4QrvPPbALXtH99fY4fhL8PKfbwzE7rFXjEk444SWYOwX8XJobbzwv6KYu2JmEzaVU8r7kQ
KFW5KONIRdc42mMRgJ5kareYRe7aGWLzzeoO+t+EAKpHN+ZG5gfvQVBfWavLZhK2t3bcnJ19uQpx
MGlp2pSqyWIUDIcaPSzypuCwRTkeayg1mrkYnDsdblYvpbPpjrSNRiXPPBNUMV+u2XwGq18RHNQj
KNim74oyyK7W3fiGEnUEe7pKrnPj3aVK3OcxSIBP9GDskel8WiMXYYfUFaEkx+OXRNg8PDeNN9x0
Ns7B71BKlR9nSjcq+0rPzhRWyVkdzik0lNQCzkqd5Y/xiCQGd1fD4z9LoMB4ReDJAINFzAuD5dZl
lYUwmgTCzlPjdBzfBK0VAVKKLv7Y6mhiyRdAUVLP49T67sjZ5zGjjRt0Ctp/GkeQVy+bkajtFCj1
zkesHvdxQrUj3vbWA37kksM+Ji9ZA61IJHfEwriDDoSeeWSdoXqR/fPi0vDJFKtBbkFBB+3kg0nk
c1UO5FSjwJaAYE7U6/0Jr4CwRFWLh/EyFooQ45mRcREMKXxHGkZ0VctY6gYPeXwmCv0naG3M4EUn
hlKj9t77HvCJX3/0djRrF7gn7/4NgsANoHW+M2+4o0SLhOjbQfuSDy73KWs4Nf3Q2jgGkmMqtqaP
0OMyUoer5UySTDkLUvicuyUoP4d96AoUCW8UCZ9u1O5bbSOGtmX0GKzfeYNJxSMQAEgVOv7PeD2X
Ccr+zwlWB1stA6nd0VH50eW9y3qKKAEFV+DCXB/ziQSPGiDw5UuNiOftXqiQnYPwCxYyV5z/RgOM
a4vsqn4im47RZeX0kyG6As7JxROh/6RHoFhevI/y5levdQ3oG31UfybeozvSZ/2KGwc83+u2OMSp
ZHhMjMCm/VDPFUGKaUmju79sxd7pOv8lSltPunt2u91bmm6i33j53dPkXeFswRnMpFitaKiZJQ6+
TMDbtqUdNBm1SId6MNcRJ7KnGMJkGfxJPcr8nQdLWxGSP+1MWHp5DrHYXfrvR7rZxhCXE2DJI6E+
Jmi8Trrgd3YZ7EjD1YJshKjZbSEPKe1es5C4+et3LZvtdI72pHMxEVXrRX7wSNl8uxv0Kx0ZHlry
l4Elz+7iMgRYeOu4OHsvVCSgXq7ft0KKroc7Q+g232OrA1D794KQe/Nd6fjWGa7ofIlaCbNmssdD
qiuhgA2D+3w28+q6mJfkJW2B7NlYhTRg9x/QCxhqWBWZs6jnIUcj7GZTYeem8iU7rkK0/zAdXXvt
FogcsgY+ogXT1kBh2uiX2r1qEqQbR9dob3M2giXSWzwirw/8TEKC7wBM0Z3muMcNqN1rtg0p7zyu
TBM4nyMjbK+kL1JfCRh0zL9KtcsuzfaqWjGBj/zcpacuRfHzBzmkHQzT5X81PH3M0xD3BpyzxafC
rRt6/1SF8l7k6yjt2M9dK+kiPVKFN4o4hslq5atk4IwtgEp6hlDVD+RyUB1Q3SbPz22oXSD8jIrt
7o68ZkbXq5Wo5rT0FRHJiU1S8uWrqicmfXQvFd1GmQeb1v0bQ1TkNZ6LUl3yk8t4NQwE+A/cxRqt
nW7OZy3fwGA5Lz9ebMFu5daE6pDeeQECPhy04yfanIVz6vibEg9nA9vK3aDQKZUISwHUff0jV8Pc
QQfDNqQe8bIQuRf88ej9ird0Ur7VNLVCHVxFRYotWK/elzM06jDNL4sRb9pvov+eI2aL2CBv7Foh
0TW/dDSEA01NaoretZot43asu9/a3CO+7wRhgLF512V0Q+CBQILPSLcIAfrDR5s4wZuTqcRobZG5
Xl2Jg5rE9DUJ5aV1J+sOmFOu9sy5tDG2h6AUQCj58ES3RDpHixnvhFGasSbxQlQjC85yGegapq1q
QEZYO1jiRVjMDOGLqGMGjES2CzIThrUIFv8Uank8pNupR2j2j5na4J7uLXo3kVzYGNexS61Mu6FM
us73KO4i1L2cQbnjcu23xt2jJhqpKJ3qKhK5xaeW789dU/KGU1zf8lykp1CMOlUsMUeqvoFZMp47
+sDBsifNAZoj9OSEnWdUNQPf+pCsQT9kmpAIRe62SJc39k9luWDiE2w2YVlsCmWkHt/XW7+5DQL4
TZZe0CAqdkxYtHdqkszGnQgJ1VFFdgTlzMuGIc60Kays/SKsAcNGagkWcBJfi0u/3DryeEJu+njv
ta6eiyNHchAcRZZGULEQm2Hcoce1kFXTi2VXXEE90snewS4Co6UsV5BOZ8n3XQJwdbjrs7Ijz2/u
xlFb9NshmEcVW4eyij/b5sJ2ZIILlZeyCmCrD0oZaMmvzqvbKexIGZLxZB/HD+CVEpMaT0lUS08r
/LJa3UCWg1ztN0no4QxmLZYYZxMvv2oeufZL4kZyww3jzSl+QJEnUK547UDYZ49lUky+pbLMLPPn
AVi4FY2ivGVyIPGAuM/QJsnIV7ffxN83XGMcgEpv8RR+B93d0n7/dQM1N189TMAtyqSnw4c1Gc4m
LPsrXVRieDIY0mEEVfnoG0JQLX2Q2/EXIeSBwvDDaj2xZ4bgvrdLBTAAF9d/iy+qsxYVYSSgHQI3
O03MVB1ypu4Oj8wo5FBP1JX+N+/7SZgHDAYXWJog5UAmiJGLu3QWTj9e63rL4s/M3nW4+KnQgux3
BCx7VdH4VcCvdFwGDYesZrq60nUkEZAcroleX9UlyS8Z9QblV7Tfr8l7c2VDdJLqsbBTMVCpbH0a
mLE0rDydPnWax6wtDny/kX3a4iVSiR0a37ei2vU5f0hCINRPinOfKOF8c43Tc3j7wL4wsfXKflct
yIlKQEhX6yew31k4LsBcvcg9CLEbSYX2vjr3rHFsbEu7+wvox671fHlDrchDg8m2lABlXAhf6Bv6
6JpBw7tZysaWOtRUfIczLfB8EwGT+0q2F2Q3tLHj5OqKkIulekfflViCHhMax05AbTTLWkZxwyh+
hQhtzz8X4a/QbkOTCxHexgdInx45Ipy5tpQyugujURWf1rAimL2hc2CzzLaeomdhe29ifRv65dKJ
e3o89zLpLAliKVQ9xICj3ivGp88LWrzDrP6PlpBxrVAnSUmQE0GSLDs4fiKByhKMlbzywRsAZ8Rl
TQ5Ev/DjMrnnmFW5yxz5WvuQsSAI24LdsGc1PjiXzpxDiByuU6FrwlxfoLnG8qjm/LUn45uEjKDA
+sVLOKIke4iUXcp6GFDJQ0zgS9MR5hdqQ3TTL/XOuSGKCgfgk2Mm4UmNvIRvtG8PqjCuQUS6dHbd
INGzs+f1q/CLlOFEkuAV3gZrSepXS+/kC3IRh3eO5HgwaCzks543jdup2PWFYrHy7W9P01Q92980
bbfymrzkrk7KsBaGGkbgqE0g3OkyJtBjy8iA9Ky1D4FVhIYmdH1T08aS0x38S8K1I4Hm3fnP3iik
UU+4YpfxdYeQFJrHdtWvsX5TL47ODPZPnnNTnhVIbvO0aodrz6OPTrrXZDZ2r93pT6RVfNkCK+hT
AoXACBK38Pel5byGGS936HALSAAjbADt8tKCoac/y5qvy9pNC3fDyPeBb9Gl4u8/xM7vTlpy/4oz
pKuSKOZaSd2xcw+rHEXAhSlpMblCuRR8NTh5bMQYjHECV/M/9b5JweABNsv6vX/cgbkHw+kop71M
1V7dAem1oPVKid9M7BzsSjPoebODm8TeeDZqU26GBQRPHOzwEzT6/6Wuu4sKDrxNTFpMhyOqcw01
NmQo0zK9BZy5X7YW/9rm7magC712edHoypUtmQ1tlU4nFHMsIylaor9MbDHjhqJ3QHa4tMzgYTEU
aynO2Wi94kTr1OtwCKnAtkB/tTJK4fDzykuuk/CHE7ui+INUmARVn6Vvb+KXQGtgcmYwyVIKNZT0
v3D4eJH8hc6BOzVrtXQCjgL9EzsRHt1MN/3kPxQSmDkdVY3J4pBuw2bUs6Xs3HQ84qwOZiTwqu2O
7B9IhgMRgeMQTl6u3zWSYyxxfJtSEMMWbFqGeGewGz9Nzt9+FZRNtuGhImo586XHZoIGflGF8RJk
k2klVnwKvZUE8KvFHds3mpIKZqhOTW4GMWZmS940Ur1H0osiHOrkirPYQ4wlKkSdpMYqPiit0Tm3
SSWWvONkMivMKx462UlaelxqYnDOaQpbPLjbw9cjZIBGg2Q1LuZOXfmlzIA1HT0NpWetkF8Jgyt4
fog4dawd1/rRL7LPWLBZxngWVxp75w2z763GM2fheon0ZGWxmBZuo8y2B7CSqUn5jCqmOgwwcM9W
69nWEITo0mY2sbusjaZ4xUkA3gv/qtZnlp4whYWSQU326p0Q3Zw7npc3jI76AetlIaxvshqqsWPl
cTlE0kiFQrjtpXe5HE5h0gtkW+APaPKV0gnVBFZVi3jFSmtXtYVfkKXdZO9+66ug+szIgePni2jj
lith2jyTDGaWKItgBxhntGNk+aO+IfTZ7MSR38wjX3EubpraC+xjT+/wDtjhKY4bDKcGnnqtbUBZ
Lo2zeVX15yZ5aIaJBfDuXM2EEi5Jywp9wGSSJIN0HnDSRKDOigPRP6g+GGh0UYBOUENDaX7Czecn
sWppvtDh91JNqYdqC9ZG4tioP1sd+RjlCNvEvlR7rGvIe/EXCo1Y5csH5nUIOz+GVwF1WCPxbzFR
4nJfDFS4mApuebkVRM7tw3f+CZrG+Po8XhWcpfc6rHz0WCFQLyVXyddaeHIxNKKVv+5ZWCOaAZfv
JUPoaaKMF61khP45VCHp45LJ0FGXFYXZnF48gh98u6EfJYVJYhAY0ZoL9+rSKjzw3UZzqbb7IBnK
7kFrSNamMo5dwGvSTJvjj5fpuRDDglAkVluiTsZ61s0s8EJc/61y3xXbncPWFH/0eGer8q10XZXV
8YfNlTRWqVFMxcyDVd75pL7lNmagHW5EonfVZoguizlTmYHd4N6Dwr8k7tZkEustqsccVDhn64S/
wmIVg8zb4/WM6QMmCIXOOUqAJeCajSP90VDEI9yrt5Zz8e8mQe/+zp6Iq2v6wgMyoRmn3XQEErnd
ZAChkxOuoZiDVs6+lcItZiFnJXLeZDaGMwAYMvG42x/+CsoE0PeMcI/XPpao6pZRIAzv6YLFoY4r
MDe995A0uNnxBEsVmw/MOir88bDrEr7AZWvW7dMe9ND3XUJ6xJ7YR6o40PDZzXVLAhSmF6QTarKF
Fux4IJdBNd6jqDldsP80OOhvdzfLbFvw5YMeKdoOsLM2CzIjGuRrBJXe4zHsx8Y9jFZBbaiBhA9U
/N+tY2vVAYDegsxCE/ZWJDf5+ZPLFVGp0oZQ3ziYSLKqP04IoNAbxToFDLHekniWeEH1gyPZBR67
TZziyP0kFs28nPp+ipVOZ8Zt76YBCalqcc8f6lCuNXN3cgqkP+28GgC8wI00QoeqH17DynRDSLTm
D3QETRtZZVjtBXy0DakuEdL4udE8KrhxTwXNUQpbxRl+iskII7kPMORFZ2ue9RHtJa/anfwu+8KI
BlBxka1UKyilKDeCWHnViwEeGapKFLJf/IJ0S+tAadUP7EUIaVJJ3MNl+7Bg0qBJBCNUTkJw0W1l
a6lG0Fwc1egV5KGOYAo+gSkZX7+qHcAhFh5If7gMlOwDKBRQhGtxL4o7Qr59CQ4ddmBz6D8S2gTy
rrHGTLUJWoKIZGD+E2lpndIobslGStJpGMOZDxEa9TpjmlRk2Fwuzi6aOFQpyybr9PgcRYcV4XG9
RjW8JWEDkN/T8YLw3ctoPlT+CurqVkkiCDemRlOMvY1d5WvwFSIIwG6jPvWLuRix5xfN3Rk6y4Cv
L8di8n4hxJm/42WADldQ/Pfc4kVP4RYNfJJN7DHAVrL0VAVKyVoHybFK5WT8l2etdDyvMqwZYFyy
6l9ndDFKe18HTr6NLzHWo1uDkxs+tx0osqWMFlwvC2Zy2xjXVaxfJRtNPG+U26Hn3EsgAwgaqsr+
11RXHj/K0VKV+BdeFNSiav6rWHBk3NZJcjhj02lQBeFrTFHxrHZ4d1D3hTGFsG0ggAMMM7LYGabQ
nCt0sF19VOJe98gl52tKlT0UqK/EX1E38wCmHSkpXaUKeTLmWSVF9F7Ux0gmLVVp6MvC5pwNb4k3
4TjbdAK9p5mfysp0bt5BkKM4F+e398HpZNoQJhirmQbPCim4IwWb47ziAMhovKfVfnghXo0i7UBv
zTbP2jaM6OY9/x8F50OMCi2tJz+tBZqmt1kzkWWJIViNUxn5sPjVxW1aIILwsYxrXGZrFkN9lsIp
1+JirGFlbai8/6I59pGr+2v9MPVI/13UrQBh7Q5ckp2s/If+sEvmohqCzctSSOkyz8RS06G3QJX2
COYdyOp7ZpAx/Fp0EAm4Vh4mQ5sbOuoorPHx4i4i+jOGTYiJcCbpBCNf3yv67g82gTdjVJeceV2P
ZbbG492hiGMA53nbKpt8xpugjwgbNVQ3+VhAvUpaYirQPxqiOEX+MRmK/po+ato4jyPY71xMCydj
sT0pakewFuIFIhjPeadNOCTOjDVil12kd/viLRDcRpKEU6DQzG074d2yB0g+Gp9caqgNI5+5Bq9B
fxNKLNCB7CMtRibDIpU0co/wWpFYvoR1tjR8vxAXKNE70AquuuAYn/bwNg+S28DBPOmNHj55LYvp
Z3uz56J7qJzzDWv+HLtUt2I0gJB/C/+fAEc5jg5i8aaDe5f7BP4OKKVVzidkcH4Z1vpxJQ9NXQY1
lK95xereon3iG1zWrcDZZv2Ywa6J6O1+wkHM18dnhmqUpmfqhfiCctlh/usL3rYroOED8XXjhqak
kixrxxnEHXOkkVvRt/1PdtqR9yKEZMbhVVvtfEvJPSP1HUuIiM54fX9EG1jxbiOmuBEOCOk+f0jO
alxD96/dXWPA6PEoTGHLZQjbM2WfklQUibPP72GjsgiEtGNtj8NGBRfCNsgj+2/wG1df0UqSaG61
Pb13vRMJQkOValNWKV4o7kQiFJTa5R7WwyrNwVt9ZHwdhl63fvvHiRLX+gipEbLivPH3ZH5+Qd/Y
HOlVPt/s0QpdSk5dXbb9YvjXfMJmNU40balXNnLGzNjZ/zPejEjezaYOnqGyJfEosS+YxYcaRU/I
bO8O2Gf0xZc2StbPn/IOIb3i+MFGlnhL9k8ZziKj2FSNpgzcjAXzmtK9BSXX6JPCFE4u2vXPrqpr
VqrvAvV74rtOMeXtcnP7ZlgWSL6UmUUCjHDSwZdKhwDzmyc0SaMG0+KBOPzCTTlo+MZ/a5S+9fHt
GwR0PBSAqoGOYJWA3ttuj4Ko7NBQZLSnuEwjeJOxQMIaazlwUnybwjP50qwrD5SSjN0KfV+HtbeO
MdJCNNCYkwPYc1QrSfRzkWXxWS9uVXHNGqINmLMcWNg6uoeyoKDMzbaO+FWe3RX1RLMpCf0xSZo5
/1byOiaoifcuH+iYNYZrMrw1/IQPAYlRX3MwRbxopabR/tUC+vgv8vx4YdkxX7CzsXSnuM+LNGXe
ZjYt+AEPR298npj/A8qioQ6se9A31JLuDQOrPexYSVv+dTXKj4DPgvLc7dFwrJR6VSUCeMttcXv2
QkX/frfhcnmcCYs24lSWt9SrhskdkM0tS0xlOIBH2ZoccokR6vJtUtU54bC5A/cmlv5FZfyM2fdP
ZufcofBHNVPa8ygwZ+3xOHCg7C9msG4ogd2jy6V56dfAzpWO0aVtStVk9QKT1sSTG2hj8MpRuulx
FQTrEP5682O9dp1/9TP/fASMjRIu9UAugzXLEO5f+q/1L05ZaCHsRSXcVR6s+6pGmbuJNPhBLWnU
Hkq9HvT3KoOQqBQlAwBu2qVeJ9b4WrdS0OU7viCt6rJnkTaNC4yofYm30LA3GSFnbACX2hFVTOj+
9BZHwpFQxwOW32a31KJqR/lOPONmTOC8NEVDSQM/R5DnFxp4Q4Jk/lMw8GuVnaT89r4dRSrOVfFX
rFiapkyIs7+dfoQjRG78+oxCKVBE2eMwycMnThhRpKyBlhaRCfMUK7Ij7h7g//kK+Sdj62fQeBHJ
id+ALtB6t4KhTfQ4MlCiw4rEOZ3vswr/zG8q8bEwOkdXrPKu1dgsQUFFWomfhjNczJm/h30/C4Rv
jFtXi6fsY3rYH1WD2sOU0U46XNGxhhvnCpXrFt5BGuTKk9x5JNi+prhRzB3qiFHWAjrZD4q0oiB2
d2h1O4NIgbnSB33QhJNzhlXu7fj4MGIaj6LULeOmYlLQpJh/qLuLz2xZBv8DRW0GSn3vM+9z7X3R
Dadvl0QHRdtHflLx2ZqFN6y8Sp1LyLzmm2X+RcbI8+9ocOGAhw1UzK0gJiOfz9fUuEP72OA5dZg0
GbAJ4PUVkrIApXRXo0B7P9EkMga7hj3W5T4FAkw8lW6SOC5UOBUXzTjxPIQVBdFqviA6bvdjV3iq
RlVK5LXZOq1jXNzsGAyYgdRzcw0pgysyqD5PVIw5MKfrQZISg7dccNlYHErnHueBJPSOAR1r+65W
1r40PjRtD++/g8RdfGdbs/4z5CBEW614RChGftaaLYwAZwv+WlEOFLY6grLa4yJK97ZzPagRf6Sq
W7woSJgcYjS9cQ26mB6JzTrOjYvndXpFgOV3vBWc9lL9CAxMbtIwdJzOOOyvH0iOjF/0/drO7Y3E
UetMFdWXBKbFLWrR5RYVuROhD+gIZZ56kxB0aGCvMOYU39bL6ZkHuiU2/zabbS01SVzyr7erQIV4
GeU6NVH6OejYQoW8CWjDwm13IQO0pEf0jZtan4HLNVOyKh90CP0NXio/uVI4Xzdz6MgKt5HIYCGU
zO7bqM31obCPArHMq0XSe4wI/OtHE1dB3vObO3+4f5xgzUSsyg0nnzVgndjJ+PpdS5i89e1S3bTJ
26W9ZEWTw1eKXo/qyJJdq2sfyjyw9dDXxj28GOi5Ie/CMPC2HfXEFC+3i2bXgDT85YAfZy2KAEd8
C/y7tmzINaaF2vKSeFFSJ2zwiQ4+dm34iN85ik0SCUd+e9JDrlMNlVeIUe6tTWk7Ym6Gzstbq1rs
nqpkaaGl+dtnR6Fev4ahenqowAH9gDW5zIOT+r36D4lqpzapGzthahOY2ZwNOhWGiS3kW1Z2wFWz
f5SjVR1M68fDBznXMcd8OXhvBvNd0k64wBGGgrRuv8zhi0sqc1tZ+WjNKY6S4iyIQSq2EBjzgoDX
IgEtZtQrBVFnoAniTvhZee9HsKm3/5XH0RPS4KayHe3bgha3UlwLH/65/XdcTV1yNJfPSyqK2PVh
cBjFQXwXrz0C2B5EMBGET3JH38NTHS8iU1GTRvMO6J0B3JbEsVCTPEsR3P3m/pJDuTdle7ddbJBT
TLBIlU6PzDr35Ph9TNoL38GkaybdQAuHhwbSXQfYYPBEOVxejKVPkvAfbTSauvL9qdYGkkBqDLhH
S6y/9FluOuTzPaHs+O9oI2QLCkS7JUUgPv74Xqpf4rsTK/lWgWW72MvOj9v6feZfY61k1ng0dQGj
5yer9f83Cp7t6uOeiwQnguRzT3V2E/z7UWj8E52ORcblOz+TgLVRER0w655Z/aGyRLePItR9eLuC
YX7eSn8b9ysT5aBdYZ77ELLa2cO7fWWI3vLdlawx2JEUT9BPo8wHLZpSqlh2aFKKayNQZfOEKRW8
PZCTuofTDOTgkq4cHVlbx5ZyotJEvBJ7I24kLjxyboXmS8WoceX14/8PwmmUiNWi+iH6Y5idKTrt
MO2v3zTAxhTVr1CPZ5tVhUeiaVQTp0fIJIc9TTF5UTq8e9+WZFWHcJIPS/KFeag0xJET3zK3AI1k
KpAQLikEPd7akPA+Tyo8FIdzWJ5GCgWHyvm7YptlLXUwz+PVgqKVXtYWWghGnfBepOwb2Q9qFyEC
go7yPUlhlc4dshAER9DtX/e+Abh8fxaws1kALmvt5KA6t508g7s9ltZSh8dVaqR4akVc14ekQj5+
UFJ+Ue8qHIsmW6Ajg3Ri6wf3jNauEir8UyxtbCk7hhu/dUw9xFmf1BVJjexI5eeO7TaE63B2FtpF
6XhNlqb5kfG/AccCzb3LwbEdWgAbgqxMEWN3tuWllD+QsgcX1BiauxiV01FGoDpugNY8UBjExoWr
5sLuAWWRquidw2f27gq8aRkcy0/eRIRDZH8NcRaqy99rV8utb0h6iFXEjcoBq9O7apWmctsFD27Y
tLvmM1pSasxgPruKOOIpCCBDLaq+tug2SE/AOFmHA3ayiViSx9Cl4mcRtL1tP60o+8HHPNraGir3
3llu9LaHYd6owI43NA0qRr4gaQt1PBG8kb0wnGLTcsPwMoPgzn2jtUd1bZN8AX0L8h2ARZruxbAV
nG1MCi3L8sGhiPzsZ3mvixalM8X0DNqr/t0hmFx98NqLPOZksozv6pLsioMGYg5PtaoiDoZGjEE1
3kS8C2fMDxBqrQS6c4VGICFNp0bbtbxlKW1nJvCvXQSDjXfH03HLVfNg/sdkFur8SulmKanMHvaf
/YGrbfjXZhdQnDpP1UYPSFLNUUAJPknenpirbMO1GHGVA+UOcsW+X7/9FVYy8pICB1MfK7FAfWnA
TivtKtBXnmxxaAJCaW5SV87lyxExSn/0cwaOomOY3ZNTaxyKN60Zbn9i5dk8gDQS8+fTS6c7p4l+
9gwj5TP2orfIPYYoIYdsLadhq4fT1kpSk4URn5an/nbPYbXtsQ1QgoTOUaQuM4PJj2QJC1j5co6n
XukTgezexVLodhEKCc2rPGfnSBq9f+Isqqxgeg/CO7GsAOsVfZW1ZyFtvB+vPkkzN4BMkhp7XDI/
Q3lal4P63+ZwN6B84jNK/LpTmTAVyJgdJOYOAC1uVSZvqIIRDXOW9GgZXtxTuN8gNU4BwxztX+jZ
q9yLoIIz0vOXNEeMY07NXX44iDow6L3DbJB2LleMExBrgEKDUSfzSRAfeVASX6FL8ksV140og1jD
m+zK+PW4OGfZHKBvAjeDkeoSv5tnkXTaEpb/SgGrDippiboAHCBihjqJjEWC1vLjVYN6wjCMIt/s
KfRUJxiGZzSpKbVbNiHCHduZrisK91dEN5svyiWcI0aIL4pzyqzgG0L4zoOnqRSwo7ccE8v/oYRz
5L9alNpd+438tkcHugpZ+GqT42XHhMd6TXQ/qY7gsmUHsWrdGMvdqL25oYf2PWPHRtWAyFbUj0IB
h69NzR50bgM5R7kxWWf0OltTqNoHsYqdc/UJLvKZ6nVI7JTlSJMFFsYOJ9gMkkudRkIcQkWB1em4
ueA5X2MBggC1phLZoVXtTusp1WBlTxS+lEeK1NuCxR8zO/SWfTad3ZYQF9bN9vZOduFifdv5Shjv
JOoPNOvPFfZ4HBeiQFZCr458YaLYx+lX4VMhnk8zLTWrpBwrhf8XDFEXtts5CrPcTQVaKt1XqbHZ
3Quv85UopTmOekH7FYckr6kBFvTiNFWDllEudzbsCLyxa8XdhD1+IVHNK9HYF7oLOnVs7+AwO0bn
eId3KOeG1H8FXT2zxMtbes4gk++Qo/C+RVONxIU7Xp1USR+UHyzBN3utev8WBDLq+XyJtOq/KT3J
Rb2db/QH4gZpfHegYj7O8OacXvoHtyKKsl75A7kzcyzsgIh3wfx3kP7FpOWKd8hhk6LbBRubwqtK
wKJTETJMp0REhXH7VNORGIrJ2bpTYRduBBycVZboOvugcChAIR1l3REWtu1Fw8m3ETIwaN7shs+9
xnCdGsUBLcTPjUwZkFu/xMIsrUlmwhEsDb6K/5INF/J9oYFuQZi4Gz0KPmzMTxKcmjWjOUl8toBd
cTKlqXWbf4mlfAQfj+kFGWC4ZT0bmjFoSgnkz4uSHkWwUKO908Of21aIBht1WJz4jF+wGIFxxya5
OF+C4CVO+KGBJx71hp72CVIRfrcotALSaFX2pGav8eLn9eBoSKOk7skBp8/dm1j7UpcqBAV3fM4X
mA1w4Ha6vFwOQxBz0kKHWwe5p6qpyr0neKGdQU6BspdAW3dGP0TtI8XWdZvEk9EBj9OXpxzjQWXM
Ah1kVgbfFN3IWq8an+UJl/GiHHa9JG9mAloDVq4qRsvwYImTFi9buE7WTKayJLqrmZH4mQZuZRVS
nVLrdJJu8irX9jvBUvNYSZxuy/7/ZHhXF6Bk2N5i+Ub88FWogYysFOhPRtX2ypdcsXv5WsfrLlvF
06CbOAjwVB8943WV2g9KHokqxaTnCRnt235k9d8B4NthGBDyVnhJO0Zqc+NuTEDZ/rLLcNVxuxo1
HFmAx48z5HfKEKkgTGX9/KSwaHZij3QSVvEA5yb7jVxiL+8xmnnRWyxrVlsvrFCSRiutIfrfmH0m
tgZNpE6PO+6r/sbOVOlgt0pExbRRUx8AJ3yGIdbe7skOPv4nor5KuYnB/koSvHAYgbmi0vnmnZbo
or4RdlhsXfFAjHT6pqFGCpXGonFuBzTx2SOTvY5yDITsQq5/uUVJA1K0Sm6fY3szJCwYHCyNvJFB
ed5o9BbScaRKzPvXUpvFyafgIa7+tHRx9h4qwYqkAzv/ZlZWrXPSETBeu+pHAy6qK+hS6tm+J7qI
m21wFkBisZ2XZi1NhrDeVK8rSyAi4HStPuSO16rfCm+Vo2IDz7ttiIpzVxR/kErOcvjdagKZCmpI
xJgBx72YQKAJ2227wsunIePp8EMB8ayX5U516knqb/lqRtdczJ1GWOHewnTYkewiNGqLBwpz44xb
wgIWev+ArBjdUnPvRyCPhVIqgYorV4HpaAk3GeMDZe2ZSg0Zjzys14etGiLRlS8u4TizEGABT+f/
NYnyhEhy6tDcFMQz+tV746ia53VnqI1jr1503Mf2mwPqHZXW9y3tG4HqtOsmWWVv59+6d5DszBsd
6swNfE0i+42r5WWnR+OjaFiKIQ6P7kJlVVslynLp493P46cYWbWSTS8Z2hmhnOR0AH7ThRln2R0o
/1kZV+PBybBPM1MUNMj0RlRC/7W+pGz9DBf7H4x+pYsrHmI4G9ymWRpP9M4ZFbOnFQ6yBOH4G93p
yKJp/lHxDwj6+nnVW1pQizEQf0gYbqk553bYLnTuM+gtH40CISHkFZG8tFa/rRFKV6zAieH41gZz
2RFIpiM6+4RgoIG+HhIBfL5tmW0WDFfCZx7b++OUsQ8SQ9YUYogcmSZVY4hBojfjCjCEpNVBjUPq
X2qcm7fOp+0sSGX+VUxmtwUqV+m0+tajudhuDhRd16XLSH3t0aLF/iZDZfs9+/8unu4EzM02rNj0
zeuzk2jDkM1gFFd1QaBpruBveRencj00byanaMpFId4vtii2m1zhofaRz7N8dxxsyBd9ujwmLVLd
CKK6vBhgQCL3tMoMAQGMmDCw07iKTj+JakHeQYK+cfCCVyxiVDjCqqlxG9AQ3dSbIgxMjxL4MBKh
cDmW/7NQQ5BHtK8i207fAGIyCIZV+rMrXp4pIxiZrVUXV3KZvyThuOCD8Bpt2ynlUMuZkJIiVnDD
c36lhd2KTJdb/0KhGkHe5cEQE/M5qhgDT7OjJf1Hs0ugtbWgj/KABG1gUjfoKHsmsxEGb3QPFa2+
c426FMkca6oYRDejl39o270qGZl0DwspawTYre5Ec+jcNeBtt50r1rmJ6ioIwJZJ2s8apOr18azq
2X5amSkHpENuueNfq4cyMLKfuPl1pW7TpLX0bus+Az2Gt9ZIbKRGP0YpY6C9SytFocH0fZN5vy3o
3ft0xxrd1yDsC1LAeG1AKyQATcfeEPNsPCmrHfFh6rFK+ezsmsRo70RmshhyIqJ8X6MY3fqpR+ZL
9ByaMKasHKoPYXHCkYSy6CThcBNjMRcWbv4PSrPL01u89/3qStiHnI6Ptoq/IvGJu/NdUJLMMIeP
0AgP7yIocWXE9XcaY0/sYncUCZsSlsPCQrSELdbc7ZW6w0b/ca6S70GlrbcZ/W9SeN5ONg0GeMI0
hU+xBMepLa1hbAX6qBw7smJkFPTupYw2Mn+YHtE7IkqMNVXDVlg1t7l8GiYlqkdK7mEKCTLdo/N0
rVnDkQuO8YIcey6Mr1118E12r50xwv0bdXUorUeOPakeQ0EyD5cOOSv45B4eYrO9N89qG5nA6yE8
hh+Q8aam/VGXppHQMXdjG3dw3FVDSFcmsDd6HN9IImJn1DlJ5WPS37pOQ95e4KI/sU4ZMTmaT9gy
YSV9XwABW8QhWxXeMFbCEwPqFBtbH3gaceTP9Knuh4MC4mZHUXLs6wNy0h5vLLDfShl9/AaKw8oB
YVg13TJXvjdzbqG6ejKI2S6aJg8PjdeFLd+nRpmWM+7c6sGKdFTSeR9YWpNfbgvWENLcWnqmJKIE
Y9keu7a13cOjfeqbaL//0H+/ha7xYlyaMWMQtBYaIavk0fi1A2Nknn4gcjtPmKT5mrti5ini8Ulr
/ddaZV2NHT7poQUr9xIxs4/3DTZ2KJkviWP3SakPCo7zd92ZvmxinEHssWi6Q05eaEWb0ekaaCY9
6Ceqo18EBdDGqDM87gMXGY8387qcKCvaAwPD50szG/r8cU2R9E6aBU+zwTMBnK1WWRVX4PZBJ6/p
V1KxWenbV1kzE1lnZqLTWwTf+5Z5fpDeqzs5xE+W/OwdYQ4dy3C4M9W4MS8/XrhhXzAH5TfidDyQ
uNbREL6q/dmzCJ1h83KtS74DBhmlYU7h0YKawXTmWr8T9LbcUe/xpWIJ6znE0/yJulqpnzKhwHa/
ddBTwE2rn4hVS25rxBm3h0o1ZBzP/DvVv4AlsQQKDEov5HlwJlXq8Ij5f19OLugmhrQVFvdYCryG
rQzu8uXSnybPHfFUjgn/OTeT2qC1APq1RI5j9pZAIoSCvxs66YwzuKbwXfzKc3fyaqSLd0rZlfm7
0NbCYJEzWIuJIckKcPvfrDTtXo2dvzCadhF6gy3x5PIw+jLctDHYZ6HeDPpRgp3Z6dWPq7DWjf/t
DYlyZxsMFfMoWbaaXfRJaMIPKaWQRhxHdN4dKnsFk75k+i1cSCXwGy59c1oqP0SLYF4BgqHqgcCL
wk+FtaVmL/gyn8uTuuN4sIAXwFOpgxjE+j3Yc6qRcqxNgyZOcWFwcm5tepDorfsNs1WfpfPhH9vf
ihmw5tvC403J43jG4T6DZcCS4++tHVF6tChLppxwAnKTCE2za2Qlw4zbuMBFG2vu1p02HRIELaJ4
wtATJXGw169o+YHTUPaut3jDgtUn0GBRa+XNgiLcYY7roInBcthpdPtvZimWj0z4cV/QnlmhN1BS
b0CcydLwgBgVtbQNatVtNltIehSXxl9iE1yO8HsSWjk04H71lgwMTFRZkXy8cq5UwKsf9Ps+vHEh
vLKmew3rBJqXt9pQFaA7Re09+SNojtSZ/8T2Wkh9Ju+EIVheomseqfPj+33NDyoXIzfYpobhAhwY
V/VcMJ+M2/sESURHxtOIs+zphdTWyd3NfwlmVJKGAqiec9eX+CONpG3YM97bGELUL1e7Exhi6w9r
8/I4lBRA6IZvQHUvf/T3SrVD2V4r63Gg7sBbkttBeuwJxytd2GXRLdKODf+XaNORoOw78sQ/yj87
deaMkdPziqRHBBoujC8GpuS5WJFQ86fBB+SC8OYm44fFggRuW3wDWeHHSZhHKZy0qtbeQzJbdBSw
Ixqo4Gx9BtbjpL6VOb9mb5bNC1zusH8jp4peS14AX5+iPNolv15LtCEtKzJGhGMnX/28yrCn51TJ
ItSpTFwZbvYTiQ0qBWPWFeD/O2JinRVi2s+Yj3Eg0ujl7D9qXPiIgFPFcM+JD8Qh9f4tURPdxi3/
lH8TceTr5pxugVj3Hr/bJxWQja6IS0e6HODh6VyrKmMRhjbjdeDNR+ZoTlXDqFZRmdX3VqdAJ4uB
T/2ydZ3aQE5/FbYCbhd9xc1ixiGSBurzLu8YyFXDGr26s1jgrCDPs4Tin4tMUUf72mjQZSoncN0Y
N0Ajeiv15TZuyp3fg+cnv8w6DSn6KJXDLINHtvpRsxhvkuD60cN+xpMsAbmvTGF1f2nZ86QuXH27
VLTnHAr5UcQSD6wr8pcenPpZzM3ktPRmZ55cryTpKqLMFhUow3WZAPXYUUtkvRUXqfjDSxxjGhrl
k8lZbsrkmIuCqvkTOsNNLNEzGGUEuWikc46py1s+tmsZCuVZUvRqBHyToCfrb0JzDJHxsKc4lKgn
0Dqr9EvlZUYRI3rzOiD8x38GGaOADRxy4W3yK4iLZ6QorK9Xe4EZTBvTNjKaJAcbQzTT6SilXekg
3c43AJg2n9/MkYuffEUZHPQA+cyaiA4ZsO53VjEX2Y4hv3BjeIukm9VIgfREZapRGlUi8vwDecWo
uci8htVVC8ozuK6e1WNNlZEmc9Y5ooGecQK++mbRxPmuEJCkuGVl3as2s+4+h1t8EvIu1frILmLJ
EGKD0enJ3wIjGrGSn2EMXjwUX70XoPnvJKr7FCdQvCFhUjULcc+bQF19c5nL+HP4HY6fo1qtHaGI
y8fLOLQSbhIKKKKAawyUls8QDVekGLczahMbGDT37ILFpWwNLhnL8pNl6FTEGQN6MRlmU3k0v1I8
Kk/sUGfHn0P8H2dLpuquCBIp5u519ZdwvZ7xBUaORuBiJ2SptQp19QdYKvPdUwRuCdkh+mRASjPI
xgYSCRG4Qj/jf53LJAqcJgFhmxYrArlumz5V9W7x6RUYRZFIEZsuSpivFCx3KkqxTCKwtDjsJIAX
dt480NLAmfMuPdYckxmUkoNR84uTi440Z2PTQ/qsexA3V6SCSp9gnrYu5a/p9PswOb63LA8FO0iw
dXhNBjf+1d1R4eANkWKreAgtLiMllpXE3XhP7Ziy0ZUcli4teuVoTnK+n11whnQQO5O9n2EIW+10
4Y4VOKuNRoPwHqx2uymIaIhG7ziI8RnK7cRS48IgfpiDdwZ1aO2lW9ygXRIn3DkxI3ZgBufKAqnx
DmotIAlQA5yJJE56Q13jeLV9M0mLE2MSoKZyBY96/uD0d7yuQoi9V1rpZ7sNEfORslZrJb/4F2w3
dJiEXMEN6ZeZkyTAGprfRJDq4Dn5etJbQYznt0tV6pgkzySetvh9T8hGD1YfHs+11ynzn7ogECP8
E7Fz07ASMMM2hzrvsq0Ja0NAe9pxkWO35MKRNjsG/eIxLHcIFo4CXojYmw7wwAMYckM/yM6U7+6v
mj6/Ev6H129FB5UTLLC7aNGWVYiALcZo2nlEHQFV9r6hWBeLtPdVzKopF8ed7yr6flB0sRoinqw5
rs4MLWVjqEr+ZOrEkOtTsJmb24To7Rm7Z/NQnqbF/zOSCNX6m9hXXwENJ4hMDQ6fjF5IFf08YnRC
c89Ln/kdBovSfdASH5/pMvdW0eAYLQkT8EKTlwJQNIH4E/LngdYiZoe+urklpFIkq+nsmW1OH3vZ
qH/TS18ed5yZsXHakomp0uZ00lq0pfUAsAejDaCD8f6n4NlLjf56t0smu3ODjP7gRPcBxoDYACmJ
tVC8aGXnWjnkT0kicLrCRIverNpI+VtOA88hBxdscStqme07AH5Q3q0+V5tHb9tcxWLdnqSNIo2W
7w8qexCBCZa2sISqO8i3sREZgqrtmBir1aGl1+dGbDB8P1YSc1fQSFfvN2m4ZwmJ0m34FidzwFCl
N5OXf+TsoRqPrd586d4cfujfRYehD3PBRbz99XLF9sRUTmMS8+FGlITtVvHvp5NtHTHC2+LVqqZh
0ZBI38H/Fh8AJWIpDzmiiqzyFpIp54jEIUdyACNbL1ql/G9Gqq9j2jXbLcb85AvPGjhZy+xUrDhK
23P+Xt6m3dLobLPRmTjU584rWa1RxIcdtZLKbjBV9YcHukxSExqQbVw3f1xRKMXQDzQeBr5XI8V5
SQrwBd+VNR/nK2s/nNG3hwkAfGVDUkbhIcuCM/YSbCCHFcZlZlJYJxZYESlf7dgyazCjjfPiBbUJ
wdfCGHwNE+PXirthvZlY30FFQyXPI7ZcEi+xLnjmvJPDwyQe1bYTzBfyb5kzcdJBvJYOCizwQL1M
GNSZ7XWXTwKebySTecUBnBM2Z9B5AITSbI3FvkLV1cp7ikoJpXKppS1gzyTfzcEbEJ52YkhQvuTX
LuQkEDJ2dyuXcRDZb6jhUGxUwHTMuthw5wwa4MsXZ/iARAU8qYcyfbnNWMfjG51dypXO4CVKGt8M
NdH8trrgM9dogoTUwHkymfqTmk+nZPpgTHeCVxzCNawzmKnihmBZjdVIZeTjeeHW7SjaTL3XkRYW
CrUNXlL3DoqqTuBk0hWXU9azPpwbAkvpMsWKuV8nQLKlvLt4QL2MbJx1JBsz4CtKbTbxwQ3NNMzO
ifQl7LBJrXsRwR/J3BO0+bTQfiVt72EzKYDVsFZd3zFkJfW32C+G2/W+h7prfDfRrwxm/lZYy5ri
q361cXZ4pWcvGPOB5UPexrPHCf4c83ZMv8TCxe0lnDlnhKSdCMBxepCgxUwVZd34H6qIjmrfkXw1
kE8Uxjkcyt4DpWKjR0B0E20WAPAtEB1Dhk+8jMAnSa+UsoAbyG8bjXjjw2ar9sVqFHPYLWOy30C2
4qEQ+XmSWPitodel93fRMdm/uaUDYSX4lJv3keCDyfiTrQQt6RlDsIj7QRtZgXf/vMrRpsLd5VlB
SoGhJsdIQe2LRlMS/u8kvZh+REnhbbcpQgDh/hRb5DIFoEpbsOG6nqIb5cfPutv0sJbzE67ruiST
rgEoVn7iAonB3xD4TWQxHIDR/uit1Z8zK//NLGY8hVyNhFaRzmEkp8cdpnb2aBENyf+YN/5X9Mbs
7a7rOLL6bqHOM5P8ZIu/HjwkfIRKsxbSZVDhfN3uYJ6+3d2cKGvM8IaRP5FxlqewfFFlKlzMstUR
ISVfSf7YWtn3KjyyYLyqev0OrT7WZA9B5HB9so3i4WvSapGSWyieoDU26LHNFthwDT0ek+ZcFgJJ
dwYZ/cI9iar6N1T4JG+w4hcy+EJ25wCF8P9BEEhU35+Y45yLIH3MX4Kib/rSOqvN9Z4VyZlGmuFK
BO5yCOKRed2++16dnJ0pLRY6WcgYIm0EIvz0Suz+3w/41WBqe7R0Dwy3+iu0ThfI3E56ysufQUDk
idEfvJXjjYD2YRFBi9iRD5YJmO9BWGtmXPUCfUmCZCpF5VSRk/YuPrFNNT4VzUAgfxlNBLMSnFFi
f9QzlJxPOH1gh/PIHsDc1nzKdX3HyBl07EBDwA36hbZX13tXLVhb4py8HKBck0S41hG9c8LfQQO+
Nv3UgIsfZY/oecQfe9k+C2KAPpNVaRSLU578XZypQbUl7o37QKoZpdagx9oFOLgf+Ya8AdlFCOzT
lOGNtPe01sVBhrFaD5/89X1vHlIRbAk6sAFg+wYg/PiUlFoN73HRSF9jaBrARZwRwS9Ro71w1n2Z
CY2nn42zLECImzGGWls8B0NjRx0w1N8b+cWrkO9Uo6mHGQh2nitKCZUQMy4sN/ueDgq04oxoUyu3
5Gbo/eOm3OnpMXRHe8WyySK00CwUX9IKla0C4hVSSWt5SxNszlk4uYSSeO6ejVYNerezasyXhGZe
gtAD3hkCKZf1/9uBfxmwA+J+omeXJhqo3qsmydNF7Ktte5yjQXqsT1ogBiWkrITAb9f9qdDuRHSK
6T95JmktMi1diHj3eOnFpJeLcs3TtemdJQZupaLW9DY4bOHF96FMDkmRvCxYc1eEIP0qJReoIyBn
v/D7sLsszWnNWg+oJMPktkf/3OWA6V5eUvOxtmF5toGwBHvQnDmC5iHQRRvZyds2X5Dp8/KQ92K2
YCFxIbeL4b5V4dbUP34VDYiAJRbkIH2WzDuiiAs8+xCSmM7fhG7KpzDOX3PSw0kDClkn+10zq/zZ
UL8LQ+uLcIuozwaYjxljT9ug3PYD3Nk5Efqs10v6lBb0U4dJ7XnWKw3pna5AC9GSnscSWzNwIwtI
bsJvhvPJm0HWJg78LZJxgXgVPjNZV2oRN97Xv5huZu03VfDZtyEEG4VNaYybpqLJviOpoM3aiFzy
pcy5fEpV0VNy3mzRhvhOn5ey/3smNzzg3hEP3ShRR+cKUMBa44jGJ9vlBJT85gNVAKLGGTtUWgBT
GhOX/Uk2bNqqRcdtLERS6okQc/lyNztsGChAFTS3nT/mtcYuXbUGltct9ldn0UrNnAtzLtSb/bWu
bEv/0qGfQPcoryJHVtKiIMWlSpARNu5WqqX9Le6+CHtLww8hsLezQ7RrWL0+06ts6oV5qtPdNoFh
/KR2M62wlYSAkziPGE/qw29CfrT7kR2dG7TmFK7DF4o0WNgQ79v7L0UZgElloymlNnw+wu8wpJtv
8WXXyfbUycfjxxjDVCkvH1s5xaogD8hpYU3WLDYi2vRwJvS248I0Kw+qp+0hgV4SRHRaUf5AHAer
I0aLoiR6nfzyUj05IWtUs7OETt7/oxBheaKEWZwrA1mXPIAM/st+9p77685TNgzkHOcSiG1J4Cz+
lM0N8aWd0jeeLew4Ewa0RJ4iAR9ceyw4ipzRmcqsm+B5pntAlGv8WpF1ubmwA2ad6u5G+pc2sqT1
zd2UryeWDUDdsGor6h5UWc/yzkHX+Lx3+5wfHRTPXzsBenMmBN3T8zPW/ANXNNnOhDz5Q1O18oWj
Ht4IiLYQExqNCSTwkphBsNO2M2/6pkMGCjYVVGxbGWng7KUcSXfTikg5hPAD1nF8Vmg5KUQZuCF7
utem9kCYQ2CMFsuUA5VC0Wbn0zaJckiImMZQu+oyaLsiZXbyfaPq0KyVR3jSyX7FbzVRTjm07qku
9AKodjDX+EwXkg+fdMxBsWKdSoufduiPR6S4mnNvjCfd2JdWSkpXJwDj2u68R0QLn19Nqh7+eM1R
FfvSeshYqAgEoPHrMZv7Odcbgvz3wPoIl3BXX/zjefV4dej2cScqvnkYIyeLOCENsrzz9Yu/Tute
ubGbusACu0Ko94vshDgQ5Qk7wE+zo2PVFGm4W5LR6EpcYBA9EO3rZcck7gfXqd/x1ygaP7/JRmyo
zD/N9fYAuoecDHn6Zhg8PCIbbHZqccve99zmfICV3clPB7l3fdfyuB0xJI+bHe1qqzr+VOaQ3LmR
BEjhYPdLYBy6AiKYCH2VNq5JVqCAnDuTj61GoaLsUgen5XjLXXyi4oRP6fAK5lVajgvoAKGW3zds
ZCY4taHzKOruZWVwHj3AmR3M1eBva6Qtf0DCF3sWr/37qGmkDwN4vxg7NopDAXGjrK3v2twaKSft
qw8CyBzO53vG13mGjZ4t59Es58s/MEK2hp3ZMALHOg1vc3H/3pwUmXpEXMRffNUl/nfyhnsq1eu7
xcpYanekHq4pY4ITaj73/hYgdQxx6f21TM4EZkcqBQg5INe5qrJRVPXKtyQZZfnWZHWQ7nADVlE3
1ZtGmUDLaWm+KdM9XwlzNhNbWiU4hys+xGC6JhvBIWaVo0qHxaKjLcChD+eTg6xvfRgGMzj6kYqH
J94lrMuiBQABXLVLzdX02R+k4/ngUyfYZoVCNZ1WDq0iMk5Jp1IQVv5HkxUDpmufX7IHhu/XWWye
d7KhFWhrdMyrpc8V8aNPXOY7IHvQwgPfJ3479cVT28Fjy7lqLJzW9EmL7YLmtRFF9HbSApcMMoiA
7G3Rt0chMiYEEZTOPSQh3IjoXImKOoRQyME00rKPKEI6n+8Qqo/n2G2X5WQmGHM5U1vfUyGFUqH2
O/ITBdhnbbjLWO+JUXdm64eK6f99dRbRQTmu3BB9RN4kJONtBOoSNpzAWYwO1qnjcJJcSxhUxJXP
jqDORmupWYCOc+vnk5kADSyZJtHv7kxyxtXCcGsKLPz5lT7lSeA/IzOJyvXKHm+5+JM19IsDWVpZ
f0KZcHZf4VUNk8dX2zF18q4MkqYTMf9+KeWdvqqAuf5hJ3fYGp0gQ9u01gxxWTYDb6YW/+6AVYqV
sQtaz1pa7q2W5PF6FeCVxZsbyM68Gx7tZBI2uxQkZowGlJ2q/z+uvLux44hpek9Mplcxb0O0gJOo
4oFpJt/PY8Iu8hDdv6kYczZQOaF1xd3n1sOMoebe6bRZ5+jLiZ72X0OPq+joayz2EfHvE2PK1cYy
Y8/YylaEAshoey+WJMqXQXqii/5m5w0qNoWTG7bN5NL2qC3xKGVOOY+QUogD3LmK7qAkfHCILr89
mZcTyllqFFhf7bUOEsIwM8ntjuQ4Vwtm5vt940Jaz/ineBg4xgxGwt4y6oDjJLbqeyy3a0FLUrfM
oOH2qlgrlKia4nHE18YZiuQjE5trqpVN/6uCRnUuzAE+1TxHn1ji3lv4pyPL7HFWLpgjCN/Iaofw
ETZ2SKUk9Ba8igEO9kbTAktlkGG4gwp6CbN+bf2U+cRFEjE0Rj2qwu8geic9khpnpUDTMUCFMmJS
8daioCYpUwYW6HlTX5ZMymXIVjYFpJlxCs1Wk+t6fhKxDvhyaljVLZtkFbP0BnIDRON7xaJ/dPuc
l3RVu/dVjcLYkwzHIc9nl890PammGw57m7vNV5ow3JJNL4Eb4u04+975PBzjVGkohRITVOqFhspj
inOZHhIyuHzlqn7y2HoWeIdm//vvSCOrNRkC+7G71wQTpKYasDmVIkL3B+vQDrOMiAXqBF7RqxGe
fxFkYxu9dxAI5hv2y1UfRHK/JBo/xt6fYW45OJzKdf8tQQeEjbwjx4qY7MwkbUHIXCCT+FrFVuKH
5vBsJ1AvruiuIFY3/gVzEZ30Z90V41nvvBD2RJZYd/1RsHtQp00zRLFv5ZPoqOuKQAW1xNf6n7+D
ztHQh51ijSJPPabUCXcIS8uDrxoq7QufQw1pnVmz4tDPJ34Gj4q9Ab+JXWGCVbnhwqqsteg51NNQ
MUoxm/DY2RhBbo6yyG4JB3+9OiFhXsK7Lotafd8z1Rfe3+ruOuU1W5sBLFW3ffwDt4bMPptNBvTq
tWARx4x0mZ1Np5m1sGZzU/LqSY2SZsgs9J2Sma44Gx76Bh9E4JkIcyMrateROCv3ARAh53xoeVKA
r2mA/NGL7/XXvFsHf5GeFF0j3/nhrF7yEFtDPQu3MPgFV+8IcsQ8sywmOY5EFwYxjRLQNsMuz3mc
qdKbBOE0uM73nH4E8Ih0QOfZvVK8IjlixbS5Y67n3hU3KQWT3W8ViiSduuRRi16oUDmVhpoVaflC
VFRYQYgQSN0ZwOmgPW/PBPWsrBmaq/Muu9wOJ0iaGVpvE+OabTu0uqgso1Vu55fJEPnyp533YUGI
TgWqs9phGBj00gAeeCrOFradzkLLpOcDwXzQjP9Pvy/7o7/Sc0Mx6v1A2Okoweu44p84PZem292j
VLVq9bQm4KO2IeXp+Srp69OgeCVXbMg2u/qPg/jji8Ti6BJsJ7X3Vd0Lx3Ch51N9UVDMQfX3M0IP
FXXA8yYihhuDMAcUyfDPqA+LtTYDyH1S3BmV1xAw5jDZWFdyo8zbR8k+gAhjpAYCux+stFiResXA
Iq6Lxqd/G8OEPuo1yNZc1ck5ZwZUC1I4nRWzojALxOAOj/+yfYnmYvgb01JTavHlRSdJudmT19mX
veIM8L5o6Ia1TrtpMdGCzIkDha9G29Y776Ara0uKv7lllneebbCFoaSsrf1pwjVSU6PtNiF0x6i8
U6sF6xjfWhSDxhJGzhb3xk2ynCGT5sY8ROaqnF1uqhEZO2zYYf3a47GE+kTy74zGJ5AEJzojtXeC
SK8b75sJUz1YEtKjlNbU7R0AdI9DiA2S4ubQLqOaiUcTAc19XF1iex7yNgcvygBnrNUtx8JuaUhq
vEgoXXZAdNrL4qn11CeERYSRhgTWwVHBEHT4jBtAGDY4UMzlHzV8DQ7mhbHI7cIhuiQgW+f6C6Cb
bhFfhOWtO16Ss6ZQ7cJYciyMdoTBT5TFglq8hGPoF0HOyjqTmo8sIGeypmQ0doywnxPxA0ndtL1V
DGO24ze2KSFu4RHv9geWRmxxLczY46vP/wuMaiFVCRbXpOeU3rR8YDR6K8ZMxlwcC69VG4aa/WVj
uY2l+OATGWindQQT9GR909+nPwPUFVzxUVK5nRCMf3uTZLIqr7qUKe453PyaGNHeKRB8kI4U//gj
+d8YUvGnUZjrRbobN3rgRlp6LIUTRM2WzfJsyTDGeitFnp2QlTH/BQVmJMfF2VllI3vMTc6XgOhQ
D5wtH99X9pg25LaXXv51prSzcaD3E0omf1SsWYpV6D41lQg1LQrkX9aN2urilb8Duvsg0cpU6TuG
HwMd366I4FyEf2qdSORMbMS/I9Htyom+Fmgv8CO7XoFj6zsrHCn62ikEStdDHQYx8anaP107iBZG
ZbupiYwajKQ93s0JgLOe7cZ33UbZVKZz4lweOcv7qOnGcqZJVeyeO+IePuiPY5gKgZzssASVbAlz
G7HIo1cUoN6lvTU69xF+26e7iuulqxCYnC9q+yLvQmFmRVk/6QtI73OtC6y+QEqKB649e1vVLRt5
LXUO0J6KsMWEGL79rkraTCQKfDvfyIfbmKP4CqGcYBfk3x5309eHKDWiuSiurK0rkZA+wb3RvDnZ
hM08K+UqwDwaUikbPLupEgi5aN5PlptoM6JbaTp/CNj/QovjlwqVpnMy9DQzBEBaaVzLGv82eDva
O4owFVFdxQYuTT8eX2DN9qS/Ccjo7SivhhZ8OPi+DEgmPtwT2H6VC5Zujgk5249H07FDe5m+xwpn
ELk5Ge2cAnm6wbxjv4riOB7hMERbLQORNu+6r5sIFp3yqDciQpzhBwyrN4oM+7PS6rBZCD9NHWsY
MepBW5pa9fj7c1S8s21DjQLsWHfxnNuajVm/VsrxOwMS+GZ8dv6/txmbi3L/RdZz343d4smhAtWT
lS8+zZs3leIekLiM1X7vDs1oHLzGVlyKNceRtscFJg3zDYnNeGTFGSFypMbtbcfDy+UA01fvIV+x
hHONM3yQsjPQD82CbBjmTBJtvW8Mcx/UVCqXnqdffr2wRml9p4aDroyBd47T9nJ8gmBHQR2lIxoE
vIsZHUE4sQacoAcKpyk4964gShD69BnKzZKaa1nwKCrHDht2wEZtLCuP8Y93rPNgFSJOSGKazS1x
jiNFyyijWUYaZ3NKcRdYJPDK0OWLzeKoXMJHlUKphVSb1x0oucRW2TvXd46OAsXj8M5lokK615xW
12E6feV8fC+fORDxnKJqK5whoNE7OLh+0bQy321cUsaCuYHfLdBSS5JUjnKtLPV3bCNN2yzqTFUH
jIrPlsB6lYgnOCjgu0BtJcMOeVGExcqrxuPPLOJ5TkDCAAI6f6XB1EX7ETKzFAZcgiKBOphklPZL
kwaKhhOHCvAkufe5W0Nr4AOHnwEhYG2w4MbCxoxG8s1JkyEjU9qAmyE0nBL1Nx9CZgizts3GVZ9j
Lz5qPeMEvl0mHYlshP+9xj1yyHEvILmpHEzjJipQBoZGLD/FAp2Z3QyQTSN2oQqR4+ahPbO5Ru2a
aUqITynUt5HavO+OD0a2xTigXObCXJ8mMv9KqNl0WZQ72RnUJk9d32ayohyQIEOhlUEJ5ODVDED/
WiLB/kCQAuby/l4/0FD2IcIf3Vg+BmGrhujApSJWjtBFQGyBCvsT89AxGSgGgnHsvOfHbJGS96yb
VTh+sTPB6VlqTcRu2FWz+EVazakqwtODbZw3CTA34pwb/5bD9Yt3VoiiO66fFxzz29CANFMWQOaJ
3d8eaa7uYWKAeULP/n1j5piBvX2HWWxtytY5l8iCFHlXH8KcyQFTYNOgwtxsoaGlxr5E74kawT2K
ZjvhEJ1aThKOyGnTI35EftFjueuSJocoyfkFHVqkjjjQ8ouBtlAcLZEpDrN9SZK6A1ip5O53z1PZ
KBw5TaKcz4pVk5/AEK2b5V9bV0zqq/etU7mPLjJFebOKmRgwEhB5bZZqzeD+xl8GjgI9s8KRw+2h
RB+qYXdWd+jOjnrRlVGSm24X9EigeY98W6c8PmgkLbtEcujLDHtPSXeBEAFKSlZS69LTQwA1LgTt
r4dk7Bwkrgx7RXkRNJBK+iaE4IAJ7t5S/pcgbX4MTp0LeQd3J/Am0JQq3JKazJwTKq+BOdkbNzX3
OAY9e2NgiRWdSGG6JRfKNEy/ZafC5ukdzj73hEvMExVYjIyBvDpbGQQJGSXwhmuwpdwvra39G1RV
zMpzv6PoQCW0PDd2XrcgYyKuEC1OS6LCe8Kj8CWn0tdrRuanuKWD8wNitr48m4RZofNZcnyhUrqI
UoWG1+cRRauEGFFIy8nNtbqTX60VRIEFTdg2j2Ul0SXvrjd07kGrqE+kQCk04QUqf/RqOOU8oe3K
BgdZCLuAvRPHIHlX2hnJlXYOqDFE9SGuDG4Dj7wNt36dfOla/DAjr7kQSRbpny9tziXz0/5Fg0OA
frhbnFXD7Qbmjx7QcxwsDApTpKoLoIn9JhtW1UfoXPnYLEB0PuUMg5I6aWhout6DeknVviv5ZWHc
HZoni71dY2B6IsIEeRHW+R96CYjGOnEZFNVuU3qGNPEsuWsfY8sDfI3Esxg87fT3eTEsFn5KxB7i
CaqbSbf9Jr47zv585jhBe8xn5zovNMKEdjhbEVuoeCwSMc4CoX/jjjZYJEFW9T9bDOPG8DbLNkl2
YpxsF0jyOtKjIceY9DrbuH8b1DXp3m7+TyHvtQ5Dd4ie6i7g4J6qpUBaP1CGD1FpLofekkb0P/15
iHuVO6CeWCPJftLoJc+pi8oQxpN1Hp9nsuJZoVuHYg6vCIuwLn5TG+DONx4xTVjnYz13eb3fpyDe
Mpyl7YPGKNlQTu1pwZvAMtkmasXo8uk3Sj7aqUW5STs0MWW86ImZpPB8xPTSd29tCVR/y/Ja+FOy
vkFicjuzRdjkpcbhXaCPPqDGg64a3uiLwXDURnVnDBVZ6GMNoev7v+O7ZXuKgyJ40v3swhFPv3u0
jfLncDHz/OkwK6I1C2R9XRyZTxiEE1K0HkSzn4Q7qbsUe6VLYkfhynLwDeNCSO2AXUI2rQ5dNV63
XQwlweSK0GXPxiz+Xm1ToNkm7kMUGNa5UERcUsFg0C8Jz1STyweZsJLR2YpfJAMGtxOh4KEVEpyd
IdNwU/gsMl2rhNPepCpdcSUr5Nfk1mK/bgoQK1f2DVTeyuWowP6kbgpPEaCKRpey2GNQ6DdqMxFn
6Er9Mu5fgF0cmscfozhQpLeRLTymzNEb4HUHZTeZMQETdvcYtd+JgEe2eey13xkMgi8UlUJQ58YL
VfpYrhe3l2FKZz6WSFSpLRbFfjGUE3ZVpkjgsJmVYTLJbje1IGtl3fZUgxt2C4R7JmRuxSUFSZsA
lLe1ITwPu+Ro7gN75aRztKIve3qUR+decluZk13cYXa2MFAC+hHBWK7FnX5coJXa+W9uxQSb93NZ
nZd+2wnBmApIea1b1sxG+FNCEAmspKkxuU6bePQuRrzLSMGUFNa9D555BkeCx+S6fH6xIeuHy8GV
6pjhb/QGwKI4eiICp5M5xMHLSNWgcLBUaYe29FrrlY7qt+oCY6LXzL37ZranJVtRwL/mTcYfzMfO
ByvpYdd1yBLlrA43A+LXqmegUVf+XiZIAsL/ILNUjhKLo4rmf4EAm7GufWqXFPoK7Wop/WQr3sPR
hWnEYmA4/CDI4R6pARxwWq28MKnixF91UWbtqKvz/qAZZJGjqnikP/C8mu6d5ogFDCVzt0liT1ON
JVreFT0W8cwtOPl6JMaobJrGsNN31YRTee/Ok/oe49s4lGbQxEhaDdv/zQW5Nn2YKc/8A8BcHx1/
p/EToFRa2KZDpzkO6FEqL6dKRqAcwqufDy3u7vW0AU2W/aim3+9J+TcLxD7xb/KaeKFvE5yIkGqr
uQJUHWfa9q+PEGKM6NfrhNz1JMrSus0ZnJXlQh8ApfOypd7k/4WBAog5p9YWsSWJ776SXenTldEC
5QA3j8x8T9sqNUD4m/iDCeNv4+Xuv5rJIDwSiuGUkTmr49uGeRZJ6x+qgerw4wcgWfa6JdwINTUQ
y2vGxpXJBiAey2OVvS8q99KrhtrNed5f9WPop32wrmS/qCloiNBwKBVBWnlcHgmDbWudcoGnirt5
lV6RLZFX3UuIzmJTN+LCv+WrjznGStA3wZcbqCooKncrPUFkmVLb5bBv6DOm38/Di5Nla7jZdeAz
0Z/GjX2u3Bmw5tsyYVuRqJbEJjAjNuRdpL/pTotpe4zgBksY4LNUj7ROR09cNT+f06ESPAYnrF90
0GCMlSDG8kIfxjKHM67xontLeV8ViRem277i+bWZSHJdoyuYjWAjd+6zz1usd/diUmy8xXP39GOe
/QV83wwOP2Gv3JGKH990w0ytWp+QXIm8wXsJZfClIjf7oYccbMzK90eryFXxxfFarAXOw8STu4L0
wGMebJOerJDYAqZ9rLFBGndb2TBRAdlOcufih2ebkddCMrb0mgA8jAmGzuRgxMaMy/C0IlhHvExk
xDFv76OjK5v/wQsKcdT8BKMUJZ9olUdB+wcs5rZ8atB0Gwp7R0mJ+nnR/UGfxJreQsOlsgyxmuB+
fL+W+aayh2Ko3jxWzZyixAZav5BQs23WurO1N1ZQQ54jDfMcwKjMZ3LKJhmKqQc7osyu0KkRA6+z
yXLd8SHu8upafePIBtdNxBlYy9v949VS3HWO5Szh5tsy4irlfbMrh3ubn/Z5wcSDXoYoPFEyFIJZ
Zr/wWYBzqYbrv4zCNj2flH8DZJzd7fwa/vZHckEHnE0vCGBNZcW9J3R7tYGGdnTQOsm4lvVF3DbU
ufFj3LpJngM2vu/w0V7Z9JF/x4nFG0nhgqHN75jaC8Db3XG1YV32zhtiuIQ4x7tkdoG5Ljgud50v
iXNwmuYCeFXL6fLVu3F8Yl0uVYguMi8cL6Alr9HWmoBqF/uyrBmIk+byT0Nyokuxd63QaA6kUxRb
8oQwJ69MkSNGMc79pXjWTiEwKRI2+gfhp4Gw3eGyrYQa5+Z3jCTZgeoDhfVTQqJdxHwIAlEJUlPA
oleNfmKQVS+iH9Rr3eNlunFZQyPuY+A5pbhLFJPQ7vW1ZL10tzzxs3ZagkE1j4XBRuXvDXabt+iX
wdMMnZe8A7bOzHznSMVrCjbQ/IGZTcuaF1VBI5IpUEFTDAzJDxPPmPD1Zp/OL7awN9rNpkpBB9yP
QdvgWf2EDqsR/DtA2RE72x6o5rVHYp9r6V491EeTQJHy4TZ9D+FYXTwIAYCih0Xx4+kF5UlHO63e
cUbK+9WKxVcsr/8N6f68CmVT+E4+JgXq5PkaxcCEE4K4lfKha70zLkICmejBVJCX//9Apa1dkn5G
gG0SobgwHFFOrrP82ld8RmhkrJqU10TNgkExYXDe5Wd5R7xKSr4VMQSR+ewsNqWE1psoGeOVfK7g
vtVOes/MfsB2f6KB4oZqCWKBt5Q4Oqvji1zvbAcyTCD188JVF8NzIeb0yoD9MzwyKJJIz0dDuzgY
OGNkYsfiYYx82+W+Ub5WcLvtVhtL/U/x1bWF/0N3AonLZzH77tYC5lxPUzgmL3tRw131uCw+i1RE
223gGzIpOL8P92KPHghirGLQ+o1M5cstb29SeUBh7oThohwsr4Amd0Ljfr5st5e8ZTmypUs7XXT5
WdXWJxHwppF8i51kvE1Yhs3utGOvLr3w2f3u8gm8rWD5JywW9Sz2idC5mofENH3kL+8Wad6Oc/qc
NAPWKxwFBgpN5rKHJLWgQYNWw/2kf7VQXI3KL4PFjzWIHl1oXykcdW530o1zPy4Li1NaEFx+rS7w
usqooyL7X+tzRW6NQUhQKSKviymvY0MMXTB/WMbO3ztPosVykON9no6d0i4Qk4Rp4jadXNfV1EGK
gsgwh5efWk2GvwC8L3E2oK0m1sW7tbzmM4qlxRS7mwFOY9Bxd0e1BlNErLY8abVczg0PO1Em4Zzy
jg5AUHrBFTU2luY5LF53TfQJqxqO3aCdQLyrVgWGE8TrPk+LkAhDLk5eIduY7g1/jRqG6vLHk+eP
19aWA7hgRJPHo95DucIj8sl5LTIxtzk1+x69jY14PR1gc03rxXUPSWwDYDpACxa/xFH5Hbp2M9Hg
nWQuSZaP5QEKdH1TD3ajbJJstF0e+v6aWzMVAIHftnuCYOsjl6DpJLXIxFzo5v6JVJIapp6c5R8h
f1tLp5I1d1LMznJBkgPq62PSyWJQZLriOomhR+/Wolp0kX0DkcPnWGYaelCWPv28GPaDTDTRiCM3
nHGCJB7UGKvou7W0OSvE4fzHUTO7QSFxXGwoQf09udtZIz0+bbkOeApYVqos8nIKvOMyd47A7Tj1
TAJfJ7ihnA6HsOqfHhIJ9El7z2KW7k910xiC7oPA/ik5H6kG9jg63i2W6UVx6h/fp71aYmjSQFSP
SAHc7w6IP1cM895X9XAqN5iCeyYGwe8+7oKHOLXOY7EDl4phoYguh2O+nrzOVkQl9mbeNQx2lH0w
7FVunuT8WYCg8M8BbUP/vVEVTdhCeJWljqdSk6n0qp09nbQciyScz2ktZED1h02sF7y2AkcfyHKX
690JTCtWiFVWtKiDXxcPYPIp0MUnhuJ/M/h0dk1W5awxW9F+Iwz9za1Iwn124cqRIgoJnYC3AmmS
jgH3aUr9a4ClOlC9km6BpRN77GOlD1JXP1+VB5bGMygdNt9g0WhkQ/eoa17FxIbTof0vZFsY/vbc
1fxE6F01cgMsfvqsiiIej5SdTL23OEiD+hu6lR+qcycJXfSRCIswxnNmJkwlcs7LHAPL6APeFWe5
kML0asGx0DLmxzIqAaANz+IjRcOVt7Q2Q7uEbGyTdJJu5dNgFISYgnSpymSXx4zqNF/A06RAdx7q
6Af0mOFXpVBpr646UYt3Qxl9+iLxduxFQlaqENeUFEiKzKcGFGfzEdNcdYO+TP2/f5FnpYXsaaXv
t9uueBphnOGyF5k9Bv9q0rALpcIWPZgkz3NPWalQZhgKtbDT3OYebZHklRLs3wlf8DuKepiKj1+k
VCq4G5t0Ilj554adHJTI2eEZEs4OkL+sI/6bfU1EvjC5u222IepGZtQkPyZEXmyBs792WzVTQLQE
ri/6Y1Y5tgtDYjuqG7IslV84MTCWF9NRXpApC6VlGswHE77Vyu0NkxXpLYt+VBvHnDXWHKsqJTdO
61uf0IQcSkfEZihs7neTMpcRrpgtw5hsVoDPMG4IatPDk0YDVB9eUq083qsgmdpH+qeh9HSaLTpl
VI1qPO3lKtdXHZc3lB0k02j61F3EZonexgNW40fQgyBlFHHpihpG2I3thgv4n+x6GY292HPE2Aob
2/n1S45LWUo0LKaXpI662+qygEHjwsOJS8cvoFmg1j1l6aNl2fcPL93X4+2gn21khH5vDnN9M5l0
YBPKo7dSo+CXXgQRTSXci0UYA/5qgbqt8+Ggoh2Cn5EZ9X51FEnG7H/bt0qPcK0huizA+zgYat+N
RkGrrs4xh9hGUl5Fp5XQ/OkjCccrOg6BSElgy6Ym/K0PkZykAsPzZmtGXk3S7KNTSKtt0O9vjA63
nfhheF2R47Ts8MobLOfyAqxQOuOYt/9PND5rSX4Rsn8WIlLLSVcJdUXav8TgylwwWbE3qAPsMuRX
C2lQuExSJvt5t18+RUP8gwpLdaiaRCGomVuDhAVJ7OXrczqevtyrOjop9VOYN9sPb5dbmSd4N0B8
QCt28zzxQ3ZyvOmcF8fhJydXaWxuuEVVx1UvCDbCQkPoBwwd9UIasth5/kQjbhSUIogV/tzaTWTN
2nFY/PEhLdbhbT4AX90oq4nBpr48jDsZkXgj1NpdE6FbbWWeJ/bibi8miiwCAkxQEyRN2lZ/8CVm
uusSck3eVKWVvtwfjUG8UEjtT2+9NGsf5FvuV+Y9N6ZeAHf7v9FBHkBCKB2YjMlW55fhQno2JEY3
rcZPd5hEAyqODZ6PKrJaFuW3Tt/vN1I15FYJeB/+hLZT/Rs0UMmDf3u2U+ukKC1+JcIGKeFWX75b
BQ+FXpPN0Soc5K5O/mwFmDY3LX6vqdQ3zvFQGyFWmF5cM8q+55tZbdNlcJlbLe0xt2KN4MoidHe6
Ub/fdbIRRfYHE0aWh1bAx+PSyBf5A5RjR0STpA25EKGYqFfuv24oAGBXkGk3BIsRIFbIsMSRhB97
NCG3OzbgK4O/UJka6KoTst+lN2nep8h5VCkvnv7WFqNgKW+NPtPAOrhnTtmDjIgaA4iCCi70p3hb
HC2w7sWywm6FZ7JmgcIV9K5ymV3NqKQ2gePx0SqR50L6928L6Uyt94ny7cmy61zw3Gijswcncpk8
Ll/+8cQh+95M0oxWZlZL8mHmrsNYjO1QdkPMzaSTtk+g6CjpvciI/GSbfNID/yHxMnSDHvRjY4Q/
qnPMyLrBk/o/F8LP0bOql3SPLyyh3v2WAPPI12Ts0+GhmoAapfoRZYUBcBGGgtTh3EXyijqZdsIi
HbocTHC+KnCPsA0r++8OgH8PFc1WCLtkkNIv9z61CBBYOTTwe0R/dS+Zzt2Fqrs1zqbHa1eI7U3p
AU8MgPSssQlIdhcEc8EfblF9h3SK3Nvd3MAx5w9AzNNWBwLxZgxCSSwzlMKj1lSBgsnNZOq7cTbu
6yXhwhTbDNNEpqCr7CD3CVkHbYs2RSDGW4/75D/LQ1Lhjhsjy6I4rlozOJY53z5r/9v1BMBBN7Ip
nxlYjG+yjfcCpZoP0oLGPApfOCBBegKaZum/HSH3WzK56jrBogQ7jY0zgTsCcmR38TnUVOiaGzAX
Qh8L/BLZ46lUleDAXs9Wk0Meyt3lMD0jPwxQJJXKRwwqWDix0fOcpLA+RXolEBuTW2exqFopE3fv
oh+caIYB6+wVqlNGugOtDt9WXqsUV1DP4eVrvGxA3Zp5x8L0Igezwe5Et6yMNn7eBmqNe6FJU2nb
/jy2gcbszwncPSf/fIb95GmU16iwyD6LP440MLBDkqRLsjxFULz1t1PQjPpxyly4Fne9PjHKjSzf
sF6vPy/Y3gpvxKqBFPsZZwGeBst9L6MS6o8t/1cdupKDnyLLU6lApwbPujFUI43Jowz47waOqZjm
K7HmFBhWWQMo+2uT5i0zfCMBFPtGaWH5jeJm34YTnTakspeM8/0QPRanIFGhSy5XHjBqwcUW3JB1
fpN4xlCbE4QdRveq2rIC0vDBka8hDlt8Nb6ofbZCisJD5JJn5FdzpYHNqH2w3loZM9/kBzpS2ME0
wj3cfYD/5OlQG4TzDtHXGPy0HjuTmRTaUjnxj/lz7uuZDzP29kv9TXwlP05lApT5tR0TT7BPVhIm
VYiKSDTaX/QVit59VcZUYUB9DA9xKfIjKfsiRtzxcWa2ZJcYtTXHmaDRVSZMj7V/vM0fRotEZLcq
mZ+q99G+MWGIMz7a9dlO7XVI5HakXbH/A8hcXx5PgTaMYsWa+1UIdZGjzSrEdQCaeyLswGZ9Rcp/
imvmUri/G/vjPyCQ/YTl2bJoa6FAGxGcsmzY7jZWRiEilTk1/YtRD7jWNclptdmPmZC8xsHUVM3L
irU/Zz6kZzK4pSnZFBkTr3pZqCqJVPOjZw17avXP9AYgeKWry3ueJvBYTdYkvqtMMUp+9RcD0GRW
7sOK5+jAsu82P2Wiz0ljBfLD2sfKcPKmp1pTkIMAe0QKTlruzsVPrt2SiC8RE8YgXQCih3nJEu0a
4UCgwCOxf5a3ng7vy/rh13jrjYPnIdUdRPYS6o79zY8nKLJywkkznypq4qIdvBrnbFWNkFHmrUpu
k5E5V2GUijd8X32QfH+sg/+jCOeEAPcYc4nuCNCPZtk880cZcVEVAV7Lyatnqa7wgpFWcp2aJzJh
CZTwGMoQWCcEl8ZF8oIQFlmrfwgCjmAPSoaVt6ZafQjaFoaVhTe72N5S1MKfHMtAkAEgibgKKMPU
zBTAXQMumTdZZGUqNrJJn3SRzCY5tPm4DIR4SRuSVelzdA0ZkfZpDGGLzDbrns0piF1im3diQNl+
Ubb62iF4+mIFgGEleGwD7kwK1M4vO4yhgOTTBkV21Xhxe6TocgG/WNuIcA2FcDr/ZG/AxBcdJh53
cMvgmfHxGWMkmnZNCdeqE6GCkieSVCfQNjNeCj2QrVjWGaQd/vhvp2AhV6NGj4800VbUl+QTKv29
4g8yJ8JgOALb7YB/nDYF400N02gqXFg0mDpDCWzVqq9MOcIMAeGerlbV2pzjvx3a4BwiQqF9qu9j
QrxOQVUbalEBzAjVU11wgfEK7kJTv913Bo+/A+mKKWrLDXcg3o2hDKISGIyKbO562ukNtlTMkSa4
LBJbu2HU3W+XX/A8joUnOg1G0CqY8/o97Bzv0bRAFB+NmuDmpCF3HMYEI0G6SZPDaJQScyf0wGsA
TSsnr5KlcPlzqgYcfVSo7xC02U5NlVrJpOX1ydwrAiN8h1o3C3Ly70rUIGAx9CyL177yk5Yba2My
EehPVcgZxo5QFbqrUE5I51WDXNNeJ+tbCloqnkO4E1Yz4xbl9vFB4vsIsU64TkeH9gZ9Y2zU30zv
N/Ol13YsUpOMOCyiQWd7FJIX0BjXHKr+4yBJ1nN7l1INixt0YNESYHn18jmsM9RERqxyLYLhDywJ
S6UOkZiQEorLFPW/GAEpKaThx+HrDh24cMEDn/GULvp3jZzerdUSoJ0LQXxLGdIm9RZjPad8G0MX
IDuLpv0NOr16jkyGC6lDAreuVzwwBawRvOVcGPnGpVFWNKREtU7QXGR3/6zjH4FOXhfXHqt1k4Cn
C1u8xYdsjFpFllmPHkCDgKh0/xqzRiUEQAC5cFBR0pk69soobl6HPZ5BGIbYik5rHUuwZ81ovsQm
oqxasO2k7eAoPB7cUJHRv7b/UZIaHs+5pyEHWJ3jYln2GE6+6XRkYfo1MNVVBMPSWknqk+enjExa
u8NVtvxEmGznIYdW5ZPJVBxD5brOKYUGUjRTjzweQcJIwSkNpDBqoH8/LfemzROh9Y2rZ204NPDZ
Qkos3jSBb7rM96IZjH3XYb17IHFu04NQn+VYtETpXolq+jqaDvDk1klv/FjVg443xee1d4TPlIjc
NOwO4i9NrkCC01+yN9JdBbXRsdiMqc2BXg7pioZPYuiaSHe5j+OmwPcFboVz2Jff7orlDYSw3R9p
9dig1hdZSlpJYGBiLPLHLy2TRnG8+GjoBEYXDqc6Pd8snixdRrHsRBhPw3w5fXjEU86tTXHL68gH
7gMZkwVVF2ECnvQZIMa1GkeYccoV3ysD1B2oU598hoLcFuQagNypTOEgbVFEfdTC9Iikr/N9R8p7
QS6KpzkfjA3l7FgHFSfv8GQtIarHg6OlaQq9IKpxfKGavJQ4AuOvrnSpbsay/edEAB/GT7ZHL+0e
eHnt2ponLHajel6O92bgju5Va148cxjAXx2r45Gdu0CWjaHMZ5dY1TYF9X9aiWRGtA+UaTvGLo6W
iWZOtFPyvM92Pimfb3l5eHjN052ADxFc8WQVRGmaWjHJYbsx7b2slUUEjv2nmQjG7mKm4ZQ1gbtN
5m/bpOdFimO2bUGeMNQ5lRdrjMzeaF2TyAvtJwRcu8I3dlDuTcvttscInUCytbRvV6p4W9sk3J6l
KyyQmNh9aEFzqflnv6QlcIboeNYfyarAX1xYrKVuYDGwXYfClB4RDbYU3oYia1ZeyoqjTaORvPga
2E+/WsHJCdvjvuQ6+Qk4Y6h4071EsMcbWOsyTH3x3Mjyi5MAAjYolHqBt1wdu4z0YR73ed1xUCdQ
gBT1BQd+ZeQLUvh0jVLdHmVsu2qRKdloSTnmzqNDjZxCQMjwS6B7ezng4qK0H2Rj6I7Lqvajp7Cb
TSvpnCck+1lurHkRAWPuo1lIFSpQafkeqPalM7audkZHNFjokukdpPzeDFerUMFo36rNE89rHa0p
2rK/2SiY1W0N+0Tyc33jGdZeDj6dh8MLRg8QLzr7nQQKJRKhdV7sxm+9wz+w043O2bDPorO+TtGf
nnh4wxJJa5+KDq8JrLNlYXAMGz8ocs+KT6OuMvM6O9XE4LWMn1Lh5vDJnsKUltYr0A+2KCM6cHM5
8uRTuK27XZy2cMpzzwYfaqWH1OcixEmvDQ+NaQ6Tt6TJ3qKioAtIW1JX8DqKIVSfK5CwVy664fVL
yrjH/SdIwI/2+PzReT4UKhUGA0Moirrhm1/PdgtUdRGLZokXZaJU8wNrDPoadc55WFnjiigSqDeD
Xa2sNzqsb4j/T8ngk2nCBDFGo5UBdh8QCJOfM6Msy5WNkGyXZYz/RacMIpY6ZuaNxqcVcqa07083
hs3ZFuKESvBYDCpdqEl/HR2hsjXQRG720g5Q+cKllJmREnZkyuaV7c2rMxlZpFROZiaNk70VVdbB
B8B9KjegrrrxdFkJvvwfWtOZ1pY3lRwArKmoxaYM/6Tf4zVsSUwKKaXmIS7SYpyCAqS/XNoBNtc/
CMlOSa0HhU8zg2i6bUAW1Ll7zQLcjecniKVRyCxjMLkJ2cBlRNIOM058448eS+/ugVlPc7y4irLL
GT2B7Pi/gmWx06OWXZZIo9ly+x/bD/Oxqi1CM/UJKYYXX1lVR0dCDPdyeMmr7235RZ4ah3E6v+m5
arMCmHdMpVFmWAPa+CaUIBz3xjLOW+cBCSw9XsHmroCPnqx2hOU+ySb8JGHVuezu8FPAhhRJKY0p
jlEG5Vk7GcgSsEObNuKq5+o5Nuq/VNCVIH+hjKyYtxkLEnI7jo9G3iL3hHwYVzSMm8o3hQwHgy8h
G5IujyjZv+i7ClD3BGbh1n+wthRvEFNlI/oxvxJR+gUqbDOQPSF9yEolHRug+0Ie/TlzDU96Qqlz
D2fS1b4onOTTpJOoM4wXlbOEHygYgHHdKil7d0oXpcUaxrCTRFGcIqpY2w9jsamboESKJhPlWoY7
TfvUPFx/VsVMpvoCFviHG1iz9p7H7CKZ2guc9/Z0kPqthoUWaEgStjN4dWQPQLXl9DWbviYFG9Vc
Wp2CGNMYFHUH5kv0GjMcevGx0oRdB8dBt/IxL7PMk9IFMqg4dJ62GcZjt/4HhQrCJskuWeUyUxIs
QgRDfj6WnRwpXi8dKIWtjn8wH2IFnAco4ondJBQTfnt2GWNaN7gDfZYD39iVOxLJfj0ypWAY0ltH
P3oW90q8by9z1bobj8WwaCMqEo3nWRsSUlZPygdabDd1MmqNHzypfDPvMWJzI5RbmYnPlj1vuJMD
KBDT2jx8R8YSi5SJ8diIIq2ff29YWkBhFp/esnsFaFTzq3x/JVDl3lpSOEhn8j6629NRdF8S3hin
bZxg/W9u3VOMF2z3YiYmxJSqVBD4Dbvijf5Yj3QGMkV5V3qHyKopVxTVDIxlaRTtY6qgCGzGs823
qK5oidL/R31AKZGx+umt2h64lRARDLZibH03ZtgSbLVGhMgHPHKwqGxjNpSWIborEnGCMc9VTqxV
NE4kc8znAgzcNSRWU0G37rUBBDgxIf83EhuMXVUbHohTSQ5hDfNdK8PVHk9I1PIjXnrEJlWhk7m8
fnJGQ2u2Xgnh52eixeCvehuTwylIcl/7CcUVYQVF2Ui0IUw1qnz14leJthFQP+d/gS6vmZk+UIEg
env/B7EO3g9I62RSDDkPRXMGKy9qmIBSUclN2CJtReXMb0kCDUpmZYTwnILP421fa5GLDjzqEymQ
WZtA+4GdvEklJPf+tqqqlOavyi/nD7dzbYBStuZunJvTv/k3P+40Ol7sitIV0VCL5TvMmCLzE/QH
a+TdqFSKrfQ/RFWmBwRG7QFe6VsfHXAkuftekvIyJPU0PR3wSPNK1pIHniTPqZTTzpEb5MixAEvx
IoHC5q8d7qWf8hDsabUsvbN06+qezdvrTyDlbNRojwM6HRVncs9RpH8u1XQMrkdrlGggdrhjkhQp
NMyyyUIAzDzDZc4sr/97CHiGPPT8GBbaWfyIKXAWXjUGEnfULoZBIEZCSyN0JjgvwfoRfBzJj8Yp
/rrRCMQClr54ItnX8/8SUdmWpjysrCTZawCq7FfokNgKYmHfb05sy5ZL47pbQ0cexXabfbXz6zJr
5GV7QUGO4VfMNwfu5ICM/lnpxbVGsQwXudZhIIekD36MeDGhbpzgKykQmu0mCcjI5CV/X9dF0I3p
xs6ENT7j+oPhKLY19NeZDMg/b+8fUsfuqziAO6wXQ7QKjb46+2+Jfx4PEwp6JcIMpDD8OXOWwLNx
EO8IqLYdJ86iA30fQdz1z8abZbGSCZ8EzaKIDO3XhPPOJLDWWIRFYNUjerTt2FGrPexAFGEKM9YT
AIq1lA0ZBfDO8ySTMwrKqXA0YLweSabxpp/AKGmfNZBGJeSmqfUdR3jKE8+eP6elA5ekI/ucs1Z3
f3IaYsLEBIpXAnAOwF3EG53y463MOaIEXijGOX8kcY4Cd6HPqIYjclt/6aaWq7TMai4CWbc4DjNm
pTlZH4G+Rfl0PECNbaXK/0Oo/bT480qEFttsov3AKFj7uvBjDe8zh3AXyJfsQxS+rGK//mlt+RQF
+f1e5V1v3em6JHM+YnTqXRjjERY1vsVAp+f0cNHStIZ4iaGE9F+Jr+eG3FxEuHvl3NnoSkPnFYgj
wVkFodX3Z7Axa853zBuLi6D61baMeIvxrvhSgOgiInzYecEcpFWvn72/nPef77qAuI+NHHTmftE/
5PPxWDTJDYx1TZ04kUmlbT+QjXOok/nGwjXYlU3aQCrWZ1eMkPYtQqcOTsdUU+X7RbqXzYiDe9eI
Qyf0hIyEJAuHRy3H+DK880ps9XzIRXcRE4+quONCbNWhUR8sj3oMKsr3UTfyhFL9rjG0KeeiuTj9
JPMRK5CAUYlUWRt+vGwqALjtd0K+WMpk78+2k4+5bdaEhfoJfyuZHIyzJoFVRRXHhIl/AZGaYYZu
WqSC/DbDe8Fy+A9HIqARJjc7pB4FXswvdCaWvrYbAno0v3RnRWUVIGMeEMRzCE2o4bWPGatGjZGk
tAofvGCygPXSX6Lobf1BIl1s47oRMbHLRy7xAFAUGpCNZ95lqGBOodxNZqc1E/TAH/X2UBHeFypB
V3XBjq4/TIEoQd612Ugt64erG+PspJD0wvtzdUCHVuzG6TICs/5B9/icPG5Arey6ylBIW2Bq56tj
XGSTsa5YmcI+hQRVX3b4Fb/8i4sODonZj+6rRsh+eG96RrFMS0DzAJs8nouDj5WLuwfFXI+Hz64B
VyJb9yIxEXLNfuJLA+mTOqlBJjqDKe34/dPevLcGeSWTGMCyBHnbmQKBlD1yM/p6P8BVwLw4dWxe
IZSZlrGxj+YrELcqdUg1dZsVkE7zn7DUFxpVdhQmEvDHfZD1Vb/Vm2MnWi2Xa4K/gbOk8/+f3Qqr
dQXC62NXA8xcmCF0Odzl535b72gpnIl6R/06qWD6gZjAS/pt1moh2L6+HsNWbeOmIsAMjVJNeojb
aIOnkdGKyzP/EcDtbzK7fsMD6LUZyupXBoZ2FWoA+fhWVuxOFBD9HSKNhBgkZLmXq+Cz5bMpJxr3
3pPRVKISl7Yd59pkQDb2sboXcdDrKpg0QTCmJozefXYx0lkW8CD7PG4UnYwQUcf1qWiOUgJ+fQ2D
InjIs3xmVmklleoH3Yu617Kb2pfKBDKyyosn3P88T9iETq2+liPLFZyQsljLR1P669/eBzylvCqd
rMmgFiiaVnirJyre+0RsVCT/DS4Llse/sWfZ9nbwNHdqcvlv/0+psovYKqZng1M7PWO5lyVOtmbs
6kmlhefe4RwFSCT8DS2Vhh/m8eiiAM3Rp9IgrN0riCJWVBScm1f9dBVBXmWrzN0C/3QCuyGgBTeN
6HB6i98a73Ao35e2KgwVPEFkyI8VFkFIcuw+o76NReFZyO3Kmu4cvcRZy4EW2EjsgUsvcAb/3wgD
2ohIhsG1LfSCf5YuduJtHt+3BWXX8Xv+9iJinTC9POTX0XdrAautICkvkHhhh4r3uvViRe2wtSFv
tYp1x5bTcdJpSUb2eZeSckYHYw39eg1J7mSS7GJwJ9Qyx44qjZHAR27FonlR7lPEcg2lRNz8xakK
sEpR8dPtSeb2F56ciieT8PrSsLXLAknKLyfQNXSiGGxpHWgRrcU+1qptYfdxmJ+OD0rZ26lxQMgV
RXnmpz1kmxJFiDtWyUkMAp2sYaMVJYEmFdYj0D6XGF01BatmVPN0tNsjrmmOQyKV3PRfx3wZGcqL
Bjew3q7iG4HkWsxp/6FIZsRgHvP8JKSdhP+Ic+cOKdOcxpMPoYwkN5VSSaDJFtQSQCvo37D4E1rB
CMUtIwY+0cE/zEhsQItoJtWbSD1uH72gZcAJ+w23qBoWWGcR3eUE95zu8rUzgIYYh2urjvVQmppj
A3Xsevk+Tvp3Mk1j1IZPl/NmJ2QmdX/PNeRGO+FoVig5WbOq7AzfftzraYLiZZz5yurEnU3rn48n
rD38uMnTn6hQFlrn3ueUHAJcTAJ/VNTlJcKr3bcvJzoAHfySwihQe4wCuM9GX7BqYv+noJ5L7xtD
9bibI4N7Tv8eU4Jb0xk6uT+qe5C02r9cN6dHerOJmie5XcgPs5HwcEgqLrR22KVk9eVYYOg6RB+6
frFn1+K7V0q5lvSD9Rh3Iqk23xwVDxD91k90nE6btNy+DjnKFJA1joAo3kUpKNuFjFbTbxoU2SEp
85u9eAka5GxBeAMQhoXmRbearHS0/AcE2OUe7SemR8VdvQ96CVHI4wcmWv7eDf8T51luogHE0Uu2
6U7kG6gBpeanEp9EnCex1fq0qyim7GQE+xOyhgQ3JPULNoShZI5YKmOEl902B+68prJHTi6UiVI1
IQrTSDUwN9wXZ0Z6uxoMC+4tNgO24/blixHE3oMpcAK1/5vegGtlEAEB04feWWTLmcmp6sh3n5qB
FTID+zivO1l+2Uei4070HOu3ZN0nmFDN0l468ucvtY2iWkgZG1M2Rx6hjLZQ+wka14fYseVajPJa
DyMFbIJMcRmi3AC5HLTHiBHLlmleXCRiBd8q9VwcR2ztvLavQcxldpJZdrBAwIiSH/NjD53/IvZN
XM5nGemt4J/VNG/kQBhFgAUNARDHoq2PW6C9MqoOOOrqtjSBi1LdjKVo2QT+OONOBh8mwCOW7ZPG
Ca/623aCgqnQbquz+PeP2k6UxYO+X+dOroqx/wbaj6l+uZ/0SR+I9VOE20VjlOjOWVHGeJiWK/XW
+V5Zram/Uj7NxtWWO8NuynyDq9uNOPIWzJu7W9k9OYCEFy4UwEAB5PYDfahuUWOaJS3Xldp2EMfh
TCb0gBrP8jRyoqFnv3RR6uTu1H9SNsHacRaEnsqrj96zKVlwY29VXEziB3u49yljqlnCF8Pp2HPE
SZ2i1a8gUYvDCvgHEc5xeVQ9PEJHfBqk5EEkdM6tiwAPfivvuY962bvdO5paW0ac5QWLxeEl7D9A
Yq7NwEmJuOnbf1Kqc1gcGPOZK3Fd9eCmruLLCrylZ91X1qjz9qdEPrKH6ra5sdFoipjtfU+v8Hq0
ZGbIFK/DzqjTiRgsYIekdzj17D1bFqyB9kIa8xT++8GZcBr5a8bCHr76RFhVBi8o8EZ+jD8lYTy4
2vKIHlVxc/hIn95ZIrcrYouNuSIvgfONBdE//KZ0Xq8q3UrGkR2otf2VZP4ckhDDoK1lVRLOsOO+
d69HYds1ml1Z8C5HG0bndq9dwaljqnEDg3I3TQ4hfJjIZGNnIEBHAf1Bvi1Hns6JplX4H2W6iK+q
dC5mr4seZto20aUNZXrW2FwpZS112PVyZOyOwhDlzsQeTsdac/j9F2qtgzIyx+JlXW0S8+9bf8jV
wj/bTXMjj3BcSCuQDOmvyULLtOZ3j06xNSVysmrWB2ZZEfxkCM9ERohZLfdTwBWoJlGwi/pzlt05
5ByXyLlFNCq0KvoBZ/YXqHiQzqYMcrUc7PDDbIQ9BrTp+1hpGtf5/wES03Ceh8HFW5S+IJlLQ1N0
K12jdV7rp+/NsWVklIVtlwOykJrSUkVXB8KHYP4Lv+pTdyBbIWucS7bwpd0hU3PYRt1uBootKNay
Wy++ad+H4/HLd1+P/G5VL4doU0HGd09ZWYtg3PWIRNVMhwqxc1EDzEjPzoV0opCbtrNa8vjYPcLL
ve6mQEYVYarT8rpunU/uDjZw3+hGj2redVE85YL1zVZJU3AGktUOvaDJmz+hApO53EGL3pBsNNJs
HJ8+POrkpnufHkgKqmQSbWKcIMWDtTEAZSiNUQqgSgX3HT5a7xJBBPNmmGmfgA1bTJNG1tI6KYZZ
pDWbI5x64f3CX7hq5Drxn3Cu/PFGYzU7eGbTknfd/8GFYSr/3L0L8Z2/dsO/FPb0xY78SK0YQG76
Nd+IYWdaPo9zGEuSeS+6e9nvf9TrGE8IS7x0IUR+xMAsxi9tDLYbMJMx0XEeWr63XMaPir3HY3w4
WQXsnD+qok8DiPdrGNhXJZTIiCsq2VpQXHt47xNe4ZXm4ol4VE4eO5xtP2+h3U2EskVfjLuO+AyD
RH+gG+cXm1MK2efBep9UuI9VBlRVRuoytWxARpb/BBcx6oRNJkvQvpl/PLX6kfvM82QT5V0XS3Sj
ECbZHvX0pconFq+givm54G4JZL54g3SePRNUieKHC0A6ET2DoF+NF5aOD2F+Z7zJlQHJISlAfXPj
GlEhIEucPL6dzAQcu/SNCqNZrg+AQ/VYkfygQwzVcz4Q7s7LGdNCjBVcDkThbuzG+vfE//N2nOxO
7zCZUZpdWxOkGJR47WspqAiaIyUwcOy1idceQS+2PcngNLnsfF/QBjK+/vIifePi8xaiNjrV2EBY
Qmeaeqhclu+rsVddg/84vVBlLnnPIGwMhRqKLfihkCQ5MFobN0cCka628l6uAcYxqCIePmwRKPE/
Wlwyilf3liXY5mk6rBsP2kTobkxwHK8eS9KVcf86s4FjdPuyXUGZ7gxp3JzCcGUyNw/9ruzp4dyD
LnCpODmJqQeDZZMa/TgSnhDhiWfrupcJmOxkI2ZYJFk7+nZR1DqpScpMLfJXO/BHC4g2t3IN5ivG
Y/2HjznCb6DJ7/vToymdUBv2QDwS6TwNgMujGASSnzXLf2EqDWsI4FQGMHVQIky3ggQJBZGlSJ3f
WGSBro3TIukeQM8XTkzvA6drJNvb+tMFANKzVSGxBw0cnr6UDJMHT9d14xkigT0i9SacT2BMmeYk
0nqToD54JYYKQrRrvTCgRZc/2p3XKmJZ5oCW6DPd35WHW/K+0aEtC8AMBQuOFpgsQJt02HUGki6v
WGtgO11zNZ3bh+I/wbnT7KIiVOFjVKGPBhBz604L985E8pZYkDWlxpDHyA38d6C3KroF78MzHmoN
nKCvF9e5/xOdOmYGtoFLLqLzPNN7E7348i1ymhhIPojfgelHgkBI4ialUwjYnE0KeYtMWGF+VybV
ck3ncdFhoXC8/F59B0OY+z+Jh5IrcCtrGTQlVYLH/6j9davE41NeVd8a/co+mG5QGC4TeojiH7mN
vuoS3dyqV631+px3Cd6Cwax3nWSI652TBUN3yXttS1bz0wKTH45Wv4Tn2yOL6hUwDlDypauVIZN+
p/JLjY/7iL40jHk/q/G8lVRwn6oiMGj8vwQyEYzpi+WEUHJciZs1vXo4TULJfxIRJ9L+vChsKnvc
+2k99py9HkVANPolwQesjHhycuMe8glPhWb37CIhICe+Eyb/SAcYIH1nhOoWcTN28hIfrDA6JOt8
hFIU8Cft41DznSHprKZGNU19pdcbo42zDmXuLLbObxa22yLWsaT4176ZWtZVvq8ym8T38uA/mODE
BH/r6f3Xn7cAXmJGynvRRwDMkiAahMkNUiCJYqsz2XSA6k2BXZpmuszW8qaioY1NqvgVETk/LIYY
rwaazK01IfstNXe2+RdnCdvwZROMt8ovTOn81Q3rdF27BmgxWWPx9bq3PMpIMu/Uk00oFYTAYXmG
vaZc9NNPjotmvhWZ+8quc3BLpuI6NvYZq3SW/Os1qOMegV3JQn294hQdqFDYx54fQU9+kYsOiIHh
RVt1trGIS6hqyqSIBODBjNce4XgRvLgAiPRhiipBAOZm4VHz04H3Ooa0Tpqemo5BaQVTCdAP1MmW
/lXOVN7WJU1I6I2D4X9TYKrqgGcQ3VwNapVPrtY/pCAQKEB4Tq+LLkalmD1uOCJDqPes86UTW3ZV
7uGkclSheKJHY1Yc5oCEYXRiUuCWzqT8eixoIsGr4iOvfpvL7YvQPmgqc3FQLROhmbLfBlgMr+py
xm28lhll6dXpdhARObqMkJbFvxs7qtBSgfB7o41MlhWZBPi9Sxm/eMea22kw/ENhifoWSvQmMFpA
RO7OHmWV3+QXbg4toV6wrEkdIt2Byz59y11Uqr5l0VRr0QgySc860cW2oOtQuWg8SpI8NWz2V/CY
VfPFKi/KTji770IZIWV+cc6TfKKnLQeOntAHFLpXj8ApJ6wTY/vl1PCmOPrE/5oV5X72dev7cxVz
+7fWae8w24Ig1+TToALdgYVennQCKY72Essig3ThTARzTEmMrhriIqPuOBxmdkeJRTf6ocggq39T
/aVzeQplOk1bGSxOR+7qEfgf0nbIRaePsjgYnIiK6Rjcz1jcbw+f0iF5HAsnhpC831vP23szaMyI
6u0fof5cbplwEI6ePjXEBGT5/YmEggkRE0JCzhHXGFYdz3uhvsTNXrXejftLF762mTsyPYylwKoG
V3cG3W+L2zJlDKAsePvEU9P/5LlPpvZSTLyaJSkokoVvlcMUFO360Hfc007+nFKDd8MFWA4QGLIw
RQtGjP6WabtNVsbnFa44cy4JH7PXtGdIZX27t8MoQOzWv9GV8TaZZ6iW4/yCW+Xcn4RQpSGbPTja
RwV7iaV5+8Je5IwwQAW/nAnVBWqBRBscG+BBBslVAAnkUvldj/pxQhe2hW6Hg9Sh46ELGZJ8/2wE
I8AKBsvYk382QOT7Wo5378GH5o6bWY/oTDKIjam8BoDEQipsNAItM7zrW/WkLJuIf8fUxG7NZaoL
B0UMTBsnfnDj26Ch2gIJrVugfvLFxta3JHE/nxzGxuWZ0/2OCQ2QiVz1R7wLVaQRaKMw+prFers2
QKcMRDRfLXwVQpmhu7wdd3rxBHireCtGRQdf9DdGoDK+JFGuZUBFrOM/tm7HHpm6ytVb96muC/6Z
6bt6adTCjgS0jSuyJpYbw/O71tiypgOGySqQ7iF9KmyUfoDOI0sin732nur3GI1zFcBz0n2JMbip
rEZE/trT0xMgba0ktF9o3gOhxJ6DvDOsnlU6WG41ciK7EjdaluVOYK/myo3eKIXbbMCcjYZi1TCg
wrQJrBJmYREArVwcFPQndwSXFj+gGp/Gdsx1J0i1qsmOmk0W01tQNmzQjikHPOaJagstZ6ZgBxDg
pVUzkJF0qG4E50UWavkT0QwzylvHPEcV7MLidNU/WE5IEje+z5VQRsva1NJRdCSugqmXUJmH1Kn3
lOr60RNqoNpGT9xYx1Vnfbj9K9TVx31lWewqm97GVdDK3/0RfRCDRQ39ucIs+EzvMJgBgC14tWf5
K65U1X5HmyZnslygD2hV1qVVQQsHipfVY+I3QU1zvJx0Re7TLkDS/VAWtsnvLPiX6f8qy38sFSNM
8BinBxab+JtbiP6fzaiNIFghKmsPtsa2tiY56yrkozRPmDWWFcVMEfwdxZIm8pKPk4d8B+LsHsBO
Gip+99K9xzs6LKzOgOYdyDSne6J/Hd8T83y8W/1JmKmpue+S6wcARxdLQZ/8o1HgSBhm269N/kdb
sKvDoFx/gBzzerbduxdBbYLkAdoJri1EIbWH4WH/v2kUY4UFy5qhmZvF1UV5M066DFLn3ah69sO0
GlRCgVgS4vXPvQO20pgiv433HzXgLSpUTrUz945X81ZqqM3sgK0dgtYBiaqN6jMmCZCYPG7PXcHT
p9J9Dbn/fwIIxPFm65vsWrRTYI+RKMgGkDOHU7k2hifEMWEJLyBncVd3K7M4vE8H7dc0sVxkbDyh
IL8YZgXijyvUHlbMTkEeRUGo8uoRz9D2E3nO6tM3w76x/6bAJ/dDAFrtyZ4DaqxCBtCLfBc+6MOy
JBdQxWvmwvddeNfR2CwQEoW18sryEDPSya/evaVoeyCC2ow+WD3ADxQGVNR30RJO7sr/EMALwpfS
nldy464qqExrxsqB8dl7OFHMWZwq2TPtfcbimO9P3jiJubBY9DrvH3waKvMqn08tsKbGgaa+oKr3
O5GdO4YNU7AcTQa6ysOQTUlD6UHBephMnCGmYzePyiQRi2VxiucBOvfLkCFOaXUSnDDefgkUN2X4
NEc5/Pqwav1m9AiygUo7xq/l8Untc1gk/zfYSUAJs5B9upFpvubaqlxiHcuEdZ5cZqF4QjFE+B1O
AaITvbx2fOqv9pTdAvUvZVt047kc9KuKYWq/N2phEFeozG4kjVPn2AcXZRjjZDcTJvjIYN4SO3s1
lF5GKtFZupAeGYs0DDmzcAEPX+JZMxi0sjxEAIWz5m/7eZeHQ5JNpIbqLAx3trTUZMuKkY+FqkGF
i6T+Tc/eSo1VBSoQ2Z9w51MGqwHmysYVOTqJU2bjDj0TIHM+xjlM/z6/GE//9z3+yOLRbvD7lq2L
yu7QpXYp0+Rk1WMshMGuZaJArdTdTN6L8w1YG++gd/T4gxdh9TFGbya9+eBFiOSjzg2NVb/dOVsN
NvGM4wUnPtMTCPJM/WzVvs/LQy1CMtoQABfbEykfD+IrFzXBiKqBn+M7x3VfuSXGzt24BifW6Stn
EnrscNv6DC258MLMQ3PLQ5FwJyP5dj86vaSZduVNisam44YgJJ/TnsQ8Km11I0IdNyzRF5Z/OVSw
x5gcNX9moo11WWxFLVWdWvesVh5eqwM03uwoA0DnWfmfCZjgOu90/XsLImkIR5CUAlnVZtkNO1HC
s6ybaKte19OhDFeKanWqzX1i3BZTX37KCO19g95WL2zEMyRxhne0WZa/179XR9FNC1i0I95N30A5
aM+TSIXYiDm64IDdI/IX9f4p+RD+rO9HHpRGtTrH9AQycGgDH1nUVstQypIsYpTKPRopwtoAbuZL
7aYRwinEKI2DT5LGcwx9qmzviSOlljqCFDHpImkrzqdc/1H4vJxnnD6Risx3fHzCUx0f/3qfgQ16
Uj4oBcGQ65wyA56e5J80oTGRjEZILS1WUKaqvHpiPHJI0xHt9ycO8ZSztzHBEFXoBORSzK/EMiML
r4EwH1J0f8+Wrji2Jimn2WeY2lNvsu+14dEFm51NoOKMIM/Dwj5nZixd+65QzFa6pmJFaZAPX8gD
hho4dO1+T6aS4gltsTtDAm9wVcB3yc0FASRxwNMB4TW5xU2bx54EkprhA8nhp3CMskUIq0cAmirP
jgjaOkQ5iqRzcKk6O6xNAXri4gxkzMSntxiDU/88O0/wRZZudFTeHpi4Ef92t0srwLLsNglatzfF
Mlc51DQa93up8VlyPEDAG1jFOhaM64B4pm5rAkFdtLn0NgTzPkvu7bIR+fNT7lw5+pYGHAsXxDNc
mxxKc0s0H+6pME30C3UI5UT4nR2m11KSARmQb0M5UYfq8ZV3OeGKMro90k0soQn+aylaxIUq1nQb
ADNygYsmOv9i9xOBbHSEYqRfA3y6ht8y6QE1AKsNkYEs5xIskOl2RaJGkFBZ4uQ9xVJaxGMCBlqJ
2HLqyekT7LIgfLZMAk9+ssYR47GkA3+4wbF9X/EVM5gaj1b6AsGKBbXmZNSFzMJOMos1W7tXA1ty
c7JF1oBo6X4821plt6UnsePvSTPdp0sPzT1LwN3bTHnuBYHvWfIWgUxe7UzKuShm9zBa92VSzdGZ
GGsvSJiFmlJpDZGmzTfkjWM7AL1sgoiNeJSQfmMU813hhvcrm50ZTJxPp1ZL7oSD8kG397r/uWvV
VkZ0bMQgOpsyFAQrjbM0Orvcq3arWAqRYKOVZ9UZ2klic4cpjXy1hCkyysU+yXHIFV/KGoOTMQRZ
tEvNvUOZZblTmt7MnENG0GZqhXmw9gtq6Utl4DN1KwQvIYVo11B9L0Lri1DvlHnHNTHlcaXIt6c5
RpCotfyFDjyFBMWfKQpqGdRzTwwiF45C8b9wMmkG6QQRmzMSPAkdizlZuYdK197TyAzbcfTQ/7qc
eKQvc/aI4QdmFo6rv0kPhY/vRqePGJm/U2HWCW93aL/Rs3Xc1T0831OXYt7cuXdtM8VtiKtfaoKT
jcuS2JZn3djjmHWtGkM0ATblSeYtEv9gb3nrsJG5DR44P577ih/ZHNpQL5+HJM9E2cw2UO5Pa+1f
h3r1HKGyxaiJo/6M2aHKIvVlYwI2wF7mnpFN2wJ833aL8LS3YygDcCMhBIkClBYopf1N8cEJ3esI
ap2X3TAsVlLMhNpco+tzORJADSSg4VrW3TqcpX0nkvWct0SM1uApK4Vt/+xmY9DaS0auCDvO2uGL
mA9iONR/q2AX2kkPO98bE+gg7FXyKlsng5fqzG72sNGn0bS3xOAe98NJsnGf4iGmOSTiFwcNsXKw
+BVb6aiWi68mdWBxrFyP845RKLK8/mKuXqmGdQqkGQKXJ5qKuq7h2/FE/1ivMvC/Vb8h2xLEzTWv
1Y88U758hqiMhsvQ+gPVWPvpkDlPRJ9TMytdfCdE7+UB2CBeSWu22Ias/MZ5hnONJoVnRXL9Wiuo
SxYTgYb61zaFhUUHRn2oHZ5sqNzvDWSc0JRFP4GeV8nOd4CNkQizAxol9f9AAqW2kmZ6KQVZv5vQ
Vamwftg/F1CAjNXPIZJT42w4W8p4lUEhPOvwjE1Pl16rIixOuOaRMcWbCYIjcgRJPzgAwgJfAZVZ
pdgLvXoEuSx/uAnxmWSq/KMqkxs6bxYxgJ7NWdTkCVx/gW9cgfzcmgIEPt8d7GX2bM0nfLCeLHsn
uyaFw2/R1TF2C6il75hRPjA6UcC3/hVH2MIX3iC5vHKqwL93ZOK7dMNyA2P8E3K/g+w0CHWtH/DO
wYHPL6G1bTmM3v99oTrb+HAXV865lFlpnZi4QvJtUhqx4IsZdHOxo70hoHaMLqhDkEy8xlHVYpTx
nO6EP7bfCJIxw9+dB4L6zj1IEO8K/2lS2ckpjOK4ps1mI7cVAMOsCWYbpVGi5OYEHpp7K0jTMPZ3
XursiL1y0cEw78ZUI1c/wmM9M6b6O2H41RHu8FrNSidWqCYgxSBS+/+JwBn4FhRob8NQ0Y3R8V0a
bULMfuD2Txl6kfJy4dd4sYgOZbpAL5Y8hSs1DHs6FeYddrpWEa/QWbLsh43Z9nBJ1oC1dIfn80Vp
vqFhZLCh10FOyoyZwZ3ATgZQ7kWgC5maJxengeDSCW48wvhugJhrysh2d1+Vc3CosOlg2Kvu2+Gw
rAZpK1s5frM3NAcceXssONZQfgTbPmGp23KvROn+P/Awx+5PWyHRIJChzpAg08ktEPjP1JRoRRdo
p8aKZH/TFF/x60jWMmompEMZXC1VpbQihee2Jf6syuuvZ3T2Rw2NcwAsvSgzN72BQxXUoh4ymgvE
QPsdJc0Q4EHfBLIEwrzmi20o4Otiske0Q3jZ56G/OQy0fdLhGPrNwE6KtYClznRkVWgoj5DXWxo0
HzgFXvlF4Q+IauGsPRZZwRGoZoTqRib3v9e8tLJti7GS6g1gEyKH0gE9RbmS8BeEOsVeNqPXsYRQ
3k9hR9KH3o2/zN5kXKn6dRAUFWaUUx1+l82gmBiqeajM95/heOxe3kTXkQDGxwZZaJnqkoXXlv23
1uf0UUi+8smkGS3vbPzfUpJmsNs7nkMxx0++/WjthIqO4ct52uQ6xTKuWGtkERE7sMHdhd85vv52
fgDLbOZALKNRK3R10MAtpK+MWoY/ct9OHSgYpEoC0sad/Vkq+4KBj/ZMVLnegvhKZIbszPtrTgB1
azQy6v3v6ihXU8Bpsbz5Qq/13+bGnFP7dJNrRevu2tZ+v+FO0Hyph6zfBjtdw2l3pqvG4o3yhnWT
1tSmWVXY56lKPgaQhJcPU4pw3jRuEoHSvlSEPEUAz9gkWDNbc4716CGt/XCX8JUl4j0+bouZl9Aj
trdd++SO9d48LcMWNO2fOWYS+WPRVMQEnM6UUZR+SMMdEYnOv/PypKzEZToPRUOgQUH7f8A7f+ku
1qvbTCorzUq2dIfv3VUuwQMVWIRveU+2HJJ+NqC9UVsH25iRkfAADmOB2+YMbvLsSEs5res8H3ka
PciO5I0LinqbSUtoXraFRl8ZIQxRqNjNLD+ab4Iu0f6JZ5JLWL440G0VNtm87V7VEmR8c+aFkL9Y
W3wVNl5Rv34hlEdSov2MHHuwGTT3SJy3yFwdeaT1NqkFMHh2Pph3tXXxTzdM08pJyXhKLguTt28o
wJIA3Ughxfmo4YiNoBscz39bMEsutc2/mRLfYI6xM4b2zIAYeugRm4qgi+F+NadBSb7BfveZq7Mb
+o7Y2hpZWxpoHXmpEd8r8nGrUvG8JLOk7w1DI7ohfQ2EIQKM5jbGUYYglc/aTGJUn300+cInO/aG
PROS6xnEdqLOXkj9GtpnTB7LXAeM3a5F+H2i8MgaOW1QmIuSclV5boNJX0JP+xZOeT8leTqx1Oop
nhjCKYItNrGt/vWmgVBntISuUwiDrEz6epR1QdXiNIcBVi8nWw8W2tErKNYAvE4CnlWO+jJdkCnn
3OT3D9PVjbzho0suluyiZCrEbJdRMvxEGXOck+Z3rdWm5b6/PLSqGuf73A2U+JTQf2t0AouLJBfe
pBzw8VWP5j0ZwVmGxJA87gnQE7GLnOkPlrsNy5dN9kbGBV64xZsoJHp7mytKcOdd3cZQQP8zInIo
HKhGT9as0Ax3ZjhYRMzaxoP/OEn7/ASprNDFsd2KBDIEGobvsygmE+oNdSXy2GvVlo8dEk30KC9t
SvZcPfD8DHxgIr0449wQ1CjkTxG3zsU2swYCfEwDTmqKY2dkBveXOEufJUfCTjKTPk03WbNEXTj6
YGJm0uYUNn5U3KeCQ0sFbu/zz+BHF4vgBubKPfutbQQTxDx212GrTujXiuBG9OpjPHDTb0PriDqo
BilVrmudze7A6qnG3JxR8MWMYyPjG9nE0MjSH9RgGqSONMJ39Nb4DTJEHx9HeKGJQQ4GczoQqxNH
TqsYS4yrGV4/dsYBl+7j6SkhPx9Sfi9ze8UOzEXFsFKrNhVqMyj8bVBXFieLt9Ta0ZuXRT2QckpG
qwTn3BUmo663a7kDToiI6T1CFWSmKnhMiYO4H+cgk4RXlcSsFF5/hp4Q0O8yECjTvdkXma66CNzM
HtN2BuB0Ejw/6dDVao1mSSPrTzX3oxE6Rs1owYt/KJowNd1KRL75xE0hVKLlpubiOZIV5031/IV2
7auPgD+ph682EXwbkSsMotwBVC6/J1DS3oMyMIkhW3XuONcCM7dhdocrMa9TVqCq20cb5Km1UGp/
AbdRc/XqLDvKE7o0nugBwELXdbH5/CJxDnVAMqh8kx7pnp0f00JHKiM6ywEQW13BHEvP7BXBvXbk
SwvDMHYwaAY/AOYnDR0JeEGdJrBnKIjD0NAA/cxnkakDcXUaeEABOSGjuIbvsvcsW8HNnFkA/nhd
j+kAQudgiSh/au4fXJq8g5o2HdSgfcmbLMqlV9KEaA6Isq6IItivVY6is+8t03p+lOx8JuCtVl2g
9G4HVObVEmLoHnfHkq4Kpzt4buaGWb2Lmh0LNKHr6g66EcDvTcaN6K9RUGDWTkQegv0KN/btbc0G
v9stiFQM7ZoCD93KfPJJynHpNrnCk/AGL6nfbi/O0U9v0BWTOV1ZX/ln36ohXY5Tn5JIpmnmldS/
gzdAg9aloOljpTaGpoGzDHkRLGMZpLHb4NQJktwSw1jkiE0ESm+k2PBPKwLHk3gCYcGjUNo6YSd3
3z7SfnJ4GmycfPL0M2YYPaW/YRAAaUAIK9Eyzbgy6eLbY6z3sIL4vOkb6SCR4YJNYFdse/f1P1CW
vEEQdZ2FosFKVSEZ7P75opHIP5gJd2hEz8ak01/sldqazOcvqiI0va1wNXxudXKrIJQocTEQ53rs
1dSgzOzL5QDQJlGLA67Tni7x1QKu46GbPkFwhjs+uEWH23WHcHEGd8damKHzmzH91tjKrd4BM5Hz
TGIGa6we0okajK64Bc8qN5qmMJybvVIzjWkdXysCdefoUaADFUQbohskzwVdMK+EIQ0ZzR2rAX4t
IgAClUGoo9jcnF1AVa8KVo0vNaQ8O5MU/apu9JzdT0S7fqdkXk/GsG6BaCfKVjGi8qG0Tm0kBxOr
+UhScie3ndkVupew67+dtRoQsBlWvRWg0nrYukZxCcKtmoUxqJ03yOxctVXodn8kYl3gNGF3W9R0
j7RinrggJxe1lxSThzF12DHvoCchkobdtseb9qY1g1DpyU6RaWSQcDytFxdaRfZtjKSOvL8y6zz3
Kq5WQzToynlxHz6l+MsTZA/sgpq6wyodLCNZRKKR+0Oh0hLZqvmboAY7q4rER7Q6XzmbilX0v8tu
Jiq73aaatwyq1X3XeOQDLjjTrpvXjbSwKyGwnxb4/WxOPWJoGjYgtuftBSm3rvu/exfG36hcdyKw
qm5CXOXyjZQPE/Ktqt0ad00jZ9lHbe3IHzlY/8bZMj88ySepGCudosjc6NEpHdhzADpGbddyrikL
Y9nMub1jDX8ACMp8T8vkQckdmgiFiZLOvQNSfv2dryTS3R9YbbeKB5rGXUAzJf+3d5RGI5ossLDl
1CZMgycAU5pmcrCAhb/khZ16JBNFNC84QoQUEqLVcx2AimEP+i/qHdXj6m3nYzeNQAe9NX0snr2U
GZkiZ/rZIxHkv1ER2uAhaVLQfdWhgM8uW+wDlje84nkW08dlD1prUWBxEZ+4u+SzNxcCfVcf51ao
zamh5EA7U+wiPANNKjkflMgfHBO9+wZWG6XqzWJbbgpw254tfUxdPdlxSj4MFtU0fe7+QuYvcqxs
mVLNLTOoOc7TrAgjYUebijWAOA+fsm8b4Fj9xZtIdOmwDJhZuRiEeOY2Mv6gNa3DBDBYhsAwEBYN
9TqtcK4nKHi29ZZaESN0NvFhI2xS8SO57f9eLFIUm0Gsao/deRtGEPQllV+UzMBaI5R69OVc5wqA
mLn7sjzDhLMAw4OTev1yMvZ1PXYh0uSAZ9WVUB0m8VgAkUVMy4626E3xT8vdU2xYTGWWM3esVjH1
/HTIt860fB9PmgJK+vx+KsRXTd/Cegc+IkmG5JZwqtFf1cJQTyVM82NxM517/YkT0N34CAXiHUo6
aoaTYjzlvnX/330lLIq+okmGVIl9WSzuUGFqklodioUCtwLoffPcqZ9G69FTPhGAc/6UGu18afYO
+vpcsinROl5IpydiI7b8o9hSMYNAdLJo4eN9hlgrndPtiy2UnSAFFM5g1Pam9RZRGRI2w1R/4mqC
sxnF4EiutPA87dYV3IuqexXR4ICvuTtCREawjf8UudYJ01tePQNWjYQ7iFQ3He4n6aqQ38CY/nfC
1B4JMNk26Arnii6WQo4XX6ZbE/6hT7YECCj6at31iHrCSQcjWQQ0QfOVhQz5ER9k4rBb6uWf7czR
wxu7Yp6y0Ac4py0xSJXXfsZyvdWu7NxSXlitG9CyhPlsvAppjP8/hxfGH+sAALd8j+RfD0JXChEj
CHzMB4vhPHQBz7b5s2tVJ5OFUSLuRLv+FM6yJHigLLa7E2krvpSbpKY7ximl7nCit4FXUnq4CTEF
982HBd70ye6UcXXfkrkLEEI3HJuzIeybqfDEBmobS8OhhnEhOsQvbekEtFzy25kf1/gqTP0PuAHM
ErSeH+bAfrhd1LDRbczWwtl9XKKvkovJqCJ7lL8iVNcIkkxJ3e94Y9gOBntt9Ia8IRR1LuElM15B
0zR37DbUpShEKGo+ie5b7Aw+cSe0sQBBgoFaEuAbELArQfaTvIWp9qNDqe7tuZX6Tseqb5pPOQ38
iv0i0XKxabjMJ54jFbnGZ/4oo2gFF06TTI4uXCaQYE67b6hm2GneOeHFJjHGmr1cxYX+JydtsDu8
7FFgP5pODxV7pUaEm8PfP7qeLPwpTeavzoIh58OBHlEyMV9Lfyq19/IUyOebK4ekKlaRgHF32/NA
QloODHTXIUZ861LjfEIlWB3eAv7HTcG6wisRX0BjmTvvV01zwG0NW86ClXJei3S4xLGozhY4nUVQ
lvuOLCli0xhn1q+fmwr/DhO6+nslGPEsgKiPns+37cwPmXIULJfM/1PI72W/rkv5QEqeOf7cxfGG
rzXfpqwZte+dmgU3RPZd88Y3Q9HiZmPoQ8gzF4Y7uxoJxlsYk1HYQAsaINz0na7M1dBbfeoO7B5B
VUzF4oai36h4bI7+u0UwGzcDOGqxA2lMxIHBRQ+Ad83stckmClueYf3haTU44uoJCyFNX70qOjZ3
fgN7UNUEPvHCWdSFDBEayL7PPyL7V5GPylF2VR6aIyFtlw4kG/6lMavOrZvOFTFXso5H36ruY0ql
s75Fv4aSdcMS6mobiVqRYQHOG7kfM2p8XkkWQMw9e9fSNhtaDAiEtF2fNoNDmOtmXpN/qkHh2PBc
Xju0T9zmcA+x6fSfXX9AxE0WprPVbD3nYRAASTtMeHUKGMPVVfoHAmP+J3rlzi2eYqiMjfyIncTx
fSbwS10oe1YoCsgzLqLyurUZd2pB/EEn7pc2ym/WkqZF33Fkh4C6nmOgv3LnOeScwcC7Z6U4WTyA
QWNCMFh9pNZisu2X1wGrv6mhSGXPaJlUwtMZ/X/b2tdP7zNd/U1IsxyReAA2p/UgAA1alMHxLYWh
MYZyv+odU0qUrmEdEp4kAgMQWtledlHmpVxlEOZQuJR6VOmypzr/U5zP6rY5mVf2bchj1/FuqnLT
cdp1EnBEKNe/h6asa/0oSCK2Sn7wJuXH/rloJBJLrgSQ6ls3j1oxzaMGhvpAYjL0VWIOMsIcr7lD
6hHzpBgeHVhXuAWI6LBWVsu0BrI+JjJAFNtYxnm7EXW3Wuc22O+Z1MSqseDw3x8T8ExhRhQaKDtn
/skglydNLpINz4VkpImP0h83RvmXW9Haf3HZEBqmT+hfqQ9yweAMKiqILBPFBuiA3N6hY92axSVZ
PUlbJ88zCA3t57RMwt9ClAjG6ZKYMODTyyEtSQ/XnuotuGWjIwl3XOqaE+siHlvgs5ZB81C4VCYk
HMe01eKoLcsPpqI0QkAyKCr5UBrWttWCWArTNEv17cL6k/sk0SOeBM6xqVmBq+L2Be9ssh5LJpfO
EODtJlVFmk+catf1EdMIyvGHwbTrjT+AmMpwTXKYgBcuD/fmc53Epw3hqnwxJSWWxWFOsa7WvQSq
uOxOssR7nSmmvnHp5aNNuYfFcKwmGqRi+7jtrt7fFnDOTAzPQJYdoOyIfHgGWJk9z+t7O2qW+Fyy
5As7xVBzrqrQ2ECVZkQn07pQjaCyPwE7NCkWqyIL1fsbC/bdyWnCVHBNE7D4LAIXTnHVCKBkue4r
+5oYHCP/zRWLXGAYWuTTyoQuvJcaLvmgUhdiTJSXoG/D2uGuoQau6rKETuECJg1LBCpiiIdSZWnq
YN15jPSjsq3EZH/f0IQllKyIpBfdSgnmkWzMdt017Nlgp3q2frg1ppG1Co++J0c0FY7S7uWt9rr5
5s4lrCF+XcNGs0m/2Fqxt+4zD4PKkbDQJ/uXaeNxmwpro/7FKUVVZW4uZ0dEVVzvF5lCPAFdu5RH
DcFRsfcxtDmJsaKecK8sycqrCTOn8QSIGJKGGpNbfpr2CDY4h3qUmnKWn0XxWt3bceOTPm/m7X6e
4TTpqjoiCLBP4k9DVAZtrbQnTaAdRvFlXuK4BTyqI9/kQ/JY+OqVVAhEIomuDJLrZPY86jT3Ohzm
ZOZpq1qsH7emPIthE5F3pBKtaCau0jvB2D1MqxiTzaggmdt5QPxpV8uWkLsEruwXth4irQTHav7j
INri20F/SRi5yYRofZkML/STmpplnlHK80l8H+GRuKbIKZXKNch/BKiL8x7A5hUgpL1n1UwviWeI
flinC4qsbCjex0h5J+ldGOX6frbhIpge/zi4OBsPXkVJ7cRox3vaD1epwnlBVu8amS2XcFMjckUy
i19OkL6yMr+LqOpqxYDJwfyf0hNqfUvZeExddIe0dqlQkTP2R4GeuP1DOzRvU2BX0j6/PgpwER/B
adDg2L3llTKMVWAUtkZIU1k5HeXrlk5rDA6ebbfnjHLqc+6sK1bspit7V1wTr84UxpvPmPCSzLld
W7mx7gHne7YYrB3+E2Sk88j7H8Ax2RNcjmewwUukZFrPBp5Z2teP+qTkZOHISaVRNg9AmYmhKP7b
fKZpe6BEDQ8IJPXIJu1SNH2HZ9CjVUue8im/4TCCeyTWxBdSjYd+khwFk3ARgVTqC5209ZUz307i
0nwLSJTQ6waN2JwF1aNQfgw9T0UUoOONxBh6VAgH0nICbEXSpGQmC0u54lZSOzu4aYIgiBKvcxHK
ZtiUBGfvEUv2JOHsyPlcWngmtzNdaHMbb1IxOvDxhcFjgqQttouX5+jtPUjx4gwr9dfvWfs8ApIZ
9wK4N7DieqqXZJC68rLAVEPCYTXfsJ0+heYef1o7a2mTvoQjESFvTtJHQyaW7IMIY+zyKwgaTVUl
+BQpYKGFoXsVPrlfd/AXE+hnqEYsnueowld3bOMyEKyH2zC28fY7R32Ih5pIv2NwgNTGojjw7A5S
jfxa5pc+LsX9J8Vj0mgegx2mhPEfT9xVbVvGu1pPup+iKxaRHWUZx8m8YksnDWI9ktkh0WRpErNE
eef75D3V/4M1LVtUVZ3oW0zkgeesuicoXlfBaUBuY7rVGF7oM0+Aph3NUdtMqVsd3SVX/3itjDHg
dvOiADXIukVle2NU+KTCERXY1v19C2N3kHKNPXlcbZfSEBU4mwJWQHSP19/aI8N6r0EUAmZg2MuB
VQ5amrggHCX97Br5atpoZD/Sz0XzQyG0pVkWLXAGAOAEEi2jNpAlS60pMrqG7hqXx50Wo0p2JH0V
WeAjYp56NGGKHQkoCNez1NVr65NaoOXIV3BbfduUSyA3io65GQYdawWjg8ovF5RZA61JyWrH/fBk
zx/gtgVHbKH/Xyt7rYmm6i7FgV3kup3JJ00SnXGk2VLdhY+R6bC4WGbbbnJ/ZwoSKRSzlcqHAVN5
DRIVnII3jJWm3vEYeD0wVvkzsaF/l6u7ZuBMm8sg/XVqnAJhJe6dw33O5TSr5o+wZqGA9DX41jQk
4DU2gYDQqE/9uVKq8yKahWsLoLlgRgYUDojzaE59NpmhCe7rWCbi2qWwfn4WvL9KeKyx0f/HyK8Q
3HR6Zj4uRupChLfkEwM1P6mlp85ZLCiJkz4/vRAfUtsSyJvGt/gMrjHpZeJktUdyCLWo89695VKm
XF9waq+6j1dWi4ooYWn7LjU8g24CyORikbJjEFafK9DKKQ56gQMQ/fuNskTr68j1BFs/ycVRG/TU
4fz7d1rDLavHZOFWyJp29/qTqc14XI5aDzo5PV/4Etie2vwlSC7p7YbNeeb+xqZwZXgpqyNj69oY
qXY+cZaWy/S43fwiaqCcBoXdpzCxXLetZFXLmp00O03lITTFfzfqCDKuh09239m50sN1bUeyuCr/
WlvXw2GLZRopW1yaK3G21FRWMjaawHd2ccEbGcQpJPH7XrzBKoXwPnZqQpA/alFm8DdEFC4u2K27
NoouQIul2xne7P6lzCrzIerXAUR9LOzwkqUKtwm8zPnXePOePlKyAE+uiY0/c3yT4Fm9cLzdThjw
qntvVg0PdodctfVwWdM32IyeWToNCak9i2tfS3EO6KYUvdgUs7W8dcLBgk4dFShftqbE4eWvoP56
vdI8t7AIJnqf2o4RnzocUfZHwYz8Fg6hMQJl6HvMRs0kI4xehz6hf0WUKV3dKRae3u+L2T9ggP7z
QGBRTnO9J6l26E03bTWogbzah0pTi761J3umxWn6wfhI/9bTTgWcr3/iG0rjM9rrOcY5ppJMXo77
luPooyNFju3WCMJnF5L/YX+IeBBcRXG8Exnxo2h8/ncufs2QvyC6GX+jvzqHGH5+gRAPfMma4r9p
k4MdBXahc+t7el7pGsuJZE86hmwBqIqDvfu2rQ7K9tSxf2bAGcbwiXQP1fRgd6idaenezQtVqb+a
9ApVgNdQF36RoGrfQw9exK2eWTllZIFnSuMA9MkhoS1q/jYR3hx2UaFYN4PH//xevWG/zIp0rSSr
sT3NP5np/WMCPeCWaQ18s2TkRbBPvBxbevUjn+IXKZNHDiEGSgk5A/QZfoVIl0zwLbcduk08lV0R
hUu1gn3KZ/OOxdDHvhnpt1EdyGmgxQcHX3dz9ZoLzsN/VjT+f2althJej55XMMho6vKcr6V54ioz
U1QJz8uDsYnPG4OKpLMV0muj3SvCjwoA/R+KrlFPQsBjCS6+239PEfvKpWD+1eVbQ1yqt3z84i0s
UOPUNhPNipO6a/P4qvfl5UUChv6GClRDm8ryU+baqLst2DqumD+HIPlN8SLy1JtmDsPsPWSG7SRI
Tmw/hzOrDAhMgDdvIu3+WFGdq0hvI9h8IVefMPPveZpal1SYSlfX2BziXTdXP308kL6yqaqMAY4C
006fo90CB45pV9JXTW+X/6/jJ0aE3tLE0/LVELNT6EpWoOvIYoHTgkYgccquLBrSr2l10EXe+UoL
8BuvDnbaAlcaPXUwd5nhGWCf076AT4tLbvvv+G4OcYI/ycBVD+VITjruVQNAN+XbV9+EKsUXcrX8
Mj0nt5nibG3MMazhgDVWrMdcZKvtR8QPhZNazJcM63mD/cN8G+3vBNBN45Ie+VDDbtpw/eYTDZbv
BHcpdDpwCahGvuyClSVSsMxfqNmbA7OfCZx8sJgzbv28BahYe+DhkZWYwxleKWJZ5YPCQ2B7qHgF
MXzc417O2Bd5LxFUcDpgZdP3L/hX1ia8Q8ayJM8rS9deQ33OjMP8pybhboT2feLWYTDuWwmO6QDa
0r1oOjK5ZaEVOU0RzZA3U5Zv2GSgM8nOWwf3tYFLyuzVSxIXYrdfZGkjJi89GcVF1ljSIoOQcXqt
h8KlGMOf3bbSbX8Ru+BJGEkWK2fKf5kmBwGmVGbzSCnwpt9pWvBbutqRQdwB5ZDCjRemjO59CJzE
2HgtFSncJavb5+CSSeaPJI5EgukNkXQwpKBSAcdmaVKEsiRfMGngJn7KYJwSw6ow3qfC2tF6NDAj
lmM60q1Sg2Qmxn4n8vB/tU3qcSI9gmZPLa5w6SpOoPe363iw50B4FH6vyAdPqEaM8Xqp9+GiaeYH
OEHgZgTB4Kch+S9iOt01Pzqdkbc/oaMj7FVm/cbpuU9mNQiKXp8pUvvyLvPKE2oMXFHSPdncOsL9
qtvPZl0SFJIaXaNiJE0XSOabHY/XGjQ8N5VAdwuW38Slg4tdL4fMWbG8DLxCvgGJucLoSqHdNICc
hfpyce9Ke2+Xb0QgwHNVASvfxAPYFf+u0A1U/1SDNrP0dUm4iXuqv8GDOMfPWGN6fAqhfjz7dQB/
VkL71HZhvN4y871eU6h8PNsAmKpELRnybxRcMdusPTA138+GOPMNqQbiNbKA4lr6xSE3Xc+Slabe
XfptanxZH4jMYFSeCQHmTl2kn6N0t4a2mJZ2JvjVLr79MZMA+2vtDRt6Cmcj75wd9SZlDtP86Sf/
3CWC2tOF5++wSM/AFAXLFFV4Gi2r8j8rnKnn31hOodxADQNS7xUzZ3LCKBLSQg46TrPOA9JXoF0M
FrocpbQsn/m1SSTKSxTFquGYDZIeo5RvC/8S9AyG573/nFQlO0uyqnDQ/R17q6jICMnz4K1YqfCd
p08pelbRjhZ+aVdzi909ZLAPrIO1YLHSFkx6ro5q9sAhn/6FEvBNgI/fWa3568SVxg+mo3z0wmnW
ycNoW04LeAO1vVBOUQzxVCVO/rvvTzOOQw+heorILc0MpQkuc+p31JH5xGGIW1nxrDUlnYno6rs3
TVwDnge5jgaUOikk3tYnI527NkSm+4apyFrpWiqB2nQxGWQLNc1LIQuPBLF320zVDmjPkuMNlRT7
KNlsvxoBsCCGRlcO5A/B0yNy/YNO9+rfbdRfVvck2zo5KG6d/XIYPulm3cirQ1k6jUI2b6W99wk8
0jwoq7sJms0I8CqnKAp8reakM6v1fiWK+wTxt/aWggFLDBiInNEmN+/fnF2avz6YOLpcj/T6OYEd
GRMvoB4INKyVEwdk2lXdXYYhdlYxieblXR30vlIHjtpsdurf/ySwODnCN/rm3S6jJYlQzK2QxZyQ
rVnrAhvWp4IvYaetTi4rl1xKfC/FMG3NeNapMsvn+naF5cGeHeaOVyLqy5cy2UFoI118ApmI2ahS
5TvTTiL41j+F3UUgsgEvVexCz1DBQThyxdC19sLaZkDR0NDofzwNOjXei7kQUMxfJxt87Fh+LtWz
DrvPPCXO1irmHtriXr9zXtckIETeXWdHPAaNrcw9UViaEzOdGDAJZfhi0qBh2zuR1ntHFc0mzAdd
04qcBeo498D4Ab+vVwsQPLpkIKEOtFIa4cy96edJPxDV93AGXYOFd394bscDk+vXKy9Hv3+sIiDy
FK5iZiJZLWXOVtByc7WkwrLeF4d0R/e8b7AN9Q839G6AvGSKxqpYTlW16nwLqBmJW0xxXiIHI1gp
HfP+F0WqoYr/LXZ1VbKBh+hSB6bY3NPOIO+HoLWe6R4mjTfmQZ40SRiIgNS0tHyOEjnMBWhWEH3v
q/hPFAYTSVzylPunperPoSkzbU5qKWqL0JNPrnem8PkufQkqd+WkZTJmK2UHuymIf//9+dqeNMcR
k5e1P851h3zY+pkR08de0P96KI8xStQYKAZr/P+ZqNFeyT+D7duMUPal216jnG0Z7jxgs6nx0cGB
k7UcxKXO5SjoMvdlicDJYs1Zy1KM5T9AfN/AENi6eG213ygIDcISbR9gZSypA4xT08XYtuWooun8
aYwj/R/2n8S6G14NF0Y+ZsbY0P9eGjabpQi0dksdK98yoLILaPtEki/IRuXhwOLuDWUXXV/u67Qq
9Wu5aejKGxtW3xcqb9M5/d5ZaxJqDXnQ8ay0QwqipWEJ5dpJMouXQdufokvragUco0TxsPVoBlwK
jS+PBMmtgwRe/i0lieDCrXrxXA+BczbfcMgpC0vhQL0rJIC9X0iX7zRqBR+DMD18y42W4SWqmi/b
pODM77PjQqJ1AOO/4i9+1pgpWFqjOFbQ8S26baOrd//SRGY+xRMZTlr4s2XZyWBUqMsy+ZPya/Yn
LhMrDEiVCqeVIvJPTfaE5OPt8P2qB5vMFsF3/c0D8XA6c1GIG491PPQYcIIOn5JwFEEvRuu6D9BN
PY2Ynv4OpogLbWesIhs8+YP4yTWiA5VshTaUdaDpflonJ5F83nUToi7liZm4sDc+u3eDFQVsHGxS
/zPqE2DbtsqSggQ7GeeEWw+HLq/cIcMEd8n8+uNaxgExaQ9GauJrwZQflg93PekXvRSdIO7bVEOV
6198F5IuznEoDZ4B+nt1pg8cRsUP70b4wSNq7CVqTvP4iP0rygtGZjsVuYwfDsdaHt141TJakXZs
2XooVzqcvZvOHw1c1OCFmZHTz0PjC2jIat14+VsY7g6XP9tufsuy+Qgr9Srmt2zixyakl9ARI/og
4v6vukRGvLqsamex+JFkRVyP9cXGIgA5JFiL8i3Hrua8iqJ0vWOBh/DOqeTWmLDoXv8YU+TB+oU7
QZUAXiKL+70w+ptmcAvEXr8Wu2q5g5Iem6znE4UpqFid83NBwctG0ZfQy/AZ8JuW1G5lUL2a7Sxy
gGLGsaLHvZapd/EFTnP5c3d6VuE7up6shTZrfTnZdXFMQc+9jJg22GuOc4N6R8C1GOUS/45rKH2g
uwquWG7L8NRoukRgwxPfifGEZnsSv5mVQCQR6zIT/vo7kdRIhx1E0FLP8E3nMh/x52SUElAax9FD
OP/GCM91nPOfcDCNbaDeRBkxjv0Rq8ccJGhLs/9+3rIfMSbqJDKPs9cDAdzFr0j6uWOWvWW6Rxn+
oZSi8BInZSYpxJwa2IS5X0kJf5gj9PF3hZI3E2s7quBLSxV15srQb1SAD/1Qhn/0rKkxUkYQdfBS
JujWckuQJrScSd2zdHkg83Yb05unvzlv5zKpHI/CNa+0JGGG8cPN2pam97lm8M2e/jf2O+bqgY3m
qZKDpwvEKrmZlyhg5w7QRiaZPflTAsNxTYbwgX+MKJACvhN6fzncBOK1wJteZ+zHhQN2lN+sw/22
guZZ154JHUhc0Vaywjw/6rNyqxjk7TYDbWmjKdNsrltpxFcPfJc5s7toPAB3Zavv3fhGnv4Qb8ZZ
EBDkAacn7xWUIIEAhrdqLhEzsazE4N8Z76nYSJ7sWxXjam6C5vaXDY2Vo+dM+2TVEH8DkE5Le3MP
Joo2qq9m4B0+fE23OWilkJ5W6FYHNEYEn66aSNWaYopr5GJck8vl/Ei141F7q8xhTtBYx7B9PuMG
q09xsNRZw74nLcy5Iy0lrzokyJgUvLiCwCfjYMVKhAHQzPuInApiYQzfGXxuEKb2dYcisDu526xI
3ZMIbMbIUTP03bwRfF/45xPQNBoLrmF0mKKgv9rIYrgJWj6kHZs/+S4bPGtKgWqTE5xG5gu5drkw
UTeKZ0Xh/ep5zzWnPvfZ439jC7Fl08S4HT+8qKdPUoyjbNi9r66lkT00Fpn2R6+c1jvEe3YvmCy2
qnfx1eoGPMzk19nOFtgrYzaHncw2PjZnG7hEtHthBBqdfFIK900h3z4pA2/R9ecbcuVasuf1p+G6
6XpuWjzTyJHUHVEjjUjJNBU7F5IAQ3f4rE9Z/lQxoGnFgBcwrn3hshgHUa5qu54sFcfSwasgzgwp
yZ4o9llFpfV7S4I7hZRNiKKF/IXrhswCnjVKpBYN/V4UzLbUP+lrbyNPw7eHMej9w06HrX4+eRzR
Lg1f/aKjCtJyPZZDrtFMueQMJbGHkm9k8JpR6f7xSK81mzHEWa4qOmKiwYscPzn0CrfWBqZXRTnM
NplIjlBSM1dTSTGVa/WLKIwT+TOyESelpxxqIRj+2M5rvC6VCO75zy9GQ5vpFdlxNk54KnfWnxNN
+cT5ScqSTyoj3ZPzJD7Zg3kCTfZ+JX6rHdQlyNdb2hEc5qXVXpL3GsWY97JB4Dr3zSbr6ZhiaT3y
kwrghRkDTa6STkpFy3plGSsnHZCZAyY2tUXDIhrj6BMdn0HoniDsbc30sNrvjIXeEbVjOtZq4ey8
kAqL2Mbg/OL8Xsu6YTNzwULk4zXqy0SxacbrkBXhEhvaQnS16hx4j0lBufNq2O9YaKyFGbmPvAH4
fbbH4uhmwLwKd1DOC8AMcrOjeRVgl5gV33VryA5QpPz3gGazAf7kTLYRzIHlyTHVC8gE5WP2zIxA
tQX4Y5p70lnyRUD6aOfKTCdLK9IX5wp3fLBXDVxr9z/hb+caRPhRzPKimSjnT/DAymUozpXohFHw
vjU5T3ehsI6gIcX1ahpLVu8P4ufgs46+4B+Ym2BQUhP484K5rUPyLofMT9ME3tENX9jvuqCFlOT1
DTpYfImyYGr/Kw9Fkw+BY1OKY09BR8MhocX80x2WBMb+nFXjZ09ulsrfImSm8NmLpSJwoMOCDrlK
ue8+p/X/5PCnbT6XzhFv7MVWw/QgdB3NTspVcaDjhjfCEKK3ocgEeO6xqc5irLO5+GN5iXrn3gGw
Efon9EVmp6N3JzEWFTSgvtmN8v7+vfz9ID5kho0xC21kb8beLjF5Om6FTHdQRTJmZZXS7DvUk6SY
wwWlYvmahU6zCoPOM4W1UQjLstqySZB9VdDljY10kMsKvXGRUSzR3FnSlr89WGZcmj/Qzz56/FFs
UbhwZqtHF6T3soUCVyNzcisDTcuWrseREGtDXkNfWjQiPoXb8sWAxBgI0l4kFC8v7mBm652C99yV
01fJdVe2ZOzFCnfxKR7NDv3NnmzYWsCwOuZE4wynwJWFpxn2nxZ05rvU2bsMN90QhROpVfxaCaW6
wWAkMzrzOuerUnBAAch71+oTMmXJYZh8KUBSqZ5LmT6QQEOqF5w5pBl6rFVCtsbK0pZqepjrZrl3
HeGjVIIFXLLcy/B4TjsscF5wow2tuzQYd6NZKPWfyTPYtEvf1bNU2fyt7Yko1yJNzwxlEeGMotap
sHBSB2t1rqE5B0lIk05dMjtmW6Sbxa0OQMZlC+Q27vvCYGOPUZgflF7bcddXZSXvsGLaGMjOr1DB
f16xTpxdrebtnqAQ1k6Lr/GFdpm6ES3wWHbKaXExMKK7HSOu4yG+swX5YS22/IjxxutQsAx+nnJJ
f4HMcgQYdU4BSBAlDZGokEYKf+Dp1S3CqWxXBf6JamjXmfjxnk4GthXLhoKqPtde3Qj6Ho3lKX/T
WvKcAGRnmbIwXl2KSYmUEg8l/UxBVwtJC7PGM1BJ9zfPelmEfy0zjT05ZNti1EMHu5R8sGCz7tkd
iu+Ju+QyHoJbcrd0yH13AaIShj4nIZvUBc4739MWFl/qqDZ9PpPtD9Ogy20z8WoEdS1L2LNuA79C
ypu3UnRATExxNAPApQDMntndq0UMYcGfW+24KoY0NSWPObQ+1RIKnYFFB+7qp10Bd3sipfkT/COe
d4/wKs7S6+WV4ejkD88PSJabawJvFcuFhqnTqbyIpkRARIS0F9MZqUN9N6s6ZyUVauh5uSwUcGCN
tSNft5mrAkhGErV8Md9jDC17RetnoY9NnDVHvLrWjaU9bqbTx6fF9m88ONYt5V/3gfOrTkl7W7TT
FtMxJ3HPBSem8BViIkff04NWraNSA+oiLhY88fQ8TNeKuZ2T5kN0FbUCViispJAR9XT4pYkF/DB8
/exRu1fKg227gIl9og3RcV0nMR2eQrxGIlmePC2Hbq+YHSTZ8y2qXukGXqpZuhNOdQZBognHEoUg
7OcBesvLnk9rKc8kQlY052y0PE9CzqK3erAKuI7erG9WlcgMXtTQR5xavKWfiqIl9DHHco5lQueY
WHBYA32d+ybCE83PRtS9CDhS4ksgX++uWAwKrHY1GI4PkCBQFwRS7iO0ojPmI1xWFYAzH0AqkYJz
On6j2xFR5ValGNT/stDMCv1GUhT5MK4cwMAP3XdQKHoACedy/pW3QOKEtCDYnlL7YP4Bg5KfjGa6
MjVsbczXeiLKs2DJfrS7hu8axxkwGTKm8OcZ5M1FDW8h322VkQRAMwBOz4Nms7tzINFYoaTBGdZ6
lOFAzAhL3oP0c50H2PG3tual6/GivCmET1y8GoSzXiQE7VcFjEZnqHIgmK1YJrrTDJ8gamtZx5XS
g0RBmsRCd+d5VEgNX7V0AT71uZl5MSI2Yci1QUfQ7T39D+FcxyJDqviNyqlaHv9goAMRhHOMBzK1
RnNHcUon7DjYoNEerKP/6GCHDKqypmlmms/QsTVFkH8b7ty4rj1QRdVMVodolYM/D/wPUyntA7r8
p6W5PwDZpoXbcmzA1I7dWHvQkQw224jRXC6YUiPizyMDJIxVhwhIlKdkOZlIZT9dBgyTpJzOKvBV
jea3gQEWUO/NlVpH2Al9HaUcpy9BZ7qeLe9Lkcul7znZx2BTkwGWao/MmaFw1FKvqUnxfjS257+s
d0UXVKnmoQKehXIJLEX1+E7g3dq19cvZssEpjJq+hacF5aEKyCF+4EXHY/aX5UJPg7vaX2l1bZt7
eCUofj3HRFHa0KlRcQfRNjviID0+QWBV2sck9nCLcgH1gjcUku8pbcMfgcjNkj5J+hNb2LcJIWgi
Dxxqsev6YNA08YBM75NePiLpjny4t2fhdUSBCYeAQUHVqo1SMR6eRuGeK/zdCJy0ddZ6eUDWmvRT
zjXLSGb+9u4qqFRNDfwjl7ks6tUFgPnX1DiJaf/HS3IQ+eXVJ3F1X2fpk3tL8hf0VjjWsHXhD0R2
qFgqNtpUU5iMskHGS1j3VD4kR6XK1FfEyJV2Ta236cnbxwZNiVXYwcHMua8BbOC+sV613hc6rcev
dL4tuH4CAb99RJgvA5vV/odlEaWpR/vpPdxx198BbvBMT7v/B/Er7sLar3Iy62DfEM+tET82Qgqw
ZwFlqI7TX+sNYOKx9MAJq1VrBRVtNfVaXARfxw7MhCnhCGzlk7qnQ71qtW3mPIbZrX2aMOGt4LkT
U+3Nh0JS9EYkjcDttS16+qU21Cb8T/DnqgE1MY+f6ginh3G93AEEff9hwakjgdaIRkXQbtyYimEm
l0mxOORGDhyjghw7q4bIVOMVxJy49RuoChKFLvRikRCWbsBbrB/pRK/i3vzbrbDc0dMYKq3l2H3z
fa2wPjTnnwJBe49gR+8H4LZ3J3FKmnCDztfD4RAIop7LEH4CQKsYvY5bSgh+hAW+drjlyn4BzjYt
H3qRjAVkCPU8Rd4x8FqGo1akB+rqaPqkBCuqja6nx3/ryWjSGkgfwW8/9e2qmNl2VBGRZwsnzQUO
QyylXyk31RTG9H1Qg2rcls/cdnI6IK/skiObA1UoqXEHxlBXIEKsDfmgNTMWRKtyIk4QThwSQ/Xq
9kN3aLd6+uMWw2AlDgbldXzq3+vgJ/8svShVzSFtTu2DeKN4LC++3KneOJVHX3LfYsSayx7oXxsi
1emJMhGaMzrCdQZVeWSUEikV7zG5cVrHnl0Bt8ei06u2wZZRmgSj3gCuF7pwg2efJFfB2DO4jF7A
WwYX6y92fPxxjIa+cwTJwgcbYk/xl79yCJhifYmTJcZfzIZO+0N68YNyx6N9tFl/JpZFEJzEqU/o
sVBoBJ0euANO6D707PY13VlYctY8FyAtoCBlfr70tP4clavF43ZMEiTFauGQDW1p0cmbhawWf35f
eKpBD0giZqQd2TGyzoG0RS3TdDslgVCewCwx303b8DmHgL1uvwfnieOndShdiLunQ/c450NeTRu1
OEQvzq1735CRIqiMrYvCgCx27RTxLie7mj6FlcW4C0njyw6YezcStvbp1wk6cFCmOZCGyos4UXLQ
23lk8JOrok5o3l+GvmP9+i/IE0/mvnpPVq2QDydUeeljYfVgLV4fhmtO1nqgcwXRw6+kvXZMTyv3
45zGnkU1UMz+QO9g72f1Ak/fBH1UKfO0lb4P7oVVJ+mVRlytcUy11wj/hxA3Adxn++lEs7Mq3Vbw
8QyPyqj0bKD/DJOxf+133qdJkZFSt1wXanMNJK0+ajKu9LhajWiZrMetNyuMEE+bLVlBNpxNNaYh
bX5ZnOp6NXTwQAIkutbIRNv0dh+bgP9jEwVKthOcRCa1P5LC5yMZtkD9azmLVK+WnAsMDeS3tX9o
CP9fullmPTbJlXQKJFGyoxi62m3VthG7MHAzt5Lg0GE590vK3E83pdf2W4vlIJiHAedQaLff26W8
J3XkVWMflppvic9KOLHD5RPeGhAKGXODQmJOkK8vOd/x4XJpvs8cXVPU0RoBDfSw6P68HYCYFp9n
Jiys5VujzUfSRk9AAfR7Qh1dz6SSYFfIE0rPe4B9CyYrslxyeEIoPyzkP70rsrrhpqxkqULvEJfB
lKExhq7ZKVzc5u35aUzUIceBbvCYhkR7cFgx8hJhfSUOq78YGfVuZaqxsS3TWn6PkgrOjKwlpz4X
XPCxLUanma8ivSLs1xHBKRDyBQQ2rTXUYTmB0vk39pHpgKmkFEjXFXDNyuiow8Gj10hcip2bpJZ0
U1ZSi11xGr3tAxKtu9SstT2lgGn1iJSLl0WOv5qyjUqGt4roaQFImP/88K5ER12Neci6XXbE37sZ
CYw5CwY0SqMgt83Oqbu58QOSr50Uqi+95OHIMfgxI6qOrRpj0Yyt+CxcGtgQCGW7Xn+PvshNfNv/
D4quh5k94IOeraIQn9tipiqpqFAanzDNuqKrmdmng+AwtWC+wV3xrsAEbgpyD8LcpM+F0P8yCM2D
N1fX3t9s+saP3uoV7FVtemQiQrnUdgl4uzQ/J1nCDbWMK0c5xE0bg3mAWvmDcEb9m/llgzT4rj2d
a2AZoKRBUPF74m1tpv/hfll79a/qkb473l4T6zYCL9c4sQyHfX/ZLpGYfwJ7oFoiuc2TtLG+HtkQ
GRapXRcfmLOrr/edypwjCfEDs75YU8Ykcly6SyQyrbEzilOi/ID96PD0DvtgPAXg/m2+2+0tkVfR
zwiV/YCroxqk262QCrKljrJ+mnDmwYUyRJPWNSF/uw7Y+tFS0e3JOoew0BO7/7Pz4tqgQORkJnCm
wDEKndqqkVoADADG5/LjjfHFRBlllE0u/l99n/MChXumQn96+ugdaqhGk1Sj/VkOhsi6ajDa8v4H
rjkit1ALgM0fScpzw+06g/15cowYJLV2+Bt2+kaYoG45mws4C+htuQuJRsbWR+H821DzqbyNAkhK
eCWYpTFFRDTKl/yveGCAoXtCpx2Xqif+kUcpWD1YaDnUw0Fh5Xc4ejVU49dfKvkQuPpbySfJnGtR
3fnPiUxGlop6BgpmYOw2pNVeWQIMdmrZ/VZVDAry/Vr7bpOlQdjolvuZ0+X/29/IoAcbaCt/RBgA
WDUBDFyxlDuDmtWMScGDoTpY+WxP71LlAMSFuOVg5nHa8JtCxKgElR9A4hmwEgoVHsO3YAZ+la7W
+YXj0c7eL/Hjd/lEE8tAORmEtcqQF8T8stCGBmUINV023sHpY1WouQwErd+p53t479Gb0ttuMvhb
SQnx1pZbvc+bOUw4i5Gl3cMFP77jI/r+X12ynRG6cU+vinL1JRcYOeQEN56r3bANBE7UD8hDN8Di
UCfbVE3U8J5baO/OoJqZ5fhBjdgLyCSP8TnXyiDIwKcnjpaCk3mq7BXqMmyY1oeVW1SCf8pxnP14
QdOVhozms1uc2FswVTEesRhrWCTDV7u8Kg4PJKPJyW6RinsIy5U8EtZafFky5ToT23DsjS0w5r3d
g3AO4pF5agjF/nB6c0AvSBIYuzeIOD83RAlwCi7u2k+1q8b7eXEDMNQsMotxSNiNy5/4+66x2GCy
8RR7KwNS1H3kPoIEr1L5JHegYX/EOxHmHjCA6rZ8EO7QBaJYfLJlrM0k38xn/f09HjM8pHiWkhkI
KCp/is9gnqMkp5TTOt0DQQzhcQ16ujRA65DElvWy81X7q2A7YPVEFKMiiiIyhFq4S/blCPaxExIr
FbeXck0nUeltAPYYFk0RwR36F9g7zRTh9T552L1YqBCh8oI5JCYipBUhu9O082IkZwAqaMY4FnHm
Vi6JgX0Xls2zE7LwAInr5vsJk1VlUolBHcjwUR+X52EsrsZA/L863LE7Lrpfx9SwLip6/3lLESfX
19qq7qIAvbZf9yN6Y42uSH4ou0IUmJf5B08Nb7FzmnUx2B3KxXWpAnzb6O89cUSdKNf+/Nn8brfB
1kl5prgI3Ot7aiKNcEpeKUJPT4HLwpsqRKfEKoGl/O2/JVHByRAHf+ELL78YVFMi/1K7lE09kZYD
sCKIsk/9GNHZIxYQV8lHDvgJmrfxYpP1fSqqRrJVrbBa7iQ9PLtc3rAl3KBMaaa565/27aHiviu8
p7G8n7zE25+Aigb4cCJtiV0eJvGjy20eXFoSaP54iBSBGI0OkZxJ+gzqQgc/2VCNFniW4dSItMmv
G2/uBQBZhI5snRJGZo8+bkyJjLcNrSAIaYJnp26nWZpn2JTujRf8uMzeA6ENVvj7r+M/vv83uhKT
OTU7J26KDIY394XWQNXPNBAjw0G0qkweuBlF5iWUGEztShZKppsNifZHkK1m2qRrTq27nwKEw3Ds
MRvvOMRGFego4OB9KdbKRJ5rbhgY7HhVc9wrMBSYs7Xjgo3XZyG8PaagkA9gaw1vHW1nOp3CAijO
gO6RPc08Qr4AySj1f3GWIJecHQp+1vh38t1pIZWPqQ68fOUI9gsObilEsD2gKVHtrI+29e77Yrh+
dc4oAwJynw/799IdxX7aV3BPYy1W5s/VYucTF6rr+MIdXmoYFbO2vBYNqx7v/TLPasXNMK7LVe4d
Sfka2VbMOWbEdbJJ0pbDfhFF+b1rsHve+nBK6lIArakNUaLXW7WMySOcG31sRbFqlQfkZ09hu+46
0YcjTgs0YzG7qZgCaQrHwQBvYsg1IX93yyrDmJqYDkGPbJ2/V+iRP0ZIsuhmUTaxWva02eFywowE
BQwjnQKkIicXOToxiY9AWn28K6dNbUFpPP0Q0u2kuw8TL9xDp1A2WJYFxoUXXw1Nt5PKV+Ch+h6q
cqf2hneLNkrmu91zkXPrpgZWmatoKXtctn6TciXDGyxRDlOQjcnHcm+axb5dpVhwTrYYfIRSqdyd
YtUMYnI5yhiIGKTU0Pm79xK4YMEN8A6qWPZ6zt+gKIJLDKfdmvYxiJ2aB2E5WF8kv2QsFnhKi/0Y
6Aq2NuByRxqe2Wm66Yy9rirnaEL9QlRUMH6//9vYQO3gPeklecZ9xwLnBKnzdIjwjGoJa5loJ5jE
WYUvdqVfYFX3LkmqlRAz807M8HtsRC3g1QMhwpjFUl8jIV9EE62V5SqoK/LlueGJct5ALAEJhkib
XojCF4ovQ0dCUGqTr0BuiJs1XJFcx6hLSytMhy4X5M7aKtWClGCKA06c7FxmRlJgLQ3NC9bLHaj+
rAE33pIQtA01vB8h+bl7ihLYjQ4UeYYzu3Bh3kwO5d2NXN7K/aKJRlJ8qSMbjqT+ccb3B3vvNGZ1
t+30fdiavxzF60uvE1mwt5/CLD7SKs9y+njiZ7kXn7bgpN+k1mhoKj7aPUJg+zJuA9uK+ycSoBBC
8D4DKxiKJEPXcRwZX6Y2y5bH6WKooCXWMEST5woXiDssEIRGAW2zlOwEnp9nDj8gbYaJjHKa5OXn
Gzz0qZM459ip9HqkWE8mjs7ToS4/tX5EN6KrhZ3X3PYXzcZSrPu3rU3FpzMIFWtGDHY0QenR93S1
QOzUj3b2mO+jsw/jkSOipfKaXMV98lD7WfoAS7msfALewuXeIl2t+2TXVJ0S7Cf/R1/u0lA5ngKm
rkHF1NsrnLBXUl9obJBqSM7N4uIGiYO3BwdrVUjPfz9TR+gB915YX/4S6+zTWrdo8KIVMTNgI82o
xPOylWZuBlwstezY+/C0KVYpHf0HWoREAxIjTiOxaR0PVA/eCY3mPILnP3yjjyjNZ3CU68ZAdasH
UT4c992FjZbbTe8QAKHSsB29WCCruEkn6IY8Glk9v6noDNbXZTD1D1dfBWmSZYHFK6iCnUbElWCl
5qQJCZZ/iVOBZd2HwQwyQLyfPFROFEuDT2ThTnoLC72tXCDgSrT35Qir9narkEy7xyjI5Sl4cO7I
LoqsZXpxhCWvYE/oLTk3IWk2Xn4B0dyG+879RzMUHPmNiH83yw4ryPTmMIx/HFwnoJBWRL/L6TD0
0YlZ67DwrRu7iSNwxOkBdwOLVT65UYUTXqQ//5Z0d42AgxQO/noq6YbBvr7jvIt5HGv2a+Pkbmpv
S8y3bl1PxnB47zWht+DLqIuq0Jr4SXGWgJiIAme23GSQ1XprJYzxjmtUq/xIwYw19DGuKHYvFh+v
Utrv0eoH83YLMTq+7484gfssYszkfiqhRdPnV0xmCjKHCcVFZVN8wl6vI1e0GQorHOpSk4Z+LCSL
Kehox1SPsiUb6Cn51Bg1nRY6AOcYzxEHE8AsKwwsZbONXkb1tF9QmpgbQueBUSQjKNrduLX6fkZK
jQGF5aeZ6vNwtzdemJiLRe3/MlP4EB0Mxc0m5XZ8KcvGaory6R1sKGlvEpoAo3bZPZ/LmkXS/3tQ
Lu44YXB5WsUOQmZh2OmB+Bar10shvr7yBzDR36NbVXwF47mTMjsxeyJAXg622KwJK1VXaDqn1GxV
+JBU8oUwGh5KYiWOFTpqtgU/vtvyXWNTKZxaYftfx9rW6FH7r8zq5Ur4Xw6tAUdfOldNDlUiuV5R
y89ehBBzM2MmT9ya+scpapnII42uu1IZUkmutQasaAGYoDbyLmoo8yg6bvnrNWuKLG8sYfr/7Dnt
m6PZ7znhFGeEwT4QE1RRVWOZrgJm6EBIvcBOTt2yIIBpZwO2Wa0JJdZfhEbmHCfA05ap+t8yA6E3
8hCqigGZMx/RRA5NzbThwc7TBwBMt9VATBinRV0yeGMxEi9zSxU06QmwpE3jI3Skyp+sCBX18miW
o8Vv4YjwVZNTsvjDbRhG5KVhV5YZM5gqYNVWH4jLsWxjSGbhWSNA00jlZP29eSJq7hnMdP2iRB4j
Fmo3+DriHpKj9C1SSt9gQ+T+uZKDNNGYvFAwNakZqDDloXjSsqeJFDFsWINxJPoRppCfJxKLFldX
1iolmicDoTGq2wh2cjeGl8cJz03zEZR5+kmKUeLN0CCo9EgdjXFZ/4iY7tPw1SD+6taFVJmKDG48
JzFN1VKc11iSe4NdjZJtibvtssHHL26sfl1CAuNxyE3q0Eh8pS1Ac8yDCC4tzA+V4mJ+60per7qc
kmvYfYvywxpbYhDmdADUXEIChVfSs8GsfXGwis4QY3Sw6hZ0o9P83Hk41lGN+e+0Lxym2NAJNSvz
OYb16DkAk3rzb0xgapUpi2uejQSoEQLsqW02OcdS4QPb8W+i2AvT9PCdk8/3NxenhmOa2saX8zcd
+Z6S6BcPFe3mKhfzFdJAJG6xG4SFWuruvTFUX1zxlgJ7cFbwgGWxafhdCRfVdWoGW80IfSN0Oaxj
4VlWQlipQ0Tfli8B738hqAZ2ODaMebw8QiIR8c6b2o88ccSq8rFaY85sISNmUWFWSqp/wMSmBIsW
HnpwTT/jXA8JoWDEaabzGi4r/6VqbBE7+3DbSC0oUdKHhMyPVLKgimORA1lUEr9DFN6x4xbi4bib
6Yg1ZpI+SM3R6o+lnHUiy9WQR0kJXzUKJAWeiaxP5e8BATaQru+Ft1nO5pQvvaZwBvQLKXc6bB9z
y2lnpNe5mcAOb/uNpa4Ypc1lbrFj2PD6SoS+CwcxylzFaqktXeC9CbcH0XmcX68hGJvSmGwosTlu
mAfy4nOMsmfZDILpuofZVRKZ95Cvz/bdjqFeqQGWf2IgqHjf+GQhN8ZqNoBsv81Xd6ZhSJdvkCgI
96qrZY2VLPX+m/wwLa/RTwqzNsEF/x/sNzolPR19HX3wvV4WkUXq3uMLKKkc8yIW7/G4+f7N248v
ouSPtYKQZ4UVE78tJXKwnuXRkoQJrfq4xIcYXmqqmO4tIiPsbjyOd51DPcdvsXHNGlHB5O8XVoRn
GCQsBWPZlkAKHxupwg1kN/y/BgYmrBPlSrr81ZhpZwBn5IH+nigXqDJkIzIdHufq48gExwpeu2iQ
Z8w/SkmJyJRUCszadtJjnnbOHWgZp0L0pQuK9SSbgeJ80V6SxPimdZDr68Ct3gjSN0C15fbQJuDJ
dukVEqoIwZSHOCBxmlDBbCnLjlIePHgx77XBnj3RM7bMMhD052KBg46GBeIw9qYtY/CFTwz7RtR6
ln4jm9zDwBwBrH0+29XIb7n+w2wgbb7xHiAeIPnrR1kTU6sCWVktjO/5pNzi0mxu2V8etUXNhr44
cbVSv8/0r0t6a8w5k0uD7TdnVj5mb+dikbegu8UORGaxJtME4XjhEv7zOz82nwEi8raAxyt/1UvK
x/L8wE3+CLmUO5jRJXnTu026T8Y9EObq3viQOq/Bjj6JMCKqN+QGzk9WBIeNxSclCCyMdiHN2ylY
0WRAbxEKy6HqDBYIuKCP5ofXrnFD+VG5Rn862AuWnFINjPuTEUTg+6fHtBp1m7CRHWRkp/83x3VJ
zcf8co51AqSLSh9W8GK89+ASXx8+Jayh23uEyOlF4Nxg5rv+F9sRDX0vjYtfKRftXTZc2xMp69RT
11HmM2qfNusZ6m257YmLcGA94BaYlPzHUeTSoirlmMG/ptZBSlIZ8sbXg5cfk9O+dnHTyzrZhTNW
pBND+fLzeuZoXxkFqGxvz6rZYZ5r2e+UJIapBPNqm6sjjVF1p48bqn5Y3BT7sQJHWp47omS/ZEy+
l5J5QMvdE2D0w0YeX6QsD0DZ1vMqzeEvoC9a2txBsMfyS+ojaTYmfutak+rV6r2c3gnIh94Y7IFv
pOBC0AdDh9l7dRC7vWe/6FfmFdjDhYDosOXC4/KfpTrU2MwSTRG0R3Fm2fExIYCCQGGjWJFJ0tUx
cI+eIPjEz8aspJavTTQuuUVbZFNaMSczA8+/Zyp2pOamkH0hUGr/+sE6vUXM+96qD1VvjxClY8oq
BD+PGo2Yk8hgh5ehs+ZZXMS76aZ6sVf+U4LHJ2zW4Px7HPADXPcS0UyTSQwpwlMxK2t+VHsrh2rt
vABzv3OueR6h0n2u3XMMZRAyA0/TDSCW1et6Ycys8YHOKLjqRjzWwshHx1x0S74kuGejy4cuXSSz
w7OMBxyoJNR0o2RSt1rtjDhvnG12et5OzV5/The7jSXI9EATbXQGUBRhqaDDig3wsYuAejeTwOtz
26cO0xxkbZncS7DLvWPGTxn/79osJ7wyR+UvxfAOOBGXCluQlJqQpNtl7xZ1QK6YyW9ttwrpgubn
jtbVLg2z6kJfKs8r6C6O7ELD3hJcPENa4Rbmuodtq7TsAuL9PhGK/ynepTXjTm8CmTSq4uxe5x0Q
1NPzwUylrat28r9oPuS0aLQ4+ibzTHV7xD+547QZ6cPZA/ZYvq7ZU7hrgT3mAz9tmTtSv8OD+ww1
c7nou8/WmE1caCahyla5P6KuHlD9mTAO10eoYQhRzCF4DXjSunC5mraU91/zmDv/M28z4sJzq1Cd
Ntq7hrQFWSPCngC5skbpI4zjhmHuim2TZZSs4B9v/lf3ybS888FQIpmkpiZTGyHVewRBBCL4g/n5
6+YFBAP+A7cFrYeyqS44ABuwQJZZMiwFOaCniIh8rRHc29L5IeNYwiTSUeIWLllhBGJ5BIWTO8um
ZU6Qt3l6MYclxq2xFrPIHIx5mszE2eQAgQgvDnPf3HX+ABPkEk+R4Jo3Ac9vexQ5Of0BrbiqO7dw
dKyGJCVP8V924mzT9wiGmfV6N6thMl8GNWgaIsY/sQXAUMdYwz7p/W5iy8FqW6gtOhJWQd1OMczi
chlMGe+Vca5AThfbLWsiGNbRykUgWgiJ2SRwP3VfeXSBhqAB+q+Xf1FnykhLQ7vzaR8ojNCoawPU
8TZJICd/JElTkz96ruxoGghyFI3GL2vgt8GtADKIE6/2Bbw3xhJ1RYoBEp9OA3gYkqxbFDTjK4Ma
N+hwvVkrwu3AntH/15fKiT8pqp167yU1Iym/fCiq/wryFb8gPXi0Uy1KcD3PrQPmaJ8FXJjZ2+DM
z9VKXNIBqOxVtG6tJl8/Zmo9opMhp95ZOS08d7jK1S/MHfJoas+LR/a2l7yBiZ5JEn642RjxI+bk
s4aujhHO4/FOPPDHmogTVjf/4U5obKc/vpqR4tg+oBAOSW+gnYpLlDbo8plu0k0Ou9SpoyGV17W9
i+OebONVZR3meQTNfoLcL02KTMJKPpgwTDKwM0UJ1+H4CAPc9ItHysOqp4s+hOYsbd4LFy9l2jWV
SXJszfAbil6EJTkzfJR2EHDxMAvhgz6TcdPv8kFjYSegCTnIr1VrAUd+Z5GfJgnTpp5DMUer7+M5
OgCbMsIoBFTJzjKFRMukVb399Va3u91ArFAbjtQhLMvDd5I3hJA8qajM4MYt6AyDBbCTpV6OI3GT
w957NfXkcipg6LsjVM39LsMub5cZR3ydltXREDkDN/gjQ3BNhYOgYr5pv/AiNhK5ODcJMrapKMVV
fA+KJGnRFwux8SIbIyoOcwAQ9ADaS+Y5j1uVIKiDBe/7W7AtscE1QZZROjcTGtKCIMVrs4kEmTfC
2mxtnU/vyHKxmyDL5QWzc6uME4y0ubgGJ5Dw4Mqx5Nru9xIY3geCKKW9cSvmRNN97wDO2wKqK/24
V4FHY8mwK74Y/EBSqv96CR66myCLjfjEIm0tICAtMkN2W7Ic3ny7jZLwrIEQf71UJ6y2E+DWGwBx
oeILql2hOlinM2asZF+eRjOixuF8PhfUBaD3NAAtB/h1sxNms5W4NG0uHCuC1qbgV9X1UBOFIDwI
PYzU8JY9YLpEWwRQxgI/kbQWmuvtLKJIeoktAKmGG6mdfC54JagIR1gY6jOjHiRKMoNLIXWqFd+Q
LGH1/CxKvRpEz/xbt7MirZzv/COv8Ly45Uo7YhawKFZ/6siW3yBAxSqi0YPzF/Ddlv5U35esIbrw
+sv30Pv0GHXsYVnHqSBwpSXG0rdJzTw3zCSpsfG+QnT0MxKXMzADh4KmeT33zCPZ/1F5QG5Xq41A
aGOmel/6YP2JzDv6sneDEym80tI/eWHzcKZc4pJiX33GFQhZQaCX/rvSPkr1y+UIJlrkmJTqfLRe
XizOWkMAj76vogUrk632JwKt+4UjFmWxycY+n/C8NQCnZw+BcwmxzBDU+VVPfzqdrMSaVV3ICwZL
Ix+tQ0iQUCgPBTEjKsZ2+tn8YrYWTAuoPCuaiwshN9oN4pSrOVnXyxQTKRMu6bNlV1Z13kJf7ZvG
Yb22OyW/n26Yh2hgIv+eDV/NGzjIvI1m53kvVjWwvqQqui6qdYEJcKfh3N4L3b7Z/cvxHaaVxnUd
ikDAlMenz8d31+TQaP3H1qyn47h2cdnGQUQYbmnkd19WANW/JvKqB9Yrahn59ISJSCidR6/1dEj/
Cs9rK0KJSs42u/9X4NLcVFJ4HgO8Fq66PylDSuNOSaf9CaKsK/fuiGMBro0j8QD+FMm8CagCxmKV
YUjnCrOBlqJ/JP+K9E3EdNHjJ0pNqxT32gFBsF3K+eWqU2ZKxEls66EXmOEjqjDkSA9bjPUEvMUP
pQNM1RQ/34489M7E2QotpKyRE7gJZimH49iJgV4zV6VozoIQfQxw0NVwrMNmrDsE6Bp3VZWS1/Kt
ogh8AXJlPzDvIR6UwJpVZgpe7bvpD9E7XD3FBw4oo4ztCgNTSHf64PGe4+bbVnORNh21ySEAlZgP
v/zvcwqyg8bv3sUAav3wxum2Pxy9Xrg/Ivi83B3CxtHo0H/q6mw1iFAPPASnbr4sM101LqjYjsSU
Cz/BftF8JHDdeVGqbgNjTS4S+GFQwnO/5rrqtMe9vi3RTJOw/1anbu6kMz7COS7ZmMx2+zZCVMgo
67pLNbgbhCVdyejPMcjHu02cKKKVDG3YrCXrE8qj1Q5PkMFPG/Rx9w4uAEs96DS1fgIdWjDzDBfh
0mz8wQ5c7jafLldQeMOlMpzJ4Fl3c0Nk6CtlhF4sSJnqLLY5LZ3MBFuVPmCZVQES0MRQ67so2McI
ltor6GHG2ey5+L4PUt4wxYv8g/WB+IA35SeFuTHpWWzOLGdqejwd3hb1qn/ewXZUyn90W8GM4n31
g1boCU2uT4tKMKdxw3xpxnnNDg7bI3IoZ8her5RWYTLCfzlheghmC4sZMvYCU5FBT7e2PMrsOuss
3rgoXSa/wt8j6QDht0SO3rO6Lp9tHAdqOMQm+rLhIL/O9G5qF9MXhUKlryc8fM3vB8ecZqfqGFcW
qZN1LEuRrp365Uy5IvcWqJYmJnX2Ql4AlBxDBzi5CEoco1lphNPDx7TbU6OnHGOOcI4yTovI4o1s
ygWCALH2N1v5U8ixsXWHEY19aOrA8enZBgdpb7mxc+R3Hk4CQwN5/FfLNuPEkSFEEWHmRDkMOKoZ
FUUQhCmB2gaiV33Cg4XqPlxLzXic3GCyDbCNTlw/taDPGYAXEmYnF3AFQkeTv3gHDaG6RbyG/slN
oeHwdpizkdsxJcmZ3AwfdKqr/7dCEmrFAItx7ZEqvV20aJuXxg82+4yIdu4ItABTHjg62kxNM/B1
NLfRnS9h52O+9EILYseP7072OrKLvX8JsSm69iAB5hiP7OuQXnAEWZ+7RAIbPnHO8w/RCRi7a2LJ
Py5S/rGDNgX7r+tfiNGCxQrlAH5aBb8fNhkLs1FrYfIHhLbwNBcbeMAwoPkWqZbfJgMa1NBCot+Y
gdvQ3KTJpztr7ibFDWm/Pp/cbstPcqCFYVNAVGCKUGvXZ0h6VuAmlOaZdrRe9KD3lg9lM1cH114j
QKHf6IqERJNUmvX7K4Xeodr19lNaGrecUxkutyQMwlOLKc0o+qb4ktmILwcdwAErhzwMAF7h9XxH
Neyogfkv2gMg88nVo5yHCCDtpQeAfqPMg95bbcn6M1uQ3YKhJQOOvS7VbQ5e+kWplqF0WITYhiN9
8Rt5WbOFkf85M/obuBw7yI90h2m42RA1CNE50W/kTiQoGQika6jY3riLwu4KHo9RapaNBxwXPkRH
asD1Di+rgHI8lAa6xSy95zjKgRqcd/zWuC6ObahZpXGZX7D+J7z4afKmzYz8j5MsCCzdPJ5Hnp5K
GKUN2qAWHZ7SCliXABdXvS61H+/TZlB0nptnfInepJGRRI9m/L95OrejJXef8/hruEJLwAKvO8aw
DHGDjObmSuHdOpvKedZIXEAl9sxnks7epyza1mNCf5pewpgsQuOK2itgQ4jLqE0t2A78ospO7Kkr
HmdgpvsKTI8c/YHh58ZOQ8el2paYAniGXiEmVGmw36M/ul+FrtuhErXJSTJcsvQRXbsU9xidOT9A
KhSHN8/BHGaJkU61EM3ZYCuY8ZO9BGEQGCy/Sci15C55e0KhyaJRyn1oSTqZGmWC0rT/CUVBtPNX
KW6MxGs6YTyu90lNOBHhlo5UfT/ESIi4jGPzVyHl8C3tN9/edf3cqlV8O0aqpNgVesz+MLB2V68m
Ri3K4YerXsrpidMTo2+l0zVlitQoEAxVw/8Wd86vQ4X0KzvCi9U2hPyBK5BUEIplcOdeTG1fTDD3
hObQql/N1ih4Atns/ix0zSeZOa00ZSOyBCZn0WxYyEXfk5IWtocZqSvuuD0z1QGYI/YPqkaGYx9D
ppOYOLQczseZRJ3avnLs5n6nLv8hiewkYSq09+8AwYIWeKI6bSJYCQKC2nJxR0Xl0ylKtwKLiSQ7
OR7womIlOa4vle/qoX+V+HvqsNXWKjNB9cfBAY9ykMCVd9e1ukCcbcPe0FKrfMPiZrIe1o2tjzWr
51lgq5YwFY6bYScpXuqUFPCerHFkJnpzxymUGxoUK+C0XZSF9/RndhBRLkGZM85afJR+UYFbaxSA
sqHxxJ31BjJa5e6tK6l7ervWAMa3EI/vxoiB2w/RpnVrdBT95cFaB15NpkIzSZT9BPMMfXMJC8Lx
8KQzJEuRmUqxLSHdruO4EMce8TBfqeIq7x40gsUP4gUYXEWLdt4WbH+4qiVePJx9ACyU1APpMPQs
VpjZ5ePLbcVvJNz6lUYUapd6ZryP9+1vpJRPTgSl0QdEryZ4PD7po7zD6N7UhmWd8sLQjDl4qOTF
6ywEuCR7BqPa6gfhZG7cdZPuWD45xhGDbzAx1DkKZlxdq7rrN4Ba1RPahWyeCc3EkhS6d11isduD
sS2KbOglMc9mRp2M85UbdOD06mYvqgIKzUakqHUdCG+BTflC/JWf6pI7QghNzaH1D9LscE+/N4w1
XB10/yltK7hXDTYYTdOutpBK2aPDGihJb2257W+fqUdNvnRzqPr+5sUocELzataQ9I+/k5nLpzN4
mHJ3USJ6oytZtIRuRpwhWde19RhTyqHan5rcYhcZW5kdRPrs8Wu5Y+vCArg1vFcFUgNw9/XbJOUT
Oq71NXVPYPeL703+qoX8L7Po7DGM2A6RzfRNjao/Ac/wZF1t+C9p33FGyJ7AKMMflEKK6C+xViMy
eRswPHKtjSTTu4itwtOn8CSs59qmhoTiH8mjnfX29gKhnqM70S5F7pqPmBtACHoRaH3aTzL05yQ9
3QieNEOLvxhcbEEEJiiXlRFy/sbISDobFWO2FhUPNOxAr31QVDsDCqeAcKtuyw/r96B2kT6ClLDo
tWDnfDKQjNaBBMNiJPOaROS9x9mp5mBdcqQ+MJgdeOEYZYoKDQ9ooN7jVSTYGW1gPiSbUO7Ggc3V
rULJXxn0VpJgZygG9wBVeneKneACuruBiPfjXpjFuc05oZCJgudacDlrDWnUQ8eGxM606V477OZm
KrglDHDCAB8c2d2BOJJ+IUZEOIAr9KMWHCi4/UI+as3ZJP86+3gWKDByYDv83Ya8Wjkol2UvEhQz
OmaaMdsSAZ6Oxe0eUwzsCIvLFmAOyyp7rY1ZRzPAZzn9c03u2aSFlxMOdzTpR7ERwV4XSIZn6jFz
rY9dZwC4qe/FIn6+RvN5tESZHEbTiTidsLnWkgka1khw4bRTX0T7IKGuvIZxNrYtKd31+3b0shko
J/gaWmIIJkGMFcf0OAiqAdneOdytqKPe/3FgmGOqW6jwbw4CdXYg8SRSbhXNSMakmGgNh/guCFtI
e32rs7g7L6IlVj32MJbQBfipM+JTgQblKCUEYvo0HGceF4D0uHgtgjAmIX6RPNaUnpFSBgZBwzhT
dt8Ivgr20BsZcpiGLZVRkGeUhWJC21oSJBxAbpC5Z0yByn2CmRw42NJ+yh22umHWFb0EKVDvSOAH
XXY2I1yRADxgjStESEyrrifN8FOY58WGRD5tU4BXxanZ0ly4Ko+KXoVYXLE2RYkZ0hJWAYX6b0gm
lZPbNSK5qE5Rr4lAQfBdRIWHar11Qhq2giwNvEX3z1/NQxSeJfjy5YK61ZUQeH1i4FXMjhHaZcBE
6vZOHYrxcZ7wicwhGmX9ap8F1eaNTPF7lz3UKjzRc62mELhLyCd+IdXEQoT9dW2yW/Cfqdh5Q6HL
SpmZQLvwiSC06x1iAQDMG8qsVN/BAnSS5GnFPSBVJ2hQOBV76i5hLrBz9CqlewuLP5NeCmjOKCY8
uIBdUhciMzKYJEgwKe9HhwDb4GMV0w8g+l/1rLK6k9rTkIX+lxf9opeVa1HPHn5yuhb9UoG0PklT
RETScLg0GdW5XPDgI4JeY5eHddkWJJJpjJS/PF5pfPoHLgv8aiNkX4IT+RJ43PzBFPdi34I3UKhS
fllSRS4HFRimUcPj222FhciLUz9IHZ8KRCaCe0K95iaV1yhRdKsfq/w9pSMNHplKYb9yeyB1dzX4
9REG5DXtBeMGWW2v8YsWU3Gkfu9vIPxT2qfJPc4IEeQhtf3k6Ew/rsxqkOq7ikLYyOsfEXYbwjVc
VV62VF8Q8TySzLt6NQ14z7mnY4cEMmSm+9fGdqcHQ5R/LplcKP60krZJTc5NyRFEDtiEbGG4PjAG
PcM0JLL1I4n6k0dFZsF/p6nD0tKy5ZAgBXzxMhvzSSJxhKFW5oRnsdlMJ94bMOi/EQ3BuOviOXP3
CQErLblZ7RGgCKY8CFDevkZ7duVMpymLt6CTHQI3CJaTfw8uJ5dijBjBbbQNJ3ybRUYnNCxvo/G6
VuX61roBS+tl711m5oKDHq49yXyS6fj+TLRHH22dcWHFcAPlqk7vNLCJb2pATa1xaLELRLWZ0+P6
Fx+hleyBf3OVgUkdMJEaN4FiNMY/CK4qlVkTY/7EX27DW78z12+j8v+ItRxkBUUtNd2TLggSmJVi
8IYapYLN9bxg3mMBGQcxWsQXTcCT3fbLkWhaj+Oxzvy32mH73o1gROnG9818eu/D+Gm761mvz7FW
T0bmrpW1HFRvQoLvTwxOzxmH7O1EFcWgUNJbrCO3EYT9Z2gc3prS+1BKwXbx4o3uUZ5ZKrmSIfch
3bOHmxGNx46CeY6QsJaOaOGf6cH7NFejOYsgMAVnlAjEGP26aQk6AJKYVPHMMdsLvUXKmusXWAzg
z/lOS+IxV77VRbhEfrytvq67Rbd0qGxefq72k1YdOTQTdWHN1YuQQx3W7CzAXjHAQTdcwHXJiYoF
FpDzgSz6buACGA1az9NuLt+Os64BL8gOij/n2zXXViBHxzsATByfFGyj7CaeuvecSsYC6Z/BcOHf
PMDt3xUOwGBj9vZZ1wsG+hOc/Xm5zSiDGeP3jypd6IbMmSjXeK/FVv3NkJ/QLZZ721XH6CAUysV2
4Z4Opt3MP8D5JKsLzTUaR3SUYSU9mR3K9C2YcwbV56uNoWN1AlKk1Ov4p2ajfCusQN5M80JELuQG
M0WHbHjCmTw4pF8nTQkGwR89zqWPcqAaEUMPNleC9+SDqql9nzieaDmsj9FbvRNkkOpDI7m0uWFc
wT9DXjZ4sY7w9HDI0D2R2GIbXIsJI5bzz84PtWt5hipvPZIg6JZU8AZcbh06rnzkOWWoUXgmMKEG
0bdMtjNqjt99Es7X9qdoTt/9cV8HZDRG7zEqyceMjJXbsVEmD7Hujpr81mnh2GB7HYYQboJOzuc+
z6DpkhUy/a6MMPI6M2UHTKZoBCzEnO0gl9asbohf8f2MJqHIQsAweKlyYL1E7X9DQibUFCC+0bQL
OPeVwJ7g3uaTNNNf4wLVsSIVAiKR6PVt9d0U1SraNOBu0P8SGpehAmgADsaNW8Kq9QSIOiYyIxAh
GYtp38sXeqz9ETkmxNxyjou4XI80K9tKD50YAUNCyGaDAMYZFFMNCi9BV/ScmzbWY2rD0iByjQ5n
zrqrTKkRktlvm4T+lnrT0Liwu10qj+837+bxnzdbd2jddJHxZYRi6wHtWJyXzRdyNKOPvbDfNmqX
eUQmI9fOyxgjSowWpiSN/xNtPM5M9Lhj6if9LGxGm+t6fWsEn0QyRy2CK3A2pxnA8gTKIsI2ulUq
bFFPzNHfe+x/OFELzWiaPv7wTF8Ap9LiLRHHB7f72dgGZQuLIDXxvNN9s3ARSl57g710ntuRDM1Z
jvNKnyPIuv8Uivrlqh9+AlWho1arfUJlgKM+cHJHDu+WwiPCJDTvHWICkw06jk7V7qDzGyyn2uMn
IXbAgekWUSonIfkTHjd0/FcAVorxpz6c46Z8l8y1DJMYgjubFIvc2YAM4Q7iFxUxJH4f8b8=
`pragma protect end_protected

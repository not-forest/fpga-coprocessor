-- coproc_soft_cpu.vhd

-- Generated using ACDS version 24.1 1077

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity coproc_soft_cpu is
	port (
		i_clk_clk                                                    : in    std_logic := '0'; --        i_clk.clk
		i_clr_reset_n                                                : in    std_logic := '0'; --        i_clr.reset_n
		o_dbg_reset_reset                                            : out   std_logic;        --  o_dbg_reset.reset
		o_spi_export_mosi_to_the_spislave_inst_for_spichain          : in    std_logic := '0'; -- o_spi_export.mosi_to_the_spislave_inst_for_spichain
		o_spi_export_nss_to_the_spislave_inst_for_spichain           : in    std_logic := '0'; --             .nss_to_the_spislave_inst_for_spichain
		o_spi_export_miso_to_and_from_the_spislave_inst_for_spichain : inout std_logic := '0'; --             .miso_to_and_from_the_spislave_inst_for_spichain
		o_spi_export_sclk_to_the_spislave_inst_for_spichain          : in    std_logic := '0'  --             .sclk_to_the_spislave_inst_for_spichain
	);
end entity coproc_soft_cpu;

architecture rtl of coproc_soft_cpu is
	component coproc_soft_cpu_CPU is
		port (
			clk                               : in  std_logic                     := 'X';             -- clk
			reset_reset                       : in  std_logic                     := 'X';             -- reset
			platform_irq_rx_irq               : in  std_logic_vector(15 downto 0) := (others => 'X'); -- irq
			ndm_reset_in_reset                : in  std_logic                     := 'X';             -- reset
			timer_sw_agent_address            : in  std_logic_vector(5 downto 0)  := (others => 'X'); -- address
			timer_sw_agent_byteenable         : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			timer_sw_agent_read               : in  std_logic                     := 'X';             -- read
			timer_sw_agent_readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			timer_sw_agent_write              : in  std_logic                     := 'X';             -- write
			timer_sw_agent_writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			timer_sw_agent_waitrequest        : out std_logic;                                        -- waitrequest
			timer_sw_agent_readdatavalid      : out std_logic;                                        -- readdatavalid
			instruction_manager_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			instruction_manager_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			instruction_manager_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			instruction_manager_response      : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			instruction_manager_address       : out std_logic_vector(31 downto 0);                    -- address
			instruction_manager_read          : out std_logic;                                        -- read
			data_manager_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			data_manager_waitrequest          : in  std_logic                     := 'X';             -- waitrequest
			data_manager_readdatavalid        : in  std_logic                     := 'X';             -- readdatavalid
			data_manager_response             : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- response
			data_manager_address              : out std_logic_vector(31 downto 0);                    -- address
			data_manager_read                 : out std_logic;                                        -- read
			data_manager_write                : out std_logic;                                        -- write
			data_manager_writedata            : out std_logic_vector(31 downto 0);                    -- writedata
			data_manager_byteenable           : out std_logic_vector(3 downto 0);                     -- byteenable
			data_manager_writeresponsevalid   : in  std_logic                     := 'X';             -- writeresponsevalid
			dm_agent_address                  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- address
			dm_agent_read                     : in  std_logic                     := 'X';             -- read
			dm_agent_readdata                 : out std_logic_vector(31 downto 0);                    -- readdata
			dm_agent_write                    : in  std_logic                     := 'X';             -- write
			dm_agent_writedata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dm_agent_waitrequest              : out std_logic;                                        -- waitrequest
			dm_agent_readdatavalid            : out std_logic;                                        -- readdatavalid
			dbg_reset_out_reset               : out std_logic                                         -- reset
		);
	end component coproc_soft_cpu_CPU;

	component altera_avalon_jtag_uart is
		generic (
			readBufferDepth            : integer := 64;
			readIRQThreshold           : integer := 8;
			useRegistersForReadBuffer  : boolean := false;
			useRegistersForWriteBuffer : boolean := false;
			writeBufferDepth           : integer := 64;
			writeIRQThreshold          : integer := 8;
			printingMethod             : boolean := false;
			FIFO_WIDTH                 : integer := 8;
			WR_WIDTHU                  : integer := 0;
			RD_WIDTHU                  : integer := 0;
			write_le                   : string  := """ON""";
			read_le                    : string  := """ON""";
			HEX_WRITE_DEPTH_STR        : integer := 64;
			HEX_READ_DEPTH_STR         : integer := 64;
			legacySignalAllow          : boolean := true
		);
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component altera_avalon_jtag_uart;

	component SPISlaveToAvalonMasterBridge is
		port (
			clk                                                                    : in    std_logic                     := 'X';             -- clk
			reset_n                                                                : in    std_logic                     := 'X';             -- reset_n
			mosi_to_the_spislave_inst_for_spichain                                 : in    std_logic                     := 'X';             -- export
			nss_to_the_spislave_inst_for_spichain                                  : in    std_logic                     := 'X';             -- export
			miso_to_and_from_the_spislave_inst_for_spichain                        : inout std_logic                     := 'X';             -- export
			sclk_to_the_spislave_inst_for_spichain                                 : in    std_logic                     := 'X';             -- export
			address_from_the_altera_avalon_packets_to_master_inst_for_spichain     : out   std_logic_vector(31 downto 0);                    -- address
			byteenable_from_the_altera_avalon_packets_to_master_inst_for_spichain  : out   std_logic_vector(3 downto 0);                     -- byteenable
			read_from_the_altera_avalon_packets_to_master_inst_for_spichain        : out   std_logic;                                        -- read
			readdata_to_the_altera_avalon_packets_to_master_inst_for_spichain      : in    std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			readdatavalid_to_the_altera_avalon_packets_to_master_inst_for_spichain : in    std_logic                     := 'X';             -- readdatavalid
			waitrequest_to_the_altera_avalon_packets_to_master_inst_for_spichain   : in    std_logic                     := 'X';             -- waitrequest
			write_from_the_altera_avalon_packets_to_master_inst_for_spichain       : out   std_logic;                                        -- write
			writedata_from_the_altera_avalon_packets_to_master_inst_for_spichain   : out   std_logic_vector(31 downto 0)                     -- writedata
		);
	end component SPISlaveToAvalonMasterBridge;

	component coproc_soft_cpu_SRAM is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(12 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component coproc_soft_cpu_SRAM;

	component coproc_soft_cpu_mm_interconnect_0 is
		port (
			CLK_clk_clk                               : in  std_logic                     := 'X';             -- clk
			SPI_clk_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			CPU_data_manager_address                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			CPU_data_manager_waitrequest              : out std_logic;                                        -- waitrequest
			CPU_data_manager_byteenable               : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			CPU_data_manager_read                     : in  std_logic                     := 'X';             -- read
			CPU_data_manager_readdata                 : out std_logic_vector(31 downto 0);                    -- readdata
			CPU_data_manager_readdatavalid            : out std_logic;                                        -- readdatavalid
			CPU_data_manager_write                    : in  std_logic                     := 'X';             -- write
			CPU_data_manager_writedata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			CPU_data_manager_response                 : out std_logic_vector(1 downto 0);                     -- response
			CPU_data_manager_writeresponsevalid       : out std_logic;                                        -- writeresponsevalid
			CPU_instruction_manager_address           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			CPU_instruction_manager_waitrequest       : out std_logic;                                        -- waitrequest
			CPU_instruction_manager_read              : in  std_logic                     := 'X';             -- read
			CPU_instruction_manager_readdata          : out std_logic_vector(31 downto 0);                    -- readdata
			CPU_instruction_manager_readdatavalid     : out std_logic;                                        -- readdatavalid
			CPU_instruction_manager_response          : out std_logic_vector(1 downto 0);                     -- response
			SPI_avalon_master_address                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			SPI_avalon_master_waitrequest             : out std_logic;                                        -- waitrequest
			SPI_avalon_master_byteenable              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			SPI_avalon_master_read                    : in  std_logic                     := 'X';             -- read
			SPI_avalon_master_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			SPI_avalon_master_readdatavalid           : out std_logic;                                        -- readdatavalid
			SPI_avalon_master_write                   : in  std_logic                     := 'X';             -- write
			SPI_avalon_master_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			CPU_dm_agent_address                      : out std_logic_vector(15 downto 0);                    -- address
			CPU_dm_agent_write                        : out std_logic;                                        -- write
			CPU_dm_agent_read                         : out std_logic;                                        -- read
			CPU_dm_agent_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			CPU_dm_agent_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			CPU_dm_agent_readdatavalid                : in  std_logic                     := 'X';             -- readdatavalid
			CPU_dm_agent_waitrequest                  : in  std_logic                     := 'X';             -- waitrequest
			CPU_timer_sw_agent_address                : out std_logic_vector(5 downto 0);                     -- address
			CPU_timer_sw_agent_write                  : out std_logic;                                        -- write
			CPU_timer_sw_agent_read                   : out std_logic;                                        -- read
			CPU_timer_sw_agent_readdata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			CPU_timer_sw_agent_writedata              : out std_logic_vector(31 downto 0);                    -- writedata
			CPU_timer_sw_agent_byteenable             : out std_logic_vector(3 downto 0);                     -- byteenable
			CPU_timer_sw_agent_readdatavalid          : in  std_logic                     := 'X';             -- readdatavalid
			CPU_timer_sw_agent_waitrequest            : in  std_logic                     := 'X';             -- waitrequest
			DEBUG_JTAG_avalon_jtag_slave_address      : out std_logic_vector(0 downto 0);                     -- address
			DEBUG_JTAG_avalon_jtag_slave_write        : out std_logic;                                        -- write
			DEBUG_JTAG_avalon_jtag_slave_read         : out std_logic;                                        -- read
			DEBUG_JTAG_avalon_jtag_slave_readdata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			DEBUG_JTAG_avalon_jtag_slave_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			DEBUG_JTAG_avalon_jtag_slave_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			DEBUG_JTAG_avalon_jtag_slave_chipselect   : out std_logic;                                        -- chipselect
			SRAM_s1_address                           : out std_logic_vector(12 downto 0);                    -- address
			SRAM_s1_write                             : out std_logic;                                        -- write
			SRAM_s1_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			SRAM_s1_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			SRAM_s1_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			SRAM_s1_chipselect                        : out std_logic;                                        -- chipselect
			SRAM_s1_clken                             : out std_logic                                         -- clken
		);
	end component coproc_soft_cpu_mm_interconnect_0;

	component coproc_soft_cpu_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(15 downto 0)         -- irq
		);
	end component coproc_soft_cpu_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal spi_avalon_master_readdata                                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:SPI_avalon_master_readdata -> SPI:readdata_to_the_altera_avalon_packets_to_master_inst_for_spichain
	signal spi_avalon_master_waitrequest                                  : std_logic;                     -- mm_interconnect_0:SPI_avalon_master_waitrequest -> SPI:waitrequest_to_the_altera_avalon_packets_to_master_inst_for_spichain
	signal spi_avalon_master_address                                      : std_logic_vector(31 downto 0); -- SPI:address_from_the_altera_avalon_packets_to_master_inst_for_spichain -> mm_interconnect_0:SPI_avalon_master_address
	signal spi_avalon_master_byteenable                                   : std_logic_vector(3 downto 0);  -- SPI:byteenable_from_the_altera_avalon_packets_to_master_inst_for_spichain -> mm_interconnect_0:SPI_avalon_master_byteenable
	signal spi_avalon_master_read                                         : std_logic;                     -- SPI:read_from_the_altera_avalon_packets_to_master_inst_for_spichain -> mm_interconnect_0:SPI_avalon_master_read
	signal spi_avalon_master_readdatavalid                                : std_logic;                     -- mm_interconnect_0:SPI_avalon_master_readdatavalid -> SPI:readdatavalid_to_the_altera_avalon_packets_to_master_inst_for_spichain
	signal spi_avalon_master_write                                        : std_logic;                     -- SPI:write_from_the_altera_avalon_packets_to_master_inst_for_spichain -> mm_interconnect_0:SPI_avalon_master_write
	signal spi_avalon_master_writedata                                    : std_logic_vector(31 downto 0); -- SPI:writedata_from_the_altera_avalon_packets_to_master_inst_for_spichain -> mm_interconnect_0:SPI_avalon_master_writedata
	signal cpu_data_manager_readdata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_data_manager_readdata -> CPU:data_manager_readdata
	signal cpu_data_manager_waitrequest                                   : std_logic;                     -- mm_interconnect_0:CPU_data_manager_waitrequest -> CPU:data_manager_waitrequest
	signal cpu_data_manager_address                                       : std_logic_vector(31 downto 0); -- CPU:data_manager_address -> mm_interconnect_0:CPU_data_manager_address
	signal cpu_data_manager_read                                          : std_logic;                     -- CPU:data_manager_read -> mm_interconnect_0:CPU_data_manager_read
	signal cpu_data_manager_byteenable                                    : std_logic_vector(3 downto 0);  -- CPU:data_manager_byteenable -> mm_interconnect_0:CPU_data_manager_byteenable
	signal cpu_data_manager_readdatavalid                                 : std_logic;                     -- mm_interconnect_0:CPU_data_manager_readdatavalid -> CPU:data_manager_readdatavalid
	signal cpu_data_manager_response                                      : std_logic_vector(1 downto 0);  -- mm_interconnect_0:CPU_data_manager_response -> CPU:data_manager_response
	signal cpu_data_manager_write                                         : std_logic;                     -- CPU:data_manager_write -> mm_interconnect_0:CPU_data_manager_write
	signal cpu_data_manager_writedata                                     : std_logic_vector(31 downto 0); -- CPU:data_manager_writedata -> mm_interconnect_0:CPU_data_manager_writedata
	signal cpu_data_manager_writeresponsevalid                            : std_logic;                     -- mm_interconnect_0:CPU_data_manager_writeresponsevalid -> CPU:data_manager_writeresponsevalid
	signal cpu_instruction_manager_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_instruction_manager_readdata -> CPU:instruction_manager_readdata
	signal cpu_instruction_manager_waitrequest                            : std_logic;                     -- mm_interconnect_0:CPU_instruction_manager_waitrequest -> CPU:instruction_manager_waitrequest
	signal cpu_instruction_manager_address                                : std_logic_vector(31 downto 0); -- CPU:instruction_manager_address -> mm_interconnect_0:CPU_instruction_manager_address
	signal cpu_instruction_manager_read                                   : std_logic;                     -- CPU:instruction_manager_read -> mm_interconnect_0:CPU_instruction_manager_read
	signal cpu_instruction_manager_readdatavalid                          : std_logic;                     -- mm_interconnect_0:CPU_instruction_manager_readdatavalid -> CPU:instruction_manager_readdatavalid
	signal cpu_instruction_manager_response                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:CPU_instruction_manager_response -> CPU:instruction_manager_response
	signal mm_interconnect_0_sram_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:SRAM_s1_chipselect -> SRAM:chipselect
	signal mm_interconnect_0_sram_s1_readdata                             : std_logic_vector(31 downto 0); -- SRAM:readdata -> mm_interconnect_0:SRAM_s1_readdata
	signal mm_interconnect_0_sram_s1_address                              : std_logic_vector(12 downto 0); -- mm_interconnect_0:SRAM_s1_address -> SRAM:address
	signal mm_interconnect_0_sram_s1_byteenable                           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:SRAM_s1_byteenable -> SRAM:byteenable
	signal mm_interconnect_0_sram_s1_write                                : std_logic;                     -- mm_interconnect_0:SRAM_s1_write -> SRAM:write
	signal mm_interconnect_0_sram_s1_writedata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:SRAM_s1_writedata -> SRAM:writedata
	signal mm_interconnect_0_sram_s1_clken                                : std_logic;                     -- mm_interconnect_0:SRAM_s1_clken -> SRAM:clken
	signal mm_interconnect_0_cpu_dm_agent_readdata                        : std_logic_vector(31 downto 0); -- CPU:dm_agent_readdata -> mm_interconnect_0:CPU_dm_agent_readdata
	signal mm_interconnect_0_cpu_dm_agent_waitrequest                     : std_logic;                     -- CPU:dm_agent_waitrequest -> mm_interconnect_0:CPU_dm_agent_waitrequest
	signal mm_interconnect_0_cpu_dm_agent_address                         : std_logic_vector(15 downto 0); -- mm_interconnect_0:CPU_dm_agent_address -> CPU:dm_agent_address
	signal mm_interconnect_0_cpu_dm_agent_read                            : std_logic;                     -- mm_interconnect_0:CPU_dm_agent_read -> CPU:dm_agent_read
	signal mm_interconnect_0_cpu_dm_agent_readdatavalid                   : std_logic;                     -- CPU:dm_agent_readdatavalid -> mm_interconnect_0:CPU_dm_agent_readdatavalid
	signal mm_interconnect_0_cpu_dm_agent_write                           : std_logic;                     -- mm_interconnect_0:CPU_dm_agent_write -> CPU:dm_agent_write
	signal mm_interconnect_0_cpu_dm_agent_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_dm_agent_writedata -> CPU:dm_agent_writedata
	signal mm_interconnect_0_debug_jtag_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:DEBUG_JTAG_avalon_jtag_slave_chipselect -> DEBUG_JTAG:av_chipselect
	signal mm_interconnect_0_debug_jtag_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- DEBUG_JTAG:av_readdata -> mm_interconnect_0:DEBUG_JTAG_avalon_jtag_slave_readdata
	signal mm_interconnect_0_debug_jtag_avalon_jtag_slave_waitrequest     : std_logic;                     -- DEBUG_JTAG:av_waitrequest -> mm_interconnect_0:DEBUG_JTAG_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_debug_jtag_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:DEBUG_JTAG_avalon_jtag_slave_address -> DEBUG_JTAG:av_address
	signal mm_interconnect_0_debug_jtag_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:DEBUG_JTAG_avalon_jtag_slave_read -> mm_interconnect_0_debug_jtag_avalon_jtag_slave_read:in
	signal mm_interconnect_0_debug_jtag_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:DEBUG_JTAG_avalon_jtag_slave_write -> mm_interconnect_0_debug_jtag_avalon_jtag_slave_write:in
	signal mm_interconnect_0_debug_jtag_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:DEBUG_JTAG_avalon_jtag_slave_writedata -> DEBUG_JTAG:av_writedata
	signal mm_interconnect_0_cpu_timer_sw_agent_readdata                  : std_logic_vector(31 downto 0); -- CPU:timer_sw_agent_readdata -> mm_interconnect_0:CPU_timer_sw_agent_readdata
	signal mm_interconnect_0_cpu_timer_sw_agent_waitrequest               : std_logic;                     -- CPU:timer_sw_agent_waitrequest -> mm_interconnect_0:CPU_timer_sw_agent_waitrequest
	signal mm_interconnect_0_cpu_timer_sw_agent_address                   : std_logic_vector(5 downto 0);  -- mm_interconnect_0:CPU_timer_sw_agent_address -> CPU:timer_sw_agent_address
	signal mm_interconnect_0_cpu_timer_sw_agent_read                      : std_logic;                     -- mm_interconnect_0:CPU_timer_sw_agent_read -> CPU:timer_sw_agent_read
	signal mm_interconnect_0_cpu_timer_sw_agent_byteenable                : std_logic_vector(3 downto 0);  -- mm_interconnect_0:CPU_timer_sw_agent_byteenable -> CPU:timer_sw_agent_byteenable
	signal mm_interconnect_0_cpu_timer_sw_agent_readdatavalid             : std_logic;                     -- CPU:timer_sw_agent_readdatavalid -> mm_interconnect_0:CPU_timer_sw_agent_readdatavalid
	signal mm_interconnect_0_cpu_timer_sw_agent_write                     : std_logic;                     -- mm_interconnect_0:CPU_timer_sw_agent_write -> CPU:timer_sw_agent_write
	signal mm_interconnect_0_cpu_timer_sw_agent_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_timer_sw_agent_writedata -> CPU:timer_sw_agent_writedata
	signal irq_mapper_receiver0_irq                                       : std_logic;                     -- DEBUG_JTAG:av_irq -> irq_mapper:receiver0_irq
	signal cpu_platform_irq_rx_irq                                        : std_logic_vector(15 downto 0); -- irq_mapper:sender_irq -> CPU:platform_irq_rx_irq
	signal rst_controller_reset_out_reset                                 : std_logic;                     -- rst_controller:reset_out -> [CPU:ndm_reset_in_reset, CPU:reset_reset, SRAM:reset, irq_mapper:reset, mm_interconnect_0:SPI_clk_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                             : std_logic;                     -- rst_controller:reset_req -> [SRAM:reset_req, rst_translator:reset_req_in]
	signal i_clr_reset_n_ports_inv                                        : std_logic;                     -- i_clr_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_debug_jtag_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_debug_jtag_avalon_jtag_slave_read:inv -> DEBUG_JTAG:av_read_n
	signal mm_interconnect_0_debug_jtag_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_debug_jtag_avalon_jtag_slave_write:inv -> DEBUG_JTAG:av_write_n
	signal rst_controller_reset_out_reset_ports_inv                       : std_logic;                     -- rst_controller_reset_out_reset:inv -> [DEBUG_JTAG:rst_n, SPI:reset_n]

begin

	cpu : component coproc_soft_cpu_CPU
		port map (
			clk                               => i_clk_clk,                                          --                 clk.clk
			reset_reset                       => rst_controller_reset_out_reset,                     --               reset.reset
			platform_irq_rx_irq               => cpu_platform_irq_rx_irq,                            --     platform_irq_rx.irq
			ndm_reset_in_reset                => rst_controller_reset_out_reset,                     --        ndm_reset_in.reset
			timer_sw_agent_address            => mm_interconnect_0_cpu_timer_sw_agent_address,       --      timer_sw_agent.address
			timer_sw_agent_byteenable         => mm_interconnect_0_cpu_timer_sw_agent_byteenable,    --                    .byteenable
			timer_sw_agent_read               => mm_interconnect_0_cpu_timer_sw_agent_read,          --                    .read
			timer_sw_agent_readdata           => mm_interconnect_0_cpu_timer_sw_agent_readdata,      --                    .readdata
			timer_sw_agent_write              => mm_interconnect_0_cpu_timer_sw_agent_write,         --                    .write
			timer_sw_agent_writedata          => mm_interconnect_0_cpu_timer_sw_agent_writedata,     --                    .writedata
			timer_sw_agent_waitrequest        => mm_interconnect_0_cpu_timer_sw_agent_waitrequest,   --                    .waitrequest
			timer_sw_agent_readdatavalid      => mm_interconnect_0_cpu_timer_sw_agent_readdatavalid, --                    .readdatavalid
			instruction_manager_readdata      => cpu_instruction_manager_readdata,                   -- instruction_manager.readdata
			instruction_manager_waitrequest   => cpu_instruction_manager_waitrequest,                --                    .waitrequest
			instruction_manager_readdatavalid => cpu_instruction_manager_readdatavalid,              --                    .readdatavalid
			instruction_manager_response      => cpu_instruction_manager_response,                   --                    .response
			instruction_manager_address       => cpu_instruction_manager_address,                    --                    .address
			instruction_manager_read          => cpu_instruction_manager_read,                       --                    .read
			data_manager_readdata             => cpu_data_manager_readdata,                          --        data_manager.readdata
			data_manager_waitrequest          => cpu_data_manager_waitrequest,                       --                    .waitrequest
			data_manager_readdatavalid        => cpu_data_manager_readdatavalid,                     --                    .readdatavalid
			data_manager_response             => cpu_data_manager_response,                          --                    .response
			data_manager_address              => cpu_data_manager_address,                           --                    .address
			data_manager_read                 => cpu_data_manager_read,                              --                    .read
			data_manager_write                => cpu_data_manager_write,                             --                    .write
			data_manager_writedata            => cpu_data_manager_writedata,                         --                    .writedata
			data_manager_byteenable           => cpu_data_manager_byteenable,                        --                    .byteenable
			data_manager_writeresponsevalid   => cpu_data_manager_writeresponsevalid,                --                    .writeresponsevalid
			dm_agent_address                  => mm_interconnect_0_cpu_dm_agent_address,             --            dm_agent.address
			dm_agent_read                     => mm_interconnect_0_cpu_dm_agent_read,                --                    .read
			dm_agent_readdata                 => mm_interconnect_0_cpu_dm_agent_readdata,            --                    .readdata
			dm_agent_write                    => mm_interconnect_0_cpu_dm_agent_write,               --                    .write
			dm_agent_writedata                => mm_interconnect_0_cpu_dm_agent_writedata,           --                    .writedata
			dm_agent_waitrequest              => mm_interconnect_0_cpu_dm_agent_waitrequest,         --                    .waitrequest
			dm_agent_readdatavalid            => mm_interconnect_0_cpu_dm_agent_readdatavalid,       --                    .readdatavalid
			dbg_reset_out_reset               => o_dbg_reset_reset                                   --       dbg_reset_out.reset
		);

	debug_jtag : component altera_avalon_jtag_uart
		generic map (
			readBufferDepth            => 64,
			readIRQThreshold           => 8,
			useRegistersForReadBuffer  => false,
			useRegistersForWriteBuffer => false,
			writeBufferDepth           => 64,
			writeIRQThreshold          => 8,
			printingMethod             => false,
			FIFO_WIDTH                 => 8,
			WR_WIDTHU                  => 6,
			RD_WIDTHU                  => 6,
			write_le                   => "ON",
			read_le                    => "ON",
			HEX_WRITE_DEPTH_STR        => 64,
			HEX_READ_DEPTH_STR         => 64,
			legacySignalAllow          => false
		)
		port map (
			clk            => i_clk_clk,                                                      --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                       --             reset.reset_n
			av_chipselect  => mm_interconnect_0_debug_jtag_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_debug_jtag_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_debug_jtag_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_debug_jtag_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_debug_jtag_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_debug_jtag_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_debug_jtag_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                        --               irq.irq
		);

	spi : component SPISlaveToAvalonMasterBridge
		port map (
			clk                                                                    => i_clk_clk,                                                    --           clk.clk
			reset_n                                                                => rst_controller_reset_out_reset_ports_inv,                     --     clk_reset.reset_n
			mosi_to_the_spislave_inst_for_spichain                                 => o_spi_export_mosi_to_the_spislave_inst_for_spichain,          --      export_0.export
			nss_to_the_spislave_inst_for_spichain                                  => o_spi_export_nss_to_the_spislave_inst_for_spichain,           --              .export
			miso_to_and_from_the_spislave_inst_for_spichain                        => o_spi_export_miso_to_and_from_the_spislave_inst_for_spichain, --              .export
			sclk_to_the_spislave_inst_for_spichain                                 => o_spi_export_sclk_to_the_spislave_inst_for_spichain,          --              .export
			address_from_the_altera_avalon_packets_to_master_inst_for_spichain     => spi_avalon_master_address,                                    -- avalon_master.address
			byteenable_from_the_altera_avalon_packets_to_master_inst_for_spichain  => spi_avalon_master_byteenable,                                 --              .byteenable
			read_from_the_altera_avalon_packets_to_master_inst_for_spichain        => spi_avalon_master_read,                                       --              .read
			readdata_to_the_altera_avalon_packets_to_master_inst_for_spichain      => spi_avalon_master_readdata,                                   --              .readdata
			readdatavalid_to_the_altera_avalon_packets_to_master_inst_for_spichain => spi_avalon_master_readdatavalid,                              --              .readdatavalid
			waitrequest_to_the_altera_avalon_packets_to_master_inst_for_spichain   => spi_avalon_master_waitrequest,                                --              .waitrequest
			write_from_the_altera_avalon_packets_to_master_inst_for_spichain       => spi_avalon_master_write,                                      --              .write
			writedata_from_the_altera_avalon_packets_to_master_inst_for_spichain   => spi_avalon_master_writedata                                   --              .writedata
		);

	sram : component coproc_soft_cpu_SRAM
		port map (
			clk        => i_clk_clk,                            --   clk1.clk
			address    => mm_interconnect_0_sram_s1_address,    --     s1.address
			clken      => mm_interconnect_0_sram_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_sram_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_sram_s1_write,      --       .write
			readdata   => mm_interconnect_0_sram_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_sram_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_sram_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,       -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,   --       .reset_req
			freeze     => '0'                                   -- (terminated)
		);

	mm_interconnect_0 : component coproc_soft_cpu_mm_interconnect_0
		port map (
			CLK_clk_clk                               => i_clk_clk,                                                  --                             CLK_clk.clk
			SPI_clk_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                             -- SPI_clk_reset_reset_bridge_in_reset.reset
			CPU_data_manager_address                  => cpu_data_manager_address,                                   --                    CPU_data_manager.address
			CPU_data_manager_waitrequest              => cpu_data_manager_waitrequest,                               --                                    .waitrequest
			CPU_data_manager_byteenable               => cpu_data_manager_byteenable,                                --                                    .byteenable
			CPU_data_manager_read                     => cpu_data_manager_read,                                      --                                    .read
			CPU_data_manager_readdata                 => cpu_data_manager_readdata,                                  --                                    .readdata
			CPU_data_manager_readdatavalid            => cpu_data_manager_readdatavalid,                             --                                    .readdatavalid
			CPU_data_manager_write                    => cpu_data_manager_write,                                     --                                    .write
			CPU_data_manager_writedata                => cpu_data_manager_writedata,                                 --                                    .writedata
			CPU_data_manager_response                 => cpu_data_manager_response,                                  --                                    .response
			CPU_data_manager_writeresponsevalid       => cpu_data_manager_writeresponsevalid,                        --                                    .writeresponsevalid
			CPU_instruction_manager_address           => cpu_instruction_manager_address,                            --             CPU_instruction_manager.address
			CPU_instruction_manager_waitrequest       => cpu_instruction_manager_waitrequest,                        --                                    .waitrequest
			CPU_instruction_manager_read              => cpu_instruction_manager_read,                               --                                    .read
			CPU_instruction_manager_readdata          => cpu_instruction_manager_readdata,                           --                                    .readdata
			CPU_instruction_manager_readdatavalid     => cpu_instruction_manager_readdatavalid,                      --                                    .readdatavalid
			CPU_instruction_manager_response          => cpu_instruction_manager_response,                           --                                    .response
			SPI_avalon_master_address                 => spi_avalon_master_address,                                  --                   SPI_avalon_master.address
			SPI_avalon_master_waitrequest             => spi_avalon_master_waitrequest,                              --                                    .waitrequest
			SPI_avalon_master_byteenable              => spi_avalon_master_byteenable,                               --                                    .byteenable
			SPI_avalon_master_read                    => spi_avalon_master_read,                                     --                                    .read
			SPI_avalon_master_readdata                => spi_avalon_master_readdata,                                 --                                    .readdata
			SPI_avalon_master_readdatavalid           => spi_avalon_master_readdatavalid,                            --                                    .readdatavalid
			SPI_avalon_master_write                   => spi_avalon_master_write,                                    --                                    .write
			SPI_avalon_master_writedata               => spi_avalon_master_writedata,                                --                                    .writedata
			CPU_dm_agent_address                      => mm_interconnect_0_cpu_dm_agent_address,                     --                        CPU_dm_agent.address
			CPU_dm_agent_write                        => mm_interconnect_0_cpu_dm_agent_write,                       --                                    .write
			CPU_dm_agent_read                         => mm_interconnect_0_cpu_dm_agent_read,                        --                                    .read
			CPU_dm_agent_readdata                     => mm_interconnect_0_cpu_dm_agent_readdata,                    --                                    .readdata
			CPU_dm_agent_writedata                    => mm_interconnect_0_cpu_dm_agent_writedata,                   --                                    .writedata
			CPU_dm_agent_readdatavalid                => mm_interconnect_0_cpu_dm_agent_readdatavalid,               --                                    .readdatavalid
			CPU_dm_agent_waitrequest                  => mm_interconnect_0_cpu_dm_agent_waitrequest,                 --                                    .waitrequest
			CPU_timer_sw_agent_address                => mm_interconnect_0_cpu_timer_sw_agent_address,               --                  CPU_timer_sw_agent.address
			CPU_timer_sw_agent_write                  => mm_interconnect_0_cpu_timer_sw_agent_write,                 --                                    .write
			CPU_timer_sw_agent_read                   => mm_interconnect_0_cpu_timer_sw_agent_read,                  --                                    .read
			CPU_timer_sw_agent_readdata               => mm_interconnect_0_cpu_timer_sw_agent_readdata,              --                                    .readdata
			CPU_timer_sw_agent_writedata              => mm_interconnect_0_cpu_timer_sw_agent_writedata,             --                                    .writedata
			CPU_timer_sw_agent_byteenable             => mm_interconnect_0_cpu_timer_sw_agent_byteenable,            --                                    .byteenable
			CPU_timer_sw_agent_readdatavalid          => mm_interconnect_0_cpu_timer_sw_agent_readdatavalid,         --                                    .readdatavalid
			CPU_timer_sw_agent_waitrequest            => mm_interconnect_0_cpu_timer_sw_agent_waitrequest,           --                                    .waitrequest
			DEBUG_JTAG_avalon_jtag_slave_address      => mm_interconnect_0_debug_jtag_avalon_jtag_slave_address,     --        DEBUG_JTAG_avalon_jtag_slave.address
			DEBUG_JTAG_avalon_jtag_slave_write        => mm_interconnect_0_debug_jtag_avalon_jtag_slave_write,       --                                    .write
			DEBUG_JTAG_avalon_jtag_slave_read         => mm_interconnect_0_debug_jtag_avalon_jtag_slave_read,        --                                    .read
			DEBUG_JTAG_avalon_jtag_slave_readdata     => mm_interconnect_0_debug_jtag_avalon_jtag_slave_readdata,    --                                    .readdata
			DEBUG_JTAG_avalon_jtag_slave_writedata    => mm_interconnect_0_debug_jtag_avalon_jtag_slave_writedata,   --                                    .writedata
			DEBUG_JTAG_avalon_jtag_slave_waitrequest  => mm_interconnect_0_debug_jtag_avalon_jtag_slave_waitrequest, --                                    .waitrequest
			DEBUG_JTAG_avalon_jtag_slave_chipselect   => mm_interconnect_0_debug_jtag_avalon_jtag_slave_chipselect,  --                                    .chipselect
			SRAM_s1_address                           => mm_interconnect_0_sram_s1_address,                          --                             SRAM_s1.address
			SRAM_s1_write                             => mm_interconnect_0_sram_s1_write,                            --                                    .write
			SRAM_s1_readdata                          => mm_interconnect_0_sram_s1_readdata,                         --                                    .readdata
			SRAM_s1_writedata                         => mm_interconnect_0_sram_s1_writedata,                        --                                    .writedata
			SRAM_s1_byteenable                        => mm_interconnect_0_sram_s1_byteenable,                       --                                    .byteenable
			SRAM_s1_chipselect                        => mm_interconnect_0_sram_s1_chipselect,                       --                                    .chipselect
			SRAM_s1_clken                             => mm_interconnect_0_sram_s1_clken                             --                                    .clken
		);

	irq_mapper : component coproc_soft_cpu_irq_mapper
		port map (
			clk           => i_clk_clk,                      --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			sender_irq    => cpu_platform_irq_rx_irq         --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => i_clr_reset_n_ports_inv,            -- reset_in0.reset
			clk            => i_clk_clk,                          --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	i_clr_reset_n_ports_inv <= not i_clr_reset_n;

	mm_interconnect_0_debug_jtag_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_debug_jtag_avalon_jtag_slave_read;

	mm_interconnect_0_debug_jtag_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_debug_jtag_avalon_jtag_slave_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of coproc_soft_cpu

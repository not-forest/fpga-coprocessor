`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Q65PmUsbrFI207RC7M5ELo63LI+SOX2SIwDeyzUW5h/KGfVSdhTVXAyhQwBWMwAM
dbuVUTdom4PsB0SFaJfxpW3hYYdElBo2ghFvxRgyfCc1jaMtOkTNdy+19g0yB98j
LbwoaucknpuNSYzlW0QykWTBIFkTx9aqrX2gTk6lTBo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 15536)
j+QbVtKO00fhNHLGKVWTzxmCdChZcHusUz8mbpJR9GHrXClhxUft5at1C+KGS2Ag
bK9A4abjBDsrDysqytCy3KqYszMb2QaOeazCGReybmSw/HESOFI3ToFEG8rmgvQ5
OZQ6E3KCitu3lvYkvHYI9hJbYDjflhYNlG3p9g/o3pY0IOxOPbX1eP7osVVRAleM
aSOCD+h2VfxLZn68AOItRPwvHJa2jutg/8qNnM8InkY0Ayrr//DRQuIyBue/YvUL
ci8nBYsmJfBCFPNSuI71iLcl7EkFQRM2oloE7vciBrS5URefTcLvvIfDPwzemAkk
XfQIxEXruOD3Bpthoydza/ryVvSC3DbdPs/j9NsVi2aSiJhQE9nqJrJPcsOFMKpV
5S59QX1MveIcJoeIZlug+6/+cagzcU9iYxKn8jLOq8XSiJbVvzme+LbWPCpLUjD9
gHH93fsPa6nb7k0PyND5zGd+L75HNc8NV+5J0OlQ7CRjAgLq9LtJKh+OpIuybWUv
Ql2O3E9X1Sxql3jo5MDmylS6AOwFTjZPM4EmobgJMFeoBGq+EUfwDD7e+qj4JE1d
GdtmmMhvhdgW7XZAqq22mMiMKD9x63C5904apcDjfYS6MGr1uNevlkDiLrnaY71e
sk+6bl2Ny21PkRRRl0k7dHVKDbmgtMIM+RVvHWb8YBtTKl4Ti8aK/ZF8OIsrSZju
mjZ2ExmCSRjID8GxvBs5DhMjfPc+0VXPYRZ2IfJ0i/p9gCV6DGM8wNUE7ftcWJRI
W0Tkic6Ip1koQYCiL0XY7pszn4osx3RK/U7RGit9ksgf/MTQEg9vqtBfZAWvQYo1
V9wHy4407FAql00JD5JLA/P4XzH8yTup3i67WaRQh2KDmCl4jVPuYOLBBpiiIsez
M0hURdx+zokYS9kvXCDiV9ZKT51iFGKWU/ts0vb49CbNzq9tQZdDSgxf7P6M9hbe
8hbbbA81nRk7WedNRAoW93mSWM0W5MK7elSJHhYcG1nbvhsbS90WXTI8QfRsNdBq
kJYrSWCtzNe3uLczwFNU+jLAKyU7Q9JM1Z2j11bm8asazEvBP3/s4l0C/lz9uqdk
FWEGhheb5+TekXTfj7z+2NqRQKVkbyH8tDxXqQJajWNdbFU189eC9UzWYsBIdo0S
74Da5/gygxpUJKxTNmN8gThtK7ABa+83Uqn+wdXBEsAiKbUF4ywezTFyxXA3Dzqz
gLS1/sJSkkl7NLFNyKJOUdbj7QwoPVuYBsIFI8M0ljvKvCgrMXxvzRgL411IjBeJ
gKGCO2eUfo974kFzwya6z+V7UVBkxCKD8Xyi1zRsDIzX4me4ov2VKiHbcf5oJb05
B+Q1blqngIZUVLQ1EjXGLlhFyyJVjE/RcU+vHMu8sExa4VowBcSxt8h3UNY1Gcrx
nmK0NYCHLcJNAfpqQAR9o9E/lC0EF+CyY++tErieuoZcXH3hH6EgwEXVNH0rC4Xb
EWacXkmyhX5AWGFI3DXNC4H8JHNOM9xpJ0FNEtv9vckuafMsGCE/sWGNEbl+F9fD
82cDhA9PpHXEb09lIS6UnoSF+djsQmei7P9x57XlfakvEZyP1Nba9Jw/P4B1TeNZ
JXDcMX2avpyy8jKxLwTfEk14svtOBnwi4SE5S8hwaOuAHv2fA/V1UjAdsl2lNrVw
G8b+MjCnDk0HrqPUT0bDsABg3WhlbzNx7DZL0+0WpD8BiFuIkSwMV4DAoy1t+f84
t3YuF/GZRgrcvjzs8I8YRVktBeiWia/j9pl9y/Z3JRYkkbFG7EggJE8RVWI6NRST
e9PHab2TeZ0jzltOTI/Dm5C8dq4R3DfMcK4wb9Oz3zKaVV/g70H1LlQ5JRHg0ciX
7Wo5RXmAHcpyN2wohYPgunHfST5HQnhSbDAGF5T2WrgebA3EdeW7wDHTH2ah1a0t
nTmWowcIjpar/qMB/vb2C7N7zud8DfmGOhuY6iocQsGa9knKq21eJSg0X8KPhPDh
9jkUy+eRGliCCXZbTpfAT6OXN8aMrdQs5cgA5WK0v1DEXXiqh/M9HXPVAcZHHZN9
Jwhj/jfqCF82oyMkJ3zkx/w+/XXedSCcSCj0mlhnUhmuR5SDpDj7BDK+cFeS2yNe
ivqF/Jbog7LmpfBqqefqna/nLv3Z/qpMbXgiubn1ubGy9vz9xPjx1AwWKBe2Unrh
VwARGRjx5bXZwy7XOCi0XsM48UZ0joEX1j+CTIGuKaeCsV0D4vocFkEghFqmo80J
dkg0Tc/RR4hX4/XzRVtljpsaXCeAZ15y1ygph9Ua1Vev6U8Rz0eUNeiXjqbyPXqW
sPzSztiUltFnSqEWkYrvqA7iUnnsjGSp4w5yTOuZR8Rjmd1uF7eGFaXlBoLMs4Hz
dAcP1vcC3EFkuRGiirR+LpQikuJAXqzGFmB4ckQ5gkiDaDbciESmekyqb7/hjXQz
unpq7XPVKhEk70FWi5NPZdDVseuQqXrcQwe1VwC3Yh1Su8VF+0h8/EORsfimLApT
lTdSAKa+cO1ISVApOL+U/RaW3OPEobIXBosSbDQQUYUpMukAHjP2jC082SStOH/y
V8Qo2R25Yxgzon+81hqIIsqbS4XftEf6pcDEtXUmYuQR5NxKs48i4BBa2MgfKjUP
ONCMxE+d73jA8oTVTDfcK64V17jRlsjmMtOs8yf/iHVJE69eUeT4MTYvbyxp0x39
4cFDioh0aOwLUHMtaVeKgdlo21HMjIrDgKEcQ7RVVCDhUmlQxUqIrBLg3+lLPN9U
seqn1RQ6xlM69bvNZqaRv0SSziL98pmHpZDNwZD8K2EaeQhGFwkzVYWMrIQMJW1n
p8/OEvhBvSMogvEKr481hB26A8GHp3q9HyWEEvLbiXDO05wJsAScv/Qx2xb2BEO1
knWGOCOhI7JKtTPgTC1QKPEyGyn2ZBSQCSKQsILakvhmMa4xnVrd7pmW8ZyFmJXk
3QSmk/viTAS28kpH3Nv9Hi3PdRP6eUOO4z4DpPeXtij/MiUsnUHxaVcOMALlJplS
X2eSe0cJqMp9aEIYaqAstY0XPEAsqV8CrYymCtqqPANSm7i7wHChASN+y34GTmM7
RZOllYdL+AZewExdzhQAKg6KRiLRPv+1grCrnke6Rjxj0l8mo2LusxMaP1xoOgGr
XF0D5lipb9uJEsfnoXbeho/vnTqp/9M+iINUOW3QvUuGzX8JeUfDGh9aaXE2yTrF
loyhECRczxxJpokPxaCFwuQyPO2c1W08FICUszcIf14ZjJpZN0gG8zkCj0fshY4y
X0ZW0J2Io8LgwZr9KtcMq3YgLHgDp1H1jNeESpghWkW3WhXAdpUsfpcfOXsoqMxR
ALvPRivY0pUhQOQLgrCtb4n16UOR7Fs/vHXMBWjkCYAZ/Qgk1v/MLw37WE8w0KfF
JAf6dMbJ82uh+4AIncGtieZpy4f25K84/qdmFR8GUYV9jW35W0ExmkXCyE1YQ6y3
XZIzeO6Gk+rxUJQuWXHrl4R/Jj9QyYw/WsOdOlHw/KIvpmWt7q0tUnZu1MkiNE7K
JrUeRhiQ/lWX5vw+8BD6ucmeo7qaS6OVQ9bw68dJ6SGxW3izROHc4v6spms2NU04
c1UYi7xRm/Zer8LGvBRN4f+nG6arHFq5AcR8z4c/K2+9g+VlEIHMgpsuYVNWwUM0
WthZWI3eJGjna7whV92QAIPWbXj1Aqg1R90Jq0SWmZRj7g5zsZYRBOenNn1SaegY
T7IAhpiLn9A84oaEnTx3HkEKPh2aklo1kgc+CAvlsGsBmWDR+AneAbXkmA1uuxFC
BRJiP22bA+3QMVcp1QfJBeIYopOUhAF+z/ZXLuuRtttNwJwRnmLzgufZNUtWxG16
uEXP/oh5apigRY8mWWRciT8DQe0qpfOmSE/qF+kudKXoYbmAgMuJPnD9/MKpwOtE
Fn5HfIn0hvjGeIpONOGuTT1/ZDCE/rCw0pD3jtdjIWaCgGV0O4vunv18+zfGBXDw
KHNcEtsVtHdTelkrUyigyMzotYsMdWq2ajEMwt4o0kZCSmsmtA1wShp6JFAb5iXB
DhRHxHmx5EyBk5dFVmu3xs5aCVW2ZEUCse6OcZpFzfbzK0u6YIJfRzvgnM358fA2
yJmhFMdds5mfk+8KHR8EZLcBElXC2lQ3MKSzrWqFhiv2JJvDgQjwuicG9apYixRn
l9fWMwJui+MjEdicYkopWMTy4npWiejWn4qP8XM2oKjcU3SWmacaOLDaRr26fv64
ED9EW5J4S7wPqkukfdjsqTyRM+jBg/aAGHkpkmqecWtN/ixru3CHDkWdrFIkmOcv
ZrwyH7FCeEgugylmpP3sLzdeKFmtZKz0E5AHzLI1QB/6DiKnaCnak0fyrB76h03K
+tu5vlby327UpW3xvp0uSghlVD/mMtkG+F9tXI/zqWAwglqYFEOC+/ikNsfl664V
nnu1V7mjIxN5T/UhJgu4nECvBizXJH5NS3uBxwz0Pw2KLdV3pZelRG91hOYr3Qc4
dJ5gUqjLIQS3ZBeYsDMKHLjQ09TXoMHLaRE4YXtBzvcQ+c1ilKqMeOD4JYq5aotX
gEYj/zKSC7vzV7R2/grCnTzR+gFFy18avzNsU3eajwfxfbzz156kl3TU8072k/3v
Axrrq5We9LpNy69Q21dRXuH6QEypV2jgDdiXTRKInBmPa5uwLGZHOXKjbX7g7lCn
XtScIkBXPYKiG4G+enyA/AahePiZqqeHgpntOujqjbZxaetBaNdD6kF3DEH9zEsL
MX5qgf52zN9BV57ZUO4buN86CDqUsLaJhi/1vRrs4X0KK7Y/8e/CpvILaJ5gdf8F
un35gllTjzlMr8+yFe2ZoYaGkX3DpaYsKlHjBQuT6xzsvDPIFeISLMsJFK3sdZED
XZiij4cA9l9yQx9AchnoBT4scffCB5E2YjVveQPthUTFxKImgzERukSjnh9zuFBK
VpVrDG3b4815yt8NzH02TuXZhkp4YBiWq7BwtU297+8oXcxGyM/6GOkt8Yqhy8Fs
iaGeEsBe7jQwl/Kw7S4pW0rDxE4uuJ3Pw2v03uWa9Dje8tesQdzlKYfxwv7PIB5z
oofHhZUep/f1HutWj1EXQght/s7qPK46H+Rm0Wwdc5wsoknMAmMYHqlfefiob678
EqL6ZMKht7QNNjoORNKjj7k3vJhuj7IN1LVcImHhtyht8Rf2iDXbesOvyiqc5DUv
8SA24FxXlCPiLQR6BNkgy0O30PYlPpXhqFesC2sZ8vIdJaGf1kGDxyfNi1BCnvOS
u9n1M9f8Y5pEwF4N1gWShbz8GyUqdHd7jyUrrhaTtZfdc8a/GY7kx1ebbPCDteQ4
J0iqsWGJoeQ9f7Pq1/+0OyWZ0AJ2AHlVETFntLzX2CmbmFEBRDRCBHK3Se8Fvlea
UeI3JYQoWqNBnADzVXs1D4hwftPEw+yDnQxIxz2/dM0GpPL86lMNBfCBnzrTLGv4
HK1yXw+NBxo0wrzm0hKcR3HCuYNVoCG3jZlgYUST0s/21l7VhcBCxeEZTZCIl6tl
KmugVw8fCu8d27FHy8Y7ihR3uVOG8SMu+H2MGmYP//PDakBuvGaw/Yx16S071unB
4GyUILP6isQHEcVJhBy/5Xz8kvJWZpBzO9EDZG1G0Ik2t3HN8iHJ1dszgjkxBqWz
1meCdNEhbBmoCd6bW+JHU05AaW4HnHcrwQ0DMEPtRmloSVcUSrE5X6SSr4g0nt1s
8S6F6x1x4sAkm1NGQkTtKzV+7Ysby0a3py/ni6cc6gE7MUd/ojKDahTIfhKuZVtE
3LRtjoWiIQK5dI+3yQKxPHZ5lJ3yaJc4FGtzkEc3kyNQLn0X/crzYTi3J8EiH7RZ
tfnlsV6Tp/YBOIlypVxt3KnBQIw24PzeipRRFYHDviChed9lH7rAeKx6J10yQ4Si
NqCL4eMP0avUAkFuBZfGyCFTcsU16qzOmP01nhChfJK061lABOOb7xRVlsvcwM4q
3/hQgU5C49zSf/6ua27DVt+PfV6kboXh5wQu2dWD4I0EelyYLY4rKPpG8svtfYGf
cNLzccJ0/h14DOiNF3oWYuHgyFlpnRDrciXkY2MSpXAo/vDZ/NchOqEM/V+eDw3T
EGhR9182LmEbXlgKKVLFjG1yS+UEDCjJ2ZRxft0TM8nIQoSf1ANzxRqBhF3GJrBD
K2tALOBirJSgwoeeiGgsEU7EDtgWfeEvsOftLVa4a6OizkkZBEnz1ZQazf7O+WAP
phfTueXbQyvuiv0RianEMrbZlTqpWwqPddolkf9Qi62ul/SISp1Bm000LJMO3Voy
2iV+j5lplAaZ4Ihb8lAqW5suCo8+ydcrH9e2ouHvwM+sUbz/VfTMdM+EjwYDio08
m/qZxS8X7+ODqzsmw+uirqb9QZcxo+C0B2u0CLwTeB7gE3sJoKkfolTJbKVvMQjW
LFkP5+G4ViWf7PJiUePolvSaNK+zh1SUOV4MOF0UHq9kQT7jhJK/4IYn1+lzIUSH
LQF0g7YGpdtJG5CaOlxoxZU4MDwV17QQTZaarHXu6ISUIk7Smi+R0dy11JOg320D
ixgw0VYZE1sFqUwIjfMv8lYmy6K9KCZC0esnMmxHR4u4nPR0jkKZK8GAQgR5rust
N90eJzaX40PRIUZKm4Vz6WRpLdVZojbnaOqaCB69OvHY1IEDWzFQQuU1U4KMuGL3
PQDI+xG0uij2ApUFRcYXO2tTk2h5cAAlY85DujOWNSRCguQTj1s9cyE3uvJ9CEEF
k10i6xcfvchdCPt7uD2f+8d6gp1tNQ2A1QkHE15IbRhAB1dBLLHNDQ0WMzifNdRo
MXbP1xaa52xMc1P/fqzLqwWrFzNUNzvquxAX3BjBff1pT1d6QW1hKtDWjtSc/JFI
k1uPsLTZAedVgz3baOzJtEDMOk0e45cI/1NTUVGm1/o3Urv3OoAfPG17nHZz+kD9
vIkIsFPuNFp2SjvQ87CHq4axVqqnPQsZwwJX/FkD7WBBpwApSOcq1EsTYF1DrEqO
xDSOISRyZmu2eMNpvQD7sOfO9BhbYd7+28gc87mxUu+RbwoojnHi7m97e3Wiu8pQ
G0mpegqZ43NeW+sywDiuihLuWPleVTUQUW7vAHR7P1yPHhEAFoSejjw7vT/KbMp1
emGeosjd+vO71UaeP4OuJ10LAzlCsIdnt6vtCgzTc23fJn18//Yhg2pUPATVmyEM
wigwuYWDRo8AOs9YVyrVQ+FN8dRZ8g8O1SW8xJkzK3rtMu9mrFkJ5XCd14oV953w
cb1Kf02IngReqnwBa9hRoA5Bx3/BNDTN9nbEmFMeUJmDA+lmw6I/Z5G91wqqgfvT
sGVWjqRzUV6fpGJ2rfQ130DF/zoeZtnhjFKmJke+TrQv7mEm/vSFciyuPF7c/wER
whiBBQ/PMMjFUW8+9vvJxvnlHNPZvz4tNMZYCoHBqDb7BI1y53XzaVw071v7tend
EP4tuKSizYFBC/f0/1li4K8e418C5Sr0fn2AYtM8s06bfo/ee8MEFR4FgaeA1m/N
7KIGYhnUerBXQXWrnPPV3ga/JGGcIQJSl90IR6n2ubP+26Yp/mKpy7tLxb1ikH+5
Le6DrpWyIuRX/j7cm8q9cNSXVGFdUlitdrmKhrT8Y/02kQLN+nrrLQL050YKZ8gw
nSBQUKZZEEt3TwGk40gaN3YNWVAYxomty90Aocn+O/wWYSerGNqxb68dXmAQjcgo
zf8ULnPSf+PXGh6OlQlLyXMySLWKiy8i9yFoC6ypEc90dn08KIPXN2RdZPuN2Jgq
ZGqyGhbiaqP+3Ts4GDy/+4q4K8jJEVqVkvrWKz1ckHfBV+mjSI1OS7d5ORBNlH2u
hQoCikAdhYGxAGrvxbxdQ2VQTDSaGHjEvJ0WCfnIw2ssIcdjTc/DsxY1GUQ5wj03
SBBkDk1+K3IJkJUZoRpOsVnHDaFttwf0+Px5w1FOHE9klV/ug75KC8DA6bWTXlhH
L3yAs/7RF0bH9+lVtdPZDPD6GdZLayeeVA+eCnYJUgFIoeDUmNTXNk/3j4w+Ezec
2TN3u0MLxii9Bhqy4/rGiUJl3Kei/k6PBdPpeJp2+fTy3kLNq5EVEt3+bgDkPeEf
octOezAI8hPXuN+lgg63Y/b7NCxrd7RvoWAXDDxPpcYr8P3vLW5SW5MH5LB82RKA
kJmtvt4Jfzbxd8IHkkuS+mphuhciJDAwBojW22K00+8farKoU41dJ9KKCBiXG8qb
xhQkVIIjGfAFuUEh21nnzxJftPVgCW7Af9ZKRggDArxUAhs8rq0Rz47B5XcMpo8n
RQKS1VcAF1BuS/EgyK7x+WYLhOSbOrxbmxI7R7uMdgt5P0ruidnJLZH/XDYBeUiY
aydY4fI4pEzzzVZD+S/7X27GS8w+CL4rBQ8u+hdRAOea229pw12hxnxQ24DaovkK
U6EMDmOk0OsamLRno5+oOxJTldgCnNg9uZ8MW5Jc+SuXEVozg7UlCLglJ8mW34nj
4WT8EpcUL6doej8QqmYyjVEVhO8MZ+kGbEilxA0CVWo70FKbK6Ji53+2vDW3OBL9
oD2Q+OpHMxH1SPTZW/BbxDYxgOua10/VVoIkKPhr5QQdyP7NqYIt9WfBB3AMtMVe
VUVsoz0Acscfcte0amtPU4faMBm/YXTgq7KZa/txMcy0HPikouCX2JqekJWC369Z
ThMQWwpk1oalm7gSUEueQ1HW2YnaeAvwXGUd8wjEJ9Sv4pkpp4s6nZRkryF0XOmJ
sbmlPq0sGMuQ9hzFqmb8abFc2E/9FBLOShwv/XCQJvXZmysOsPs3FKYYavAEzbw1
QIbFYJvSRmMVMzZ6ZE9U0oZYknfpsSQGMg/MNL4tfWcXT+EUIckyjFPiT2QO4ZZA
yxZLOQeX0f77Ch+URUKHeIYozNgdlodiSj64tqyoZ/QPJwZMynsOhogrrfEBFX27
1c00gmdv5CkLXp2P8xzKj0W5EnhwUbwAzi6QCflO3vRcIEki6WHuPSj33NJr/X6q
8Fimhun7UABpaunZyVOx2eCbUPMDmj6TOicrPQ4/rR4CfKaZ+Ye9Ej6smdqPBse8
BEbWcNyDXHFNl2eRajck3UgleMsLcO0yE5di9W0ysVyy8Isnq5mSMwzXn/JVwgKM
VndxO+5X+QIDlDZgcF6D7+PM5zSkjUbtq8vfccRs+vmrA98myStBjUP1G43GWaPf
n6x4Kc74yfSfriCXHuX10vxpl9wCIHyZu3pdi8mt2Fsjd7SGvomLU/AKr6k32NZr
Rok7YAwJvGZnPd6+g32QUgyJ8b61QDRjvcYb/t73/LnyBA2e04tX1unFaowtddiL
lXb3EA/4/UA0lvAuEFT2Yka1bDzNol70TfL3bhlDkHFqtpqlyZ36PO4i9j4ZCFwR
ibCuI7IrXpA79IrlsPfjS5fkzOw48gyD+yy1XDr6kkZaWLJk5veCP7UYIe/TWJD7
84awa8q+n0Ru/4PttpsBAeE1B+92x+qDHZq00qnXORudnmpos6ewvG7iS5Yipa7P
xUkE8oR24CHZs/iddhEP0IHihm2l0uq3Ojc+0Ke9eIqS0IM8yUBmQD8LxqCB1E//
tTvW4p27FINDJwvHlZHku8qMvDCaoFZ7wH0yLF9Z+ueepPIUHKVEhuDRN57nYp96
PcSU2ZhPvtwSSK/rdUunjHVN4/QFE2Lnk6W30ptyH6l74Vm3xkgAENtAcKRneX/V
UCxLyg/Pliopk4Fbg9MS1TJCNasr6exBcl9wxV04PUnxUxi+nfDQernE4RUVFCXo
DJjPaq7K/0TXhRwxZPG+rerT2eb2z7geZB6QWwFdrTkTq35gzywW8JByCU59rGE+
dVBqgPJLgM+uxl8lyqW9i0EmO8CasCCqTHSlrO1u1TXxsCKmTwn1N7y2y9pCdaD/
CfdJ1wumMD9w54fW2jNkNtQIyMfMx4i+obOetKEAglsP3+beIrwYMKAa89tyYa2V
WD/dxJO9Hcti1ZetOoQfllGjstd6QbF+Q3vsnpXI/VjnVmgY/Niu8Tfdox2F38lc
OJxnlVooH8Nyk8VoelS364V3CDvzQ+4RQyrv3U/I8PX7DhUql/fDBkgA9gmp7yQF
80bOjmtasVB5CQlFCkLQqk03gUylB5Dc8GHH2A7BAhUAwNfhPNEFYoLpT7jL+CeG
6d+2GOIAVa9H2npXfxAbO7o1erbJ0dxd4V86LzVO0C/3BKRe/XjvDK2ZZ0obaYFa
XPu4iseJ8qY8sfvZ4nipCb0kua2VfeuCwpZm3swd8cMNG8QWJga+kwbM+11VMspc
wgTG0ngzu5mCtr3QJyjWQ29TRWnYn+UIr9bjxLMN7293YjKD/4LbKtpKUoap3k5k
wBPO0Lb3j/087eP9b7D2G9XUhybUVITsdOhbI7CKqPDEGl9W4IcmOfQIRtzsUYBa
3tNwmDBZ6fCQoirQUQFBRsVIts+XdxmcB4M/onnSRxh2rK9C1XT/yKt8mfVdgd7W
FByW9lLa+Z/6dg7NQh163DFyb6ugntISDRJn69yXXZd/I1LQNtkYL77VmB8yURs/
B2VaXhE657TlgbfHjTbVjLTQKZUX1WXK/yS4gJPT9OJPzB4mwpURWSuOBWpwxrjz
2zrUfIC1q8OujJWppR05NLg2vtNzr3tXMYdfWm/CVpZMIu/uGTSPNNFFVZBo0QzE
u0xKFinvgPxqEFAvJ88sWai366lcxBTbd4F/Y5kh3S0ZtuEUJlYdWH5e63milAEO
AZOJ7eHZf6aSD9A6dk9HbFmL4VZbCj5Bboo2Vge+U49gDZz3u5L0F0Z5fdDzWk4C
xjGP/DZBrLf7iClpncHO9AV+eJmSbf5pUTz4UrkQXFB8DXDWKiGOHFxhrLqZI3uN
+iBUXy1tPwnw0paJ0QRYdnFpZwqTjxdowzDCyE6ndU/bhlTBi/hs57ulYsMK55cA
oCZKCfDSYmSn2aTdD8RUfhhTBtDylIEWhvzrl1DUHF5bmSGKqCXvLEX/+TG9DRD6
PQAghaGq6uudnjmfOhTMXu9MzpNjwLiOzpX1DlS0xtVBAir+PliQTU6OFdDrcpq+
E/h5Eu4HzxDprMSHwN2P05CLkziFAMUkjla1HgGnaXbNLe4/NoVG1/s4ZgVO1//N
lzvkTbfHcji+JO62uBgIihWuOAc/d0KuQS6Q+cvyotcRPGFULo/0/2jwalmrvScD
qEMn3CoNnNUiJhuW7deQVb68x2DoN3sNx0Hfe1pp+fRy8T2EBcnX3GlLZXknacoN
VLJZdhNSK6caZYZnJ6hB/pItWNr/9m3yshNCgsHTjiRVH2h3JojkBiDoxAek/+ro
iGHA89NWanxpSkTETHPeBbaiqrrGbbWBkLmYD+A4k59vs+kfioVyw1snSo8CMWle
mSr1xhYgyiO85D90kpJJVUax6G39N3SXq8m4o6qbNH+nKuaXszLiM7PztUP7NL/d
/r1XhxPEMV6xLa0SGJ7RLwakzkq1mB3v7w2Dk5byiqfuU2AFozTW2IJ11HIigSTk
EDDxcQSN84bRaADSCuAs3jQBt2F7qcwgodC/iMBSDQEzgDoZ90F9vn3lJN9tfWHp
BvGIatvsEUTQI4qc9q+Jsmr6PJvhR2iVqMDEftoQU/jotBSTeo1QUtl0WJgVv293
djKYVXcTY0QbdI7fgDaY4Qg9/P+vA5DcA7yQS1bkUQd8WRPcrqhmXhyl9Ye5f1U3
BHI5HKd3AM1FPySdjSCeEd+CPsSk1jUKtE5pMck9eGy4whE8XpFTpVmCfgTu2geC
VawZm7BHFonRX1SgDxJDx6pliwDsdbnG0UOHAcSsIKHZUvIYAq7f4FUMz7uXH/v4
KGz3RNXaXnbdrEGlwfbHdiwZj92bHYsh5GzIK+8ZuKPhcnFVdYUVfUWWfaZPXvqg
ynO7ecT+1c94VzLDO9uXv88CMvKXnhQCvV/DMfZ1eQlYD5Z5D+VxzZXvpIgPsSH3
Tygnd+xCHW2h+Fq0fkVoxJgb0S8P6H0YVe7xIeeIDOgs2I/5FWYK+lXwdwsjzXTH
n3qHsqrUFTtF0duwYhc5ZsyWp5YyWyYoBDKporo6rPrOlGO1E79XZALVrLgRkdyh
Too5uPWkzBqfJ0Rf6thgUI0/0fwCAEpUTNOSo9PjAGEz7tVEtoygDOsvaa9hmW6M
f//LWpNR+f6NWB1ivhGuhfSFHGToNuYZlm+q7JTC+zp6a/AHDsolYaQlzBK/NDPb
xQgO6kmdlA4t2RvZTzCoQTOiJkHvJOSnnWon8ZDtkiOfcHboJsnMCxNFB86HjcAq
iwwOYBB47/JkofTJW3ScC5zK7e9tOZcJ3KaihvMdEfKzgsp+IdmSr1kdTW8v5v+e
26pqfxyLPnkNrAbHc6qDJNU+WjWgQ6tmt0Ucj+iGhn70aCxGogG5D2yVEaS32vX7
QX1ivSAg0RH2d6y3KkjBapHRSIWkgWDFzsgczsllgtRNWD85Pfp8fC5R6e/IBUhk
6bS9apJ8b+jwYAmDe8gRT1ZFGUgAfoan1klcWMbvyv2Ij/ly0xVU8ovRbPkXIgKY
5Zwzdhh5WzmlO0G8/3sEvmeLssbLFrCaSR+6uAraHRtO89GxqC1cmfBcErKIj3Ke
SyBzcgFPN/WagbSyV01V2eb1ersxmuHxyUAIlp8f2K57+50u4zyawMSdSovkQEBc
64FEHUZ4ckRF5bjtLxFTAnuvuXh2TPfOuxQPm+lOE28MqkwwShsMMJzPa6E/ghra
cctwZGjRzH4mdl2HBYRmixltuuJW3zoB+hImtxwmcQ0A/T46jNjzTOXDknSEHpI2
x7O2afkx3hf40dO+kFEZ2h6R4lZigvqeFu7WDn54d2+KKXB98MaIqKdOlNqRsNu9
wENZ6Ztp0EgUD34a2WON4AgNDglQmkTOnIXbNbre3azPiiU9zVIB2LgiJB9zDY7s
CuM3om/VLmL2tb2ZYa0jLxoN7Y2xpXM2nZalyHFroJGzvBBYRUaxagCXk6ueRd/Q
AqOIxec7B3rHK36NoBHlXc0PtM5jKQn5YDYfSyEsFNgWWdXPssef+p4pOE9d/rDn
hV6sw7kwhpD6fkDg4RcqTWRPT1/zSvkDIIaMSj3+/2RIjNgCWxPhz88Flqys9Ysz
I+odMwZLedcW1QqU3NQUoxFeD4cor0rV6mKiacustpJQH9tL/MKqYDT0zqQJaJ/t
/YDdenu8jvGsVXhkoUyeYgtX4Zo0GJ8zgQ1KxD4CvqoFyITceIpRkiGzVZ0ckgj5
6c4YNh+Dg3JDQU6KLQNW74oqIiKVdNZKaRZltoXuixYUIp+MSO57/xH+TyoFNC1U
Ao6W/smv973iV109/x8ouD/1sLodnvnZFXNxC6B+YZBkikHhbQTjPqltw3vMGOfV
HxWSVC4NDGfydSptXjRXw5kzXz5dtQdBntYHmGuwRWYKBcObohoaVk0cxiL4A5BV
zb+TlBvTBGZ5jV3UQoWKzEKAE4/CfombxfBEimc58UsldUJU75MEb7sRFEFVNzaW
s4MWM7/fDKtb2H62eKIWqt2+bSbkpI3X+IVuaqVBuBafd2gsmit7pXDN4F/QmThJ
b+gr5HLAeseAJakqBITOxf99nOX0de7BvjFBE1urOqIGyBgey50j3Pyyq8H97TUi
sZ9a8aay75rHb5/AkgRpBc0KyF3tI1+OG75PckkKourYrT9FHHm2UX+7bBbc8Se2
8RuQIqynxwD6TE2poE7PSJ66VKjRRetBUm1a6qt/8O3shoGDOXkpxsSw+a84Nbu0
UaTsTRGbeDnIJj+/5OL4eTTZQVKn/DzqGrutkzqQuPFqRBEcsKpSLdXn7r1CJ7kJ
Vgj199UNB1cMAkzZfmm27N0BaO7ocgi83CJV+Cfc5MA+UY8E/x3vIiBDfUyaT2yL
BZmrqQXuynYTxVYQH2UjQK0vKxulkRFZuHID1fMpjsGCIGUNLdZQ4HnDH0EWxhd+
524Czdz0Xg/5ZM0p/R6bP8/yXgj7+AAKER75oLg1fNvENDwyA19TVGiAvOzKz82p
n+x2wpnaJzDzXSpctqUE9NBGA3VzL8s4hqtiVu9KVVuZ7g+goHQBlKlatmsoxTUQ
nqCetrpnTiv0Y9HDEVM7RKQnADOhlGE83Mr7rmItVgbmkT6kG718gDC9HGsPd/ID
tTIUBVDkAgi2cQvD/0Dhxypa8LX19HOb4vuadJHsVA6vZeiU7wc3+4DHu57mb6ak
vATZSQANyyTGHpGG7SX2amMT4ir0+OCTGRBXIhlFmi+T17Ck/z6ZZquNVbAUR3QJ
64hYEUVL9a1Wnxoa7D/4HG6JH1a3MPAism+I29qJJMh94cMDq42s0+67mwSl7Pqx
lcPGZCiKjig0bMC2+LgkPqW7j8/uWQMmSowJ0/gYRw9faxzzjuWY27Qi576FgPUe
BZCE/9WHdzN7in1jClUbsGHG8hEiX/Xr4wBAzpl+e3rdVynEOWSfVG+wlJT4yEcZ
lLhiMYrrSn//a447dZGuVEA4ZiNPg1ZCbl97xBVrO3agAyErGYsQ0T7HJNpR18Nr
ehoeolBcqtq6RoY6jC0TLgSEGHPcsuiifO+FFhHGiPz4d198GIfmcZAnEljptKir
+hLqdNje/VlarhRUEZzFsfl+vxdSDHAkhHAqPCP3/QRJwgJmLdNa7S4802LRq/QI
2bBtrlFVTKLMqOLJFGv2OsHEB0NoImQ5HUubaxLzvmPM45sR/OTEUBXC2texHVRy
TttHSLU+zm6+n8xz/LPAWbZj+Drw3C3uQKVMiiila+1U/MgtnL0jXH/x1wBwsBys
VleFIdgTL6HWFiAFMbycON7CvstdxfixLpDLrTdcOj15dFT074TZqcJ1DKzp/9Vt
R2Sz2UBjoL91KnjTOX8ol8D29ocu6Qruxbo5UGUPY9lKeADvD3vLs4FLHOseYVQ9
1Op0tU80b6WVKohz3X8FxeYUBlDL4CcniKnMy1cg8HFNoubFCqfnsDj1DToq4mTk
BPJaGhexoLcW6Zu5CRV4ZCGiQ3YyICwDaHYH2NaTMcskmNU+spHiPxRmLKDxH/VZ
SouIqj6SQvLD3JwfnK3I6Rl5t1RdA3JOrV7IuR/tgHynDpEAWYSdUl2gQij+PnxL
V2APoicL5f8NadbqB4SNtKXRpywkyTv32c5+d1UhetDdZ7eR9qRpf6RTcuCjKoPP
dYaLMWzw9ZkJhQpp4a0XiRMSJVLshEn+HuYqxNT4VMR/P9/xK6hsf1oJ5ucM0G+Z
2oSh085n7D3/tGgA04k7t3uuoHIN3bpUMmlUp07WhHOYO99Gb7LMEc2htvXU+349
hpaVqfP1vcHXBOsaWPQ2ioXfB6x3SBnbs1hy+onNW7jv50Zwpu5GF5yI4INvPoNU
AuvIgbVPP5lofWL1QTOqamyrUQILRmTkJMm0VsCa/DocarH02P2aaAEnwfbKRVB7
qOZZaZFJBUWeyWwt6wuf4OdeArpSW5jkrjWi4EWmbsieb1slP0QSYH+aXyOPwFez
8oj0FWrfQ5yhBvST++pEtLnv/UlWCPkBtPxDLWCZhAeOoNhom72/y2YtV6EgLn5M
ffnF3QUGSs+S7OD/rpLjnYO3ux9KsVEfIDcRDKp5yXMO0fT9BI4Wej5ZTdJKVcnP
4PkDGI1nHx0VScB/z/+6lUM8hXLooYPLQrIg4KapKgEDeGS+wgIsicjII1V3otA/
OEEZ6nrxJeABLLeSVtM7hFFlJnZfrixh3J24/SBdx/PCd6y3QG2SCvWc7oeUWB9F
GtdfG7N4loMpEcZlcMtBDL0B+rCQf+IYo68KV3JKEgp6RVOjxiDNgDGEgGs/eGAy
lFMxqQRv8xAQHiuyykcX4fhyFr2fWf4jVIhw26anz7iCasNulixcqNjCQQhkUUDv
3sTW3O1dXonQGhWlkrkZLdotYvqHaZ4YC/BrfYQtuovIxR8oVVf2lwai19b0nJh2
1biEYEAwLn9GUIM63pggy24uaWDj7kJbM8tBuem6aBp1GbpFC054LeS8U2tSklO7
AbDt7bSoR7jP6o7+0oiBtaKLw+Y1gV4I8skDAT3z0MKYFl5X2mias3eThuoc10RF
qWgQvezp41LfDjmLaH6tunosNtsfZkk9KDYFmzvsdvy34kh6CQMMEsmmXMXhQmQ9
y/TJCWUFr0rnu3u5dHZhpKYJC1DfiYMYvqR6MInRwZ+5cytwSuKIOZ/mOCWhI+4N
xSHeypD/aaVxCfkWdW+yIZuNiFtF/QCR4MIURkR4/+s9iZhSGFAjtrk4d6Ud7L3z
ucFyFWBk8ul0VVsK0Xzxs3Pk+SxLtVVhEBC/uVlx55DdcgnOCVDtRv1e4mUfces4
dz/H8TS885KKa2myqy644Cuy2dgu1J8/3YkLi+fIQISAfR36xOmGHe7IzQ6fRKso
VxG0VxumE9hA9/i1+g85ehk7o6mFtbVbQ6QVGOKc7LgdITciW/E3tnePSic9PceA
nOuHlNNiE6vofG2uTmiFCOpCbPwiIqjc2Yn0Zs7x4/QdObifh0oIuuHL8p8+eeDL
d0NcdZTVoih2Giz7tiP3PUOg/odwcpwsAmP8zttO3h2KIPdDBvw3ZmFN98yAJA1+
Qftw4ECz2acGL1Nq5WdD1lV9YwVzsqj2hrqJ/9Notn34aVmjQBreNVZFKhgfEZVd
bhb+KiYjrL4ALgGqEy8ErsRIoSbWsm31HfSiUFW1s/pxzdnn2+Jk3EdGpysxzwVt
D36FrAZemNgBygrk/+tjd4RpLK6v9O8RfLf3w31uLr+mgIhIOwhWATkJHnIjKCo7
YrEQ1JknPBelz1U6Z5JBuI8A8Zfln7ovYuTTzBrROWvdr2i//75i6APHMmcg30ZT
/Jh5OtUi6D7aT02C5buy7VP81Jx3PQpwVeIec4EFZGNSUxVPgZcYSZqVGyh3g4Wf
mHdqJFookkMl3lmmr9w3kVfSHVoi/eOaLpHupGb7wAKA5Nx6hElEA41UjL0OWKvk
pOxGBlnJEppcWn1LLBzja+6+6BB0/T3+ObfLVPZizsk70EVXLzcqCNi7YK4+NPi6
De5qZy6pCH2XUrBJbd56sGLdhFDb6FN/hEyyc1/SwM8F+6qNeyCeXEl841/ay+ls
Aa0rCEZU+N1X5T/5gDUJzhUYmltf1dz2zyLVmWIvfXh6DC9CBAX6rAxIEm5BmJBE
VoqkA8c5uTs6L5isyYgAU4rIabgtCA+9Az16PsZ966nx0Y58M3OOUbDe9IPrTK+G
Yxleom8a1sB7Y56DNy9npWhGLt/9H4Dvy1tz3f3mF8IwKAa28sB1jpxMqpRbh8rb
qVWAR3iwTEEGg4HWjRMs4dHO3e239BOT6zkEhgkT3+YFk/gYoalaWKE2u0y4Gc/s
rqzZzAFnZjt94qOtYoD8Z8hOIv57DUZ1pW50+6M89cokcHy+b2xeLqljrm8ySf1a
R93lPfmcVmnwuvC6YgR2tIXoY6uTmfU2YcrLKOWxlQcWYv5faRTcBFEiuqbf6hoq
LYGT1hyLE6xB+iGwh7p26u/LxRSWzOjtBFk29irUbFStqzbb/eVcw2JnEZHqNjSa
9WVIFpxCiXkx72srfA4ZD/G1Se/nx6W1Y75oUFcL8YLxn7kCnHhnVa+3Iw25n1Tl
JbAqa6irr2n//xjO7+ilP7PGYX7tcsvWGflBLOJdzcKMK97oezPbvKOtpMttkYp4
u7R8rza0Qio33RsnQZmvaQCKfF1SQFlEg/y6XRh8TDdTa82Sv1OS4GKoJrcDpc9i
MNUCqlsL8EmNh+qo7oStPE6gcebOSwj1uOkBmueXZcF7R59f7ELmmu4ZXc9BPsd8
TdMB1+SPCWzoyQ2M3lQqytvzq1OQt7nxxcCXq5W4obry70ikFcgU85hrpePmDfoT
VrppkZvZxDdmAbG16J0bAn3GfV29ZD5jWQzk3BT8G2r0aes4ZTQX7Jl5e7FvCcD7
OlCg+3gv4Q32TOCp9s1QgsBX6Y/se26XnCuzHTIaYKUGeIjTeh7U2FXUAugBhs2C
vpqLuDRjrCOjvMWnDrLLF+KsNlend9QGNcl+NUxcAXy8K/wVq3B3dbZTEwfniOfY
089KvsAl4qkvqq6cWpeWfqNUp5XC7sN9TykAM9R7UhNFmb/hOoVTJza7Eu/xCzyl
4y1l5dQqk13Il086FhwNvmcbBa6xta4XMqd6zvfjzQo7enAOWGhy5QiAOlxNnyFY
hPyTXEdVEAf/c3xWl5z3sdT5TOET8xWAdYY6ofAqHZtit2l0ZqHaBS9FqLUvMAtJ
l8FyZbBUuLSG8K8Lwg79JiJ2i+KKxvivxFkWy90E1wXjKqBi896zSae9l4rolJzN
DarZ3wmWOEjmSelVtzJ1hDTnknt0wVaJgMx+NGnBhqBi4475LWbUQJItbSl4kE6L
yAF/zwB757x0GoWSshtLwV3e/3HaIn4OcrZT6Z1byY8coLBseUEoBk4Z9cqgR15v
rVBX5jEbZnTnZSRNyQ6L28JVtOpL+HULfkHapWPTGEqdsIa4SdpifYiajUyqP1Vp
rRt+fb0wBVtv92pv/xwfFn0aP1GgUGKNy1gFPVlaAwyCrZl395kWNLSm0qZL9Cd8
F1tMsBBr++OriCd72Kuo7ICLi4MP4UrboTuDb5FTeTKeKNZdKnJ7JkI3z8aKHIyU
tGxyamUcYu7/cceNUo8I8VsxWO2XinY8b6t4mtGU1vIW1HFrmluMqstYi5174J87
X5VQUnMrQLOuF9KS4YwllVc/svOHMyj+PV4Q5TgLQX+wCZdXsDBgLoIIm0cCSV88
JCjLBIpDXrG+GeAGKvsWTxAPGbnAbexQSUqkY2pAHW3JjKq1qbTxS6ixUgaxAh9g
lqwGpFa2E9bPsGWXiXMMe53m3fLrN1wknhCetY8xrJJ9jepM5h2c5Gelr/E6BPRY
ozKMNAHfoTVxvy08VVdjl8Yjbh7NtIIHeo8UYrtBd+qoirdqlVEVgzH+kCdjpFUN
OOAMTra4QUDTvsEvIdtTYlkKVrSKLIE3cAWmzuE0KIdBNyP3qqiRDL/E6BV07wis
jTYIcZrPcJtBvaOlkJigHdjvkMV+7upUNZARrd/CMLEHHisdbdkaQ/LEtbMHzhag
4+4BPTyp6+zCsChfPgt7pfpassEE5tOFM0R9OG/1V282xsE6bhfBiVpbm5YtEjHD
h0Wi9K8Hi+vIq3OBYfBTrg4LRiRjWjKb4HX7fD/5lWCDdKT2huhuDcV0JFMk3IIm
RVzrFsYh9pHf1O3F/KNVezmlSRpdiUL8mYGzwxlPoYU+Xm9nrCDnmKtX3+mpOJhe
p3lv4QV6gQ5HgIAZx2N5t+4OojYSo5I5hxPy5ccwMQzS8Hlxq7SiC+kZqHHFu4wC
72ZYP3zYslhB/lLNEE7MufQvy54BhgWHrA4tJwkzTVS+SlrfEfcjy2FctE+/YXav
AkTRU+9STxO1xC6AwKhfFTIz3JGKl9n4wG7cvJNTVnpm6spNRTvcuUkFFYDoh+8b
Ec86SUTMk9w533jpVfEOYlI2euE467LYouQfNc7fRaHdF5E8njrwC7TJAC4F8783
8GBvEAzHboS+gzFK/9zwHmIW2YzrBcASptxLodY+OBt9IN4wgTnv8el6I4k1nvzN
qCQjNNzKx8+gD/UXCCopaUqTIzZmcTNdm/IFX3nZrfLj1vfXBdtAz5CBrLw4snSk
0fzHsa7TX1Mz+a24S92V4FnIsq0yQBVbrmqv0MuO4ohvXVpMImrOPZ+Xk2/TCZJP
nDjeJBRqvYs+xUIDDKtYujPGr7QVNvAasNIb5jaeHZjYup+BUe2nr42wty19Hftx
AMSUeBggsx2ayEE20BPNr4f6f1jNn9tGUdwCeeO2lHudmfRkhpjvxgfZFExee5ZM
XCVHu94YNpIauN8WAkLeJXjRFzKUqYPQv9uVYkq7/9xbZtoee1OznaxG7+TyY1tM
uFXVYKXnQS5hgfcmdutpUWYCWOxAmD25cspAC+hbVY3+cCZEfHLhOgsIg6mi52YO
ugkiCB7xCxQwkSPAuddcu7ULxndmwSuXE40xUQX6fca6G9I4vkhaTIubRoDNpbmH
6iQE+gHdJFqiVrszMF0izijWKXmKT+Nxq6T0PtogThdqozY2bq7SSDTFCYn1gZiC
IyY99Moi+TfmxmfaaN39/V3ED6wJHvlq28TTOBEkpGqUAi73BvpKH/Lc7oC+sGna
hPxHmMFpiqdbafvXNAIUw2IjxCQ6sf7/GlFu3Lb+F/DNL3k4G23ClCI2eZZ7Qpy0
PSc1NH1jfk7ibgO984KOVOsLZOSJsYAmVo3v1QoimYgoBvVvtVbO2JgFNH3UE1xe
wV2PHAn3n1Dt5f5bp2y2JWE1Wso5Q64kNhJMC8ENIF/MZ/sAYhHwgjJE9yLkRRk0
tIsr/8VXG0KnIVxYzY5t324asB/R3YjBu7IyYcNr/s4bPwkUjkrlZRCAoZE2juHH
vPNDWV5sEZs3+DRHDhxMPtEWlwmTX+7zFq/U30knACwc/l3Q1611rbI0CAYIb6+R
lVNEdueG4XnN/GgWDnvbt1XmJdOwnY5DJ4IDhefSN3SBGJ6pv39xawq0kXT2wBeJ
mvNqEpFfxwGklP0Zwn6LAGEF4FPru6w2R5uqCVHFmjg01v/zL00lfNQbwrAzuyUN
gTX0YKhc5P8/Xn7xDi6fgg1KAHuww3lYESopYykjJ/5sohsw3P7fHSINtviilQJq
f29NTZ2rxWhXbZQMI/Vcr7Get0cAHZndMYWFaZ+N80RVuUZXlAvRjaptSqHEUS7d
Hp+Wy4QPxeBw3lRVfpeew5TmvR15mUvV9UW7FsLzUCU=
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
SGTaj0u92ox1/Tz4V0PNKQYa4lM8LIposXuxQTWvK5tHRi2nh9tftkvh4Mo4Uc0w
tKHh/Qi63i+CLk9MNOiGJeUbNyx8tZxDSWVV8IH9lmySXkvRN2Rr1EyF6OG0HTaY
vVoU1JC6btFHbdD7G85/7WBSiJQ4hr0ITkZ+xJKUWdoWO/WPBySYeEkuyDEHLHzU
lS1KhvNATQrZdYKggGnuXvzU2mPGDRLagIRkj6RZClT9YDxJq+Fl8w1wdetqdUBq
FmUkiOV3NmPithQhWnn8fGtlDbqEuy1xy1+hxOG+4z0m/D19PhMqtWhLeTt4aqRp
UAfSQDbRVHxomyWOxyePKw==
//pragma protect end_key_block
//pragma protect digest_block
rzbql+qCHySu/c2x/rLeHtMFOaM=
//pragma protect end_digest_block
//pragma protect data_block
6JvJJMsLIDT3CQQPJWR+coWnjKBXCRIaX7X4v0aL6pywCJMjia/+dqQwz55HIDhE
RPMCpk2NGFFE5yaSWNLISqcG5SMBo/xVL5XJKGNQGuaM2TSPKUAWVEJ/plv3A6sW
5xs7Dfk6rhQXHboe1yUdVEVwku6OuA4DegnrrY8US8JznHbXBwet/ygwIMHrZR9u
+D3prdfloJrx8nn71IUj7F2SyYI+HI3LnoqBoyCdgqtvQ5CYtRwMtzxPxSDycZNW
S7jqyTFWGHMOFePOIIHZxIbuOodClnRDA5/z6wh2XPk61pafYaF+ajWBK2vwgWuj
WpFa8h2TY+U1X/kRZLn4ZhyO/EY25ytrDLCqMfgQnI44McGe3LI8Q4XEAOQeUWuC
UMcgzhrZzJC9oGj5AmWrawwZRJHeZxhukTKwqX+uO+o+bHvU/b7PxMYG5KxiuNil
z+i4NnFg1ntxYN4CpdIdIkPRIlsW9Jzle00oEoLp3pVq4g2CmWmNbYm1QPwJUqRW
tuyewyvC5JlEEW3ohKr//jiyQUxAxN1VudyQsHmBRpyXr47ItmEwYm0rHrhiaXBC
X4BMb8LrOFNXo6DIpOx+K/Ui08YXXRY+ANgsrmVUtI3kI+yYw1KJ7qTddD3awpJI
1sxB65TbRp99QRPuMCbAjiforKuJfwfnNRnHWcsrk6WOhT+R/qLbjZJ8LBMnmBup
fPVPEX9jAIIhX4ChYC0GptdcSWk10o4Qp6I9I+KFvBDcydBnVrkFprJ5Cnqr/DyU
xb4sZlIUyPFRSo/duhL8NSYyYBrJJr+P6yY3MGR4DwKrD93EEAGeThMGL0dyljhA
Zme20uNHY1+2Qha9hPr8YUL3IKLbji8BFF6B72VpKEVYYClQIHAxWqqeYrliZ0Hg
d7EOohTFLOET+m6p/Vu98Iaw9mGMmZXDvTQunyMxfodvTCKwgXPiAtm0Xvoll6ko
Da0b2etlkh1Ew7iKbZWRrAfIeQ/wXpL+EcmDXXRhTJFBlDZHQjICinZEKDwWlTzv
Dm3Z58tBROrhuJmCCymZYhG8+E+cZPPzXDFuhR9zPYukFZgq6+n8UYi7DvXikvy2
rM76b+oLEtDg2+cLTf+xYBVhkm+6f99FC1KtrmeArvK4aeTWrpnAoGtwV676hDWa
ToL3rWKfLUaB9bxeD8GaCGqRnCpRZrvfajyPyyozd1/xxkOE4QkxhxlZwwxMSn1r
cvmP7Pi2lghH78RIJxU/OaPuDJH/ez3JfeSocXyE6qB4u4KSnSqfBYW5RIjqX8m/
TUTcENS9AvHwPs84TPU5Ig+bE2ASRA7/3zaQGSlTzTgj3hEk4vkTb/ZElnFp2fnj
3nZadfF0g/YigY+Mwr4gw91O9bXq+uEEe4QWjqxBfMZw0GXNuQOUihH79q9wmKD8
t0kydFGGp6kEcXvAnwOQGKvV2E1wAfqXc8be+rpnF1RvrLcS4ODCaIOAuMbrCn5Y
KTKb0bSKm4G32Xd93sECo4IpNWZxHuno2eDTBRcipekaA4LpdDmr3aPb3/BzHn+i
9t2sri3TFf04ZZXC/j3UxJ5NbG6H/60xsuf76Ycrg94xPJmoivjvMd2fKBc/7nG5
gnQUfw4p81rlIoli1QLYSh2ChPlJ+jiIOGGBm7SmQZOrTgmfvLTRjy24XkYEJ/Im
RV0tHNtYtC/VybRi/D2QOpg2q3WG8KWl7IeclEPVzJF/Z3ammrx7wvyS89NnSour
K/m/stwpOEEfUqwMlWTthk0i1aw0vQXv5U+6urV0+cT72IqO/ENqGx/x+HKZnR5w
1RyTdz57hMgBMS7urugevKAc6JTlnuytyzIWGGum/o0kl++W7NF//LBwCJb/65C1
h+HAfSw53ytjHS+umNvPdyGuMt7JqNhmkvsO2x2ADEHxOsO7rmottrYttFWGJXWt
cVGHQY8cWGuPtmcsPnaGxMHIeYnzXOB7fDnI51Wya/0vhkHG2xVo1GaAiKaNn88H
RKi18Y0JTGA09s1TwrHXCZ9Gy+PCPCtqOxVe5EkVyA4brsQtcL1PPHoC6vFpd+UQ
2fMQ49VXYdMAG2Cpn+dJYfBf8ouqC1EtuS7pG/LR7joFDELfQEjIfyPbz58Z5ULV
XqEpTn99wIsoEDjIL3wnT3nYMMqQy7ROn4KmrCHJObmT261YZ11p/YXIbKiaQ1ZU
h7xo4QzTkjNEmD0+mGu7B9+ynZyB9w5cqEzEY1nQS7ZMgHFGnrfK37fF8bxZzYZr
tMOvcTnlxD/dAVdWa7G8Ai0nkoBqftO55wzJv1dD96k62pgMc9NNDJDB8Rua8CXG
2A5G5pusfWW7xIMtwG2XLv4DqVwZNfBwAfAz/Hq1opPQYb9GvLYMMQCoXRvTh/J7
U7007HEBe/JRJm+xzOk1jhscsbngLWmMmQwubKz8D/73fjTuJo9MG/B15xWCbmrh
FQUMOOtfMcnKZDNXjywwE04hHnCRJcHgVpIhIqJz9BVAd6dtFteYm3W2AgDECjJ9
DhgBEWiVwlCDm+PmytrBNO4LhdAQgYL075o1biRpcJ6srGOP+qHH+rXaemG3hje4
ndLwDNA+MKcYttnCFavTpTItYybhKUYNu0Bqd4AMeaY2tIt0J3FvVnJSf8egzjyX
wr+cGCKtfiNzJaXBqUAkJezPhvcR3xNkK/vugTMH8fkO2H2Thllb6bnCIcmDY4Jk
wFDr8Osfsf3OBDjoWvBje8vmS/HLgBt4COBBNIgJBFEBrrfhAhMZruv6n4yHYoUU
Tw6r/3wA3jRyVZg/xOhj64vVhZTnDGmamO/xyfeWe2vhgKJH4utHPJzjzL7RQn/2
j4O3fpmscbX7Z/8qO57awnzpEXQk0R4qcbYnL5W+2GxBilBdImGfXP5gEpTGhPo3
jisihPc+nmSjXTXYzfXqTRvJ4hL4NMbS3madSAQ1vIpA8ZSnwvsafSa1AWFstPhn
2KE0Vf99c7H3MuFMv+4X7Y5L6nJ88fKbG0ciVapckx1CLVnHiSJ7swVbYAPmihde
GptN6cshlHk8GsMjiMta2C5kbXC2S62PjK/XBgrNwx0tIyJyW7X5i3Er9oU0eUWC
5JEemD0QnZI/aESy5fsQZgbTXvVYl/kg+mmd6v2th1cB9ONipy8+DMLEWCKRoMmF
Qgn09Pz5sOLt6LsU2vvO8820Y2nIIgYpUcncgZ8cXtYABOG23w1p7De1tDpeSPp5
GStJiXSoJzRpROzdvBNYEuohGnASyZXSBDPsIFD0IjUBx9rPzPbgI+jLn+FyHMGM
QhjVVYr8dFa+mfSW2oerYTi9deHrvRwf+KCoop4ylTl9rjhDhm323SPtY20HUwvt
aYbVvjp8l1jfOfauR9wv91mvjN3Op2LK5wmLIovd6b9WO9iOPZcWNhJlx6x5hI0J
AZ88KIVz0Gn41BwsvAzUj1jMM0Z3yOj8h1zVsGJ0cuXSLZ6hXbjIiRy/STNzB07T
uXHpnlsUaBCHu+pmD8NWi0H4pI6m9UuTp6MPW11k6zO37vjeP5YWpQcpCUkJ7L1u
czL4YH+/jVVz6xYcABA3+XnZbVS/BODnL7KIogAEZ4BcM3p2B05PzYPVUTLk6H44
6rN/cHVNMN9CQ+gZKNeZRXVD61P5w8/qmqPVPiGYw1H79HxVZCc/f0Hg1Gs2nUVs
rAPeKxE9ATg3SurwLDrk3ukpd7+j/W/2p/QODtb/mB0bJPaxzr1jQlzxBDmEEnca
r3wt3m+b+GuwQp9dNpwsFcIDSpe2hPzQcPa+SE5+l/GiUg89WFQTbTmulYeQ+6+w
NA0RqygnWeMJv0UIueUJw3OHevFz1DOivKBMIrQdhzxKb3s3SDhPNSMoKyw/dcqN
ccyk6bb8GfVrN0jbwezRvu4sx5GipgZjcV0vUwUqbJPISz69XYBkBj2czkUqxMBq
l2T+6tBwqlB796zTVXeSj+1bxIcwdfgtagB4Fiv76tCBErSXXeN44gBCM06OY5yF
NcJ7565Lpd4oIwB08fMDmllW/6OkGqOiTxOmnxRV3Qbe4gxfd8TlxNbEw8nEDIEB
o58KpNQNY9Yz3ljBEDtaZbs7b0wZliQoMcmZOH1mNewEONvwQfR5J+Jd551xA8wc
43Ajg1Kt53d1GrOH9R4wE0kaXsIwLoRI09IGdV4yGJ/1rlk1MBpsF++t4wlPMyG7
Dq1Iy3B1YEraL+bF2tFLJsTj+1CXgar8T1xIkeh4g8n+mH1LW1MxbRzSo2PEe/EQ
eLp+Ay1pe11vkiv8hAfmyuA9ywmS3DdTWYZ0GLWjcRNSFG+3R4m9rYS57McNTyOT
9PtoVS0uQ6ygcE5PUgI9sCtleV+rn8io9ixVtGrdeXtTQI14QrOW+dHoXCICCL+9
/xjZE3xVj7ot9scStq3HF7v5qNlQYQM0Qf09gOVyzgnI2yXC3Exb1qWE7oMFN0/u
4eRe5cMp3I/OLdh27xXzQqg2bwu3wP9Q22H58XayZcImasb2z3oo7FAjbr1B/YoS
PohUoui/4zrPAsogxzStasNB77X63cl1ohLhfZMU5iAtZcO1JYxTIuPx0UUW05Ro
prdDCCI2RSfmWdlcXdaJ2dWnJNtIgeRq5K4KyrkMQgsZiOxVmlFziSgBvTyzVaGO
MdEKQu/puQpSNx4Kb2szGipEFMdZflwGPVxMOiuJGNZOjT9nQk2/wzafXTrdrCdc
O3Kc74CyRbSYl45nynmQzDLAN3IcxejgnUVpk5ifjVY4Bj30phhwjvE7rP/7P2k3
FnAhnb+F1A6hgzPfCmpyzedHstTLuCB2T8fQ3A3/IZ04hZk+z/x9krhXUtKWB1Z1
SFHZITc3soLH3b8+LgIcJJz038eJzP1pbYmPF0t3rj8DCyOdXmkSsbQ3tPOaE2o6
L5mfsl30Fo9Z8pwMTodaJTI+GhsoDKDNkWgqyoH05HPoqZrqxUidCph4WAdGbsRv
e1h4opxj9OyDQa6DEjn01ZrJHIfnGZ7xWtZJIaFKJnMR+wUFTEAfLsRTX/N5R1WY
/4LlZ9aytej+BpYInD51+O2zJBBoqYyjT1P8PSinCFglCUt43wqlrQZdmGStAYMG
zl7p6EECXNLNF6Kk5M6zp0sxGUdCJjV7bAzwWAvecwkbjo/gy7Tfir8AiODKu6vt
XNuDVFBdYes0Ir/MxLKsZPKKvtfKGPNZoErkqRBlrGHxqYqqKNDXPINu/KdrPd/5
CGqbyeoVak3tfVvWhdqTL4j0sGY0FDKv5+xGE0iJ56It14HV36MAoOdSOkKPiG5D
sIlscd4VxM+B7jnZ1ovNtCTXcZPK1T+9YOHB4tt7KCb54NOw9OMThvfCRy+GbIWv
VsE0ufhQ/+byoGvOe8WIw+mKwnc09NhPP3GuV2qUGOwZtvL1ZAIpj/Ke4oZRILqR
OGWFpl3M941R38QmbYH/Jar+6eAfMP/m5/WkSPMeY0xgHIecqlAdvBi8FmIFcb5V
SaMlOTI+r3cqYPeRxmKPwKmOWSh8oMQLjDOxLGqXElZvc2+AZcspHsHYN4d4P9q3
b/Z9frl/YuTl2YNwi43DlYI6EInOC5/1ZDuxqY7XqxCaDoTYe0X2CGk0lhKmurh2
q94bCEjyXscEdfxkTvHvf+m8uFJ+6J9s4tdj7qcb9Q+1mvYdPrNtFRnnFAWTk6eW
xaL0OyQswCcuFVFO4pj40Tl3P7yrjClDvP9rcxlN0QhqFgJeHJDN0qeTBwGnKFc2
w3YMsSNLQ4LVuBbaEQd+QyM5yEVHnaAO5kztllDOd0BjOWktj5Po0+0rmIFHuhwM
/EOu6NjWiXk7c+nPFjWoFnqiyjECoeg4PPcJC7F8CAAyqUcnbdPTmMDWrQmh7/Qa
DKfnOKEQ0lcPo8Ntxxl/ssyzfahB3zaZaFNt9AevhfV7b8EN+sdueCDRcOPXRbCa
3EWYViO0SZLPI8zXoz05qVk0ScolpvhyJ7VBU68jOPJyJQYhd8LP3yQrtOLtheqt
KiL6x7PWMDbNd+iPy/jrou4eSkR/VPJXw52l+x3Is8PkaMbnUc0RyUhQvx4HBnbU
kpThHa0xTUfP5K8Jh5xvylzkL2XTP+RwDFDBJtuEQstiydX34H4ai5FrPajfz6DD
mdLYoHn09T+q5+zICB2BWkUjtN3e/bd/WqXDieSfcjpCrMVqG5EJD9KuNJk/u2sn
d42ZVtk483uZUS1jeM0jdrBfRUtF5Qfhra9P5O3xImh+E30AejtO5rT2FwCz6Brm
9vbNkeTIcmhIlqQfwYbEotNSGmQ8axVVzh7LTrwSYcmz1m4b1n6Ba823Yj7ehXP0
7fz5PVVVTmfZevcqWEZMJZHrUht45aGjriZKyF2/t20i87SJzG8h7oK0FepCqPGH
//pragma protect end_data_block
//pragma protect digest_block
RNfxynNX9tkpYCyA18UUYD4UYAk=
//pragma protect end_digest_block
//pragma protect end_protected

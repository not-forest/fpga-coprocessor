`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qry1XM6pVEqKeZR40VwduSlpbnqqbmMd6Pqv8GSFGm3nLaz2R9wMhPKmcPmqotIG
2bAk+u4EwxnjqNxA7mDrTiORxibiWVu65DiU5XOfiywCghrC6cFAH1Ci/2Z8P/RJ
7Gm9aHFltDf6tLMv6im02p6a58+2jzvtVnLcgS5KWBg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8672)
RsaPMqNixDStx523z+XMVhe4J93JLgvMxO75JEmnBI0SY/PEi+3LxQL7Joh6hdlH
1lxqBCYw1rXBqmBMypx4LrpePvAzBbqJU99DlDTBK9oYur1DXFTpUUolV0eibaWf
wwdhicWrmwbxPJSiTcdvxpyMZ08UdJz/OTFEwQu06S5C3PU1Jj1/guJSRxPlE9ZC
/YP9sFfBWS0O9z+a4KTlwy2x4z+1yRJhSWIXdTjjx082lE6trGCyem7oLYmVpGhx
mRnoeNo/9sEfQRi6PWeas0HgKm9Oee4HDAAwHoFIVDxT9GSiu8g7Vky2vmBifOjw
Za4A0aDy5jAOjs8goX1OiWRDKVHM+0gg4Skm6+XjZPG+KQYyCtk4D1jtKokfadCr
xrQOPkT1wouoOVpMsB07GHBWYw93tNN9I+uDtRWJosgLDBvPSfON7jvN/LJOAGtp
jR5MKfvHs2PVkPLy6kaytzC6MWVAn8zguHkUM3ExZXmjR1w8nT44kDvrZsvEK7K0
wTp1kVkD3vJuzk0ieNDLQfii7az/yKYFEy0WDCon5na2USmcgfqDUW4eXNL/Fp0D
aNXzMOEUIeVqC/AwLqfEaFl2T3k3mF74usivnwoWVMsJOyD+05QAs+FP1Mr+g508
Y0NqLSCmWU2E+aM+1rbVPDOY7w58nj9Rt2Sj31s+T8+82r/kTBvfgpnUjn7TGPgJ
a8ZtkD34nhAobZq3O0M0mijeaCdcV7GoAA+oqLPwRgeQf5/pb2sqGxqNHc0vcLxG
n07/iXgQiMDdj1YA4CH10OizgS1EtEA18YUJieB78/ACa4RMyL5GhDl+DMTldiTQ
KSiNDqtIML7elGkPkMBEMXwrumyzYhhoXU9nq3MaHdmzJgX6aEBKA8jbrlJxX9k+
cKbai+d1Nkp3l6YsSn8wMMvS15vqtmLyxTiRrgye7FU6YTZ0NTvBEfzwA7fNeAHX
QOMCHdbeIW/THXEmj+rct3UXsBbzUJ9bXnHuCW0lbjWh8y1xaKwkFuqogmqUWZqU
0S1hMZ5OnsKXZKTy7iW/Yj+zPaJ13+MizW7IrdOkYKlDeoKFzBnh+OsextU7xrDN
1wBAPM8zd73kLVNSlHgBU336eyZ91cb7akuzsrWFWft+yt8/jCz/SnLLyD3K+pKJ
YqTrnZpbLqIVcFEZgZWD0Ap4OBqSief6AEfE5hw/w36wpnZ/1BJ5MeIGXi5C4lIK
WMqpMNE4ulVpXFgagtmMMqBadfK3zZODgTSnXNhrTW0kKXW8sjbxKhHLSTnm1Ti8
VKPA3TNq2wXmswJjeq9PcBxzoyBCFjXqrvXN2IS5nHRnlYTRRukyAhBI7LhBarNv
bq8rhGSMWGMarDLNxUYi2SJlapDkHdI556eeNTuBbjfhwsLkbsG++s2Hgqhm5NsF
S7FRaTy+5AFdCsw+twp4mc5TS3CpeoC2n7PKX85g25onpEfGl4jVVWNPCfQ/XXtj
Vfe4trQeZnDyKAj1biVwU3OtcwRRWkvKEIfWyCihtJk8FgXwjI/KBKcmy+uqE7du
yI0ehpf9i+T3byVKYXHxYGA4aTYIbu1S0aKSxgBbTak5e3TCWcfOGy5d3R8QT4VZ
6R7WbGTIpn1546C/TAI5bM53OqwDsMH9gSdUf+fDHUb4PbixDeRFlZI5Y4hwBQuc
Fi+yKkJS34VvXKqSRiG18ws/Wl6/C4iVQAo3RDfGrAmMQpveXkEHUEg58lhXdc9y
nyiSH3VYxqlAHl38rT3f3Rcj48ud3GimxWTL6AZka+0VYFL5vlHS1tIjySmf1rjT
GDs4Vrbs4ApoTKLIDlE4r6o1Eo0gd1gRACt18z4Y/CF2VfOJP5KTC1giLKf8q9q/
q9S0CxukeklyIiOP2ykMbKtMN1oGwcE03iompXNO0h9ndMYCWjizm4G1H0TPMv8/
63b6MOgQSnsDGz7QdKqLGzoJXZpRZuSBSTyGgt2oPf1ZjMgNhnP4VdMeniI9yQGW
FUlThjOEpfZ7bxPgbEtiIqQM4ac7WectDOr8L2mxn/xYsi6XDyTpV+m75fQ0xBip
km/hxx0KySVeBXZg0xo2pMmikx/B/UbHaAwDjDyJo/gexVSnxt2KoWGMFZwpla2o
Y/HoZxEmLFmHB/cI0msQCEvP8Gl84OZrBHd/PgWyn89osP7IFFkxysHsc+Luhli4
t5bLVqx0qiI/TrVi4XtyxMFVrMgAPm1wXuC3XE1wPpgaIRrmZHywzV0jnXpEG4hE
Y9FiegdKAHkjgoeItwu0D+ov0kH0e9lOwWFZdFKXPLCmG6NTTqJeAz6bcIpO3fYY
YGbZRrzjcGhHq9q+6KjwKlhO/09nLb7mIZ41c1i4Fgzum5eAk02GochpkCynD9ZI
enLvEFl6x/NJK03BYeaM3NWRBWCHYgle9ROBQ/LsrSGpj6FTknR+QUT4nLgS3Ptq
F/i1xjJyqtJQp0B6foe5nwqW0gSlokmNCR20diSEjKylIfkhhU/JhXDseXTU5M/A
iz+V9BWvl6P8OjSD8QmHcQV1fYhhX7yx5OO97M1ZxyT4CaCbpWjpTyAEW0AyaLb2
/TITMOtNSko4HDhF9Yot2UtYzlMbQpo9ayFIbipuK/VndIJVzh6+LxaYgKuXI1aq
dW9cBZUmSUrf8mNBh8dcaIS9obFwo+sU+KvNSQ5dCzhXXiXbdWFbu+IN6rIY6ank
qfG40TVcJF7oyIV1p2laY9V8/PO1kNMZAmhkyWAnJ+k5YAPD5tLRIMHw2oxMGTfr
1sf3LzdcOp/67FYAjfj4ShpJ92UzkWdpB3pD+B839ksUxCNo/2KqzluAz9fBr+ca
KBZo3Dcx+NdJW8HBe8WbYnUcDmffNInGMFZzVp8wzHsTXZ1D86qD8exQEFOTCyVu
Jf4iRLxc01EEuzRtfH4W0wtMMA9PVWoTyinzhn/Gw+KBPTlQxfkrBH5dG11K5Q5m
NGk7KyDF/0UcfMTSB6nan4QdZRtuvvATG6vMTt4NSy7t7nFhYD/qlxqfY/DMM7E5
vnp+lzcBddZ6BouG+GyHBIHSr32dWiF1WkEtz0nudbnilzgKGcAY8JMvUAF8BYrU
hOymiEdkNR25/CBtRzWW5menE0Xrut1RyOa3Wpge2DQTNMY8k1pb5Om1Auxb8Qk4
bCKMpwZOSpD5/lY0rlCqDdWyYX6ZkrQ6Qj4fZEqgQuf++5yacXWFLfQcy5I5mSUb
uXSQAyESJUGAMmCRCuI1M4wNuerxSPPQYYjepH6zgOLsBW5gbSittSnsA5H0tM3r
Txjphe1e53NldnllzM3Qn4/kmG5hocclWfysHTL7sDGgerq6iE8O67kHGVO3dpSj
34GkGS+TNmaOSNlDLgZV57I9ZYejPZSNmLFwHbFKHGGUK+i8oVUUN5S0ZnekZOH/
CLjVXRGRWZw5h5fT4w4e+lyaaz5nI1W/kNL1ZyyI9pfohrIK3sDIoqdCsSfDqv2Q
uc1utoKCeH2VYybfjaaqwl2Jf2lq7+1810KReIDusP+PmF08AbRY8Wm4lCJtLP6E
dG/3Ye9DFvs2wCcBfE6KvTJZ8BMIBwu6/DEELvuAbISVlpmeBVUXVvETYL4623ko
KwbeY2TgQRDV3M8vyGWjYaITbW8LQuk1TViJu8a6JmHEAdjt2dkCzxWXZOBM5KM9
bH6mRj3w2y6+RPpqOTXJnXD+tzsZvgmjdaggAfSb76X/Vuw9C9fXf62bEZiGP3Fi
QTXCI5AQShD18kM29c6eRPaScJ9FnA/iEEfvFjssjgfJecbLXBslX0zHs1LvMBhD
sSf6Mmh2xbj4i0a7N4QGcjKPJ52ymN65EIAiGy6V4JT0TdPNW5JNvDzP5LS9tRGL
mr5wIWfRZu7we3tiOSiVJhGuIQ1NLgOENN+sZDBXU4PuoCAwj0Xz62gTPYRdEsz/
N0fBTeYuIveb2CtdvBsLaw6lTD1ONud8264cD2nMwfiw4xilAWEi9kMlRVlljPiQ
FRGUOPriu1ExlSRR+dI4ZUBtUmJL79y0gdgaroU7yJuw88tc2tpQdwtBwjjg15qL
cWFWxHqHLCJYBrkyxww1s2lKtyyeaY3FXaeuL7YBbuPGwpySBbwDjhS0ca6vRw4m
+Br2dyusEG3IqQilNnUrDVbeElub4B/0mCw0ppp07TsMSrRbrMojVs04478Cvv12
cwFAD45N6ZcY9szxRapjSh4DxDV5iy6szJSTD4ZgFZsb4cY6XxdaZy2e94tIRlxH
OjBipAH0OTvq4Dxxy8u8PMbl2OTi3KpQrQ3wIfUKVT2AT+tpxWdFrojOKa4+BBjP
l5J7an2DNf+OIYtHjvpU3xdfjVoQ4b9Y4Kk8k5um2yCd/kcbjiaQ8YCNFG0rHPM4
m5jK4W4/BhlOmpg8g8C4mf50JtWQESkAMOYoHGcaR/Yq7itHPhT1qM2dIP1tF1vu
yDO+5Ybix7k4bqvh5Os3BkuPrBuifx9IIy7qdnMyKQA5VTg3j0lpQQni8aqZJdaS
YaOwPcOuvNE3iGCaSq5LEfSLYfbxRJxPCzazRv5bLlLq/eOwb/klxygRae0HPjni
4hZTp3ZjXzRIwq9GGbk4JicB0C6pqSKrftV1UbujKMUgOCMxvqVtdRMFTw89HzMD
NSzzhTKFlqk+qW0xBUeWoGHFqZ8ayigRg4W6fgFUcN5yVVSqZn90dp5HLs0ayOtX
KWbHw1M1zhx1uAieNPnhNr6AKkU5xF1q0yuu1EJzF+7dcdUjORmstgSxqHbxYy/n
fJIhLgG72tfhADciqfOWuh+pgybPc9Lply0qKKhKkB7jtYQCUI9RLlO/+eziZ5Je
PG4sx0Y6696tTGx9cmG/XIu1h8YlmFy7CXytf4WtwGzxTZxeb6SVbJv94X4GWphh
I0jaWygBhWJttuxp7B5PACxE8YcT/Uk1zOcBCXBcF9FGq1L7AgMJQ9YpK4XTb/OX
D9ongCvGefAOq7Y/iLx/sillrTXqj2lBj0KDh48UoXu534uLfqmgSgv5bEUU7JMr
FmbHQdg0C99rV1CQwvMqFd+rVFGFzueTwiCk2iKm+anqOp/QUfgpvOTmRk2ACaky
X7GRA2arTyJ2fnDWW5+i+U9isKzmb43Z1pazshQS8N7d8EiGtXgrBQCGnNp6Bad/
dgxUFKpiPLGqYBnYrJTTsa8mQVxSoLZ0V5SWGUEDl+ZWaE1eFvL28CSajJYr6uX2
p3LT2Hc7acT9ICGDygo73yDOAGA3OIo4kcq2V8TDIKtYeAr/HN8iSzgjyRCUJHcO
OmdjjqMHU90DbEw8/gZjZm47EmE3scA+Is8BndUDP/UEmsw3D4ke90hLnM/wccQ7
ijjXIJd3ho2jf/SdyE/Bt1NeEfqZxomVZsSR89rTwuxFG08b+IyH9ff9ArFYgGGM
Bf9k/QRf7npBjrrLABkZyiNr0A1jhJ3qWIoRmbxRuabTTCY8C06Wy5DYa1FSeCWY
vHfFGV1gwg/yf7qHhNgW9ZD/ox3O3JNtbzoJd0k0V6Pz8cy3XiZzkoeYNZwSjWwy
Gw45U5au66vYc7vQnIvD0eHZjX2ZhemvQhStOJugqIhoLdR/iZRWPERM90RSuiLY
bwZnmatwsBAMiUvZy/VQ/0Pp5qc2n9OOtQl2ggL5De7ztNGFwhO5DSNaK4MBA3cO
Om+8Nm+3hYd7hmDgWUrgDdoVpf3vdAhNZljJItH+BC4DTnxLT9dQm33gWxtFJTNA
XrlhH8mSwx3+GzjtLgCRESPitX6T+rxPGqCZW8+qF5I6CbH2JjU0NkuRNFDexb75
qyYWkDEi+6BV0kHRH+BKJnpSP/bjCvFWSqKEdtpcU4rIqJClyRRy1PU40vqSdMBY
ZYze8F62bLyDV3sb57nXAYEIIk4Ap6cJfZaz90Jj1vjb/7hne9b6U2kMfvXLVrKw
BiRI6kt/5KXmrNVsdhNT+sobwTNLMNv5JmG2oDyyTWOnALzzsAmaceAuBrHmvft4
UPk9BvSOat70/PfgQJIylZcMKxYhkpNVBBZNe+nReF4ABdtlUQOpCgB4izQGW/G9
E8yZA3LTVf6tFmB4VEb1Q/N8L9A+BKwRuFiBM8ZCs/wrVECHR1ZDazk7VNz582Pr
n5MfcUjHuQFneBMlQ5R6KfFN5ib1czyu5thE65zlgOlITV0WKwsZx4fVxuRLcpnq
+q0Z4WI9QRzAWLjL4KpiTgh/Lk+xsxC6F24LuNgE8iURoi/WVwhSTos3+hnAtNw7
eHX9qgPNs0VqruUVWg8oTAZPviXxGKJJzeSHNzspz7ViO9p54pncb0Bb5Eu2VCKx
7ra7R37PjjKcxc860Mmf36KuUve8hP/8JeQMNO7B1tsTPO4LP9cdC9quL0OYrnMC
cbW+4hCjjcC0NlF076KLfItYaZgq74tUvi4h90O+MjcNHe4fC1Vyw4MPEjPepvfP
FNQglBLFt9hy5dqvUjGgO+5Jmi5HpGPzUaItHtU39b0YztUHHLTflfvw1UQ7qDdi
qZT0s51fMZK+x6nClXV/ceFiLIXOFZp2WP+2rmH2bT0yVEnxVSSoYKNN2ateJ5lW
zB5sLZB4HoFW+jQ6RTyKLuxIrJcAV68p4WXBhZFhlRWiwPO1wseDQQSrot4ccNig
G9hShn0AjcKnKLAQRTfmEMzNUSZ3hL2hpFx6zTVpQCV9d6AXT6X8V3B/abpOItYy
0y5vQC8pRu6U1UqIClcb78zZKP40S3g50VpIiktpvL20PnbD0KXjxBfCay8SPVmZ
UXlYVp9UIqsyIqBHllKhuLdORhqQJ2oXoEHGs43gB1NZvEt0ChSBTxanGwstdXpF
DlMNyxHn6OMys9kp23Grk2/iEpGgSAdChOfUfbd7mwh7gNywNXWalY0CvNFGeFAY
0xODTnt5eGDejWM1R2H+ijbLJnOMEYeOb4C+SiEg1MD2SElFArs2oY6cxy9Atajr
fgWXqqmSGAR/RtilvehKACyKYe1vyAVa+MecjfP2ROd8ik6smJP8YZnkEZgSWI9l
Ep4wqaAOVpitr/cpbJ4kkdDy0zFJVcTCkMqDxeHrjbFw0jLV1w8Li8tmt+wsbm+y
fWqKStaEOOlrKSm8Z00CoQaK+m0AbyrlsmwIlEci4YTmBfWsEWdblyi4ohPYIPSe
UKtmtLREMtobAWfUuFeaf52ie/ysevTld245L3PIhfRnYwdjd8bvtLhSx3xDadEB
VOVCaOQYr2sl6IhgO/xUeNSEHMGSdsGRx09RQvtZATRJ6x4vuppatI82/sJlXGTl
tCh8Djj1YJII0M213UZi+8UHB4diGtXNv6Yb4XbXYfD61swlJtNjcgX6ypl8C8av
FVDChIYX6Hlm7eWrvdXob/SwpN/TIrLSdwA+LcXWqBD+wOgUoC6U21FEdi5ZxpNn
9pkm+QK3zHCe0mqV0yznj2GEUT3Yv6OxCGXyy8qkG1QODjb5XdGbNIEmLNoEK9L+
U4mMmyJLzZjx8hEfQ/yzeWLcSi9jcmHRi4+0qaCqmBy1UnF8qspwRlBm/curGWxh
sgGWBYSKlGCEC7tq0c54SaYiZl6Rd8BQPMnj6BeCBo6hfGNobmCUhGnAwWC/U2eO
uvrWNpK8MrQS9LMcLzn6z8I7YZG03R1OD5tcZNPhBOBIGXFz6jVkn8+yyqcqsfKA
Zgpha25T3ZBGcaWHVr3Gd2Ytm+vC46p9RnM3vYTPtLti+iq+aN4j9qSebGQwYHvx
pjgpT7PGHlVmT90s77K+VErPZd3a62zscLjl5IWCZKzPkBnpZ79+IpnWNGDXb1F4
/xs/WbMWtGzyKjjRXp3Srx2/e6cODpdElMo4/8fzBV03XiqIU5ysngJ51iWEleZW
UQ44pCOj/l1fbFQrJul2/nOEbU5Gw1+73BMndgNCNwwfTGuoSS41hOc5BgdL+TLa
ZFpdMfaGsBZSnXSQ8bKhXvPO9w9HFFa9aPGxLNnsnpYip0HpUXEXd7/LtWtxHvb4
7KcQaEvSz8bApu1JCfJuXnfVSnojKiT7MA9+7GSNJ/yjLuTOD0xxC8yjgeYSShg9
L7FM6QXmPk0O/J4PUgX+P0LRozYEYHCjOmHuqQiFuUdzF1NfzULwxVnMO0SM/mYz
tPdE92m9AKkDzZcOXOCu7XngvmiQTXhAgNJgJhe20j0JNVqSVQnyDWjjENBqLMtW
Smz3MXNGRmPMoSAJr1AEvmEya+eohoK+aSLbqG8F5h6hCw71Or5atGjkcxPmr8bV
fmJySKoBn+jpxq01NJNwS7vY6nu4XCVIz/Lule+Z+DzXovbz2glEXhGJ19NMYch7
SJUXAOHrvDIjfUrZW372c4v+TLP5+YfgkBHCyBvJFPRm7WGDP0pG7Xm3eZUtSxR4
Zq/dDsEgUNr0shqfHhEYxJJYCEf/IgZwz0lkVnp5j0VeEO8IUMTCjpxnG/dJntiy
7syCmcmIFJb5w4c8zVOmpsYwBdmI1llzwkz74ypvZI/WxC/H316B93dt5gqsYEno
a7fycQLrY78M/njN6U51Q5G0hhaxfWOklNWcokK27DqhheK9kzBbD7VYH2NvsWOm
h4bAubPZZ5sTSV32mRVqIdNQ8wW47uXTju+kYGfNabshiZ0BVBj5PYZ17Vr3jdUo
r2CIg1kXwsfoAr6ElwEutEHyY00BKjBVTNLcrCC36C+QXXmRT/xNvLxCKa/Vb4A0
o0AFTiG3flOX7UaRDQ4LsEOHb+R3O5Js01S2HhLNi+hjgAY0PD031nJxUv2o0T5S
83Ve1NhF7Se39/HmQWz0tojgxJvvAPrTJBsF8SZM8FWpXrnPFNMlmZJtsHlb15Iu
eHyfkUARCZRq2m5VZ24pXpTEfkUD2YmIFb2ikLVn3q1E3KltAzu1lmPrwmxfWga9
0kXWysYw/W0s9YKU+oyOcywK0cPXbGA6fV0e66cDgiLpoSjPG3T0/wY/vF8GqzOd
p2rOBHqChpPtfBSwr/0+9Wyf4UlxKIFfVCIj8ZUvHoAdTpAk/dytqTuW6Eocpcjs
/0BRdkk+KEKEsU9qIK6/JkBfXNdS8APRnx1DNvoNrgh/bBbG8wS/1BtvBb1OYEZJ
Xez9BrQFxwj4pHw+/NEjLqKChOtkcP4+typcrCRGtRLIPuURqOiXYmSwH11dI3K3
ay9eJPRU3XHNrbGCVT1o39JnCFjW4cWFpoXflM1219ivRSv9rcjOqQWN/L2BVM7o
ET5Jx+f10G9uhxTVw2XcsXxKN4GEzlpupJLfTzKcJ2KV76NxQhaH6EWUPpFh0g3v
tN3rKnJrMPEAa5vi630tFihwyxYG909p5Of3hfujoHO0aHGzmE8XHO6bdxBA6rjR
mCCCmwIVjJFV1pXWH2IkTe9NsON73sc8s/KAxY1Xrufal+OIlm/3SFtmhyy5FQ8v
a2ubmERMPWFupsrA9yAgwlAa9KkznUEKrwWPdt7atMME+eguGmwJnuJ44Urx/rbr
8ESwpTgBLptfIG8X6hDv0MdMZqaGCHN9bSW4hp349Tc6GYwSvaP75OJcvoaq5cVT
miGjmv+f2BYuqo6z/L7toTwb1EnXP5//M5BTYKJrTndvIpfqk4A3U8djB0OOhMl9
ax33Iwat9Cn3V7ngqSYwkrDcSuUapBVKdVPrBEvY64krX6+sxLGoqEufPUtK8OjU
PT9iUXWN1Uu9KnRifvlgKzz5qHVsNjXX9ABrH5DM/IaVNLlmXwWspkjdimLUIwTm
LnRgwxwGvun2+1b+ATHm9ZbMJV2mACtX4nD1NvaHBVVxITe4eYkafjXj1ndp6kRc
gKowKhzMn+9twrJTiWtqjBrFAV0T0m58Xirau8PsJR0j/BV87qQJMUA3UE6uylVD
188xaHW0eXlq8juJ6lk6JJCEI/vknjfnEyozyq5RwfT7+vLFCbIav2ogDgT9t29m
vO2PojyeUbWIMGTKdQUQzRD4DnBS8DnoUTOqtRJHzVQmhxUH09pIhM8w/xQfxhMB
KqmFQ+TqHFFa0a6YcLuTnISYgLCFnAd/rBWWHmmgOsJOD2A/oeVviey2y7Ilf9cB
eejm41/aZGXAIkWPAZoBc1rof63rzf3h1A4zzHNYsPHdBjWs07+zmDldD3AOW/9x
g6lVAXZSE8zDRemoYeE2M5aKkTVvZ6QJkDUsb+ZtUp5yQPm+GGNlGO9Ebve7wnel
1fxdlvujrUeDq40ObBUQ8ogaTeEy8MGXT6Zjshx2UAPjUMhp6NhaKfyMKVxK6bTv
k7XshAfbCehJ8MI6g3RwsipasxOOgtvQRSx8D2Hmby8np4QjrsfY8Gf/3Mb4AZTM
NNBWsFzevkD6djZR5MErbm77UClqyyGDc8X8OzAU4GNNdtLZ2LcC8onXoQ6EPRFD
XtloyGFB0SejegrRmuP4/RwAlqgLm42vQmoAHWAO+H0S+W0pqmUOErt+MnlhWdv8
ivo6Tb/vzHrSjxYWmO5ChjIXylPJs9ZjKa5w9AH0HpWpK3NB5wAjPecDT/vMF4a1
93FiuDkozhwYNdSpmwU4Z3U9DLbb2T72Ugga/gnz8aZukd2UKw46V9vby+TFL/bU
KfnfJPdylOfGt0qQXWmX+o44h746Nx1qA8DEhTITxbdFtVrp52/olp1VQHP/+OJ/
fi2V9GdhCdP34OBfynyjChdA5zaseQUwmGjfKJN4AH4HUN89r3Cc6IPsW1WVqG3v
bvg3uY68WNYHkSTB/i/Xkyb5SN0ddxDISZ5jnXzGbHL72QikLyxVijzeNkCfVlj6
G0SD+G07ylHv8gGAQahNUxsviKQaSL49LovqjV1D0FOE7TVWBiGQXTbYUhAy07fQ
EsnF8/wxl4S4mgnSOyX8dXsS5A+Go/IQSPQE4kBM2ra9MMmAKahxaL9zPXwhCqTo
7ibqzzrqtIHbLu1A+cCrwyT2Nxxe+EY0P/jwKWzYa+Uls3GCoWURuMGMXNFfHIJp
ND7O5kgZJO+/WoJ0k3Lx/GY2ip4dNOeif+poYQCr5Ho3apPpA+CFN2vFQ2aG7E1M
QM40IId98DCA1+8S4M4YxWnX2TUFj7pIAub2PF7CdySXXmHgcdxRoHva0EC02wth
W2Q2OJJVyDDfZU9o5vHUoOvza/KJuv20CkkHls8ToifN8anY/tFSSkcaaX5LvjFw
VFoYT0PV0BWpIyD+HfUYC1diPto8Cluch8NbOJ9QdGP5dtj55FFt87NAFZbgNnQr
gv6RPDaGtE1SbqR9gnjq3SRdszPNj7KeH1NYH8Ufb0bAsa0qOMFf6kdPHB/V+rSR
qA7yZJzk9u2aliXYM1snRDUVOi707hKoeIhWuRKGfvJiLGW2i//KxqucL03n5YJx
Xj2vjfywTGGDqugz6MeWP+m4iFPFkRjw6JGPg4iVW0iaQzD/BWd1INEscxgLnDDD
DiHjN+aP+9jsvUDElBWqhXA2vBsDf8CQf61meQT0Ai6yOejqAhpQ3ZhIl8bFvC1y
zie56GYo9HEPfFa0QTmCSQ8RYRzlsa2rTgVKeRSYy6i1rRcYox4oHkVy7jQD0euB
63ec+G143t3bxcJEch0WcmxLxL/mT6R7y/YSS1VCC1psDNPu071mBhM7AZwK9pQ1
mwysOb96iuGyJwErFKhyvivswK2fvAIwyVshe/TKMhs=
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
nwWUnV0SVhZlilONIflr7+9BgeYWMbRXKOn3NuckRehkFsjlE86goy9lPqF798eyan+7h2d7y098
Nymt572jQxZgiC59UNbUkAQ+FH9nhGZkWOh4k0xuVJBdcwISF8Hz3G//BFkIQsoIb72z3aayh6Gt
XDksLsFBXgeIzbTSp8vYabLp/USFac9UrgCqeQLz+vHpB4b5goL6ktjd1c2Mx4xvxAqhWv5wYIpG
WEgpnnqN2pfhIDEe9hNR5ysqJZ1igd0LPR3Y5g0ReiWpPeeRKovh/g+o1MO+V23dpc4Vo0x70tBH
LZUrqL0d983ymZ35CvWP9fqh5QO3QYnh8CDjYQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 4976)
tvlFzw5LPg3qbfhvcCvtEgCdQbmlRRHgSjpHyjOKYs2zFYY7gZLcbMfviB5IQ4XEaQ1I3IN5O1jP
TqFAjizEgy5FKxlWe59GadN3HBmOrdVzE197jU3PFGVehWYQpiFiX/GrcuegpVruJ15D6Uw8V0/N
AiRMkDbFU0+IErDE7PJP7PMlJTa00QWUqEIeApU5v83BlY38uQ+1qNzHJNUXBVvnDemSHsTm0DxC
rcVJUFFFGUCafsep47Hw7Im1GLD4HoppUfA+cGnHC6/frUR9oQHd9/4GLriaaJk/4+85tJ/i/Qwh
zhZW79q78q/PAXnxlK6V6DkeW6MuycGHodNdVUvkQ6gn6YgDBr/qAfcCv+0UuSy4C7DhDg92Gu5U
bP0TeDbLc62jmapRxRGUOGSgiB1goBQ2e6Ap/za+UhwTFV+gCaTdGXUqQoyxnHBRy+s+aGXKSqKb
h1z7ouTbAN60Rt5fopidDhpR2+SAnZWnNgefOhbTF8gCXJ7Iac+kUUqEN4smc2WAuWJXNM2T17Jh
c0UlPaZOFl5rq2KczE2VK/TnpNcEF0Wo1t++IYD2eHI68y7NFsSTxSOYWO1HSxXnXbpRDdI3fi9p
kX6PffFrIHoZCCP3s2ZSNSRycdhey0lNe138oTQgTiS7TQ4PsLGb5EjNRm7coTQCRk3EB8S1SVqL
esg+ekFZfH1Ya0MSZ6MrpeQZJqODi0/rrqKuw39W+TBd7xbn5JA4aTEXtiN8TINzEZun+/Htwyto
rtF6ARlzGCQSehD/gIqqgctPIYyjfS58jT7Jla8mRm1nuHfqQiKOIfM9Ck9025Ghq8GXNzRMAi7o
Tdxt5vYm3EYnCA1Mti81m2WMAzPVM+N0uLKn1rKv0bMcHoO1/P94qnPDS80BSFhv270bHhIw3rBh
lyt6RjX6bx03Ie/lD++jESjV+mEUp/dTsK/jgzg8/BI5UQywZpLjoL0H0U6jasK3U9i8z9zYrpIB
pDPdzLcymm/WJEGYCu3vV67p1bjcaQ6Ppg0hR/GtDeetJIWsYD8iB1IcwayanFQ5gZ/oYy5PbefU
ucvlr6Ew4AtnXLw71zq+gGJNpgoEdAsLTzfXbeIxhumc5knpYNEKIjblnS75JM3/JhctoVjPeQjm
S+x95C702LCgVlqRhUkV0Htfv193/LZGwXvuypEjo02FT+/mUXinqX6ntXS8hhzyZmjrUjGfBEvC
APjnSeRxvX2fhGGPUs7DHIUuGrZQy2rd1yvBYK/SB7AerJaKqiTo3nP5EYRR8D1BnustYBBGdzu1
uIuxRwVOWTerWSpxSk5CWWDvTjjMRxROtajvbRgMyl49Wm+YNDPlp8LHRjrJ/L1EGkPYVFvPc7Bv
kianz7LOpPjFtKt3t1baEQzKC8EeFjc9outFmYxADk3tVMJnrYrS0QPaK4u74Y6K+ce4wVN1WhHD
/erdwck+y+6n2nUJkF4jHdy/mJ+zSwvPseVgXqy6DAFhJpqHlu6pDJ/+AzdNWUYQjabRtf7xUuvh
4tKyXP7Li+R907viNKlLysilHX8cMBTREyNYBQkpsWUdkxYdZWqamjbVAGPIH3trzTv5JObmZTZ+
t4kUsVMqVcdeafuF70vDg75FikY7EGNgTmuCpHYXs8fXsdG3pt/uVnN+yOpXQCxqKz6f94qqy2qV
j3HfuO5CGcz2c05cHQTymIQR7SQPLEUZnmu8EqEk4MsJdxWiU9anBppVMgyF0SfPQfY1M/XcOghF
LIZ9u8RfstFv6KNapTF29sEhKQHg/8nZSD+DjA3GbL27MyKahBpEQdMCm5/CPASl228qcVw2LL5I
U4sVAa22mdn3XjOkRtiv5POKU3p1nVTYjWduTLdgpWrBwC+LwBNYKQqvBBuJ26uADn/ptF5B/Ssl
nqGr7n7EefzjyarvVA/XagzaRje+EQ5xVQ816BLDFGwI3Wn1D5Iu9dJ11C1wD+6c6b4rcfAeyNQW
wct2sy7CUxF6x1qvcvxg/C2LkD9FOVtjvqSQ7xalj7rPFx1PMJxfshG67IwFtHNYOvTZ7DC/bw3z
Iz2Z6ddZJbyGPOXTtXYgd+muynsL7eBoCBgS7FSNn1XMevHpkpzJ5sz+5YhtlW6PWjhj0FMvaEXO
w5HRegvaKnk7uZ4y4iV52TieEoRpvERhujLgNkMdw4wneXf0CKDQVR+5s3rg+RSDQXMQ+1Kjhquy
gsX1d3VkgiQrNpyfXdu6YIBm06bkYEh44u9Q2Q7L0sFVW0C6utn9e8gkwnRy+R+0sVBK1B4QQZgT
8q6FeFBkCa7LUluGrtwkTC3bQp88d7EsQsrH1WuLxUY5T1HCY2f1Op1Xuqeb+p9iEUqbf1MsiraC
VVS8dDpvSfKT0vbsE/zTXZ733tbUWLG8sOzdPGRLlFpB9G/jqWKFZCzxFSjxC4Yx/spBE1F1j3Ka
SmOkXoNQyA6S/RhuPAaRp8vKR9A5dXQsMZp6Wf8ibyDSXTeCffEQKiMT+QCyWwwWNnMQIwXy7YX7
CbppT6T3Bkjl9hdA5LLd78NiqprB7Shb1p1fmUM6yJ3OsIQ1uUwtJosAh6JGIypPzqGiANp3eFOM
dw9vTAJpofI+nBSCw9S+PmjLZvHGaINCVmmEYbvoFmoK5jwt8zFlQmIQeRpEcJpRG+XggoKjkR9m
ESdXnkRoeHwi7m1vSpYWYPIHrLW3vWAhMcA4hh0t1uBrlCnpw0g0+WrjZ8tE7ozjNGGYCAGUVyao
pAmjoKGzLmOqny70IGHOAtibcDo1IJcQ/QFqZBccTuTt21ZrZUqZrKF1LSrRIMtGxFJJXK/PtOdG
1k9+Rhc1U5RWUTKWjV5yQpyqKdB7sOyJ5c8JgYHIqF74RHZdWelgKWGo1nsztspaIszYtm7Kl8DT
Zc//nTuJq189rcuFFlKyMsQetAlp4986dwqzP0AEkwS6oD2UsBzvqx3vGZ7deib3rBcrnKpsqA0G
zpvKUyNEQ+8U3gxzYMy4ohfPvv5QATw47b/Y4tV5nkV2CgySRM0OV5noyri+x8n2gtcDcDT8Jozv
P/a+HgYXfeOVtSwhqCnU3TCQUNZHQpcUV61b9stDq9/9YM7sdffka9qI8aNYFaOLJP6orkwkWUMA
neUEm3h08iPJJfdZQNDTrWF3600K2s4uB4rDs1Lhv/Zu+f7W8w/ouhIfve8KL6ZbWOa6+JCWkI0l
WEbd8CqyAzujK1Qbr39loWGUhu/AyZWmUVoy2uaXIUmv/HRz+WhH1drP5E7pnJfZ8bBMavhKnwRC
zEEyxvSK4SBtWfNB20kPNo9XI23U/LVmVybMh/jk/sYO7bTzCxKgRDCpHcWEfe7Ebfc1qZJOdTfC
whZA1qXeU0q1/SCX48ySPSb6n05s3HiP0gvee3p8YZZQ1agAxlk1TYHRPoHERQ1JtKzNWz2RDUsO
UWIVXsuYwVrFdx7ZxtrJiQjEUfixRktSHtIosv1sYnqSQplhqm+lHFFRYpOKlHJs6WB1vk0FtGOR
KN8h88qZaYh+V2o6rKRrXRyBwGiBvmhWrrNMKyz0LFTaekZ3go31V0+ALPUjJlZXOhfazf0rwrRj
bL4aTUBUNuecu9WkIqiHBScK43Sm484FbmZ+1EpVLgoeTbKS0gZbGPw+N+l/eDe7Ihh4qEo19Nzo
X4mm3adx/XxKH54hOqHuxmhtq1g1WfyYu7w5GVaNGZrmpbjJgMBxMPMkI02Eo1fMcqY57mPRZBmG
NpyxVZAQUr8GLsted3OrINLFKUYTv86q1763lqIQPu52Q7jMz24LM0GaKwVuA7ZHG8OEvltg79ZZ
tRJqdq9wiVMOBjd0b3Ew6QyPBE8uj+sB+I+r+bWS/51B7WhReyH3pck03A7o8nnXlyNSJGAcbHxK
K19qndjYoY5vg3bb2KyOIxo7q1JxUPMUycHlTNaWxMXgOUzsvsvi+U9O3E3BNdjXOoucj3wSromE
x/l4JdNdfl1NsI9k3gNr3rzWXyVIn6nnBPT+HO+6UYbXJRc6fYpuM6bXwEGHrAkvHwfNsGMqqo34
FrJHr7FUccxsQeyVAC2GnM1moMAVyhq4Z4uf+bQfhuG0PetMC97fsCH83KCio9wauXFzni8KVdvd
5CzPfl+ne+AwhUgFo8jSJbKYcsAdFImaMxLhHtKsqjPu08zO7klK97BA7EoI4eghnWJ4t+7LsnK9
OXk9sE4oXBwMBOSKzqpuZq+Rj3kew6DbYTRy6BwJOJucDMOKHaOc5Equu03bTkI235y1Qc4lN9IJ
MQ7C76TTyl1jjPB685bj/nk2a3HJ6Jfcb+b6NwiOFO9924mDaqRY+SsEChcTOMz2GFXvKvzgPVfX
pq7S7EU1hql9uIgznrj+dsCsEVFi1205AP2V8ZXRIoD0xAKaN5fyaU2Qkgz1b5rSeShCreMsD814
ZlcOJxv9lQw6x8K2/g0hqwk5ekQ/+anVSWFNo1462iel1mOWea1fpftifJVuXeBZnjU+EudG3sDH
GgUp6CbRzC/I1VzdoIUTwI1gECY7NtYeLcxJ7dkzVn7oi5+XswB8CNDPRpHO6wj5o8vBQ5qcHICZ
naw0PdATMte3Yco+d5mOcypebd1q5wt3nYlLGsGJDJzcoGFrqa+0mkm3AVECJgU+Uloqj7PXZJfT
LI9lUQ+3/f4AR9qMBc9PzyhRug5PDTiiB7SN2/HJwv7FaFKfQp8B++JBAAITuLq3XQiUMSzukxk3
UY7PPBIduyTU30Y3aiMHZ5mRftjgac5O/qT9/kNDhRGf2MQlUAxiX3vfEMCnKPJDvI93wP0VyzZ+
phkCtUiReq5XlemTTmaDUjztswvHLk8vFQ4Rx+KAdihzQUxIupZXUakAHezctf4ox212vnQNByFE
2ujXdTNN7vCoMOUu/aananlWgpKqC3Bwhgagq8iP8yYjPsoxwT1IAqhGswX3dNeI88tfOTIUCAAk
Z2ZPQCOeVskAOBEaD+iALxVlyTX+vuDnjFNBqX/LH8vVy+KwxxGGUnKBvZ2jVzpCMw0a8uC0d8su
R85ytvqMWg3DkuA+rSKuEYl+iblhoBGLByTDJ4Bgug7HACujRQu2AotElEZi6ZwPgPzr5vJ6KuYm
vB4MaQsCcLEzSooxHicqmDn91NwVs6Hb118GjBFQGnF8ElMUB21xL/1WQmy8BfRqCdcG6NJsDQu5
eWmr1jzMvJYWW3NH/bfTcfIXO773rv+oDyuMsblrms/mnDhiM4/vfEzMJ5nV0LmnX0jsJB1WrEGD
x0iYY0otgKt+ORdM8EpCNh930ExIxm6qTe1ybxQ9EtXzvB52JwEvfkFmNzubwQh06IswNmGXUfy1
YUieI2BAddf4p5Y9sFdRU3QK2I3wZJxWiB1hs++ymtcA9w1z7iYpNM+iN3sBlWkDfn/YtjNGDhPb
4J+xsd7QQVoeakHIw07Cl9FHZzLP0pvblYM5B7JHTtycRStaHxVD+7Jsyyp/WB8V98+rWA2EpVAe
amLiM9j8hx1T2vw7Rp5j8ytnEM26gaoM7uTuqtGLwwRjP0WmhwPwU/w9FlEG1dRIdC4bDKo24n5v
WQs9KXlCUpXTu54t/bXVeC/XExSHckMvwUm7LHLqmzrcX05UvMg0ox1H+7PXvcMMvH4xfQyQRN1U
88zIRifRdu1h02prXeRb4RZFtRq4uPklKXZHBs7+cmDdRO/fh5GUHEu0igI6ULiFBku6WKCPD7G3
Fyw5CebYAK/hJX91AdBJARKdGLmkpuTcESU+X/eiK4mpFM6YOEhZR6rzYyscNo97ylP24HWucvBW
WtzrLdTP8Ldv5xr/tM20n8o4DO/za6pvh0fgaTTfnfPTGrd8Cn4tBDGAAqiog6y7KTmWizK535O8
4V7TwTEbfjro6C/6YCjQogz7ul6WX0q4CzqU3wZYP8i/LcxErk6kiqGxn5bWfb7yalOK9suQVznB
4pOhzwjACil4z83xClcTDFoiNWHMdT0q98xDuV27wazmw7oHECAgCOBjIqZf4jmIxJzyQW5GrIsC
yvfzL8JyL++pt2HKnCRtjvgHsuZOzOeZ23oE5kFsUh/CcqCeoc5wR164rJZTon3hzXWkIJo/MGdq
Q8YNdsM00EhkAwGOQK5xg6h+xiMoVFd+w1zM3UJqW/ac8lUpQLc5t2zUgzPcAnkC0IaE0w3Xq/Dd
LuXUeCST5Uq1Yaufn8Pyoz1qJEC654i6aTqTpzgAKRwQYjSmitSRYEJZ2nwtupf8QQDKHnX8Sk0/
lA80k8kjLC5y1FMidi/snki08DEt85lTeHKATNhqLUHk6sCPDf/XtZryQFlMeirVUVyyATlthU4o
bZ5OzM86wuOB1/lYdlZr7CWlIbbCSJ0ATZtzMUbiZUmdTRKup1MvJ4ov3ZK9V2LhMkf1mqOFMDXW
AZTC7u+/fUNuH9s1LOfWj0Vn/f1zjl0MWJ05/NK5lC+I5ndW7Hir8Q6qFzx7E1JXgWoKkl7SNY0i
YKbeqftXMXLdhhmtQigDvp5D9zPMdFDIfBRxX6M8vcGjNTnZMsTCJDy4IQLFuKIZATHzpTI7G4Pw
Xdo62Yv7EaBDL7YSIbtJvctFPtenHmJf4biRx2oSc5kmHo0q10Y4t6i3bzPD0jH6rJ7YfmUy4hdz
fM0MIVgi1kruZdwHDGaqsd4=
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
naA5rAFfAp43yKvC7DpoSs69MkVva8rPYAqK6iWNWK2cfFwQx2xjqkVUxS3WjEK1vAxHEkE4L6/f
W06oCi8qyQySI8Igi0EMcA7imdgTPQJPTRycGkNvELNbw334NpeKjr88pwSTmj6f6cHsc2cOrbSo
ZWuv/ckei7LMFbcMR0YaFht6g42CGNo1SF2jdE0EOZK4poAdY4poggNK0pPKw76OX1rRZHHz6j2L
rsy1BOCphANsoavOwJq9fvRcF5jwgqtyyu33J1H+iQRW3LRfeeRckZ1pElCukcjvCuGvcskhtELs
0pPQfcbTzAf83u0p3jKLVY8Wviw10vqdcpGANg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 2320)
fEwnrwk1ZiVCCeQ5TwCBHkfHQvyO9G49bTV4etEAN4KBNKAiRI5gbSyUrfzWmgHrQLcTfRWEOuH8
h1m3dN74+1E4E+/XiwDA+RRUIJnXao5ELu9YDAu01JKajxgln1x+65geSYyq0fVkF1Qrmy2KLBdN
RYeQMUmYQFRuQFdQ3/WH5q0ZEAPaCIsRpxEf5mqWs+aQFAeGFfK50zAYF10HFNoDZDNlbu3MHMWh
OREJZ2vn4oR9Zy10nMLcMrCLCyGRH7pzwVAcx6Fexq4Vg8+bn759yKGSbCTFsB2vjzxVN1GzM0UV
EliDORmY3Rz/DFECjpG0S41c4J79jC5HmIhlsn5M8Ukr7Z2ENF7om4unW2mRPmlaEQE0xGhNUoo1
UDw8FAT6JI8guKDMoZi05hyNf+HYbHtwLZCjJJOtuW/tKnnoIQ1ptNCT1hLUXEBYOdSUsu++TNv6
NIrss5g+2cq4F12wsYXCksuETLtwkbxVbCqm5m9C63Ytd7w62QwVdFgJ8eN9W1dxeQ/AFKC66c0U
w9g155oJZt0LidrKDZQ7FXebIyiPS47WFTHVHTjZcFOKz6dLGl+VhHK9ONOYjFUmYLiOSTqvGOwL
0pH4tgeOCS18s57eJ9OHeVXylFmAuhXzSVwhn6NCUeYiFFTdg/6aN6Hxrul3/97IRgXujsQG6LTU
C3Hp1n1G6EFZvAR+yKjhHDpZlD3tAFnqmzx4NR7XP6ADnhGBakIi79yEXvVCJ8jGUZjWlgaKtCt4
vBxQKanDhDuO6Z9Bv07/c8B8bA8ixzrDCMJaOVDtF1yBZJxskrrXss1/46D/OAMaVT2+Nzyo+zIV
qdMhiWDaiofQ3aWzPMb+oaRJTei0H12zE9HS9RgngkrnkWyECdqty07x8UEfgmgi8tIRUsDe+Xc3
jVxeMsihapg2ls1R8/mbAKsfevzSiDNWlsIliwFI0E1ixHlqpJzMXDDQhUDyOVsRRrQ6lZrrq7Cc
jql5yQh89LDQxnMrScMgIpWfNWwG6XnOPcfy4jrLCGbWEgnm2o7N0PMb32rcqEsPym7CtZsXUaTu
XO2DQYrVOz5b6L5x7F4PmPx9PBxGuU0+vyNOsP+tEyPzeerRhdSkC77kZXQf6MGtNkFK4oG25B8a
a8udBvSbZMrTGkwMTl8ofQQTPKMGz67ZxrwuxBxZ2kmsTmWPhPQaPpILc8v5SEfwXh9Xgd2olLA8
w/dCQDlUqSuUvao0qjZ4KqDuwiul7AW4THQ0MNNZf55URErsRj0u6V2XeQUf65231fM+h/d1WAtw
ntyZuVTlvb4LJLXfQy8ESt/ez0GjwgMCoAsziMYSMDXVq9Yz3Vul+wVBEp5B4R2pq8Up6tO3ucnc
7KQ/igZGHt+26eE+QIaYBME8d+F26lzgiVUwUxHUhgzP3EtGFZy8rWH9RxcbQr2CFnK5Ru+f9nDn
FTEVAb+yMVoAKJa4zVtHeD/tL/fKDRZJmZyFqWA71t2Ir/oZx+qTvIn2kVPBby8mdPfWLZmjE5gS
xzHUeKmvKdaP8Rd6g542J3g1ul3D/IC2A0aqyJoelNwutjw0FwzwgQRuMy4g6OhNwQAS4/i93Oa6
Q4Jb0Jsba726udjhirxTu8pgGDN0so2v7R4lu5qIrU+f20PaeD6+YGZEqg9pXPyzD3poW3IVsRiw
8LsyKZVROq7FoGDFR9TWie6bo/YMWysDiyhJn/YI6feeqZwq+pvcCnbfk/NlOoP9b/MNGwS4JD9x
cFFwr+m/JHlhxRTS6qZi9SVTAfXgfRsIRcyZ5AUzdj5VtbRoByb5inmIh/vRrd/YA8E1Z2QkWNqv
Kz+gi2DpjA7tQWEUpbYd3GhOFYtDWoCCCORl9uqA8s6qQH4ftxiIj1+V7pjwJountYOdb+9MsWu+
MYmly47S+gAH760cvNR3pgUsGfifkOgUBEaCKOunvhYysf0tBuOaGLImK7Yx1C5KxbZO4zkEW92h
+54L1UWGymDpJRx4AAjq2guZJUwcW1wFyMq41RA0tUA6A1QlThksuLjB208GsYwlUWCj6jT64bYf
ZN/5+UokPZeWoasvpcM9CJ3lBPK/A3m4lCEwHc1wGspHAPUm5pIMIBqyhvMjrZcQNdj4gV2+Nl4Y
+tIfOAabC5JESG3Bm26/O3//sHR1cwjSejSe/z905d2bAfRkkwAf2UB6qEQnFh3PYtYbdzKkUwbh
qHRx26LEVouz4XMkcwyy2IGVg9RmA6Qm1QDV6Ge29y2bxh3mQJ1ZyE+DuYkD1wAYXm23V1KFfmrd
BbcLxehAjemDFIn7LTeHx7gbNwY80jfpLHuOIzYLkfN2RiUKzsAg5ph3PxFJVWgjyOSAqMWT55B6
fCHogLWGo58b7Dxu5nzRYhRWXWBcsOQPCLd6QPglWUCb0oJaXQSC7aDMYi1UwnLNFS2X9RMUxmHU
AY0RrUGPvw0wvxMjBZqadicyWtnybTtXwqEHD5qMoVXre+xqSV+W6ln43lDK46MGljmLdu6IAiCF
tgoTkYL9gJIjAU3W+t65HX6GrkjA4q+FV+fkwdF9c4dkXF2tri9OiMhMl49+9ZQxSCXDuQhvYWtm
mtlYbapCRyru4XXWYNDJ9diqodsGgfAPBhB0pgm9MrA093tUkQ3pPlGoDBPzmlpGQCW2dwVwxggJ
MtJoiGcT+F/qinkJtzBeaAnFG+ZP/wHBrrzIcSpQsbHiuqbDmUrGAn8kOK4lvN2o4QC8SO8HZFlU
jQTXvuupVqL3mdPo3+XXv0Z+Mj7ZULQt/f60GltZOxaiDyoOWvzJj3rilBEyjEf02JnCyIH46n/T
H3SQ19t6TFITAGTOPVmWV0jx9xN3l9LVIM08PbNlM/C2Xzxgylhl40LTTy419qMQzKdiK6Ndr9ER
igE/n0bCzlAVS14XmziP27qKbe0uNDyEhAgUuIdG/ixlFjl1dSBo2SyNwARonoI2dk7NC5GaepV6
lFEbR9JV7CI6X4sMqQpyGuJikN6nZyyu8a40ZGpogofs2OE/mXh/jYF1EN/duqa3iRlIL7AuXRtY
QkHFZapiSTS6wvuQzI+kq44szDyHfgJjJUOz7+KzuD6bqqBV3RflQw==
`pragma protect end_protected

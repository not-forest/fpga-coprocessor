// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
zyuXLw1kdBwb6wKckHY9rniBM0VAw/DcKI60G/lq9ZVprulH1heJHoTNyY0rK5qP
T8ZfYXe49pXoEmv2SJ5ry/joP1tRhKLN9iYj1j2Z9hXd4zFH2U8rGaSQ9trFYJkK
52m4tjYXTWxGnTuiX4K0kvQJsUVguoNE8SwWIgn3Mjc=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 4976 )
`pragma protect data_block
FfSzzMk5c/hDaaOo/cbPK3YpgPOjX3cO4QGgMtaDv+R92W9mTG6bzJSnwNkLADlD
AqmWvxS+GH3oicoYu82zGfjrv56LMLTK2f3dFyV/I4XoCxCCOEGnXo0MnK9KqowI
rfXqFxjOOgH1tcF075F/hOpM94dQFATYFckombvZSofhmryI5wQYRHY8i33swpVP
rVvgESbU8LL5Qslrbdr1XDqsHZNuLrpSSL1KGXsJySzT83QKmniLGYvg55oz8Kgf
Ygr3jVZwFJm6vC/H0ejX6OzDA5ojp3tYFOr6BzkZims1nDBwxfHWfyG/UFdwm8+N
gBap2bAp8gtdexRWGKWaZQ3O+I5XMys93aMCWA57joWpKPWCSV7IblmhxFK5im0X
ESU/ZnlkgEapcmSMqdEfzvSDI+rWzMUY4Ot2uaQrasmK8BV5i2wjq66aNbcXREzV
28pD/d/PFJGUZoxAKrwVYpslH4Zsebv1WRuyAZgYNDIzYT8iAujT9vbpzYc+yMVO
VUEgkPvpytDVeiswYhKrMQaOTAv2VYkerim/uTYKsDpY1AzSzmLT8qSwRHpPz52k
1imSuRoiU6OHBh5azlbTUMCmPk7eDE4AfHvqBH4QdRPNNJBAfnnyixlUtv2Xg5zP
2fCwp6LTdbqHn4rgXN9RHloktL31gF0OZd1CXjiBTFFviJOd1raCnd0FvVfzBhUS
STOVxyqAkE3724BO28wWR5ZG2+7tatKjuEAwEKq0NzMOPzlQ0e1aZ4ge0stS6Xju
VosoLJqI50wfm0bKy/zNtIEMgbNPNHJEgFK0BtzsE37IsRlt7jdCBmetLL0kt+i6
pvijy8RbM5gkGhYp7+GRtlnXNCfW2/1BwzECSFNvtv/RrTj/o0eBy+RPS62ceh6H
tLAK2T8/C5c6AQ2DGK3OYWRk/uBqhps0EVaLpUQqY35LZQ0GGmkrva/T51jvbG+M
v+BmQR4xFldnIGnv6L//wYa/UUY3b4ii4mpHn86CoHejYCANQ9Jj/P/Nq9GPw6q2
RFfqUbvo8M++x72eDOsFlTt9ZK4YfFzRCK29+GgxIA5ltcySX8P09mVG2Uub9y2D
VnISb4EIL7imPbIcidkb9c8d8GKAtmNKHbD0T15mfmGyqwa7NDnnJkPxTkJsHrbh
jMTseEyJDbDglNRerMbheQBg5QN04MnbKUENMYX84tNd5awvoMW8nhxDZBnzbUCl
3ZpC3GnheHjm/zDFGK21b1oFnCdNllyVaAtT69Ft3lZqpMpQW5kGTCUO8w0ofFqk
Wxeh/Jc9KRRS3mEcFEoSgTc5C4AdJXPXKM7f039w+v1k0cLTCnFeqL9LDQIosX/+
RAUySKWZU+h2rZrpSUi6B0xTp/SVonBwhKUbiyEh0/Il6YS8rD5/tbG1Xni83uuV
ZGEb4sQdOxmOsi2TslA4qaH7H/sjQJ6prSUqO9Lsa3RtMyiMNJDuYuC594Dr+RFy
uMjCaeb1y7GNMmxplwnyC3mDWbpXvEApzonFYH59QX4aflJ+xYQYOXniei7P49Hb
T4t50oMwKDBvpbtmgoQj+KkJfLEOM1sWShcIqn2+mgesRaAtSOIPfdng5temRgXS
A0JAd5ti1Zl9+OtgcDre3agMzYZbKMOkBDOYj/k3W+bHxHFhlu3D/ztTgW+h3wdD
pe2mdDRwHFqi01Xn2z4GUsLn+rfpR5to2TrXSqWOL021uOogJU3J1sgsPbHTBXkS
R7Jb+EVuNT8qkK9WQiqV/FrRSPWtZXeOCLk0TaIEKdEzv4YWOGzeLpIz2GZrDGJm
yNUUHl059+P4IBc2/A2tTroLpR7DjnW0j7zrmrXVL7CuDZPOOt9PeQRzCoyM/UEa
jgsCgoGKqG5Z9+tF0N57KsR49gFL0adicf1lM2D9CkKiJMSdnkOQHMSXWS6I6qXH
hjI42vimsszj2Hqrh8XPHyk6AI/fBNsQnHVx5IXDiVN1sotirE3tvzDcfTLots6s
P6e44gvfUNRFQTUOBQa8C/6aHhqoX7NU4oudiqOoNEn9stAQnqPF8ZI2t0k4wBiL
a5XBcd67yAnmwwp5qWIsF0ZBhRTyp464hPqnOZlneKkqRx5OZQOmpFBalY32Feje
WVx0HchYfuBmvCHswdoCUuoXn2XfmRJvQjksUed1l/ffgflrERpnZ9lP5e4l2zpY
OljmLAzIW1gNSCfla+/Bw+UsXM4d3dT8StUl7ncWXrJn3JgNDi0poeceVPmebqxg
6SLHhbjEY3xdsHME3kLmejD2Qxum+Bm5QAKxdPhe+My75TTn9Ax1aNWt/Ejs05M0
AGzBKLKWdHl+Ere9MCzht961M1JwMyAFgeE45Vw/U3EV/M7sv8g8/C/9plHkITqR
b/0QXnwzLYIbDaq7v7p4IkNca2t8+d5vwFqX4eFFwYIqNDq/yJRSDp+0Dhtbn7WL
rFmlgr6QTuOW8uPTWpzCGnPagtQq/mi8qyRinUFe42cEVx96AcjnjmaWOGYfHL5F
9trINuVRlx0QSzIAM77Rkpt8HsDVhK104LWbD5ITCpiY0xwJSKSN4e0JuTR5ms8+
KYIiVTwOtc71MulGLHQvUey4UKe8RiiUWWf0twDoGPtvUXsD6R/A1kzntgdfPZzD
QfyRxv9G17wvo56CgJbqZQm8MfRqlfSaL9WvuadXjwoS3HTvOfSRgs301pufGqea
U71g1FG2cs2PTUS2bH6NhUwOPcnCwT0fISRsa98C5EJW82zhVUqyhuqJiCVW0tvI
63juedANNDl7WadT1ori4w5yU655/kwjaLTJ9+ra/0JCyJouK3LpzwMBQqZJaOru
YaSV0AMoT8Ujk5DMK0g2ZsciRVsw5GBG4DeafmWbGXsNZhigfaL6i855wQE8qpc6
ArmbXnX56ioXFJ8ZRePtC+KsB4g/amHfppW8aiMDGrtt9waycMIm13ZbPjBPjuEu
Fmbvzz0ZfyoRZ+Wkq7vDg3Myoo+Y3AzRXgc3oNVEFMfUT69utYOrnRaIzKO6i44v
E8YNUOTk0En7ZMHM2IMsFNeTduUxRsdYO+iRyAQdUlgBSuaQC2UherIM7f0voaaw
IrAKXaXiOg43SPI9CqXiZRx7v2YX8gDmOe/qo6bVw8yvyQzdsyy32lyV96+SB5IC
UW+ZPjBHMLhzNBeXTBej8ywX/f46fPV8C0Ob2J6aVhIIkGvaw8rrLDBn6Ou0oqQ4
BW8cTpr+6JpwXk6Q33oTGDvkSHXtXvt57Xll5qCCKPzIbxR3rA1z/ZntOmErRA1H
LMh6juaBL8+GcPoFKZ6gLiNpvqdWCT/yBoxPPJ+KaCzXCBTZZvFEtjzf1U7DGmEm
nnHmFPV5WmKfMbEbTzkICbDV3In6AI6bY9UAyxRrSOWkrWNJO5cEvh9TNCysd4Zp
acTgFeu+Rgyk2eUGvRw1k/ieaN/zefnoBYZZnM+7NHpHwmVQOxFPprKJ7IPcXzI5
FyjbC8LbyOact3BThqRYpvY86UV8ocrzRU/H6ynH2nafYIfDqyktI4UaELdSP27P
h7ZtPbfSeaL33UzNk+1FkSV47DnuIMmKyBt6Mqfuvct7eakNrwTl3K4oWuRIULt+
E4g1uNYDkw1r8UwENGgHmb97qYxdXA6HbT+IW25qM2qgtrF6CptpVoDFtFP5l3di
cymDPqfqC/4QcUosy6wo2JSKnC21Lfwm+xn9XaKRa0d/imqligsxt4BJNf9ciyUU
GTcD5KgIIUJkcmkJHzcOL+3rSG9K0v88PIlAwqdxrWEG/KxZ6yTg1XLNERTpijCS
TZi7FwhQwzwvwDxJKSsvwW8bVcG2TG/3p9rRjr0bfeAFswRimEWgi7pFH7T3q8+Z
2wPCzSu7O67eRd7bqEltiNVB420DobcRSUXSuCqYuSehZEBiiw5iRlgPu5/9MhP5
E4vRy8fWX0GOlBHHxvhv1RbD9akBk0zofR2fe1gZUuGrkq8nH+UpeKzXkh8vXEHC
i4Y/LKgZF79Mt5Go5NsI2NhPEjI6VZHhbGqC4qWMwsMIF/bDqxvn18V194VZTNNG
VO2i7S1IUvLdYfwejfjCUnksIRP46+gSucvo9iYiJc4PeuTFBzIcv6bBr8TWCPEQ
mmmT1Iiiu0AKV9LcfSZHe4xN9Z+Ruf8i1dviQz6/WOJcP4NvjhCktqBVAEXKqXfv
h0GIm0SmTaHlilQDj7iv4boe+hBMoOALyAPg/6r4FlIfQLt1GZGfuB7rd3yOZiD9
Ks1qz/U5cpcLqYYkS9hw4SaUJzC+XhB/lOKlxJ9M0ST/cGFD23R/G81TOUr0hqW0
9tlbuAb/wpoaUGhKD7F7NyTtQtI7wHDXTrow1vVb2TklJ/sk242N0HEsg3PofG+h
m2zb93zpGoe9IxcPai/faclUU8XQ0C77NzV4KMS8rPdUTPy1jTa0QYRVhd0A3i7D
zEGjNJItLypHyjs9tDMI9rDC6hw/h0ZofkaAqedB8MIOe5AMciaPsqDBdsr28slm
/SbdNhWFlo/QAO3hdo2r9GTJ4WOOse9TIRSwyh/MsKA6AvZKIonu3cbQlBmt1BVR
9//5WQahzlhZYvnSS1O8Fva6SuwIf1C5Bj+5zIbOH061vx/Cud6OoVy7qC4HY1Fw
UjkL+DKOeeF+ZiQSII6L6eGXC8Wx2pk8OUl3gNaO9yTvku4gkKbftD6yesTBpT2Q
NTvuN1TWNq9eUn4KS2G/V75vO0W4sXsuJFYNaHTgTO4S0W/kYSYnh96hX/lUsHQa
78uS9TPeZiFfT9kddZzhHI9OQ8ccRrb4gm/yTBx4KxxE08hjEidfQXJq28VS/CQp
JPuaajFIi3ECrw2vfUkl6n2vn/pKDKPoTG9o3kORPQ1Lal0BXobMkQiNW1q/0x39
np0kxMLcjxz3nwKYbQEXBWxrHplbPKmOJiPPnSQL+u04uCHj1yw5TbDXUwmnLb7T
I0YKgwGWNwH8lnYXy8I0cN2fBnzufGUsHG4B9kizZJPJYeVxX77Z5NW0cQrsysCT
rbcqZqjSWIzGiPFNN/n4qAgZjRrsAxCf98fxu5uaNkk6Z1MLqnwa83Q1paEHu28n
rcz43mtUK2wYH5VoICnVqy8h3aNXv2Fpj0REZ0GvXDale5t+OnJAth3tkYxEBjTP
w23sleahlPjwRdT5dEnxUXiYCY3T6FX/z6Fb5CbDqGzuSlBn3pNoUFUPnn58CqkZ
UVHjIoVAm0Mb9zUr8/kpZPp02+Mwf0hl0aBeF51AzUh9TIyvYWqmJZLXqPRKBe42
QE5Qux1t8HBG/j8sFdo38M0cY4iJcuUpgxfMSask82mKiq/BZIqXdoZGZWQGHgpz
0SOb2pRmVrS8s3KlsvLcOzrI4dm/E6Mc3kYV/n/leE9aFjB0h/UGH46G6RvHlesX
8qYyMW1JNUnq2QxERi29a/smNL41KZrkN+DaXzyryr04UZfwDaJuc2w3gXIWYl+U
dYRNXF9dwPsw7CqEtgVgArC/o6+agpSWojWa4uVRs9VeE1WDZElswH57dUagdLbA
0uiM/cxMR3PA+x1hEm7gOSTstThTT9+zVwvJSc/ND4GLsq1hj6sF0l9oyc6f/nDG
9NOISw6UXvTgerZ3Il669kSa/z/HssJ6qRwhHqUYoCjWfj6RqWuHNcUtnF5E1TMa
dxZHW7EImCD9/9UcerKIZR9YrU5lyaMgcN4bQ4IpxRoeHmciS4z3Od/7cOrDwHCM
6pnKHoclKqoh6rpYFKpVj7b7KQ0KYo+jJ+FNsKuWyPd9/IlgztXKBmex6pHHRrrO
CdyVhCrSLpkf+BvmHTUXGR95zTyjR/DDlRZPJKfB/Y0ydztM1UW6AkFudl/2nS0T
2/CE+89R8fArfPzA++b+NnTrnGKRuV7pt1Cyjsl3XidJaoX8a78b3DKVXEu6rd6I
wzHNZLwmv/5oJGyZ8gBLuB4xhvvFlBvWgtnm9vRP6VVqxNIw8+SIi3YMRJouYnHu
XsocrPTqx/FADtY2oEj7g9YWwiW/VhTebtEMRD9bnBYMNxtaIWO5nWwFw5AF4Fk8
WCOwdQuBxgHmN2malMSZIzz+4C6eYgLB0WacYwhthKlNekr/S4ShH8RBm8ZloKU7
R8pqCTV19IQUQMWTm/UOS61Dg3np32X3fTrZu3iYrqhIKeinuVnV3VWrnLOiRLxH
3Y0dGgMXbhsSZre/6Mh+0gqKhJZDoV9snVs5ljIqhd+lUntI2yVOht/jgtXN7QAS
d6DnAo6AmkU77hk1A6cgSckTlYToLSXA9GsoCpbSzepsu4bbV63g5p3cc78qbN2D
cUunwfH3dECm4eVYpZPc2t54qULhTp8sKYBtxBfgQKdD2CJCaWzu+gHky6Wt3Hi/
dM7prWChGypThlcmv9fjcFqieQLkECXAkKSadThhrNw8V0TtIz0DC+9ZsatRxqI/
s3JScP7BOzm+85ryn/umYCt0GECmR4NUjk+V+pjkVduXkzKQfYJ/o8ecARN06RZE
pxTA1w2oQcwavdj4Sb5IoPoZHx2oa/9qfq6sxNpPn+D2JxNJ200ywgp9TLHVdZv2
b07998L4uUiBgHkiA5+qvoYyB7W8x/BCzLGIpqiTdnj4aZkiVMrPise6J/kWEDHv
jOHGuyCs1kusSBCtHK/5Rz+Nq9pry/sVpIe9fcODqNg=

`pragma protect end_protected

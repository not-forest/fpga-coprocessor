`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
iX4ovhfWMJfI+WAA+mt8FZaH+02cRLuAGlWbTiXFml55NwOOUZQ5rsSDvYynJCo1
D8UNYbtHUjUUu3WE7yRaLw67C3n3ETzZwEvFZ2hywcSQu6BDqpHrYeGTurULXcRj
W0RV9a/io7TEl2Z23GOncx6Ek/AWasbJSOHMuwnjPs0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2176)
6CeqJLU+JxRuSOJX1yUzr8T2+3DwSYe2x4taU9RfYbEjWgDcgH6J6AEvzvTc9o75
IoXmaI4kj0TAlMOZCvXir8JAp/ouYj+fE9p3w9P8Ocku2W+Rvmw905lzjLzxjiMf
dhBReB33koaH1QrSiefMgu8fi9wO5yZc54LCbsoSAl5Re2oOZfc0W4uO6ngjWVzZ
igSqqkeBlKixK98omEPcqa6l3WU3tg7Lyg09tIJju+JpDNihpK4r9ytc+xvsrrl8
HRRu3URl3iQt9CfR1dVT3FLIFofHR1FQv+RGTAfZEQ97Sep5kSOfqzFVhNaU29bj
8spbiuOYiBymGL6oLUwhyOphJ7tdQuADtN5waKUfKhLYJ7yOSrsx14S+LWR3XcA+
xIkit0TPdcZ4bTWeHSpmF5yT3OQmgL+g7OjPCnZ+3GTLbhSwA4Ryo1amjFHFJo1Y
Xii51ADKQpFbILKmAa2f4aahIBn6u3LuU0/Atb9lVRLSfh3EqOZ/AqSJllFcXbhP
UWWkpgNuC23aNINu7tZsqPs0RPkiRX1yFIp2YF9LEZlIp8qUW5vxrbYTjAlfulxb
H+cLwSbujT/eU870ke5BD3pr1cWd5qvGDT6TM11Effbvxi7sJbf60A68StzBqtM6
I2u0Vg4au+ZHaHzbzAn19QO2lkpa4Hjf68HC/sQLbOmqBlTpb9i0OcZnl5aYYtjM
8sJOPIVJXzKzDhvBvh4T5FYoApbQ76DdTT+fX2v/BGyKkVRaRnJ1osDNiaf9Bq3o
MyNHmihrLfErEvHBrP6qe+aizsh88/XXQg05Ub5aIdAVsgfeY0dFySj/p6jdV6Gs
LGBAKTPwK+FVDbVslMDXldMQcPMBopjLkWEl9M3q+17bIgJg/OD9qqsrigO8kqlN
ykzm4FxUYPzhkEpqqi3f1mpUDr1AzoesNS4ejgRyL6DeCewSVoFtauEWovooi31M
oVIFP9+r1Jo/0j7P8V8mRh2l9KeP0y30GyX7x8M9e7NqblYucmEGSgA8blMtNoI5
R6Ym1Kku4Fje9mLDQ3R4ZPCYjhyGkfVrYS0U9U+6IOQLQZ9DwcsEeiPTVEZ9Aj5N
RuoXKIWI9864bQx+Be8JbaA1BR6ea7667O8tZPjSn+FrWd++pYCNCp70QmdCdLlD
SquqhoeqtavBLXf4/88t2wA5dU+jV1Vaq4SbPGIlTlSJjlx70bughNjKcM0e3sZP
ZCjlOplUrWUCxOP3XMFnUZBX5MSVts77LzvYeHyoMClaN+8Nm52REfK+vICgSZmI
dS+aewvuJmuPRLc4e1gk1lp2xmQAX4Wy4/15kzPhpNgAhY2HQn84635J/zFEmE46
IxVHRF2AXlGmTQx32AEFC4xTUzL/fejocCZHKNEZ0ACDiK82LZ+9R5OClLW1ia9K
nX74H3rY5/59usO7L7mmV8+ltMRW3iQTcvSDp2bJb1QbkrpbcHGw5k3Rl7VU2JdF
7zgaibb3vxuLwYMhzjOirvKqIEtYE2/rjw5e4IZkZ2kvLOXFgBg8G6ip4F5yJu+r
OJuMSsE7VBHi3Y/zV7yJ8ucPlZv+V53t3vNcPxvv5cHQ1YqH1qHmQuMOkVtFgEkh
GcbAH4087LP1F3HuUCqn7JhAbdAGyp+6pvyeUtROBdkxAIP2a1gn2LDLKQs8mJ4b
bI3ZOawH4GFDp8xBiuqXjXxZbCn0p3g4pextSiy1YbRV8upJOiv3Hb49HWFWUyXK
80hh/Hj0EZFjpU+ewYt7QDSvE1b1wx6fKRoVdr+IZf+az9SuXY9rhuQOzRMbyydx
7yz7f+U1ZPEczPzzKVtliHTFK6R/uPsSkRMpgwGwtL9DjgUKu5ZQYxshyGrIBjXk
oAKBk4YInVxsm6ml/AmpCGpvX5JFz9uVmIt50/bq+x8GFa8LrLfiSIQA99ZC0nSp
fPT2mMhVl+f1u2r7IfJtRLlbfYWog8vTKbCg6/gB23HO9ucmxPZQ7/Rv8Esri3Tr
5/nd7N2wEaxCcey5sUPVOlQ4MYpHK9iinZL9h8u8uW4Fsv2JC+/WaG6Xmrg7fasC
05c4St/LyrKvpQcfQw66SPF+c/nggW03D2JSqpWtRAOKJK8NV3mk1a4vYZb2nNR6
3KOJfrINY+C+nh9Qn+kkozadsvHiNxmtHHaqMNAinmgOo3qnbBSF2UvTtfDW70dX
up70tL4cY3YnoYRU3pD/HNZzBJGOHF6jPMAtcbfm2UzzCbj3tt3j46VaHlA/7Ymv
HzTOFzEZipCq2JXJ9GPsqUn3BZJd09agT0KMt7uClqk4oChldc/jJJ7pJMLam/CG
IRSpluSMX3aCUeZbAPwMC5sBIAP0zUMz3ctl244a+S33B3VFG19F54GyaKC03sus
SgHwgjXIKl3CLrRR5YtThlWPDmLGTq/eRcfcTx24FNjJXMn1HCNbta6Iq7swJgHQ
eDJ9drlZGJt8aXgAjmYEuXdTnsudVzksmPpnUAsQhoLopZ7l36bUfQYdHdUJilFE
rLRR0ZPQPnTPj/Kgi5Qsul28Vv8/b+nRutfnxc2Yw+RmMMzjpc0nUDW50r7TaeTt
pXNzUEBVdOze2UgTtAC9yCZkBB1HCGQmf/gLCtmb1BM4zZtzS/mKb74FHCKDjPxR
Lmio8cxOnC5ynMcJk4VuNH7qSca2pjnt/p7JNSkEYIB0y8mPIVnGCv86y5Pn0MvI
sIKXzaham0Hn0oTkvn1HMayA0glbjQHcfsxUL+GoJtTH7uYZSWYZiGobIs6Nz/q9
8cb+APxLM4HusRnkF1yL9QDa26XsyS/obNQLJNzMLIm2oFcdUt4h9NyhqYEyHhYE
WK09F7PP8nu7A7rcPoafYNVa+NIrjoyEK/GFo/U2nkXq70CLgi4JjaPXUyYSvpvi
J7viNNoc4xw0D75u1PfONQ==
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
hqqElFQSixuEVrvYSqiPUMF9WHme+9f1KThKYlRHbxrEUTpnCGRyHRNxvZoy5b37
JMPxKGUXF2O5KO4zbg9MzFcYzF0GGgy63pjitqVkvcUtniMVXtpXjgRAam8c7enz
qrcjYLJddNfvNy8Dh+KyPxZpAwJtZOoVYFGDpLTWKgQ=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 3632 )
`pragma protect data_block
vx4nrYe3h9wETgE4q7LUIt7eJeJZJRQ6AKl1RRzu34TVLdMPlRbQ0wipY8nXOGD8
h8THa2YWfvNAcDCiAhkhiOkcvYBnOLChHfCWXY1cIuSfyTFz29oFBhHRx2MGrK3+
VobvQvM+BL7nmIAYMmreiDraxgQ2lEBGSsPtipYXqIoEuXj91unl+KhhG5aWs4hC
qrUG+FkBVWZAXvEDC/UDuxdnVP8co+Ef8HQDGT5pnHd9fvS5hsDXHOylExz5BhzI
hzhoUOlGfZ5o3SbRvltbp14gKu1/1Pko4p2INgnZ3RkBaKLkPoel+0WbaPsb47fS
kdkWNKxmBXOrG4WuPAqMYG7FepLL37F9O8f+vJssXFZvI4fvc+MLUWsfgniqLYwa
roLfRS1W+1A6/Ut6OBcndgA5nEZS/ZkO7jFSGBgM2M3RdYBdvGO1/9vhPiZLv/M4
cIYle5hbGovknpilfUwsK5wYO3z6wjUfTT3dK+iyVzZjN7JJVsaL3hE6bhjd43p/
QzWrGJqs70O0eTnjmg7zabIF+4T4cLC/rb93EuBs6JWzqJkh18Z/Dn6Rg748rNol
DE4UIzRT41trXysne9bN7LlcSudFG0z8MJ74deEzQlVLKqc2v6p7Hi33O1oeMAuO
UuQXCg8Glscs6IQC9N8Y53ErQ4RmYYkyJx/6+peOYJknuxlGqCoLnmvouUNUelte
W1lpeT0zD/aGgJCjl9mGg3Uu1+l0rYkktcxdrR4WAU8SNyw1/1FoAiTxbKnpNL2H
3kHRTMBxBJTfea6hH8dVoe7nhPHJ8Oo6okA8UBPEdVm9IF+cGRdzBRkGXDVlBvoX
XmPsOsqQnKXUh3bAwjyTeomsF0aSNcEwjnqhFPBzKcdzPRjKaZGAmS7M7OUigqvC
UW4G6t7oJGPfnedpNvt6XCEYV45XpVxc3bq/53qogvhMfmdy5+QM6Dl8GqOEKdpX
ZyZUdQ1QGJtbNT0Uwh3L7Z9Li29koZO4u7OnyAFnozp4KiEv0jjZ0R8UG8V/Orjz
MLNT71dZVwk+tV7MIdFz0EvCLZFA3N2d5f4q+B26vypDfoEfnwgMz/qIPkFcU+nO
YA9n5sEWZAtZowsmvaXm/zSiq3Ie4b4TM7Nz2HAY1qOoGHRgMiR9HsJKzRNd4VEM
RXRUWh3bbXisDLbI3xxSSUEmDtRCBjLLqMZiyAoTjlluzwnyfBdpfFcCx2b3Proj
EYvgzexCOFoM/eNpDhaFIncdZSCWe+3H/AIH+Sd361+TgKisFKHplz8LPG5hyyEx
4bBevdllcHLDsKWdG4p4Qf4ffaYn/medegwski2e+xlNGxUcMhHR5s7lrdMjD9Y/
OU4Y7HC+NBVqQihe51+uHbFe0txFxC9k1lWJXJdULQAdqbsYJiLpp+xvg/1qJo2Q
nr9KhdPSusv5jey3PSPt+PZgviTc1k9I6jZdk2wXhgyYAW73/jpWFib/Ljtp/Kje
szVdZAbgVOj0398kMDOR4t6sk/6FY4jX0/l+DJlo/xDhyOXtoA/x3q/h9xs6sWsH
t5CA6hmzBKvIzDUlhULLTrjxkT7njO5+/07bWVOag97gRBlQttVYlZcdcIw6GIFD
cgnLpkTuD+9uHW21ZB6TxgOaTU3zBM1ziGz0Ch0AEwdrVsE2oCOi22gFTBi8SlH7
NrfW1b9ffVgoRtZRPyPry9udLTL2eEuOImUijK0qAcz68NgSgQZN2aqLoOFAAiML
WRJku88977gBG140tBX4AQYTw2ADIQ1bJpCyWqYyqmyQTOFXbpAiWhxHcEJd+PRy
vWY12JvM9v3CbjwoDolcp/eEdX7jkPBuRWE3RA+/cE16f67Y2i/6v/bdM0LKzCqF
YjNeWFhTZsI6VOt2fmjPA2e4/tHq+TQFmcYLJq6YzSerCYyevs0kaoidtCTf1MZG
r76jACPqeBXYTwXcO3daDs7T0psilL5myYAe6ZwB4HFnoeGe6KeP/sT5B2VIU0Kw
0KQn8TJLWIQxetKyju82WjaPmLTljd/7MrHsCmDPzeGr2o1sY1sZfTJdbN5tBE48
ZrKVeMAdH1SK2rxZC0lvJ18LuKfjY5+MPdev3s2Lt8W3ppErXdQwp1+XAl+Fe8nk
rgU9038NOEicEEwYTOwUzYNb49YZIVuNGgjEfthjHzxh9ySHWdeyKfq8mftfK9MS
SgfuXIaxuXNSrSdM3QRwFY4fpEO+fq8IHa7rcK0vYVwVg3TKwywc7Jx0ML1Z1bq/
ZWCIudRT1rv7BO1KnRwptUWb+5t3vMLF9ha1bSiNxcvICk8FO2MVyDCjDhfh+A/G
Ufxlx4C+7gXmn3zrkaQcqu5L6ASJo/lJawy7FMGkFAD8n0FAzUMypVmJnsx2eC6r
k+ZswvvV56d8eq4ah0YF64//LJWIibr27/YtDk3tOH25PMch1mlDquEZRNn1NOth
D6W1CMPI77JOLfuUDkzdTG/dWs9FdnjHCWeiWayi3DpXjl3KrOM+vvr8YrPl/YDj
YfyU6Aw4dniNesGa4wls8KXKwbTLCGS9tDFwBMWY4rN6RzZnK+Hqv1JWJzgm7+dh
2lW/yEktcuufOR2hMCxy7C+MVnFtA8Ur/49fUcPvo8osfYadMIb8toAc1J7NqJil
uv1IO9tqBjFOm1DC2vowRcPQQ18bftcRM2esdY8Onl1ahCbbNgZk7Ym/c24NAooZ
4fAiGF12H2ZwoSj8SkrbOCbEg6vUnCLjOic4dGb21hhuUbpN3kU7UI01P5s0RX+k
NLd8cUR75hzis/WS3/R03308wtXb0BAsceTGWlIWug5SZ8sOD64WSNQSVp8WOK/L
ungfF+oNLK9qbh13HeFPOZkKDcVDr/o+bR5v8mCeHUsLiSKPnBHIPyb7/gRFi4EH
6t5SFqH2gvbyPXlcgkQY2eqk946o1gz3pvieOuUBOLcYYMpcs9HhNuf5IEAEAbVx
SVVDMRtCLXklqXkSQWBi5ll/7Q9sgQnh9h8LH54Q7vgoYs8lWO03QuWYhc/GDvEW
fYE8Y7Wo83ilRsFJbsCjX2GQrNKAtV6j/Ih2+IX2oVZFmo3ZLb501f3l+AugoukX
uBcdfDS3VuzOpNSQr1Q5RzgopqmXsvyCBXnIu0lAhb7Kqmjv2QvsKWXcFhubNA/X
c+A+tz1ZQMKRHW7jcciD/btOEt6EU3RYqnC0+4pRCCegCJoSqqKDQp/QJb2nxx6n
z8P4Nqi+vmXVBRoYuynkHrVCHlQL234zUpKOuVIDUDLtFOIrRfG4lOBsdoJmZS+1
kHjbBCpIc8GRXKkdyc75fT8rsdsMQbGob9pjpzt8o8fBkq2zDWpfU/y+oqNkdgrp
/Fw7PwvmEY+qIHCgqGOFC9nfW7exj3N2ZI43UZzwWL92j+wPb/QCypmvcQlPtQ0M
JzrXjCrP1ynlcmvmhrl10enpOf1hZ3LmKzdMgfwaN0lfBDZscACupCbAHjhkkeNb
pepXm0HxJMl2a4WTOuvGhiaGkCD+6rdKJzM0wnlKqNd9MVxf7TIuk3oZplNrDxp2
xhJU8bO0d0V/5OyuYTARuuMwBRx/WqUvKyb7GYM8tqH1wGR+ox8xg0+Fn6FA4VAy
q5SHbq4Jk3ZK/RKc0IZru1pH6fxjLru3zi94tWZ1sAL76VhNVV4jbV/i5jMfo8Go
Th6D1VDMeSFxEmUDp2sWDWBgp/H/F5Y5mbAeUm/J3PZvimZNIIlKJGmxuyssGo7t
wzxiL5FtFGvBatlDHNBwvsfvLZLE3+GuAk77cbR9LO+WlEhzUJt1EY/ZMtcqO5Vz
+0/QXBh/8Ny5Luxx1u9EtNOu9ki2PWLaSAvLXj4NAJt6UiO5FhSc77mTaxQFT0rY
Ko/KUqQoveSWehLi/kZ+5i1vCNeCjTRIC1HXPgrQDJ2FCxRXhwe10ztGJ/q47VRr
pMP3BPR9AYZ1TSLetusCSAqQkH1RVuOcHM3dSYYpm5X47CTYr47EwKJsmc++qFYT
ISTYPyRS9C0+bx4dfH8m3qOOjZnVCG3F3Rz0y+OPz3w2K+lsgDDW90LqsgBbNj+T
2pv6Pb66FlXDzIKHkXnKWDkG4cor5Na/0dV/QfzcXxV2Hkp/d7W2aozn4VbHKgpJ
8orbXh36QvxclxJm4bbF/0037Pqs/9hLOo6Jgns5ig//lyLHGAmVOJIvz4CEUrUD
xZhgaSpcaiJ+ULEZyaolxecM7yDgWNL3IazFUW6XJNy2bJkE5x79YkVBR0iXAJcZ
1CtTTeyYsOqRkwG8/cmANoQ0wDF2dcAxJDE/ZPV68bnWPEPoR+CxcOmqxn+zVe4z
InHPPeKm2KoCjDVl8SzQsrKsySVRKOXuMrOQVXveBm/lsgK1jI87EQfdh8XKW3X4
lojqXGZDPudRXbvZ+mbp446ybd8XmeFqg+aalB5hYfRNz5/i4EIjf0hCjYZVhmYq
jCyIDQu3UMkSeX67KOHYSEmJqpoDE9ElEv9ZufqbfGyNbRD3GRhqfF00MYOMwIHf
ElxHB7RAa7m4+7qiuOUR5zwiDlHFXjCMihdeRf4i1Qwir7gcruLGWIMU+yMHpAid
VjNDQOU0pdH+gAt7WYg/ZRbrHxmckBnVxqqGUJ+PaD29/UtHwaCk5UV7EUrXiMXr
BX3syemtL07Z+EDPPAAU2TrsPkLeV6jFluqLHQSBqusAfHh92B+Hj0zR6GyGaRbL
zU1N1XZTNq5cKxtUqxaXXf5M4s6UEo5pwPMwRopQ8VWZyyDWuGLmkJDwkcgO5G5u
I7DODHsZeLj8RsM/W4JSUz7/FXNoC/m3CBmzn7VeBA+FLSPqkJMkf9OmhKpt4NKn
Pls8w4QaQ2MHkSG3SgMiOCg3LAwHuMR72vFie5JE/0c=

`pragma protect end_protected

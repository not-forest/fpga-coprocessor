// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
EyubLbFX5J2mydty3JDQ/JobIKuOeh9URe3+dWjB4Y8FGuVyhpCwaES0f9gSF26w
jxcUjMVvedDlW02nfP+vzYWG6lolBE2nlt0cB//O4MklHCSkp4kZ1CoDn61DGLqg
sWJsWD5LascEALQmxSAF9lPQUlfn5Xl9EUnEVZ1NmpzRAX78LZs2mnHG1MJvCX3o
ROoJH2SL3P2y2qhyZLDU2/vvH2k9tVSPmvNCY0LjJiZNg0Pxtjdj/smBc0WD5Hrg
O7JPUEfRWRP/4ryCdBsfATyp6nggvU64XBtaL9RK5jnbB5QScNRa+sOpZfWllo6D
M005gmD7/2Vx8bZPkYel6w==
//pragma protect end_key_block
//pragma protect digest_block
9Ev55aLTL6U3yyKcpB1CxYmEYp4=
//pragma protect end_digest_block
//pragma protect data_block
yK3saAyPFK4A778S7/qFmfXZWa/2LVmqWQbQY+XC4dxSfKEU0s9QYiiGcQeSB+ar
yl42U8sPPUPLxOnHv5im1/xqoOuK51LIVn31ZCsQjfEGUtWx3wHbsZ35FpO+SQlr
sQ36QARvH7wAj0U2BCQcjFIN+5S2D5+NjIEIK8mn5l7fVhNTBRtSWkoKGDPiY7f4
PyZxi4KC1rJ4gKWQX+DOK8IBNZBlsiFm+nyrc3gQqt4YwLSNjj+Aj+S0DJKnYJPT
Q7wAXIhsj/PGN2trTGFW4rbR38WbH+HTllZm+3zVGvoKTUWzBxi5djhQs0PxoWh5
nDotEvk3k0eyljxqfPwq3R4kFTJZxARQ+0K/RLJpKRJEiYGeQ6nDBJtWZbmwkOsc
xXmn3yp5GSbvZRm39l0fT5qST1KDImdzhYUjC+HThfjKRTpUyeVzRUH9kZsPlVXF
F3ZBcKaVkzKHNltMHUqojycjbwCKBYWQw8nEZAZYxG8qbBAFPrAW7o2HwXFIQ6Rr
d0KAcarF32kiw6LbvVZ51A5OLEvNUUIWcqE7qNPbkGox46FwpAMmdVuWn3g/xsyP
IHE9Oj8/52WT8Hrhrcefo/fWEA8PjLUY72gOH4iPBwQ3Kxib49Z/wnWf30TZQ0Z7
X2JfccFlacuVxR8NRnSWVUwhx3LeugIOgQWATP8DFOhy88Mbm2ptMaoK+QNDbnlg
NclCLKJ5oMHHKb7YQqcmzErE1uQaGn3wteA7VrB7Mjlgi/dvkRaq6HbekfGrSc+P
t+wCGsdZ1Zhz1Vju4WV2vk1JRhAniUYZ+XlGmijcT6qMFkXAlEjrf3BGpJVVHA4w
qKIpEK8hIKvkiyFE5sIXkaT6vfQqgTTHREoWJ2BVBGymQe58WiOkhYvnoeSMDjal
6M8Kz7qtgiImTFoKgs5RtF3o1hjA0ebOJdAARCpXNTPVyvwTd4WVkCQKN9pNg/zm
+389cANtHONu0f4nlkScwR+Nu55uH3KZXVgBpThs+MnwKplOZ53sITXEXrkyMfwh
URJ9AkVz/A0O99VPhLKpsdKjWQW0vln42Funj+UkqFqXIdtw/xsKvSgk0JN/8EQN
814TJ1MErCkRz7cj/EQI5DDlsgSnpIw7HZevUFyp88GZ/WmCU7P1iovGUuFb5E7D
SgjbVt5b5BzwOdqAZriDCxjwrwaZde+q1K6qlqQn4hWirlRymUiiULrrrGSBPoyr
RsWh3SNot8Yrw33zmn/S0KTxsN8s9bqPswqNY3JFChirjtGgMJThI6aanegkmyGv
ByTVLumUdJm8dKFOAEq4SvH5chPMRdf7RQLqtEaYY1dZCVkvS1bU1L9Dhv+soOhR
X1Tb5a1zcovtDZvtksEbQB+AxVb/IXnK1flVXYO0K8kAKFjSzDATlMkC98N9q27/
ikrLiQlfgJIHsa6fBR+tFZzktRZ2BsP6tdPlcuMqylKJfEvBq74Nme+YBluTVt7K
YpgzZVB/jEdf/2L9K5AupAacBqLg///ITdEhOvWdfG7s0ZmmqTP7jMlBq6KjnTM2
/cEmRZ5Ldminp6l0cNBhgnzxTrxnl54NPbkf790hHuFD29DSV8S/GGvfJY9onME5
TTCX65Q69oL16zWQYwppfVSb06dXG/G5pMu1LKJMvp8Jjz9C7/hUSsG8+y2mHzWu
G9txJ+qyYiAaTZi4vmVKmMX/1Hnn0cCb1y1007xMViwzeTjLOm/FSk54OI4uOYf1
BpiFDXu/2SzX0fv4kCeCVqdoFEi/+4DYSnWeGnUljn9XQLEfU9hf9gTxPSooErzK
C4lkmudbptMbkRkYxKoJ5rsGyO4jplIbHNnnjYHELIvfNPRmyBs6zeeXN05tcbdb
EK0QfFwPgnFpDrWitM/mR4kXJcCvrs8laLGIuZ+BcLPf/g8sctimRsT3gQl0UOJp
higcAFlW+vBqVyEAcIWanje+VpbUHsHHf46hqPNCwmKYVXpIbhd9tnGRHC86gQTr
xkNrm1LgwIUPl4VMNf+MtsRXkBxjqCNiuyUmzdBmW/Qa/5aHZV3HCaNfhJQ5GOAa
2Qpg7xHDYuVQj9iYOccbabza7EtjjeLXW80VufxE/hCnXc7Z55MF8qyS0e0Xq3wO
Ol4ocylqO3dDf5AMnYqlLkpq+itZT0UNqNdKUzZcmtfxi4/+En/m+98/l+HFcuMn
6RbahWKbf/KcNd+09bvPrA6I85ShBCtoicWl/9jJFmI4ORWoFinMIg4C2LDdteuX
C9tqSeKyaxrpIjmUQnhw6dPR8aZzlSsvT5q9CBlMdXWwp70LNuouJ+434DLb/ri4
t2Aw3f61yEVHzp9eYjEnPCgnyAi1vt1mvyZqgtSebLnGzY08e8SQwzMiZ4ockVpI
s1i4nNFmnfEWW5op5HLDQsiMytdd7iDUNck/NkUXdLSJy/QMa8Fn4W/bfkm+ogl6
pfsfd0keGOr0YEPUroGS4WCMVS25nRBLcPnxSBOh/vplEWoivrkZAXpBLWINUyUP
/tab57qU6ASPwyYQdjXWIOuphW1kWGRs4rkB9MtB5mWPDHV9lvJt2CJcHXulXFov
9uBMKeP2YE3vxUWGKrptaL9EwkzqPHDOCpT4nBW4Lb7l2tEhN0f6kP9bQX42InnM
e63rOJiouBLw89wROB98w5NaZ/Pv03TRyCvx6Q5mx3NRuMgqOeOEsirOlwtjsjbD
jUPdOTbDiSdrQovJm0EZfE5ge4fkP3LbudzaxladhrsE/LZt0GzXi0aR6pNuoVnb
zjp9eXBpty66RCbF0zT0verIEkPkx2AhyqZ0D6n5VNhqBZwrtNX0gAlg5KUVTy6Z
FkHLBOnZfKxbGqxHm6ncJtXBgPHPzCAzbDK7cixhIj2/TMOkezDLvCtwHs0fi+3r
L9s+APF6aCLCSnw34iYus0iXhUiWS4dwjk20zrY1VqYRppl5OAnFcqLgSm8H6jjP
waRg5xjBWwJLL9jCN+i1MmPmCFRWvYjv0N5hiL6rz8dz1Id2vIzIXfVmJiVVF6eG
yL10qYkDfsYJqGKjSmTa6L3UTXvepSYRKBgDO0pojBfC9E8m0p0EbNrfHF8GETFy
oTbeqkgdDy8f00JpSrpFyhBBZVVvE54Tx3tu1LPUij5Y4AUrVr42A6seu0OwyTnG
+sMivQiQhH8oQXb2pckzdVTJsXCXbgwZj7zdAay83q+WI5AHhZ8Fb7XUYyxbZRUo
OPKtdNiI0yfmm1OS5Z3dG2EWEIla/mkft7dH3dUcKOSca8LPBZBUEyYf3Km/httP
QEd1gmbWRndnwlZ3PFK4mJi09MpBB2s9jKya/gEFXbjGrxnDX0lO7VGbutML3+pM
sOGie44Te7Gfee6XIAhAGR8gRzwL33gX8TkCfwQccr4BJAMauNGwByVBCjtGqDAk
LaumIXw3ttr9STXC2XX9jDjJZS/tD/pFwjPFlNQMXJOnSZhPTkXxe3TzLmNKGOrb
vnv5he2UDNRSnOe4uPaH3svKg0PQ/kRljXEcqtlx90VX+8wihuRYHG1OGMXwy1Q9
GgcYKgH11rjWdGbyD0SyfP3L+XkMmqFntRGMRNOsg9SCTDQFhykKd+ZR8qlk3flZ
Sdf+1xy1bGhyd/cRt0KlCnMnOY8eT45HR0h1DZD9QEVyCIqx4NngvN88zq2rlBLN
Xh7DdjPo3PAQWvKPLTMwJxMGye4IDfCtLr2kHOI5xOFLMZBcfJ0gjAZKf+omPpLv
ozrBj/Ulyr0BfrmupHKZFaQK2VO5tPcGXgTDCTTD/V//08NaO2WXnNeqzBBaKFn/
EDwmaRnGAP8UoZwhwkHWHmAss9d6d7uPXRaWWk2nHdgU/xUpnElDqNI29KS8N0xw
Nt637xCbJLJ5ZHR9tOc+k/zkbyPqTJLSwHLu2vXO1yfOjQlof1s9hTN7n1+XJyj5
Yc9W+ybuhG2n4nZnMlcvy2N5PPoSaPoYEJAXjulL6nQNDtwjl77/MHMhu4879yRu
RYqcZlr/P0yXUwpfE5JXZ1OUVskCkEPf/GbtPpyTwSzNmcX2YbBfdlEAsi4eZoAM
qNIZlyc/XQSoGzCJcTrIoUsirHOWqBiq3oObWL2y31mVBZOX6PRx0Z+4r8L0eEhY
1SgvNpHvXr21+csl/t+0UGmMal6QjyfbKJS+ww/MR78VZzb4TJ6g4fvqwe0e+4v2
LsmhTy/Q7yVWnCevU75lXFjkiJvmy15MxNJekXxfmPeq+yDOKd0VSqVnXhR10UkW
LZmMPzw+CTW/YKp1tlwk2O+9UDPyuHtoC/86ja1kCIwnuqNxpwVdDsWRbbuPD1Zn
UsdWyNaTMEj0qiuJ3xbR0VIRcQLlO+UB6MDgXY90BZ9pLiDQkN77q5b4UCJ15V/0
JbmduHxVX8/6PhLIidhv73YawXyFY3ZZtx/YwN4Mx2v47/fgU8Ftn7W84vM3lji1
2HmfHpkCOejnGK+OL4z59Jz9EnPXDuS5HSYdMfPmy5p8M03/crXCWLRZWPFtf5Qd
3nkrv2C+ZWUX3MdXB//QW4bTisBoUJMOxlZTrhWtST9t/RRVB7B/WhIT3uRhKgPi
rpUZIrW2QqGmiiS3eCOMvewEKCGZf/BIUkB9Npk1mszqDyBp0M6egHD3sflUusEu
CQ+mk2txC4INMU8vMAWo9K1vGcBdIloE0sC6a0kUggLsp9lmR69u/jZg+rBKJhoo
QHfn/CT9cCmSzLl5miv9FUcDnzlCEhMFbV8W1AOGg7+6rPGBN0vI+7qrRHc7JEpm
6aRY22cEV19dmRtABCdHoQeqE/+0tG9oR7CPTRIK1MEBkaR6ACI5nPejcjpdTmC/
bLRdHWDoYoWwNl0/joVgT9v6QV/o5q4886LoXN6igKZ/zcdadN5YeM7pM61AJDs3
WiUcZtipv0pn3CmWgtn8sfpzoz/idmnFVCQMZwnsalX9GF8z4lqDmt2a6Z536Q+j
pSrraNkuZbEeeLvy9qcK+1TVh1PWkbeLD9F02TKCdjAC6jlEmHJzMF+hUDaSIHU8
6LBGUog5Q/Ce4H3TaoMhUdLHz5E19RfFe6ZbBkGd4e+SVOu9may8m+eLstiCBiAc
AzrNWYM9UpsQ2DpL3J6Pp/LOQxGTj01orCS54WXqrrsQnykYu6Avfna70FJr+MkG
cUxguib/yYC07Pexzf91urVO0r/jHYE8RPxc34iG2zTQj/dNVzgrTorvMl2O0gnE
NXVQLcEkLVp56np1y9caBnCNsX4KYgGpc6M+AHsc4h0mHhfBViVQFK2IfAUrNpAC
kPbNrtd4LY+6xGFiFztJiBAJsAzR04wmM4Bh0R/OyR5bM6yFYg/WLaN3Q1smDdqt
RsNK5kH48loogr3TRJwEmhD9q9ogQ1pcKfTIUFEP3oevteU+lN24aBCoFcVBf/2+
n7S/oMtjCqHwUdbjRXyMYwG2MD+iK7XIF46E55H1NuaNsY5LStfYzEasMxTHzy6+
npOWNKUtbJq3xN3lx+fzlJsyXPiaML3gWDddSYXpjAD6HtIh0l3QrT/OimWwHHH6
iH3v9UayI8qcvlZuHG4GKU+xenAXigOdt+fmAspiv5zUz+hcMObD6JNdp7SPW3/i
q8nLqzgaIjUxSmywVfwsME2B9M14uoygctjlWoi0TZgt62tZ2JDxHw++GQ92vaXz
UDCp5cElnvnpS1HihnpxBbe1LAgZsG2aGEbYPvzabzy4yJjdwK6sienE9g2xzeys
sLFujhkqOeJwMO+jdUEiLcIZTTMhvm2Gk/Ugasru+Vn3v8JQfPNdC8aAvlfTxqBF
Fbn8iOL1gipFi91bpLuZP4tytgbADNVnyJziY5tdzn7Pqu07SJafj6JmtjAoXyeM
OMglNjLpIPdDhE0D08rGESY1dKlqRY3pg/ELapLZcPZ7x7o1sSyeAMdrTEuDIcpW
MRZQTEmgKG3tYo01CGULOovmqLNQz2ppX1Oxh0uRJAS5TDye1Lq268FT+j2vPVwS
mQa3slfgPH5KwS+dzOcDaCCQCydGoK5Xuk9TWVorq3perGJ34VzH6YmiZkLeRaKQ
tC8kK755NhrmHC2toyTYcth2RH/tGg0cDACWDcHCIIv+B+qH+62+ZYaRPIFsQ7Ce
QWzf/hs/QGPVWrWd+ry41V6LyUfIClLzVjELWh0j/Jd4UALhqCvDyt9f+4f0zkt0
JXya7/fvwAaZUdo5+opchpfezDFQ0EWkFoMZkn9wOViTW6QJfB9RImCtOsRJYPVY
dZtu8YGYGimuxfKr6XoWRpXRrAOk8u/dYH5A0J0ZTNXxU7A6XT8DTz1UYduIHfWS
+tS/bZBufutMye0j6XBM+7xdOcS9Q91Kg4Wl1o6iqrVWqqJMLBZK5JUhvxLuMbWz
vgXH2podTIznBeOxErtUe0qzP93IleZj/gVGPq7nzj5+SIUAe0hQawy2W6lOlKxZ
1Zyz3tZ/l0dvABJKBaSd4fgJ5ce8sFzlsYXZUoaZ9wryhgm1N9ftjR2NxUMQN6Mp
OoVGaGcBAW3h5SOQkDIc56CY857MyZgyXce2xeblOZYV+2NQycLAFignUjWbM64u
wZPVFwPVxXJcsyTQQGEf80KsevNpTPY6hai1HxP36Fo1lMWRtmUsVQvmMPzYfEzR
icUilcNd7OunaXQH5yWcuqanSrHbwxM/l7QV6HRgU/VOSUWnk8Gh/SE7IYGrRRaW
x6B0CY1X14N6iM0IHDc6weyHF2ZvtKRRLA6mrK/4I7VC6g0U9duX6fST3FVWFogS
LdcnQEtuT0E3/8YTX7QS4byX8hRhWSy5MGOxyTSOfzFwrREzQd2z4UeDplITwoZy
q45hdZx6XlmuyAeWS/tf0TfBql0iIrQ+toE759Mjh4Fw3PCz9Q9wE6MXqx+3I8oC
1WBfvab77RtbUr1tUUjveY9+8xE6u6YK4H/7CPEyk/JvLHELSSTIINzRcvZedVPw
VSta3s9ope3PoLGPCfBIUi/l0kk4zdmP93e4ojwyR1Q0KjPyBhzrG02UKihDxZwK
R/BDqKmCL8MNXTOCJJ/3a6krQYAP53QEfOcXfVW0RDvPiVl67iVKReBXJfagnCYf
8CG09R76mC5OX86qQ3weTJbmKszsdPqOVkMhRCdYt0vpVo5GyClHdXQ5VoBMxn8l
u8mpFAetv7f0TNo0+2BlpZ9GVGxOHXr/7lbuaXQ75HkjkxBsc+kzgBItJTBo6SJW
cgoJzE5QtZLQVD4+DvY0mz/QdsbMNF8Xs/4aedMsJM4GVty404bVmiT9Lpo2IK4Q
n5yXTtQDYd3It84LPeKoLfAEQsCDNVsPqza08eLl4V1oBjGV/pWYkVRL7h3ZtBE7
ccNDEJreLCP+xnobL52DbUJhPggLWUVHXHYhqGknMOCgUNz2NwUGPjIwg83n0J5F
Uih+E8aAv+6Aa2p1No79MX6pGlHbMf/QpC4XumQRtVUG8mZs09RCDCBMXdHcD7yG
9aN9iqjYEL9m43mbcUZgbjODk2zBOVBasBhW6KcLmWnRiiEHCVAng74nvHoHpIrO
NZw61vw/aqkIhfsR7li7FTXG4/xwrfFUGxHX0gxFo+hEjUsjpld9HjYmOrlbMsdj
gaFOqfJY2Hch7H484c5xJf+c5L/u4y8+PFzoJB/AR425QsLTL/DwFO15zrsB6mPu
fO91rkc47zTC2fWYq8Y25xeUqxb/CMO2ingzHMswdHhFWBt9Mkaq3mOyl1TRxZEl
6BTfn2rYUnkn+IvhC1lpudPKPk0x//MTvZ6iHA1Va+ji0brEu9+/CooOCIQ9mrFJ
dCe0OdKdW4wE8JhWbPaLCy+mZ3P8jEM913F+30Im8B+l7o0sf3V4qW6yN1FJP3EZ
myb3gpnff47kDX+/DbcRDuhJ93VJKG1xLz7kNCNj9FFI98tk7y3nc8kVpS8ie0UL
HoLfLCVJ7d5ZDyzRNjca7PRBm4zfrkcxQi72kPBnS+MhqfHTfM7AEk7a2x0MlEgJ
L0SvAxefFNi0fbA3nx1QHLA3p32Z33OFNjxqDSh0VjQ79cr/le6jqh9tOCS4FxpW
P1sqA4LbI3cBNlfAmZtvhwJnVLNFKZLOoxNk+FIGkaPGzQp9L/CZsCVgKf7vAmqV
nghqmCKC8DwjH5357UTqCSUk3e1u2P+TKTIwPGOJ6wQIM/lZ4L7fBtY9QoFRny0a
gvGBYOTIHE+n+Lqj61MFPDyVtJ8kexPs+r4wbKv8qu2RWp+OEG+PWxM8YLIO+VcF
9fY6GyQWDyxAFcvBYCOCE19lQmyPIeiOX8gjE2P9toQKA/wet1PrQLhuGigOu8Wp
g0Ey6RYtkpRm3V7XEm03fVR60Z9A55TXsOi6/aa3JwfGZwlkqFSAJYTqPO7mhvvp
HF5d3hZAL0Y16u1JLJGP8uQZK9p4A3Ju6o+5YjhREUNJgb1GNDWVDNDeG5DO4QDl
33GPf3daRGw4z4Aj3lJt8/XAiG5dTqzm+CWpyE5OXldGjhmhlhcdwzMhXeKPOQJ/
QVCM8u9+z/Of1P5TXdgjE/Zm6nBBwNrlhZttzztfBBd6VQ2/HJlGetInPyL3jetC
mHhtoE1qpPnYUZXH7KUQypbIPY2OCkcY4+0zFrTr/gapruwiHEBxBM7Ky+w4oq48
lLD8QBzgvqLIat9/ZNwOePHTTLZj14EqNJl79wEYLJtHyGF+D0+zSJQSlJP0y7vL
soZn2uUbA9zXznrsbF9TUxXxzxS/m//Ri06FJS91jyKEHWmW9HS0v2vx8Z/Po25Q
lZpbjhL9vcvxNtww/NB200DGf4ogoudH6S6JUMcUAu/+P+OjGKbYA5oBcjWTNNIM
yjNnMd2/Hqbo9pI4ygcI7/t6YnvOTa16ZlMbLKYvX7pkbSDMaVqrNXZ6h/MtIk5m
uK960TTifs6pWyomHCIejOV4pVl3B7VR7gmAwqKDMFbGpkFV6Q9GeDtmceJg2gOd
UDjQ2wZI8Ox6rIHX+I35wEwMAz4TRsOsVmepZhWttB3fji2D0wUkOG4PBqqwuQIW
qO/13S3Qwvz01Qq6uO9t6qjEQmhmijabpUg6rMfSm8cyNDbiZZ8gNMiSy0+mXJSu
+MVQuMGWBFgTwJOcKYEP4eN6qbyDnLfeLKMeFNYmrhJUMADiJD44RTlchBM57PzV
+WKvCByYMYkw8mStnTErayrxlV4AYU2KlMyP7KU603ZErKKT3KdOTIfgmozgQumv
AVD/l6kA1vok5TXFdqcgzoyA86hp6o4Vls2uu60rhQy8MXYs6Xw69tPu3mWtNaQy
sZxIRfYRKkr8GRb+1cr59CzMZXC39rxQ36hnIpid0dyIjumm2frcmPtzRk3Nav/n
Sv9JxR22LdqTTsrkV+abamecGqIGc82oqT8CrvvLGF0oCjKnyV6W8GnES5Zc1fWP
LCAUNVNQaNTUnTCo8Lseg3EtjoVPTBlJgzVLUDtv9Gk2y8qT7kyWb5Tkf8Ke/2Dd
uY9oTuAQCdR3/1meObIFayfYQYtRsQd6/PDteH0qjBke8JwX+rXhYtPVSPWmc3y0
5mFU23Wu9e+jdYPd+tC2dAJr0x1XYIEPDQx15t645JoDiwc+VATJW6iKT3EZ2Vmw
YoLNBizV9rM9FmJ9HyVzn3MtVZNHD5YieHkR4G5EUtiFNIHd4EY4UzWAyoYb4iTZ
8tkJD3VGAYSDZaG7Qs48LUsRAk00keHQH66hx4KDtdmm5NUavsrqDD+C+hJqRTSJ
ZlFHULjHaFs73o07ee1bOMohgNycJiV9YlVa3XcIhYrUVFnebevyIPwNA2tYdOnI
GWhSP2G/V7sBSGc0hdjuh2TbHi3venWQI9IDsrC+JkE6/3BrpkkTQsTKkWMRKeky
XROO3CYkWtQ1zCn9yd7F+LO95rZQdhPg15UIMJylgaDimGrSpnCx35dLf5Z6uh38
QTVpJiCcqc5EYYG3ldT9n21DufXheUaJPyR06jSwJ5xDVtDh68PcHGjXNScgz/8Z
uWoZgg9TWzXBRqOr+tBYuJ1IOgp4z/qSMMZgGEtGv/duEWDahLvRnuIYe3RevK3f
Zlw6xNOH5813VI1ZxXPoOUfTJjRhc5ZtEDD0PE7HRSbtBnxgBCTZZ2fLa0WnV+cf
dXGlxFAXKbDQvjAn3LV/ebvJNCr4vq7d3NqaOxKe6pJhp2kMreyr9oq9AfYTHAHX
DUhP7CPm15oWkww2ZFJbzFzEqkYl6pkhaa3e13mqPXxdftIFZ9ac/tRD0E9NcYpE
VHLiqzIX6IHYkDS+BpEYZe8RfA4E/rIeRHzhk8ZPJLlEN1yqZp8uuo2vJVOb6lj1
WJ8Rsz6WE2k7iKiPSDS5yH1SB57T7jmO8z/xs2ID4qDvuDJ+JcDqMfoQ36OIsOTY
Zqp0o1gCZc36aAhvvJK3Et6jjXm8OkA4NxEAo8vV8FVpOypW5cDRTqSuEYwwBMTl
b/EopFZoNaYJV6koSG0nGcEs86IwlTadvx7sj2SWETMM5HxvkFH1/KP4Spf0rFGk
7VhBY68sO7SK7ieBw+3nl6qTo/7RmMcKO6FnVKgXiVnHp60f4HnsEF+6gzLy8Vcm
g/Vqx2aN0j2ZeJbZ65YvyJjzrp/0YGneLBh9FcifrCthRF1QAercE9a8hOX3TU9Q
69BtL1Vhor6Lc6jgdC8ZJ3nnkYYK1X/8H+bhtthmDbyNO/gXAaKYWJ9fwZOODo0A
LDGDT4uhzHybyww56+/qh25OzblX6I9FVyoGWsdr7dCuDmbXyxRphgwVXle+mRtV
MK7K2hqa+aPog47CKGNfKMXMGrjpobebdFZ0GGyYOrQMKiLFULYqq5NCJSJf6XSm
Rl4bjo/cTrdiKu0gDObOoRx7dV8NEp1YgaggW0aHgMkwADSQkkTrpYfJySaXtJos
lOqizSVJSyWJuH3xSIK7vriB1JeJWZud4kcRlEmSSqYlxbCoottS3gVSXRpridh4
K78v+1MIFwIENMFTX6mfuIE8BwCvvrQtZXjHyXu/Vs9Kv7kKXt8zw7vFZwIhvUCc
qOigE6SJU7+IH/jiX9a9bmY++RAf+nVKz/7R203kBScYc76ymmZwRtwoAzLZA268
pXW0XE5YBy9XMxC8g1CEcLlEGJvUqd5SF/7kI7vuwmVkyPWaN2MrtDovEWNTc54g
Xg1Z65VvwMN6wpXAM+/99PBzFQZUKLtSoyDUWcgj0G8mfnNdqumBE3pqXyu7sUND
gnXq65tB1PeriYj7yogSjCM78Fl4eg8zukRKmRMQqqawhZWIQC7gCtjpNxiOGQyk
G0lG9XDCeqCnelC1W/L4ILNHkCudoJvycKJHdB4EN4hysAU/PEP1Au6jkXqwIAaM
1dAVTeBChJSNX5BicP6/GEyl/TC8nSUmi1WtC0wnYb2rVHEvuo6c/VDyvkRFgu5j
WRzewqvEvOqpbopT7x7U9sHRi0syzLYFkhmYGTSN+kg99ViMYOLcDBtvZ/TEOjek
5ZQciaSCsoVXSM3e4kYAAgUaR3CW4KIyDbIUrA/SVMPsAJvl9vqSc8XX8uWC0mco
RGV275Invusexz2zsrIok31y0C1Ckdj3qUa487q2YuhWU/Vij8hV5BPuBcKMTJHL
acN76MPlFGrxGqVMMkJt39bN9kUojO3Nn1wYnwzJB7NBKqTXVVmTZc8NqfcQYIu/
CSHhbREeJqMtqPTrib9Ddzm7m2Hjk9JZEC72oiuALGuBRoCV6LhhVsIFFGHhDx27
EAf7WFgdNryq7lXt/ExzwY3gHT8mHxxqLp6zB1rzZIh4UCbJeC2pz1oYcLxGRQXg
PxSqZxMU2ulkC2m0bjyr/SfwvSFBS6RDgpLpdEPmb5C3XPAcT6cSK3pSFsdIKQry
OAhKjBC7a5D8Y4b1YzO1h+UYfXfHj4CbEZ8U6xJXqAXi0FEhD6EUA+YZ5Y4WdFh3
dxYMjGkfXOagwnLJypSawddMYuuS8S/JL2X3Wt4sNYFP3DVGZtmUjjVLew0RbT62
bMg+TL0eYCqfP+eqHq92C33h0jh+Qb7q6qsMpIFYu7M=
//pragma protect end_data_block
//pragma protect digest_block
cT+souddZwNjCg1Gteb3wHTOw7c=
//pragma protect end_digest_block
//pragma protect end_protected

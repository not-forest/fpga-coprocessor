// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
BTQVPvIQAjONtIku/aa+3kqwPMnmogl9JtKQNQDja7NQdaIKAUdg2LBlZ8/jhgsAQOZdtUmDblzp
309Rvh/ChXj6vdO0NeXejBweTrps4rim/r+Aj4dpOPr/wTERZAo0XI9c0gcRWzPtciFleDQJnIkS
t3sMHQuxqINj5KzkU028y0BaNWi8RCKuffcx65oaRixfxSofYSApgmGX3miLAdtlEImHIbin1GM3
8M5Et3EjSp+6ZyViba8KDtJbcH/Z2S2X4dR02ZmhptS2axR/2PvfCrQTGWGIGsjrrTlS2Qk/EjD8
8Jsz1kpPmxI/tdOteSlHDvskUwOTdAH9LqZMFw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 36736)
GgWJ0WKwRExnivVp2FbvAzajq1bF7s/CZTNjWkEiqRH00ZhOOBtyMvrHe75SQhG6S6bdrLDPD2Vs
YTwnrXnPbtcT5ncLSKKqiWV0WG1Fx8UZVm5Tl+lwxAppDZZcNGko0unSo1L9g5e4MmvATK54dmT/
77vSA8NM2hUgjCaTuy8CZuDxNmvtndRZE1hxB6VM7gHO3qxDjqqgvDm/PVZx0J293Re2HdC5M5LH
1nV+n66T8cIHH4+j4o3GWWGJ+v80Z3NEs5aKoTXRq15Rl0sXpZoxehSW6F7FlMP3NsXXzW+oAtUz
04VnLCtXXcNSNtepQh1JnD7h9obwSisFF1voWTZ7KER+Mb3C2krVJmpsR65iY78U0nfRDG7i+kvM
qcf7nmPOpwF0GVTEdCj7GPk+5CZYXuon1/l9sgx+s2xXCbUMWpakbACvbO18oT4IjhQmEaQgz7Zd
8+JVE9p9eRW3e7KvUzZBKXxFc5FuIlDJEPPn53nRNRY2V3Ge4oZlGFB7ZZ/lSPwNCYLnG2wJKx95
Fym703eFBk7gc1F4XtUsQbInbcxJsWEWHZD9PTNGZTfkhhXnsl7yyoXC9FAJjp0xXfHCKJeBGRdO
QgnOdw8ghIzf6I6Ie6MxR4WD1YYCdRBx/f4K0rpZlB7E3C6PavGCgqT/qrC0XbHBTE6OcC+o1x3D
o3FsW7TEGCwlYwYr2F2DJUVhPVMhgMM797tP4kADNEwF/d0CllBsKH5Yh5EKnBDYFbvxE0UWjXCY
ET3owtRkcXcToTfJMAwVXIeh/AvQH1dWBhcB37/YIL8bJ6AsbrL9JQYwmSFXtpaBwf1TZoS0BfSV
KRnTpOH7uF9BZTJaMhnben8c0k+Y5gTWyihxg3Gwm/cSpoyuB6sSkDhSdWlCs4WQCjBZ8zhWUh3d
wL130YOFpZu49o5dJoQBDHOKj0weIwJY5oNbDWDMXaTPxPlfm69gjj/NAeSbqP2c5NL0L1ZpPmZx
fvb3fjDAcb9XxGUOf2e6xvufMJBRw7lTNKln6ibJbGDX2+ADp5APHrht0ERb7Jx/7h1JQ9ENNiAz
1uVKSGp1SSnaX2pwfBAeRebAko1M7uPV9UTOlYmMRKLb+auoNGWBBJPtVsnhN04phK1w9is3DJre
DGxfgFbjaD5nvaYgCToAPpshmNvOYOYM6zXIDBF2hgBdnpRGBbiTU4oM/qnM89mIg6aITOJQhdIy
mar+6VB3efiDsEwLuaBxK10f9QLFopTY76jtac4SYnxT6jI907UauG8sRpvrrahA0KEWtVjHEH1a
Nx3M2VKW83MTZNPk2zffvsYzcUSyyU9bHR1qG8puktY/i3iuDn1E7DvyxiM7amorFt8pYR8HZz2e
deK0Wm3uWQUtGcMQDqM9t5VA93ix/YZFeBAFeZhVzbzJmOU7mJzYiK6w5DqrIetsxGnNdXkkP8OE
FHnkWaNeRtypuyLaKt8YPgiokxnZzTK392WgYOxU+j61ZGzaW+n7/q0la9Sah07D38cQ+OQWiksr
N9KnIIvgVw3Xx3RuqixIcfc9YdqtrRP+5KOP/84A1RwGOlLKlmllFlhMcru279OyZY7Rp+5pCZx0
OA8/c+INTtcXGwAdwsiufopaIwxvNAJl2RPtdnItYQPGIiGWR/kpGti1HOK+Jjt2Di4+wWoraeiG
zmkwmXIeOwYxgMoTXDjKiFemqb18yJkldjp0+/YKwLjuV6tOgLHhmQm5l9+neiUFfHmVjQ7t6qx/
DEQesajWhg+PLP41SOux7oUPCSIWYu/vD298Ncg0zuXoFE2jYH7FQmmo51WPtTuC7EpITu/xVxgp
/OF9nvR3KLMbDOeSBdeMBG1hQM66t68u1Vf/hHtTKTcPEniWIDiCMQHN+zFP3NYuPnLe2is6cHpM
I9cLpWD8DZzkxczbF7qmfnpdRQczz3BqWnJ8MNVVZpqkBCjg/3neCgMwbMFzeET9CBg/iGjnFp9h
HkwTH/t6z4c1nc3NOf23JTyEicz/O+JupDJ0g3xBPstxkgi2mx9r+e1JdHLwsSiM/jKlMZ3uJST1
G9yMuQK8KFHJqH41sVjZauJlIXPWeYa4kWsXS3x8waRBWIyGNoT+XIobGlqtA4ise3vA76sOTKUz
BCOKMt8kToKbmNHiucw87CqZNgxCdQ14C1Oyf91SZPpqrU2XsL4kaAUZsYR4p0z9mYQDRwOKSVsR
7iiC2KuBZlvWNWjK+aU5vz0odvHJCO70czKv0XTxNknMC8nwcboN6IdbW9BsOLLA1qegZNm7DQWN
HCFyOdOE0x1EOujkOck/HJ5DDuPnpKuVa69AO0vpKuX7Srt8BjsHt5lxgNmxgRhO8JA4tR8fZscE
vJ2IL69PMO1xArefW6bvKERlCa6nxw1F7vLFdmifDRg624wPZM+wYi9gtXWfbh6ZVb1inOz2kBHj
PfH/R4GBlJ7tqcW6Oqa0rYuwwa+5aA2EKBGEtJ2xCUkcI57t+DgHQ+Yvf2ENzA+yy1Z2goQ1uAIB
FDz64QWhj6kN0om3N8QT8Ih/EaCayToLcJ8S5LvGD8FyAkQ9PnfzZpuekMIAEwW+TcuxfnbQJr1p
X90CfTTQiN9wnfKWSI2HLIPahIxtDfsWdzu5birWl2vsi1j/ddc8cbj0y4bRs1C/1ouawYNNZaBZ
E3skAyFUinKN0HYYuJf3wzyglWBnpkogtT2C2XQhY4yVbAlORmwMBomobjcUHPNuQ+7ajJeqZ2uP
1I7meBOR+jKZ3TFxjKglB03/FOX9XVrnpq4EZkD+SZff8ZWY2KQ32/T96h+XNMXsSMGEOwjBrPVH
KpMUNK6gLJZeoaOc4L5NB6fA1v8tsmI7wQbOZzkSoW3mh9u0HCmpsF7lZemmjPsNQzfWVqKHx3LX
AU5Z5Rb0pzg3vyrEua+rLvGR+jQmpr18KMYmVi4ZZh9V/4wqLQ04cmQHGXmdFrUUb8qWb7dNQmkf
SXQXyfajVG00Emz2sncJb6T9cyiWvMfvzjOB8sPiqiWwzHe673wUjQR8+MgFaV0HRvgTKCjI8m/K
oyATRWEgOYEorkn/aZwTsxnDiNhNomd6Y4kRbikiKfnJvw1L7XdioyVG0h/8WsyvLA85FwTknjYX
0nXvbNNeL65u2ochbIUjtWe3yuoG21cFdSbE0jWoZi9AI9dViDyg/OaMqC+TiVZ80qkNKfKH5b5g
vpDmps/SzKPPFPvQpwel0tF95j5QDNXrjQrIn02jSE3qeveRzRp2kR5AP0p3d9UmIwmLXUWFe9zM
Guq6CLT7DEVGkdw9TA3Otzzja0oBdskVS4grTK/5d6W37AmXjHDQd3o3Vks15TruGuDXhfSB6z0n
GgK0dDCI52FqcV7kzhjhQpRjdx64mGkxAsbeBqb7eqMgGB8b8CL0jDJXsRlJ9UTAoVhwjHbb/fAk
K7auB+IpaTUeEfNHg7zALVvMl632DoPc6tOQ2g5cy1/QRlhwlbVCiolp9Bo/61k7P9Bvopr4uNT3
XHEVJNLys4/KFLScIZ6DTtCvFfk1oOVL9bFkR8ZuU6Y3P09kVEPf+noUIT1dBMychSGxeZeWDggE
jpyKnQPc+a5hKJMxJ1hoTXRHFMHO+cUmZcci43sbVpbXDgpCRIaXWYljTafUDNqiYT8E1KYmz4p7
dAZ38yPAOyoWzZZaQw8urGjV4kAezc6keU8VH/M/8SQDW/oEY84ZofcpZ4qjWWsvuv2VQtw+HfM3
EkziKmEDDYCmHnNUYRlWupn2qunKgxrXyam/X7y7LbfweJtnw/3jFoG5xlxDN1ifTTC0oCKEQBmB
l+LldF11dnGIZ8fe5xtMGWw12OuhZOVg3B6MwdswH8rrSUlvp0NfjbpVNQToutasqCeNqWYgX1SR
qHbjCjjE3l87c8kkyCgnlMa43++jupEFIbNftrIrmw8y3wqXTTFtfKehMMnUfsw5icKMXIKoRKtN
kUrFvJQcnOdylzcSk6G3BzXZRWiN8kJALj+kQQ89/1V9M7WJgTDNikEcHHFYM/D/J/8UOn+mlsCz
8sJhKOQtStdd1AiUe4Hc3dUWzrWaOhTs/xHpW1i5WWQY4AbunD4DYTpjtf5ZZfreubByP1RmKQaL
BQhmh13AG0xJixM3M/7N6dXbWscIRSZ3okgDM9UlEP2/br5Pk0KIzR9Hez6TUEmw6PRro41GNZtE
bJer3P53byHo8yxTyVYrYKRnR7bqTrOgbZq0DBzh/Ax5R0DchtsUajtfEj3XZw1KxqhxcwxTOr0U
Yt1NKrXO5ng5PViv2JEjNZG3ABj5YHJl13ym5F8ok9jbkysy1UkhQBKCAb3D5fWYm0KLg4sT0kjY
EXW9YrW7IC9sawkhK46VabPaNc8cQMCrjdrYXU8ppWDuqx2yS/Hg8bFruqDoXFW+CAPI4TAjnyLa
dRUB6UiSKX6ESpNHx7/JYrkk0bZ1F8A203IoLWv/0nbL+N5fkRdwtDRvSvKiXk1jpkJjP3j2ER43
u4+UfF+Ve+j+77xOy9zJgfwlr9/ueqBMGd651pTrmRFVmoOqygqG30xKle456yUTs2AULiyf/fMH
IMvbJ9ulgEX/GmVyo59lFoHGG2Q+IL++2tjF0AvUuHyosXU0YVBrqTGF5pD0sqG+BEDU1dWRrzHA
ji3GNvQXYxxZatMWzCIPocWwOlcCdeYjjqh0SJsPJzftrf7ag79i0gA6Cklut5ZsdW9uH3/w9bSQ
/Efn7rBOMZ9fQZ8ueOyUa03VM2XbvVtgnATtRXVOWwwukY6ObcuCFSdzXZJKAv8foOFAtHLIscGJ
gTaM7PFVxR/QdWxiDtf7paWQk5iSkW/aC7WDBkzE6hbrlz8lD7LyttnnA30lzx4ARRTct75oC1b/
yXnvDLKAC9E5p6sh++eu8CUWPec7wr/R81KAhQynSwkQ84zXkrvetezblLxWt3C2NLnsca9Aw+Ws
SXePqczhM0aW4CYTM7QVDS7C6YJODMs6Zx03ZkO7CzynitVMFDCjAzfNPvIhQGgRkoJG4G87AYGl
mmVvFsuyzhD6N6dnvA9T2ExuRFUGQa1Uz6bjNedS4wiyw8HZ8LcU4Am6scGvQtcIidEBVFiQpUZc
mfA9Xi/k4Ih8gVY70/HwU2NqY2265OdgLUJtbdymFXtRB1qZ/pgVAc3Xdiko9Sgmb0aICsBIi7Pi
wDfI0Je5N3YALuoB7LxOPsfgUTbKn2dtHuVK76a947fMGSbxTv2+9QysRTCsLybBSqjLLQIqQVbK
C+YQ45JcRdvxGeECBS9nFnGtjqlnltjM218NcFhpLzB7dLKjSFU5HkWYvGnjHimeBWOnbPcIDtuH
mDEUhucJR6YB+iKNxtsbft5HaFeB5vTrsiJaHPlKrcjuS6mw4wPenwLVgeP9nO23njLkAeNVIyIW
lu2KqVAajCN1dMGSkDoin3hNMUOOBRZWmQBB9OOWd4+KGWRmEFMkL2vPtHrBpyh7C1IeNSvS3Nre
qEDhFlBr2JwCjhYI7HxGvUANDkmHTooAg9OVGbCVoMtYY4E3T9aNdh8Zkw5bCWg+xN6kPdMTj5lO
BUU3bsuHi/5XK66A+SAtX5hPjdWso0X3eXUAySygC/GNq2jvt9UStb2lIr1gnBdyiAqKd4O3RJ8i
xBLvF//PVYixYtSf9MaA78uvKgYvdp+wwvAR1CENSg36bOVrgUF75hiq2xvkT+X5ut7gPJPBxV2V
ptnfEl5gFHY6+obJ76BxrC1bYNO9T+FVYSW/Sm57pBJIZ+9taPILW+lpUXXVszm+aXHmja5A/4mR
AlHMQWGP15xC6q6W9C3c75F64sjRoM5iKzBLRH/zvX3+Lcj6rBbCWvgkUJV2yRvylfA5EOxjcLQT
A2nx7S5UtYpKsQDggtn2Rqfvlrcxd+DAqw/u9Jg/YAzB6KhivaMdd43nXx2bPJzUAnL1zR3MfWrK
ARHyeu2hYczJ5RyP1qcs9RbJRABfytjbyzss5XA9EdWs756Ul3RBOvVw+xYB9mjxGKf6rV8AT9/R
m5/Z3/2UOyZBA24hYuUW+24UnsUtcDZXcJlPptdFzCMBeKHuTgO2tDb91yvkD1xV8YUO853mj2r+
Ga/GSiWVuXe5D6kNUMEs58HPxk2UhpocgO1HsNUbK7B8O4g3Ba+WTZR/JaX3PhB7cBfcnheDw6DG
ZpDG1VUFp+DB6zq++wAQGMsTA35OIX/CdeTooucbkhsnQI2rNl386hq3bEQD7S+xDGnVanzvGW/a
1Yc5JFdU8Imj7QaAuo5NM0AELGu0mzeBU9ZpBENz9wkK6qyxcChGa1en8nEYNYV0JTNc4D7W5BzX
GLebBtw3c/PeJmjtO4gxfwgUCuM/OT8L5KX47u3R9cbiAy6IzzEoq9zYNKlptb4PXI2umBDKdz8L
U7+Uc8UL7Iy2WnLii0+HlW44sXaq4/9uWSij/JncOI1bQZx2YT5dqp5HxL4CukSz96D11mhNhftd
4Ev4ogJwRsIavfgim4UB/VUwwKFDWsFvMtgidchyHd+Yqcvf84xzE5G4ULfaj8dBlmDDpMfnesBS
gM9YSa1aINM00r2ADH8puXWVWbeagmmMhS7NikmLQtMbd7PUlMuMBJWw4QGKNDa3xb5vpB2klttM
xEjJlmDSkaxISSDF5xnmJFpzaPL7laQHYR2nOMYgkv5e4MUAbRYRstCTc8qoYVZ14Y8bakgwJAuY
OmNrPMJ+mRNURPpYIkYsqVWiDPt9jc5zg5AroDYzt5CfQfb6Nw0jSYWcTaMyhEr1Zq/VWiMtnQiN
PUTiqelSGvSUAp6EBiTwru15BSIUvq49deArEkgUoOu7vk7v82qyvMdGt12kVzin2YBwq0KyaXx+
RuXfEDNuSdQPrjuE7+HYrY2S+7I677QFXQNnsQ5pnUdqD8ktxKvRnY/9gp1kT1c9AlO7em8AUL7D
ZnqTA0GjV7fM2B7FEm0NWDsM8pl+kO3i4AErxN+lvz6XZ0UgEjpyRFA/8CTy3nYxEzZXaGAfKqTI
rAV+0Z06ZPpa7c4r/ynat/UYdf4mE1ILthgrHH9SWEsm7M5HF9EU8oR72K9UzTwgXSqNBSI9WyuK
pMNJ9uZrhimrGSl6XIRMwUZ6Z/SG1p3S6U8I8Ut+8yD97bJwyvnovrx09PB2zPdvZWecleTv3T7U
WhYwNeUVnXN3QE24wsuXqElSdWwn1YoNJ6pNbS+0eTsnMPxmeBJU3sEtL+oqNN4H//8iOtfshzDn
roqBlXdZ1HlDSiz6Ft7BU8an0/VGMQhvZOXxj03c+9stlohpHgTqcUjsTtPIHrY5ieuvw2zSA94r
J/TgqcP6IqN82D3PHkmlc4u8ElThS0boaWuik3b07fuNgBf44y+Hbzb6B7dwDyywUBIkbKhLkOYd
q7+pk5UZIGcw6V2XWQ2pRm6kxm0mydLanMUEAVmTSAgi+S3crEev1Lv93xevWBKXKw9Li6TlWL0J
aoE5MLimf8vp2efw3lu73o6NXf64ZLvsEw36/OBCogIf12sVGbe5JIC4J+Yq6OLxdnIelhLbzpuk
IlMkUH3q3e2Z5C5OoYCFB9ofT5myuDhScilrS0HK9kB9sIHaOF5NNEzxqZK+9Qgz6iVEJlM9Y3F3
T1Y/B/VeTtSv6KRiGWQXFDEyrIvJyGW3KypjCbltKcJ4ZWSxGZ8/biR7bKHsu4iUJN9SEugGFnt7
y41rXZdcirJY4ICNxdv2LUda6BY5qpyvTU1V1AdTQ9OwoQdXqy+XuFJ1HMDlz6r9rOKtuiiifPGR
tcZua5XreFU7ef6pP9DCnnnd+aoIMtvN1NMLHJD9LhT3TcfqQsv8ciVt6AlQQ5q1lj6C+zVChczP
4gJCQntj4BvER5re7G9QgGC24mFHIZLvF41WGky7mFKI1n0h5qREQxTH/hiVClOTbl4c0TlpWEYZ
9pWvCpfaG2HkpLYKJWcaU5919VQm+NKJpk0LAZSwTmxIIlRWWeuLEd75H4qxWvY3casUD9Xzt0uZ
4FCqtLdRmmqOn/VNSv+yAGKxgUolEuG3keZlDi7c91FyZhvV+JnhnFItyi1q77qeLww0iYqCLZIm
4vOmcpgt03tmvgF7LjPADwhWDNOb4HfhYQ/VMqY22Lqd0+00KPEXl4m1ioc5gdr5k6E+W2QwqHbz
NP4FcIBqhHNdyivACXCf9x4H8djbWycdem7kLnQ9glgDao31Sca3K0FFMzYCmOS91911FoE16TBL
hUdFZrpF9AIUoot1Reh6lBYL92fOZ+zLPVZvHSBmJhkfelkn4Qmoy2vpCNw5h2MuzEczBi7XvgSv
CE/n6X22qGZYyW5iezcyJ666rPJvYUBpanK2I3c2CChXNGE015ENBdrkwpxA1kwjzC2GcVp+4xaG
perK2E/yafeebCH7TEwUTiZKtafMcF0pzJdD+jpcH12KTZTlp5V3YEtV+Vr33t7m41EqQ1/xTjYZ
b+h0Fo3ziR6RqWGyglmf3AWG76GdTLBtwSyZocSKOoYpAQE324r2t5uCkZ2q3qr7JokXpvw27TVi
olauNpNlXCSzADbuMagW3XvztKn1KRcA9EmIjzUZVb4GnJOWV+7bLBS1zQ/m9w6p9NU3OxAdNWGl
91i7D44eI2O5GdB8j6h9SXkgny/S6y4GstRksMMsS4EIJk92DjyeVwVOdwjYnSVtMEYS7qhkAI7O
NZqiJLs8iD8rJyaF2stzOSzv5LlmVur+yIkp78mSymcPI4CKaXUwRTZyohe9OOaTkqmeRa7QsffB
ZRCvIHzOsVJwoz6r/8yGyhmFQBtNul/sEQZym7fQMNrlpzAkof6bPJBPi7KZqZh2TyoEsID0+Khd
p27/E8C8ozalrKp9SuGwViqvmFva8YBcrjJ7wWs5AUwjE4Ro9spAe78WO19+Xq1KmIwngnvafkv7
IaKN0LlmzwZTNIPPddX2Qjvdgb6NRui7NwPdF8LXeghX5HTruF8YSOg4wDEETSNny7BV9LNXtQ41
MKVymA01siDTVYUYJuwLpmnCJD/PQYxr0dy+Ksw/5obatO5JoO3ovJMEOJwYaLeFOafJBJHzKagW
AllGT01dCcl947ozODgUl0ZKHFUt74q1Utrx+onXHUKvH4EtJYF6mi21hFHAf0+k/f10zsNyMrA8
2lxVXPGqjglELbtimN3d1l1ame+ZpXmkuz6XRhDclMhHv4dS7PwGLsxuzVoYU8LEBmBR87l32kc5
nIW20VjsiETtABYy+VAM/L4ovSvnDu+GM72/KN/LLq67KIPL06tq9/W+V6oPkx5oSCIl3VK4n4Bi
/A4EgVoenQYkJ/l0lciIMpobvtgABA7c9Wz8UOdopQGkZOBzksse8hYkECQpN90w5GUsDjpAMH8s
T8irDmjUD/KSTPILKt8saaONVDWPN8PJhbCXMmfZnrqW3aQ4D7U3xanzZvBmKUkE8gDIg4CUF0r/
xITi13BZiJrVjSIq0avEHDoDtRG1UAqng44gR8m8XqU0hX7QKSsSlv1Syu/TDifKabg5FQqYIiQf
1LeBM6wlDZjKQtgyoUTEh25VqL+HLlAZS+4ueQ26bt5YghqCc5vMl5nRkozPIceqPo21yrURamVj
GK962MT6tztlz4REJVJVmI6iqVBwnOZDikpIyEvXagy30jT/toWv3Fjh4CfK06ZKvxJHDl1hAXbg
mIIxYVc3QgbKcN0opS+tOVrRq2tdJeNOSASWCGoq69PbesoAwWEVwg04TvDbv02xTBEDqu/88riA
11ooXkpoYyReAFUv0r0SD76XSJ0pqiTbu98oF4MLsFTfh3gwN14laNC4tcbZDtf2KJQr5i4/181k
NknpIN6UEBGcR8WFI2K75EX7EoA8cg/NSMkf/j84QU6zrP4YJMakQVGgwncNUw3F9HHFTipl8CL/
0vdNgZ6OibpXRdmodCbhUdbsepp7Xv9AMvIccPQrZ2QH6PFItpLEBJJoJAVyUnqAmK9m8rTwT7ND
l7czsldTqY9H86SSvTZnNTqbrkLBVnKbCjAzzrN6s8vCkJbMusH7+v+++SLHcuxsuJurwMb+7Tqy
Bw4nqgmY1VY/KHImk+COoS3AzwZLdDF/q/HmJyrxepFl1iZ48sF+YglPuc75yhCnbonR0lIszXBq
6IEyYGJt0zKWbGzeDvgZh40PRIuLloFskRoII4krJUL8UE9JGWdurNr1G4stPjFQ/8M0dQ+1mFEh
VH4oq90rsffXz63DpSQ1zBGM1rMl6LByuRkK3JzN48nwrar1i4EuNYOOiPjAT+e6Kn+y8AiqkajC
FWnFN04BV5sB3SGlWC08p2AcMpsLXOlEw/WrAroKckeiZMXygD5sjk1lBwocEjONWE7/soacANzd
H4MsSoCW+oJkk1BuewM1LuT0x5A9a6SPJNZlHHR4gJlBx0T7Lh/jPXWXf6n17XcgmmoyCmQ3Aboc
suB6XhO2pr0imG8tzcVn9I0dbZt8Mryg+CXI2iFhjqr5k87377cPUvoLjOWzfC1ADfRWe8oEwQoZ
I43AVEKR5AVXBcx5YsH/PBtGZSOEH0cUVbFA78bdAriFq/JvdPhGYXhhk+W63Ne8x6mmIii3kBOC
8QlqT50T87fBfy3xngQ20tec9iVCmWCEMfOJNzwcYcnatBUiMMexNrVgQRPqLYc0oAohO+uofr2r
xbRx3yRK2cs713rBubiOKebO6dvhtMuBQM0cY38UairyaGjmoK321shRc0p8CKlN1jpUZBJ8FYMn
+okeqlqncXO8JWOdpcGthYiQVf/jPCX4vm7F7zhoeLJ1XhiAC/neHuSrDF/q+N0qZytOuF1cdgFs
esv0clmS4zbUxYLRjkVywENCLsoXuzWTkGp7ZgGoZu69pw6nbJbq2+yHvxXNzKqIgqU+15KC/pO7
GJLLGaN349G41etkNE8iDg5qUjFSpoWO/umFDtEwkmLEyb8ox7i2LdLZNAexWkpdqsb60FrhapAv
6AXGDNidcHOahwkGvbzg/qE5KhVLnLi3PwP2GKJdKPENfk6oxJUpfbqzicUDRCK62yOWTO5R7o5h
7rBTpdkiRmVtFMZdsLggSSjUiSXvrNuGzHd0Rqk+ezvmfg5BqLbzCztDZzE2XBU4hWDCB1XidsLZ
IV1/J4+830kNEg9G34RYn0oCfhA73xTrOBKNgYMK+A6UIHIy2ubt8K6btOkIrSXxuuQ111Pvs0UU
3k9mCw49wS+anxPwMsti1DFNPlyVu1S+hxLj//pcwpOeNxJXouKTB2GWn7spzLhlZLHDgb5DOnR3
UzpeR02Aik81bfpMXBzQlbc0jYm+9OB3DFU3NPo4Wlx0NqDYuexZ6Aznhi0+g/TsAce2hw1KgfJz
Pu8qZsq8mOrHo2N+F7+m8IKOoaBvmOueJfKHuG+Y0qWyvvYiloSiqDN0DKyiapH7ZXTlejHPdVLa
8IH5rb38nvqmvrj97A7Ik0upxc3gM4D/VyQDxUKAgz5Q1HZf7fc31qh0+lcynwj/5vFX9rVRx5av
/4AcasAWgoGlDX0WPlfPlapK1M4SsAD1Zzm23msPhWU7+2b4XOinvCOyVVtcoMcdjYseyXoedH71
H0u8slPLjhimIzQMzZKVsco2SGSFF+l0fdQZ+tT7Ghfiv+MvhBkFMpiWnh7w70x3Rjo4LuIyGnl6
P/KP8lD7MTxaE30tuykShQ5tkM3qY1mG8j1bHjP8gBC+Aal7blciiapJZanVuJNeFxAlfBUaKi88
Ao08oZVpfNKsj3El1BiUvhm2eSs4gTRWvQlU9xA6fQBP3noHRuoHPMFzLKvQrKTn3c006Zd33af6
4+Fi5sQzuru8PcCbO9BxqJVl2dZRureMYy/sualUKS1wTWYyWebljKJFNpegCGzczI7Pupt5XMc+
vvAPMmnNBRLkldUlr422TH71R/8+KEVHP/rZEs6sdiFh9UskQBDcdM6QkrLySRfruhlU3JnriurX
bFEAH+xM1ftjYrcHvsV/kbJQE1VycyooFO73MpQDQtM5fEgDjaK5+iH3y0vFWJqwQVR/nmGULHD2
L1VFMdbSeaQanfWlAhwHMVkkQyw/BHVAhkF2RjhqzG4OYXKUYakeRFJdGtPiDyjtk4Y4w4nssDtn
JnF4ZRiSzAamDTOvYZMs4lYGjKP6tpRDvpXDWEMZvOPLFhuXFm9x1z56jAwbWAdRdWSnarg1BIRs
iwfptTGopm+ESwGJfMRZQj3bVfRNbz2Tr04daUFkGq8e6ZeOpWr6NuMFNe3zj334jIIURk0xXU6i
YXnwi7o/ye9bPcVa9/2DnJSZ10mIoR06gtwHEV5dW4dUqfKlws0MIOXIgw/gm/5sPfsvb3+l5jbY
JJMEnVBxIYekHgaBOmoroHxJbfWJWEZnWMGkq2ZkQXtTN0zu+9tmMM1ZKXjoU2Nt4VXPMk74ypJ7
M6aMkEQkXVfpwYTfhliJSUXSOXee0cUBXakiEurHGVBISrTlWkdgQGAG0iKbJQYf7UKVeip0vxsQ
DX+O1ao4fwKFFxsY9RViXFq4d52fn/E317wN1r9z+6MO2gAtPMlkgGOOUgW3cHiytoVdQbgg4WVk
tBGFbc8J2bZfLTgRx0Yjf8NSKP8HxhNtBFv/r0r+MqBejDrx+ZhlY5CL/NHHYklhklhiT9eZuJud
Hway8bJ77chqxGVukjsSX05CQtBNzpH3WhSC4pr3hu86D9b9OVYn2MuRYplOC+VjUUQqHy/4H18A
Nh51S9R3NA4PlGSc8eHmCKjlgwFc4G2x4uUhqh3JaeV4/p4abXSsB/Q/OkF34SAFAErXC5FG3wRP
5TuKdXErRHNMBuGLcpJ+jgzfHoPArP3rXwmWQXr6lqx3PZGfnUCjwyP343wBJV5vEhJ1JQC3Mruq
SLWaJ9PzhYlD0+Cc2jC3nWjEOStfh+e9CLRBNeQgSU5/OsMO//1YO8trjppiXkYzBBxNNgU6/Pky
nnuGk00Z0gLEQyRz5+myRJEoj+4QcIX53puWiOBl7pmK1zUFcVsai9KuNbOjh/tuSif2RYS2SVd5
xWcGQce+f50ZViW/hLudSHBsw5qeSPpAODKGhQ9aaf19ckjtPH48emVgVWQmsW8KlGJfPeVzIsmn
R0aqQI/hgiaVBT+f4ADAcCHydLoAJJZZGo9GPE186QnmiVKuo9faHURDLCLG4SYa7XBBcMDDJTIV
8P42vJMrvLSPdFc8Vt8BViQyytHYJj9Ii4I8AWGc07MEYa4fMwvL+bciVhT6u/ripNM/6HVahzpn
PMBBLZS0z6VBjc0MMKnUe0HLKLGDQUkO5a0rKkZUzMz0g2Nlx5l73IWMc8LyQgclRnhecTtfkwv+
+X3x/PRqtcUsjV/eqPIj3UzQigl6WVNS2sZPw8rpXNlB8RThw+UDY3BQE7AIcbHpLc7kbY4VPzR2
RWMmJ0jYD3TDzoJd/jHk6jANP0CFbMHYdoG+EeqhxrrBFIe3xmjB+vEtPdjdO5U0a0VFMUJs7IWs
nBy23LzKFX119MlfacgaqYvJmSR/OVfO4+7OzaKp+ATvDqKs5Mk9ugiUyu1hDzTczVHtmBmxLQqe
A4dYCB6PqTxivhZdbENAQ2eSq9zSdPLf/y+4pmKgoQMLQnsZyYd84QxYb1t/4E2UMoi+uFBGwC+k
hrNxcUYdktED2HKTvO7UTI6vSc/7s20Wbz4njrxckb2FCweIAoMylTnPcH6Gxg0KI7+ah7uujZXe
5pP9ajkFfz9+R9VrD8PrVA6sx9TxP5hdlWDo94BScsDYbCUqnPbZX8+MCGGXw/XRkzPUFON5adjO
eh3uAcfLV0nz6bzJMFloTyMTwLx5Y7ycIIcOkznXkm1MtpB15l+4ewv31WK2nAyItNOtdJ9HkTnK
0jbm1UEgK7qElqpFubEeuX8PR+tNACyO/hAuwoD7AGYzJSwRbcZiEC9errNqNxVKe7M3XeYlharT
H7SuVEj+BnKvNfB9RQO6wGPOZVNy/QBHy/5DokfnEyNYr1tRrKGUdM4pAg/uQRShheirB2WYOSFx
9bTIiMixu7SK6sT3TsWo/NFJTLYQrLOBNTCFjZ+s5Qfnmw7ocPXTtFl2mAdrAVOdX8LCs49fFby4
T1Fe2cZD083FxrR7DiMkeJ1oIdg7fgFhFEO1DrQGVlnm2In7rOphxvN3gZh04DYaHKMzasLi2FY2
LCxRd7Yz43KhNPHWNYXwo3METELfqRKcdWpExbClcfXHoPAd22tymlMq7A5efurFQFjESgP/kjiP
LazFXsHSUBslk4vkT7V1PVI2w12uJpj+2dMQM5SN51ATLsoy/tnIv2aXzyNuwWEZ+dtc17siGG6X
BwECTV6VtlZxvK4AJHlJJysuTj05jgm6dlx2+mKQsBqagynN+rT2GwztPvzXn8mchOMz3xWtjzAV
38QrF/WB23o0xJn6xMYhwky9ZlrfFhTyObdr07Y7TgF+tjKL2SXOE2AJfDSzDq1meU4opdkz4dPX
2a3/S6meJXqXPS+lTSAVHcwNFAzlscp5lKO7MOS4tXpg1Yjl/NWJbErccID2SCb4M9nQ7hORXlyZ
xD8y6DWJWWb9xQSypHevEsHvbSfNQJgolmDAlWWi+T6VHxWLrn3sY4ISMAH3rlcI58iRzKF8aGWW
iJ0dI3QjMgDAUvNCX+4l05IZdxLdPxjsfRL59fc+yyj4tpHgdlcR1g3GNg1Ih02MlPosy1Ih8xdd
bsitLcijuoBQOJkMX94U4tx8wOzWTMCloD7sTZ8U28V6xAFsvpc+YgUNKBaJ4eRZpZRBbvRQ0dYG
HEOhnk226UWNWhITDxh4NYjtzKAm6FUHFXPZZOiErmXcEu1FMu/rsXdD7bGgdo57TSmg+xXFJcjg
MRIM3qHsVYeVtIVeWdwVAjKhVc5NPdFBen2QOy166T8L4ApbEJVtKHGqXZfzX1ec+JrBanTh/Olz
CBGsUYYkPix6ZN5/5RujOs9/YYSsF3Se8pDpz5HfpgaNGj7i8+HjMxy5+QmP24ypM2oREyfHT28+
pxoqbCyGSgJOV7hTEmx1/9k2MuJ2X1gqtL/nB7Kq3yFfqr25kwMbkOhxuSast5BWQQaTqDaq+kgo
dQoFSKqK2PXW2/64vCOIKbPJX//lg9uWuheEEaDkdRdqtDIMPDbeFpEuCLh1NW9JEOvzNW5FZaHi
CCeXDZMbY7yQ/RjhRZthbSd9U/u/5B+Bk6QGytv2IMIxoQLJCwHVIQJVaj9R4Su4dEPAhgykFu+f
tOAsGjSZ470zGPv7XfKWGPz8BdVhrVMyBFHK0u6+daua0dFbBld4fnQoOtja3AM9oODhj2hWdAm6
ghWYpgxTlJ4l9tAX4wA8jXy+af1T89AYGenBya3w72V8GqmNIPbgiJSZqgNCuQDpm4B7xgj919a1
SPnCoprxMyWglSKKKbkzRI7d1HF8zLbwYkKWc4/2O+gEbBlrT8XIUHycSRwQYXFMbiJ+nOXhI/5X
s8a5V04jYD5vphytTixVBhqj1GcSh/2qhuUo6OroXXZXfFCGWrywPXwY1f6UVqGPx7fzbCIqUfw0
LMtMIInZrbIkYZ0Ny/A3vy7JzTGSkClWft0shalTKmxg5C+7i3FApohDjnTU+Y7Qf9P56Ge+QKpN
i1PyBOLrnBdLtvZzZrhldKavvhTTKWvM/UzkHgL/LsXHCdrCmo0dVm11V+snAd3kskM7QVXrmmqr
8vENKa4DNtVy6CTV0AEt0cyneWRu0PW7lfmq+8QENn6fkOvrepkDtb6BZcz3MoyS8QTC9oGCGBlB
FsU7yGNYDSwh/7QxSIjAYSy6aCs9cKumYEeubuXEQ3eqT6yMu51H8PqSJSbnm9PIcivWlaCq3AbM
PrENDFGvKP8uTH7VjnH/ljc95lUGSuEiFpTiEo/G0kblj/ArU3VxS/L2TpgVUBvN7ecGodrMlQTn
y9eCtPcEmKru03IZMUXWdCHkDMRcA75khDAoAtV3+ZB/UUK/whu6fV/3TCYX/3HwZIo6fjTnZquD
Qmi/1gmpT8KQN+mChIP5t7w9UEJ+dG6njDxq5VduK6Sq5TWpNAU8wo9CqAJfx0Tgr8/3L9kvwFJT
K+xjDmaSX6Fq6pX4pA6f2KJqaYd5DJnty8Ybfmt0Ki2mU890OrCDJf4FAcd7bmIeBihoEpb9gSvl
UOvVvkVXDLMFtHnp8pNTfzGKFBK8RpkshF/kYeNVgNy9txsO4KU3eFQsUH54I5cJMZeAARYMVd6r
AogwA2AQpGjJRikMb/bwZhabSHWG7Zr225pCXN2TtX5LOmf+/vHelrsyGccDJEsGwRuTKazCBVdM
8xdB7fDIG0SBJzJ7XBOE7aqbc5WfmZR5/Cwup93o+UkG9Vtcxe0z8zZ7LqI4YYliZThFmwZjhaU3
4wO9FJvTzCzWVgkW4Yme2gCHIrPwi96F99Sk7HN218AYiun5ey9QMqxFp+JbXJkmyGwnwX8Tt4Z6
papgp2B9AaxPneNmslyBmE1UMHH59j123MclNaNTJsd7j9ghkN7C8FZunu6txuRcHN0gXMkkaq0y
oJK9zk3l+7NY9WXFxARe7mAXwvOFllKUJCaJerXRcLP+opj6ArydKNq3YPfG4L0+KsO3OBIlC6N3
I68jTzDMTeqhio2n7Z6GmpbIJuhTug0CQfs/qwlBOcJINQTi7fNjwppQJbAADGPXgOGclBa0+l7X
A9Hiz/pfSBQfSMKVy4absUBHuBWbvejBwr3e+C1R7p164dnxYZULOtZwI5rEQwjA9sEIx/n/MVJs
CTNEb36ZhFgbZsLTHeZef9vYu/BwIyHIVl/1gKKvE3MRKrm2EoMxQZYInOk75Y0ErNRAc0SNyLWe
O/C6qxk2h9YywB5gE14lhrOTg3tiEvr3kHBfS0RXwzwegWvac7acQ6Qp0nZ2lAbmZwBR7a2sHgIV
ahSr6FSjAlGgrn5O77JTqIO0gc3ozOq9jjP2aFhbIlQn7jxNe5sTrH/OfEq4dJJ2zKRI1s8BZZDt
V8BDa43WSi5Sw8hePIIPfGaKU3IsD3ZiG8vZIkcWD8iYRXRb2dy6f93DI9XVBgu0J63XGby0sm+8
a8IobTmcwmlqub2P4GNirddSsDCh6Q+ClI3szDY/GVFYLs+pQ3SdyoHqhKqbLQwG64GwrmEc1bJW
XSjRLg4Ij48Y9/cMfXMTk8cnro5sgt/05KRTnVeqw7ixyoY89C2PFozM7eFtC6ZTWsmglndu5cR/
smYiWuI8MkvRjoetIDGDomKY+H3SX+WfKgSJn+gm/9oLyNbBdH7BOUBKQSePwQjVNQQdTwubEDzu
Pkif1vGtzqvCzpFViHhGA+ysan3TXlZMrjctgaHImIycofL100IVQfQzsXIwemqPEgW2tN9P29H1
OI8d6KF6YfwwF/wlnllrkwNWxZe0GS3XtHPaBob5bY+goPXKeC3qU8k3E9pBmdSqUoKeH+VHSmIk
jGBeJJgcOVAAOGEz81kggBoTuq0FOtzUw2T1DwTSxTNhRvO8wvH+1DmJonL2IINYBHsxi8XBMNvr
QwpuZuwYKVQlMdaKQpcUF+CqYQz0yt+k/l6W/u+VKyo/kthlXxtsXGnji52Tr1c+iuK+flgd692H
7SHjqg0iKEDX1YoduB1pGsbA7w1kZC15D3xNPOq89e/h4HFu+ybZsiwLqlg8SZMMMxlCWL9omZNQ
8pvSkxaHBsFCNAWkhNqwCMMt4fwMR42kx7IDysg1k4YFpOs2qRuQPnBSBTBQUpHjEyJ+21qD4/tM
Wr0exlH72oJR1vQM/B9Q7lGD03DPhSyrYgoR031rex6yDwAliLzwRlRfsFxYFqQ+OZUBNeCjeJFq
sJhwlxY722p28RBIwtiGFHHcGtCeOHSk/m5zRzV8u/nQML0BB+JQPoWQmvY+FzYnnG3PHkU4n5Lo
irsCx9DMJ9F5HwJpGMpGXhYtpSvFXi81VjP/aa/DAQhL/mLpxPqqpTBViYdlUfgbotbVcKiH9dt0
XGcmpnAFVjmux+6jJ9lNOAjf0wjaqzCKTUdGnTe2JNVRwWycuXdqeETKW+yVrZptb4hveW7bYbwc
a2lCFbwJ2Go2FUswtSb836OFyMpeIRrysopJ96CCqNfY3RgMFg51kBHxZwbBZvzlXB/n4SPB8Ve6
W/aNm3/rLsMNGV9/KxnumC+akcvehEAAAFNIl5NjtJMg86/dIViO/8XELmjAEKeCL+Ik2HXvkmOK
M+h0olDjvARScFn2DiDS/4871IVrlmNeDytM4uKRrEmuOjf+eIXPGRVkLl4txaMNR0ZcCz1j8IdM
ImPXxzSqCra8WzvK32XNt8CZBl8H4Fnu0iwTDXgwvJ05+xUgxZMT8I6FQDJOws44uFAqhd9YQRaQ
LOndh+isdftITEgfLLn9dvI2VlKnoCGLcu8nlrbMKMSwd7/ypoIduCucKvErURNDmDiC8vMsoGQd
UonDIrPQQ2V8QNIBanKe+9ePCz9giUp3ggZKWBsL+uP1sX8Gbmd+b+l+8ainuTMmsoZCwFE47QQY
2Qh/uBznIU/3HYtvZ/QzH6+Hx58RAIvZtWrv7PXBfccwaaOuoWRyAxHs3C0UIZVWhkhvvIlGxfMC
j3YqHF59Xg+YX1b48NaKKY1G6RScs0yxIm/s6qyjlR+A9JmJk5W3mP/rY4Nj6hmnEc/f+CMG9M8E
oWk2+S2mknMVo+2L7q8iT+4r7d6nntVhZnTeTBr/UQKInbZwHFUC9trZGTeqTIj8rLzQe4tIgxKJ
AhNwDWvzl0ZiEusGz7L3e6Xikx84DbZs/ImQ2e3UiUzeVDZTm/OoB2KoUrM51bMgXzp0IliJY/K6
3HsF91vSgCiRJxuqqM/PMDPz+L8Nbn54u9JHgGB0W44p2VxfIYFQLZbgssOrm47SCyd8c/Idqpii
dnRD2CUN7omHV5nQy+p95aQPuLRXaNr1LkoQG9Ncwhspris9jBcxgQR1E8sOKqzAmxqyATkwt5Co
INEuDrWrRW6LgwKg0RvsDJ2CEzLB1Z2hboDcZnaL2ocZtzD208Vs8W2w50/Te5nDe+ok2vO3TjWL
pYoAkrNYe/FJVatQsM4UfybZM4TktHZ7KCdIU2wwGfrrIRZW66qz5/XZYTFzc3OAx/QuOvBQtveM
slmOH3Hcr/SZF3vAMNPOg4ROma2zadNMl3gTgXWFBNikxqtA6eyAT94f1Htekrkq8gcdiOpqwP6H
oAvHDFsDwlQ7WO4jJh/o5gk1BXV2M/tp2aNvS5O5nUhQ7k4XPMEr+bkM6/cRH1S/RuHNsbW+8W+O
rnFrjDwJkxmZnsy7hjvVYWh/tvH73txgVyVbNLpqjj9lZWucmvATONYJPFwp7PYw4RbhlgCMnUeo
t8/fZ7AZXYzjgydXqQU/6p5PU7jq89fDWqlL5jIQru2221vSE1wpDtd0mC1NQvPn/jgHsmY8eCtX
Lb2XM4/BnzDudOQVA4NAUstkizzd/4V7cWfv1wvWn2vciLlRodJSc1eLf8TdFC6FCEPJGmtXC9FE
106uuqlWqe6VsaKePCMxLdxlpLvohT39a1uNEv5+m5+kErX9zL/mZmoRYi0cEQ9XSz8lxPsPAA/a
0vO6w1TLYjOrg6/u7hcZypgVRL/OYp/UojV5XwBIn5L9Jrzv/+ky9bWZjnXliwBNQtYiw+xahtDI
C1GZODYn/9MlAm6M0XbVhQ988/mBWI8hf7jDF2lXlaDBGDYc9keBwcfE4SazgJ6M1V+PbyWxOiNT
tRCiLqbPZPoLel3EC1019NPEKCTwPhsKTBvULv8xXWVek45fIApfx4Zx3ReZpQK6FWwSY/d66Ka8
NKAAhTYqaLhfrvRDLxHokiNa2vKh8IBJy6695t3Kql3W0WLqvaoNNbXLl9XkMQ0Fl0ybTWP2N9AA
c6tzbKiCEs8GTT+sneQrs4zXR59yWw9wc2nzXIRxw2Kg4Ygd+2exzej7E7TZDXicKOFbCT+4shco
fY7WeLnUYQG11ibmHjuL1eWp02s/pFxBxznANxVgeI1LnHFQkyOmHJrUWvzC21cJm4Rr1E/J1vL1
HzeKXrp2eoS1cYujaYHZxuSkiWWT+g5u0FJlIP2cKLeRDb1sURPbGKSGSzGByTwxFNzu0iium+pg
vaihnQSBzF/eMYQ0v7m2AmwD6XnhO11uYEM6fwwB2/dVrrFSFgSncUnKymJlc03cL4rbJJ0XReSQ
xkp27UFJEgoPrD/mbCIpycRqPX209spC9mCQl7c+WA/6WAdqpKckMO2YRt2gUSIguu7Xd+DFtKOU
WGZiOqwbxLxXwcCu4As/UROgR8YBt29zJdoOdsBh4Ran3+WYTkuP5FDROgMqh4dWZcAJhZ20pSJY
pjvyIaxZjii26Mr5YRH8L99bt9JFyEBno8ZgTtMEQCoRzsyrKVRaBqEjeE00Xc009cvmCYo/K+tm
bZDHxT/NFhbq5QKjbVu15d0HJ7UhwLp2JGVzhEwmQ5fG72n3fTxP/6TvftBG+iM/7/AJ2GN0MiMu
ABY1VRkszl502tdI4/REndnj8Wbb8qan71K3PcxMQbN28V1Qo23Vyj6+4n5pE6PKFpHf13fEgHqf
QuwWEbkD1Z1AlvnW/raoLMw9EMnSeoCxpPSe4CluCf9kNRU/Qg5TyB1gCS2hK14Tefgcse5QggzC
RJSvfVtg3ekyTB4tdKEN6JSQoP/QH1rXv0OKrj8DFAulu1c7rD8T74WoCECvD7FXNAgPR/r8C6aO
rWnYCRAg9AAANow61CjP9yqBctTW2JxPSmAjyxyoWqvF45RkaKXpCte8LnyT2C5PCnMvtqqkdEQv
DC7yGyvTxzS4GZ4eniuYqWppKRlJYvAVSHTiyTi1vGy6gKI05Nr4G+aoCSlJDkDhtKCypxPHHmBr
4GwUxJiPMR5pkQwZGuhhXnqXTyW6LBSp6qFgkWecjaWF0i8fp9gY7jye/vuobXoxMXIxEWtDWBFQ
cuY7TEBsVfCKYxVc5OAobdHCBujfzG/nmNi00EJcCKyR2K0sS2Bs0WG5tfFx0kjL0BLpkh3+4n5A
Cr7OWidlBBK7B9sw/UfU8j2TzFLACeI9p1OsoUlyBrTy1Qg8JoA+hbo2KSpluxYCflgHKhxhIHC1
Q+2LRivO5HZR24gwa9PHSfQ5U4C4HY7Z9eNXes1O3KkQbJd0VLK5oLYIeap+02It9jXh4ItF9yfe
4wSgqvFcpfpC8a7JJj5fAkzeiZqXGqBS0nYnqk8c8YRqovDbRs+wmZguawZH6IBqXZ5xhCXAT7+x
loQgZiwTP/oGau8sb6utaNfvcwUy6svr31GAEp04moPbwkxSqzxGBEwqjl4dExk/YtN5rO0wvmYA
RHaohk4Qz/TySbsqDtFLxwITGp3j42GWg66FXbNCfZv6C56hDXaEzav3MqJUv2nnqgqcwmxh8sB9
z9+mtIPo5APjcxX+XIuZuCg4DokyfnjTTBKy/NpOLsme+J0Ap4I6QOSRckXGc0N3t+Q+RXaDHTui
Ozxi07f8IOkWoLwHRLxGnUBpLuUOsnFY+sIUbRQUY7vOdsa0M79TMYqy4sYyu8B0z18/SzUgfUVw
ksxzxJN+1vQ5dCnADhCpbjTJBUFEgtQXjUj0kwdYJ+mPGqoxdST91aNG7B6vMVElMtdysPROhc8f
lrXpjd9sUfyraA5LwZRtO4GhtC45dmc/+Yrt/YJ79SNag6MdV9+dN4iiHeOD4ULAnnXKtMgnQrmO
AU66umvYsuq6+IPUiUXkFtVTw6FM5cArjIOHdrgQ2kjtAsbVPCU1HDHBxJg+U6+hpHmlDEiAE0vj
UdqUbt83vRgQwdtY6qs3yLb2kY+O35ZiIbIYXglQXiVtuF3Qn7i/cibHMslzsG9YJtbR0qCFIv69
axL5vjUErYNRIinfXtQIxiXDctn1b85lny4f2PJLiFkA/Rw2WyAiJfbQkz7kOHmuQAizRLd5yM7u
A9ChXOmqT3UY6M+rmDQ/XbLrPBMGsIYRJZGaV4PhyeRO/OP3qSY6FIIm9B4HNjFUw9gWvZr1Fs0e
GoiMTF3SFaceNyg7QSLwErmLZIdZu7gVsUsr+B5Zc9205YGR7dkGT/cuSx4uIvm1hAhxizqRjgkq
2PfSebs9QNsVTGTnOxjC6O9jUEW1y5Oi0wXji4bVsZmx/edrqStxtHXJH0HOusqH84EIur04wLub
RkxYIaYLbaSxua8YkIdvvSMm8/gFrl8qG/qAgf0lo362jjyKiYsEjjGUuekvTjedvTRhg8jwokSp
IKmcCArL6qkrh0H81AxInUOzqsvQWq3MuVIjFZ+z5Y6pmsZM5hJXtfHH07zAsvr3YKEXdvA0Uejr
zZ8h15Rrgqe2cJNmVZclQNonFuoV8nwLYI00XKg4m7WC5XaDADIdrCkFavwJMQ8Bl1m/V2DeJDow
1crEdajV1MHYD8ivM6yc53bOZKaYk0RuLM47Pc5Yi8uD8sAMSRbmh3ZIQSW2/BfoJRfXKfOwaIcr
B9ChJTe1h4D33/zhFo0Y7GxMzYPxG35xAwU/aNvPFQz5bTL4BFVoQFUG2cnXAsrLVNgQ0Nn5e7sW
jK2w+1pEFFy9eFJ+eiP3Cod5aFVLIk+lm4SLTCkhL9TA9LkX6gOaojsx5WytgY41MVRpGTh73Nfd
6i6uXO0Q+u+MsZEZMGfgVYZ78z9wCqPTb0kt1KXeWvxU0NuLwa8UlHwKkxupdTDKtaCHDB+fcaWr
PLfrasCcaIxDiRCtVE/o3jG43AZtDwmwhmZ2kLfzl4UaYufoNRiUdrHNjBGMt7GVYI0oeka7dsQa
8dT8zOt+AfnDeA7qjRUr3fF3wEVG29EpIHbQhb7J/kb+45miAnsjmU4sbGIApA3RVD6Og2KNHWHf
nqHUtUxBtG6cyIwgimx1EmICkMa0rabG/8PIEETxH5YAgDVXqksSsoDznJ8Mnmuni6EaklnScGEY
T5xg30SBQZiyxpipCtYTNUs661LP9qDA16Ie4iQ2/9MKgDyfi41FZb0PzZxuBnt0BV6HW65xSdSr
8hmqJlv04imw6MwJ8wfQXaSv1Th3cmwCdK2gTOQbzeKHOOmyeR/FELqizvsARNvmJnKmyZ46lqjQ
LtGJNlzTEtl2Q/aQI07JRUyp9wfaTxJFKuh6jMYWUvPuaUVtkIU2EYIVw+SS1KFaTx5B2wuAtNY7
5srcPoKsOx/OxwmfJv/QnEL1Ak/2/Y4pW5VDLnWkWPzn7XLMPOnpvQ/ohC89DcSJHGbfvWb3QVzx
JrnUspUrzYeEqztv9wILw6Rje4pEA4x0aXLcTEkgkcf9Wrde8DDw44Tv/1wLjOlCoSVdtwWjFFv6
LH4Zj7SDp4VvJ5+jF6P2x03/UTzKA6FFy7PlHsDaa85Qe6NtTd2USCP8adjAA0cdbYShlDSQEUuJ
gr1pakhQE0broGX2ivvaOLXVIOzS24ej5MrnwLDIeOoF52C1IWNYODnaNHjMiBUzesnfWYyZ1W5u
u9hHv3oanKImCSoI6lGBmlg8fdmFnBg3NGv9udDxyve+PdkDfg87YWHze4kv8giE6ZUcE8eDO4jy
jI7ZIenpzV5vfqpQrO3nDviEhjIC4e1Tc7V5StLueWXAJ56ZRc9DtGhGDx0qMdcI9FHJtDivqtlH
0RICZTmaR7/rKJOVfYWiMLSy+rGpMr3vh9M5Y5Q+rK0Ahnxhht2x4rQq41Pt5OtipjWNaNiSNhvy
jyWDauHhhpuOF0/gupacwaUEqLj9wqVofLVNCn+XvEvEWTSqImAdwc1dKY9Ia3e1HZxIF1tTvg8X
4SAr9GeXxFGEnO11eEWiHI4d5sY7N2370w6j9QawZhjT7UQsfIZ1WWA/kVKLgy63iDLBDMSnU9PO
H2HeEByZBbnT7B1yItMhj2cZUZ9mU9q+w0mLwAImoejNnX0xR4kwHiXGiVJHxZLT0MN6GEQxlTjR
HCQ9WQ1N5Mx2t8YD4tzWUEljJr3X7C1nEGLErIOzMlVwfqhd8TKFKrEJ9YUWbgz0xlmhTr978DXF
+FG59Qx1vblufm3x/leysNDvzaN99/w3TvCjUlj+Xi9H2shYoRtLyKmoA8XpwpNnP6SkR83ORC65
ulNOMYniJ2qDVgk5vyoY3PcZ/cRiVP12b076URrx99QSMDRBhdpxvL8S0X0jNCWfZsNVDVkqe3no
LqsBAbXncEuOESjIVJHoJal3ya6wHh1+K1TOZNfdKwyK2DikEegHAebsSp2pAzaSFN5OD39J2GNy
rljnVojsLiyo54LrUQzj/xmPmOnDuzuGglcVH0HdRG3EwVZFbqrmnLnwOsc2JLP8sDscS0c4htAR
FwvcgGVep+o7l04iwBaXKEBHxrqi5Zxks+LhyyoFh0BgGqx6XbJwLe+Qyd92VqWP0JVtR1xx99yO
gmUveWtkXnMPq3HPKWNsx9yWDP8XYMB+biIul8uvhWzMCQgB2PhK+b5/+wuY2WDBYjk2shAsOFDR
tLJ0nuxg+AWSmVcip9QTf5g10owRgqHsftL9olApvmPDZ58DB1tcttuPqgzX7Cday5H+uvZ+18CZ
F4X+CpV5VJNFG8xX0Q1uOjBYGA+LjebJhae+n4UV+oash1tkiTTnEYF5aVCzlOTnDdC9ScLQhDu5
GpjHFbpP6Q0zp3elZ9KeQKsYYT1ESFxy/jT3JZ8tR+KKTvtGXg9lhal6Lf/NfzUn1QrRdplecz82
pSq2uxf+WL1QHDX71YlH3dWhxExthSDzOueFuPrycUNAF6+/gXCKCrEhZu0F9SVsqMNki8XcQiCZ
si4gAbYnWpn2x8CmSUSWPOAMxtRlh5Jp0KJojqM+ad/rAnAIkPhBSa8dKbk4pJT0wMwXobfaqR9L
+0Hc340lWS6R8CESG8JKoXoK+1x3srljZgkIDaTdfkq2HWo93hMe/I6FJTv+uEitJqX3f3OFbFEg
CZfNTTykPhznTpwrJKhRqrwA0rU2FbpeSYSTSMkb5A2K9QswTnitgrsnviqcDhnWldaEKW6Lb1+L
nhV7oeUpW9eZ9cTx9HzgBtoeYW/rTi8fMHpeqnzi2mM2kBgomiXWEgPA/Yat6eGgwVScbviwcvZ0
GIm707AvovQRqFxN0glSFG7Y62Po4hCqpD86e9V57J92XltONEE7RXaBBxZvrhxgoMpYTHslAuGt
2qyfZJhgh2jJtFqitGIW3zWVXkq+/bkph9nfvMG+sgYW3SRXL/Hc3f8OArouOGZXU1tDSqxytQC3
lx9RPbQeLR7V6CGjtcmeZyc9LGNpt4/3wIRuHUMdisfBPltjuiIIZw/NiCMi1fYqYkbPt6PbirM6
eM4poFPq7E0wH6Vy0uQArj2Pab3+lMCO0NN1OwM/AANb/Xo++4b+8qrTruOiBCQpCOJSw0LDuNS0
7oO+2EgtWYj9yc/NdWRN6QTE3sfq+X5Sv3ps75RHw5PYJ01WC/ae60b54jLO/k79C30yDUUBnchh
Tiu4ApG6CLBC9jyprqPZXWtts51/BRDIQu4dPuT01PJQrUSDehNHRsoEHLken3d7hHSO2G+6iN01
Gq+EbqoIMirFk/0BAPvJgCSdw79CfPx765IUIC30KzUEzMOsqCeIFZup5FyJ+SeMxe6p06uANOW3
049IVQxRZFFZBDalqbO4/ipNy3q4WwfZ9toJNN47KPUXl/CPccJQVmiv8+ZFDKyif00uJt1c4N9F
/+sB8fsEQ/HeP+xrC5vrp5OfuMace6A5BRKYgdVafMMa/GyippXr5v7jxCqE36fhWRW/qIlhGsu5
cqyuAaLQaC+CH1E4+QHu4FzbfkwQ7fyXPMPFNmpDW4o2w5NGd6EIvC1qITC2YznCHcmyEQzTRn4q
/+g8lP1eBT9srT6APorapE70mvLmQ5qsvH+fH2erTwDK6V4W5F+EJ5zh+TMs7jtSjni2Z4jTheEV
S06qI2ApnFViWCHhjQK+oZwHX8vlQoYZp8XHHhLP+aZZhERtWnSmIwwiJNHccBWYjUKvFNkkVHzw
a9zazYjjlBnZs72CFWcpk1ZW+E4dQ3uVMtPmZvzrGpwB2xZNPp3Hbia9cblAxMfGEkkomXEpl7CQ
R4Ci4WF8azcYRXbnhv9K1oW1mIJFQiP4iq+XE1PgAx4atJuwTiONgp7KyCet6htSjaDDGQ7OQzCu
vIoMcP6PhkYQO26GvIF2S+rps+SYivjUFDQBQrJMItG+coinblv3sMB6Y+7lKtI3idLv8ZWmmOGN
3ugGkTihKL+btSPQXQFU6Ee50iVJr26UmNpwxuPTVvdPTlb6kAiQYeQSizD2C+pXE167hvMSiYcR
HXsx90LIvLa5vgpLi+hMJc7IOaaDIHh12KM567CnccbaGvK61RTGBVxlsUgOaGK72xSGNQGHULwS
/wMCNOhF2Dls1yzlZzQjzGyHDdBikoUJSPCiS3gRvUHbjkDWf0BJxY7VoHDuOWvK1rRdw5aW6k6I
XW05xZYXkALmntlDGgCIQHMeK2O72emKaJOIysWYDPV4Xb7tei3daQHMylWfplM7o1ey6zWFQj6q
Wx70OLq/5pMZiN31xb3AmZeEH7r++bQqm9dF3AKRYlHkhUfwkpSdUXpTqnKc8SFdtezgpODVc1Zd
XjW95s1friA2KMHNVslNxhVSfu5mxgWut95ngTYuwjv8M5qiyUUxZTQIfD1Ic29BY1of+GUjIg/u
z0+UHW0rprRxA1p/C13iQdOYe+cTENQj7ZdCL0Ra2Hj2MwS8d3LAilC7NLEmuO3JYZpfCYeDOmnj
dM+6OKSyXwzUIAuA2T9IzFO2lY6Sxy20ko5yYMRweIJy09NSkCae3Ex3lkaffk66CSe5opGsWwY+
ihELiuQDkuaJt1JxlchNYYSWpwiQCkN+1wOHozp4CzI91uunnh4j6/MAL9lRu36CM0rkwCItoEBd
7hnvOlkQS+zbS3cz0P+HNoqXIgtD4+lo6M9NEUI+2DCIqNcz1wXzwbdeWHqyFN6tfvmlNxDrF2oT
GSv+4hE+c5na7+OrsioLjysvicDDmJ99PWh0feyHz68nay80LdD5SSg16EeSo3/szzFYGme5wEsx
lqlr0BULKS6wb/C8PQFMZVtraw196hNNMF7CBlXvKoBjZZQMb5uQiqHs/JCpOVHOwem2wdrTNBB9
Z5rup8O1J3GQ2bgFMpqVIwaMo90aChRj+tp7tO3j+6Ii5OJNg1FOoguHXt3gXVF3RNtvBzgqbQq0
N3BaTjRogMTT27IYf1Q5tNTVhjGGB69DipJiil2NSxWK/9dhckPLNsFZtsflScIQRo95WpXpdoJi
ivSFURkW+cmQXHLrkI9lqwpfispX1yQAhC3Fw8KTTM9XobZqw4uzqjQYLS9fNokxzBxhPmwRSuQP
8TlegRE9wSjXiQhZ23WoqgNRfcA2Jfxqk8Dy5FWRLjRks5+XO0kMVg9iA3aH3CWEhzRr+VlEcUMu
6NQxX7ugu3h/vWS6wc/uhyLgX+h26zDlsRZy37UVanmqACugWb+1Q18C6+/urGCkpJeU9Id4sdr/
OunkPyEpTNOSOX85zWiTqA5LEyP4HAfeEprg1iTAibL12Oc+25X+t22Gm2hZAN0I0uPV29CNSlyA
mQpsT2FlLsJj/mYggdSD57pIeM5oE7rULFMX2A70rjg2zVQh1xm+oUTiUThnLoN7AZyZ8A11tHv8
Mkzu5aDy6PuNE6RsnsQ4pc3NtaWNGUdbeynlagYat7P5NuhWmQlPyl4INIIfnxfCOnxNwSHrQrBj
P9J5L/csu9auFmgyf5StgQvpvMOAdDU3Aft8YAaOD85pi9nCihehsWNmws9vdDUuQiDTBTGf1hSc
fqc1Lbpqr8g8QBful9org1ZuhrtBt0KrPpyvcuP54kqKfAp8cNyJ1DL4fZ2ZzBfRbjMAAy68m5P8
mMIf+q8XOfkkjSxiA3EUZZR3x7hn+SHRSUatsRvIYlIHjNTkbvRxZ3/k0QVAJXg9QVVqEWXKSHyI
+0gbVENAyi1Wzi+IegnqQ125L/cGQlRUP62QFX9JtdzFwRcTjijRAVx+75++PacOOO5xopk5/9lG
BBX+5seLOV5zGMOV/riYfsBQ/PJJYSxVEaVBJKcAU2OsmPb10oypZeUjzExK/djiZ0oFexsW0S2P
6O4KKpEQn55lNFzFxrex/9Kxpl7uEdPv+g+KWaIedL9zKhGwroBO5tZPxYA8BsLdtMbAEG2KxSWE
CbEezkPBhZmphIEEfANf9shvadVZwczvoTWIiXogMQ9jjzIgybA+lCspMINLrECZ9vcFmhLa3CYW
WAp74BTtVn8nLqLBsQPcNXcECEczqNdFXOSRsIjmebDQLa+tIsvp6sDoOVTIOnygNA+sGtW9qxYo
EyTwyeA+Tp+XQVG4kh5lkgtM+VlKpx6MPJSz6aLCQ5GGm36y0J39XlV/Y35aaZA12NMGg2tOCJ9s
x1zzxzTWTnkyOPqs8yWxQgykFiRkRcvNp8VXFiltoj+eUPSbkmsffah65nYSLr4KxtnFKOpbtKMH
bErYsar3Txzf3u09HUmg6XKlsceqCbN1il+wKMkt1Vn6fxjBvgQ4R2XWRM4tK02oIzD0reaMSW+J
JfZQkQ6qLbQ53/vXOuM7ZOOjm+lB/Ux5OVPY86+MQLn0tla4OXxKiu3cTv7dzzpTebYJaMmFyFxz
5TTYVzqjyJu6oB4D60x1hgziii7VGjDE505F0UmdxGq7eU9EjzNXC7BRTRmXV87L+jNfqS0L5tz0
Zlm90em6OHCa4XuTyTONkT600zwQxIdQa4/cpFdLOAQ9F64WB0wZtd7TuUtBU5Smnu9JCsr6gWOO
7NRC1ugXMfFe2uats0E8fG94n2T00azpNOlSzkNwe09XkyGH+wB4mUkgoJKidQxLhyncs8zJWtKC
ZnoOjySFRc3XbYE96i66nplnd+zRa4Q2E8CvKLH0NOL5R6lidvopEJgtSVyq19cZfZNmEz3SXhpi
0hsSCxUJY1S3cowRn8+Iw2LZSQvJigF85LNf+vrjZ/IaHac1Y89bV0iRQF3wNqL2TfK8dt2nRHa3
+zKZkI2f58xxKU1uKZnGs4k1ao+dWjb1L5hakQHRawtEPJ5tzLVzdGvTpKzQdaNyRhUrZv0Ce9Cz
mEaBZe3YdWreWG3v7JEnjus7HrrrEmMNXg4ydHET0WiO+df4oNijeyFHGtXjmuvGDUe5HChzjbMV
SQgy556qECFdEojnPFB99LblCoaClWPgXvCPtJI/E79AaZW3uIyXVFUOmUDrmiftyrrvAh3eDtBA
6tVbFJHkw9yIdtQO4424E+rCDcUo1ODCdbr8nQVTKnEMdtRmq/QuMz4b2fBYWwKlip4qg16SJsR0
ZygQJTuwIPlpEo7gBGmDheMWYAgyMRWYFvx+oG0K2dRGdanvivtGpp9CGbHZ6dLHZKJkoIbavAP+
6buDgi49tkrabk4KzfDVWx2VO+MkzXsZS/Bipz/AZu6HmeWdlcKuJsm61MKZMivaYylmbk5Ir3hS
hf+snTgUC/90STFGC2McGkFOn0vmtx8U2k/Lvbim43FxtV+PAbm1cwihIjb2S1WZmYkYq8IYhcM2
9DafINsG2poPVQH8ZRlOv9XpVKU9qmT814reEfY1Iu0W52GzEHYM8BCQX9baGD3ZsUrJjp4sh8cy
+f7uzF6ISLAxruj2ySArsffZ0JJQD0MTptc8j9iWsfZw7EvXzX3FdIWZF9nBNw3e33ZRmJDCfAog
FTuRHO+rpxE36WpTdrQIyXzO4Wsh+USCSXNsVlNpszGof5OGvyBwOJTl4kGlfEmw9KNNb6ohM3S/
jYLMOBXW4Hfw1RSYswtfXxhQuKsOJOPD4sA9RJuBn7CfbJ/XrHK4SbzWNR7/Lu2HJp4+QCviulVj
ZX5gco4Z2+Buhlp1z+++ACFSBM+agyUBg/qTap0M8n0k8BpqMREhGEg86DJJy/LpLOqdSMpkOuEg
W0t2fCHPnojhl2MwDLgIaywWEeR67ZQY15Njt867sO8QJz71eRSQUYQMztUoHra9wDa/PjbouqTM
X07xJ5T2B9ZbcKeJNj1qxiNzqfu+bBSZ3i7AoldqquaEx8H4H/OFClnuA8KDi2TH+HQU4awTWLZ5
rObLHdyY2eXqh2pH9Vp7D7rz+u5iTzsqzhuj4QHQxhh0mzZDDC2Uv85vayvFApxKE0JVj/wJpANw
yh+owhXNrgMNv3Ynq3UIjYVPZpU9YVt3fng6uXONsm0b2XN8KszrmYgrIY9gcFO66USSHe5No1KR
uES6xANOeed8SKVEmkh1pC3v8uRpn8bug9RaOInzFHeeaVnzSMIugmHbGEydRdBc87jkAQLafWML
56nV57wOOjZ2Knyy9GE4yNM6bduczsX6GiSXfSdxPlcS//bGKYVPmIu+EJh81IR7pVTP66mIqPUk
QT3nEQ8nHPY7+Ppiaa1P0YhAhLzccGp5/LkO8Cw6F8zDqFea3sEk9Dwn9XI0K2wmjhkyNO6HzIab
HEJzUepP3D8reghCCE9RV/R8NhvLhFVGoFT0Ddk/p3EVcpC0a52lu1uPOXTIHIQxFfzq6k+Thjnx
0ZnOe1egi0BNoeAzZ3nkRZE8LSYDBmKn4ECvtv6IyBS+at4+PInI5Rl5bKDG94ONtbix9e7Dob2g
P+FtaTAcJdqPtsLBi1xphYK6C1fOxpggmkws+QkZX8siVbAhLg0dTq4XWBcroo9gPfqYZOqPtxt5
nTlyX/cOkYKhwutRdkuhXE3nTueXx7BLOHxmPCstzJ98KsjOW0zA1vBDDuCZ+9Og13zZjqRIoxeU
NBxlsgjLRVZ051vXJ/IvGohyQ3x3R8YVbp5ybyXY5dlVo00RC3w62LLMslXSWTU8to1Lo6xi8yGy
ZA27eg3b4i+pA7yTo6f/5zaHFjJRXGyQg6Jywta5Bw9j0mIZw83fpuv/c5yMPEUs/V0TYbooRWdr
AZzTwGSGSfa7yfpRLI7CCcxAnk14YwGlI9Jzeyv6JsYvGSbhvAbSCYPL/SCpus8nZfZUOjDV5P/+
OPliW59wmYsDKveqC4SKzAoaAl1qWg9qq1V5Xw6y5tPhA1kqJSA8AmHSG9Y+3EvCbtN/2QOwToZK
p6G7R2anylKH1ERI2Ew9RIQStKB8lfgY8m8lWJ3gnOQHhkmfvqsiuFuU3kDVHGyi2Wa+238iahzh
5k80zcuK5AUY2Uh5nq76lUQtTSgCsSPlFi3+R0rJQ/OpKMDChbwB+80TXYOxLxrbRWMH9HfyHghC
szFBXPBXDtZ+D6dEcOuPYUIPcG1i8Fyv78sIsIWhd3k2L17ns7Gxukt8hd++fLi+VbeSgJ4IoSct
0sgb3Ysj5mly0YVO5RiLhlmAKUQdIulJ06a5uASWasHpiGczWRPsp/co+a+lKt3uiQtsP7uCDKAK
gOayPDlyl9Gvz7Sg73+KxAFOJLTNZrBfek65RXlNdN8HaCehBIoXIG0qclALlTXLLl0+tvdnk/xv
Gr46Fw3UISU9ZTqmfflXi06iSXMsYJnrT6AnNgLng+ffY5En6qJXMdY49oLnEDWqJOtoMxguL3sS
0INiYGXFNmZTZTd9RjmsgJN8ODcxM58zllmSvoFV7ngAxX4lAI4Aw/uqIvumt5dzVghhdjJRm6kv
Yfa37f4BqZ1hhMKXFx45rYKS4YBJt11MG42dyHSqKzPtMgt3AiLCF+IsG2Ndi+ES3qWel61XwbqV
qIk1a09rl86L2W0BAzYFxB+kKiT8Z8XuN4Ygp/Gj15/3SPveYxtzcF4Q87dOMW3mVdiHi/BPTHhW
2kcp6qbBLsK7HqVTYx1UyhqVzvCMSlE9oIikjL8O/4+cpVZqqFymRrhe6xSLUtbM1Yymx6pVdFht
RySKIbGb1KCbnIAzfNOgdEz/7bmAhnm9/m9hwGRYqJedaB/st66eAr0hFmo2BiutqQ0c462vqTV+
1Y2LnJ6kh8Jx4Nu2hYjknSn3osXhlkf1bH84FBE4emZNy2EY2qxis004zjA2t5eTumnS8HVhQ8DK
TvYk6gCJ38aeZUfSvI7C2E2/V2/tBJl9vqWiNia+PL784B96JOdkCG179akGvJ8mvKkBOkJtI7wJ
yMpvBlmvPtwQ7eL1Y75eNMeM2pkfjHRdljAoHpphNeuQc+0ETAo76zojWf6E2UtRGyIXZ5IBzHdY
31wQ4qvdqrGRiaj5fr0+XEk5sSaLbH6LN/UEt43/v2E8/DcRKmwiF8ng2dA9ty9AWjZAPXHhIplL
b2ZFZHCK6ylYbTld748qDfKGrBJGwB5/4zY8xAG9FJxru8Ng0uhqqxue1emmgUK5/QACIp4Kx80U
YPMtt2SKf3t9vFt0e6PdnKhMmBe1kooEf44xNHAgxcdmlxUNyZ3TOuHaWNVuTrgfgkl84BOugzjR
HmrP6LMDKxR4xWfxTn2jQA1Rna1h+SKKzm4MD9+658fZS4/8krL2sb8SqHPZnEmm1kxZIY7wlPNn
VpqJppsrz+UdAQFZocnCelWlKxxPpLJPaBKQtI0l9rFIFarpH7e5uVyQBFW5A7Khf8nfwra6PSvE
Lz3miYZw3fKVdDL+tC14XOyNYjiPlgy+on4rSXMLpVNl4hqF1XpQ2oqWYXckOJ8qDiz4HPSDOX1G
vJK9yi2js3iHeLlaOzwKCMe4tWrFfKKix4gxfThW+2Ss0pqGQET3R5jDN6Bf52kV06RcGJLNKRkx
kvwVQm6rrGvWweXKLF6agrvWIYFm9YFTs+ZaGBjCO9tBdYGD7rG0yOoo0gHCuabbXwp97/TZk/Bg
WhkaHICFqUPqVHdQj0EDqwpDnUM12mPAYxsoIG8hcqzzd7V5EPKu9LsLhg3l6iSsduuzwPzJ3UOB
fHcuiIBiSX3fSrCo1mtey2kXIctaInQ5BHld33jAz5EIwB58dvOSIOXZIxufIlhztLf1omfdJ8Re
rR69wGJo6INE0i4pgRxEPDxSGdx/31A8eTFA58jZdfY+7GUoMe/ZtZjLKNnX5qJ7FIbkgs5LYK9c
khigEt0U1p0F3vUo93d5eeEwa/5Kz9RQHOkpiWyAUigP1c3rKVZIuGerLP/nZrRFZpR9ndhi4o+R
E5/m88xr1zuLqTfO9aCr+sg+JN0Zsy/OGnUeWx52snjGZP1/tbHgLcvAFIoiDBMGykkxdlNdz/fa
4QEnrOlSlWv0fV5tSJU/mDuz/btQHRpGXZg9LaO991FVZca7wkOhHxo7WWDjgbbobpKq9m0sxN4O
/e/V+gFC1Trb0Z0OxFitPEWyA0f/HJDMDi4Ht62ZOEP8nQt1e/eomp+SGeG0wW2u+B+5LzJJAfJa
YNgfgSBPQNgoVPm5jD3DqflfvaxHMDqCvcXH2GJRCpWV+ZFfJJUt+LNcle9EUrs5fTyb92OOZkV4
Vf+ZR5sCHovOVQBZqAc9GSJ4rMrWmEsMVU0FnhPbAqmy6SzqHvmXn1sVmwoI+bM9T/onEG2ceA7f
KGGHMaXDZ47hDVa25+eZQjZTBK47GSNZ9X05jSteKhtdo0kjrEsZnkPpQ85KzoHGfjfvFqhdNpUl
/kOYNxLrFS7WWY9hyZjFe7OLuy+Uz5GsocBWYRDmluH/9UsFrA9smpEaLf4ciFaB+5UERPef7PE+
10Lhk/jHAgMUCr1F72ATjJqCsazBbbOAz/MGnE/tQF3VU+bZ8xm8bPEpquH9kMJO8IHl57ggjQaX
/rHPLeBw3uHlYtMHIau6LNSYDA1m+UkR0OMgzMb/+AYveeQrAukp7eUUTuwKKeLr3VYqeU673ie3
pj9G3dFta+zE4s1XkHJ6scD5Ool/SAj64otm2KS1FWYVLRa+WefU0Ncrm1cYj9aJyxyIoBu228UP
yPaqox/ibpwZuvB6Uvs7ZUCJKid9g9Dfvop/WT2bnnMTRfZtkVdTw0mNJyzo7b9Y+x4zL9AzFbb0
KPvFKVKrP39yyv1+P5jSqcfgtFH62KExLtx5dHoOg9QTnqPAY82TtuDs5ZbjUlm/S35EzG2Fjkz2
euQ8PGxrghse5qj8MxjE5OmswC87x4dyLC/jGqT8GmnnGL4zovYkOvU3A/8f9wgfe/R1Ug5BN0Tg
BeE4mJfcVB+IpkrviL9hEXmpHmuCiY++TCqAWSodA+RbuUEmLPo+jG8s4t0G92ctvgnUUSaXoffM
5iI9LD5JRreG24NsC0vGkFJRa4qrAChWyLRuX32bjSpJtFmJV9VE2+ehu+9r7zSKIx5zUbLEvpNq
NGbpLkhOgLJISqkhjAQZdfSkxaJNvQGhoLGstX7Y9NiTXy5ljxQf2Cn2GpUnSy5cyakXyUR7hkh5
Mv1frllgDW46jEtyPqZFuyaQ6lAcS5NDY/Kn8TDSGVsGtsL0cUhTtMVrL9laAwOix1Ra28MLBQaH
XI1jwqszeHsHHXaQmQ55rcDef1n2mtOOL/Vwl4agDdGcBK6f8FCFTI1O7EZvAbzCcd4f+ckmHpnH
c9DJWQVXY8fRWWtlwCEHoxd6LbZq1eKUa5en85TTptFeCiLzvhJMOlAtlCyE+GWqdOa2v3Phnwvt
yo/C5XpPzuCzq8nngySlKpEh75ZTFcZWQb1gwOR6BgXvxSz9Y8CeqBT9tNk1+i71g63QzSJVJqaC
LN+tibl05NH7u/273a0zOpJdHSgLAObwQcQbje5IHAp2CZ5GSQ8G82QiO7Zou3WxjqLsLWxciCjp
aHTSfnjgNixaroZwR6UhWqB/phlkJxDtbe0ReHtaq7DvRGo0/xJX/C1ad3C1QXqQQrcvQr3BIHy4
V5CsGy5JPARPagzCCf2RdRS2KF1ylDIcCr6g7yhThVVrYKEit5ePBr0sJDexz+J6bk4Wivrm6IjE
BUnfxjZ0QLAAO5oFdju83Ds/PhZa37Uk3qkaChEBbMF2PNYF1MVfl6o4Tfw7kzndTiR2xOrHMMtv
Fn/EwPlahTkPmjKIHYnZT0HuWZzesiJ7sHTCGS/tVWMl3XoBqYpW6/YQIJC/DeYpcqvReg8mtVId
YOBPgrhFECb8mWnCtCtN5lhhz3WnFYpP7CWylfmeAy/B+2P0rXif2LeZA4oWUvKZT1QMMzN9H4RN
bKYk2ths+98kFr2Wdr5vHq1fg0fGKV567x8m/0QJiE6BARqjZMB/KO94mN5N/cNKzRnT1u5oA+Jf
4BhaDIX9TlLzlGaM8K6kfxLWB86bO3RynwRq81nSisSo+M/AN8gAVLgWcEEaWAFrQCzjJj6PmVGi
qEnZd+zNikrM3Yy9FrSs229uAL4o5VYuD2NiHNaFbuZ6CEYhNMxDYx095YQMSrv72cp7uVfpBeDy
NtA+OuygswyRoOZnnydzI2+BEakCSPqlZZuHjsFGpQ/0ygJOZSCN3TuP2B355glX6YNLb9ma2kMh
0jl/SrGv+AVRlABi6gN3Y+zpYoXZxg8yZuyB/FDRY6XGmkzeSn9HRGzumUG0MM4IfPNn3WnElVc/
Rmem4WMQ1MY96kpwgXIDQyyXGwt+iG3YLGQpRoRNlK1dTj9e2SI7FBbd3IUIWITRBkBz5u8k1HP4
9BmuKIky4KZwz/GaZiqJOI5cd1FTfdo60njNANbSvFThnaGvlIjv3+MXARRsmGRAh2rEeT3cj0vr
F4x3Q1Jr2leTNoEgC8qeiAVE/CSRgAaVCVEWANhXkZzAJdUoalLDd+MkCaC+83q8kZaWwJRgiluY
kekffJss+/LewoUDtLn4UXVh7ofCa0E5cBkK1EPSUNmxRTa2w+hVvA3nzhfvBPp6GoPVIJcgPMcI
bUBHmKMwRC+rS5c8ZU0eiWTdkDidJjpWik8TUhZA+5U4MkVpOYPzfMVXLofFlI+dCRhFBPVjQ1iG
u3z1m0yl2fy8G5hFxlc48dLciPS8dwLkRpLSFY481UO480xJmN1K9oIgBQd/taCRimAqCIX6mmIV
O39L1wuyX02AVpgzhXu89QaMh+sGhQ9wDuuZlZ4gd6IzHO3s0yRlK1WleKyTGGnFKLmjKmL6UweV
qmnQr8qJU+cskFs3DMyZ9a3EPnHmMLs5rHOkVyKrizW7zoOHpJlV3wG3nTo/Q2wloG2/MG30ZteK
l/gkhYdQtSnfgULv/v02+SSIEIl0lP//85j87dg6cGC4MVR9Y6mM4cqrQcaknFgSvBIzBIbZeBCO
0DrYfjslvQj1SUfrAuWJXaKWglcfTyzLXivPCqXK1kvokV5Ba6ES5y5l+rbiZGkQLLkN/o88TOjK
X27qbTWpHgwdy3ZdXT01MpLye3i+oArvHq2OTzV3BYvjVY3unRef+XupKHLaM8RXDqrvTV/lsKyY
YWtNPbFi5dr+MaPRlbugVghI4inEukXXq1eaw70eM0KR3tz52DkbfqS1fsCtbC5wtlOsFqqJa7sl
Ln1MiiZxTV34T2UvTzPfwZ6DSfnSgNHqd+rrfHNMJ1p3c2wS2lSyq2/O9fSPXCZ2oM0LfaW6x+ZU
3R6/6ZaOXsvvdNWkLrP5lhco3+Z2pFnSMjjPxwZhsgKJnW22W09oLzCE2V4G2pfXF9edWxQqcGZk
W28R80TM25bGDiT6Aor1kCOU0kafumNSf7aLDfD4i0/Z8syUlOpSDtP+8OW0dlbfZv7Q7k0IPFll
CRzXNgpLHUQXt7H4XhOr7nKxwkdEd8pEIQTo+H697v+sTJrI0FXNVfpXJdkbn50oayUMRuLs/h7S
nCi2h8duTKSKC7ZRKNC2PA7HZ8SbO8F+9C4yRq1u7Y00ETXVJw4ShpFMjEckI7p1GGNz7NhIapuS
6xvNCnuOBdFP4Lbf2eG8xtaYO0TXZkRyNcD9NMoOTb3U4YEBSZ44V60ORdp+I6d+9t3cpToF9lig
ANS9nhHJDylibGCDioWQReKv355ePA7gOPo8EpEedv5tZGqWZXejkyU98lXNRpBaeOJ9EZR2hqtV
o3Zj8IayMiBVt6NxgAX7tROB8/J/1i1OQrVG5T2Kt0Ut3J5XxWI8kCIuA4wQNfG6Kn0pTQvjGcXf
hekFpkeSWvYiJdEopkfkpaBI9tGIlaQzmfjmdR/jYVhcuoDTmGpkLa5eW/TfRzIGeX3kY9Vs+0Ka
GvcfqNDt7Z1J4NbdX49NR0pUgRDIXjIRVIjP8vQpin9a+C+8NB+gma1bFe/FxBW+a4sVOaToDzq6
yTvI0mURsxDKrN8tzBMZv9IfRH2JeLSDEvfRx2ONaeg9wfqKVatpIVrC5hxMRtq8yECX0JG/VMXR
qcSmfWFo8afXbePm0NPAEZB6UEqk8r5fTHTMG9cmBs8YGAp3yoXZpdwTFSjZVjqkE4ZzZgZS0Qpo
lmDrT32OTrcSIhg0rQi70vTDquP7dICyu28naFSMtSZLDLEUw+ob+Yr3/DyHIpgKk/2535skqsq+
STqdTsbEi/4xJQ4P2dmgWNR7nRuijN1jNmVy6SbzlBRtVi4Rs3p5GzGhRMp61fCgBkr+CHRwS195
/fn/ds/vjsvyE6scmf9tC0NG93GhZCR6CUuwQSIbX7mUaMG6QqALcKRP0c8Nea21G4IlRYrhSlZO
ATI2QxdAN5TRNdl2GYzuiyXXRzeWP5YWwASiZUfSwVDTavjjSelSfXCBi2vaztAYQyQOccNap54r
tNKQNT3RWMPMu4r3mXU0d3u95K1gqhODTwl0t3ukGlFW1xb1s7zQ3KtpSJmAThXX4xtDFndL76PA
gkQnUdqPZVGcVYz0pRIjE522Hzn2ZnkVtJSLAlncNtPq+zeJKwRBpNZhJ1yw51pmHVPGvfVjULFN
UrS0m5EYJdvp05iBnJFW1hlEZy+REawel6oSZzisePGvSoFGmZXyl/hJ5elbrFhVUQKioUOGYfga
h8G/9NEzAgwwgzNaw+OjTQgPHLkGaf2+9Y0BRZOcLI0Jmd0SI9PB38ErvC/Z8lRSu+6L1Th569vn
SLgdRBLW6YplQFg8e13jecZ5iJX+CpqixEwxYYJM+w+e3GJyEPM4Rru6wdNM8+GnbWRbVX/b15dY
lgRE4X90zxqIkqc+2npDOL/N1rs8+g5DQbse6PkS429Y9N2o2vBp+AuD4PkfxaPjDJY5aETk76jA
1HrJ+u5wuJ5jaPJV8o/zNqH57C4FyZElkelDjOu+reswu45Vyq7YJkCwj1OAOfUPzOaeNJEjGDpY
Fi2yYX6YIErTIZvmj5BBo0pbb4pi4Gv2gtPTbqU8cOrm6qDvqVr2iUTSOPQkK2COJUH2DCbCBTaB
YjIbkLWSRhvl75bvO+nPT75L0nmwz43hIAcTrdIA07WzBs6j6t3sa6MvrVMUXiPreKrRJh0K+bBK
/EjenH/Kr9YrRv/tCAFGz+ZEEtWEOfZrWxHcwqs1LzRkw/0ngKmHBFOX+QlDnEaqFPcKkI0UPSSc
DOGOFYkJYmZWcaiTo4bmGe7nF1wD2bTOzi9ztcSWcqxdEF3VzfwfwjuYlEgxD6p6V6H7eq3jwnxx
2IGNIJ9IUCg7trYVDXvnV9aX7Atzsd+7OaZTYoyskw0coQmkpyQjJu0wLYTT2KtB7G9B3dHBp0Uu
nNSorOVymbn3Xxpz0op3eVK0bC6xfm6ev2IOIsbWRrnX0qywZnKPOkeu8m8mvaN7aegx8FTbYDaz
YaBdaxdoCGKyJnI0fxRj43i/XY9NvBGe0gMJeGpkM09pWWb2ER2bleZCUfV0cwOT1nF89t25JoyW
g/Oy1wyS4m/TW36qSGKOqFr8bU4qsFVaIFqXBybUpkUBovs6nYaO5K+Vgtig/uCbdIS8MaxqPXeF
SzqsHCnj/tw5cODoYRRJWRO1BP2LJZIjYCHc590MuGPD0ynHNTv5PVneKukEQarqR+GacBq+wZfS
tzbt3iXHa+bbr0wrlA91hXsU0O2KEp0hHwyTEFlzw7kaAU3pJdDmaOXmJ5Ngap8ma+1jDVf8niq9
ruSRX4JOqLcAVByE9l20hS3hKC5JoiUGc9eLhwfPwv2IQs9p/nYbXPEmQG8gun/6CCKvRLlCng/d
heXBD9I26vcolHhFi5cxR5nJFRgLA0dcOt3b/vgri2QS8EvE/4tlznRWvAIO4URvAbG893IVjbA2
ApJPZjME2QUNnbgoEN3HNQlQ3NxzTd0PhX9sQ60ei8VNNsSWb5JXXQMiws7BrkJE7OT2R4ar86ky
Vp5AX1L2Mhi+e7RRDnVU1UjsSS1OEtEnJV9jGIZbcZZ5BGeFBhNnKe11c7FLLv93r+26eJSF7vTc
Z7IkRkEaA6WwFVlg504FGGSeHgLHuu+sBTw/Y6pEJw/i979NfWKemloo33Vti9BgZ6czgp6krfQd
tSyBOE0+6/aVDDDKR3A6WMZSWBe4kpPe7BI8SOty9f2asHs/SYX1/vMPDLBajACmnJjGdta+ndf5
6/H3KTGbA3TMTmFZh5XTatdppMyJUD0qyQMWSCGnOyTnBa+drMDYsPjzaXglQuIhMWWQL4at/Irz
j3S6DD9Ufvic4Q0tdXVPUpzjkyd5vUecik8gw8EOoTsRcBAHj8Y2D8HHhqmkXEJkVpEravsU2rPN
KTLDzYr6S8cxT5yj+G+9i6p/w5+Xb0re4Dmi7KjSnUCZVTpIxPKHC93Hf1w+aZA1LYorubyc/wS4
SXaX+HmR9KcnnKBQxTqtIFsxnZi/fZSBS6awEzn+v5FUB0zEk67nhVlbD/ov4fmMOgsOJNfRFvpX
hEz6ExYpvWzxsVteHNYMfk43IugywBTx2Jag9lrGf7ObTdPqVA1TsQMSE0OFWxqal6YyHllNG1qo
AWUWAUlurYr943PFuqwuxKuos8UY5hrPV0Zt9N7bdGwXIwqTSAd6CgYy8AHlE9ExqbFGYTBTfiGw
8CDUBY3ec0FDw05X/w7DEDk3gx2Xl8wp1jA5So7WLox8LyL8z51BoV+OcgAPUFETjpWAr6LGcpCY
OG6eDLVmccyW19KoqsQqJrB9pfBspJ/jTVBTKAGisLoXwk7QHx9Jt2qVcYZEmuUAXgXH/cO/l8vK
J7qTmLMvInlmOEV1Dn4v24TCO2wRGT8+zyUWWx/qyBgEmci6ws4ae88tDtqJAYgVSyCNSGMduQHP
dZOu1OrfTmEttr1g9F+lR9/fQC8RKMWP0LrmDMjjvxeMJcC/ToMP8x9UdYG3ZFy6aAYLf+nKEirp
97VwgPVA9EnZjwOYnfYNuPu7ihz3gb5JugGWieHkIyvanNVBJ24DI7UEYdBDP6cXhJVWAZyj3zYM
JO2Z04FgwZzHUoGh6XTD/dq5tNIO3OId+XnRytyqCfex/kdNdJyotNS2lrlt31Lh67+4SosgV5BJ
oziVVEKEMIO/86RkTgU7V2JliCZceE82nOFRNsBR+Sma+M5PyH6pfoVaM1L3c8/iMumQMh9knabA
a9goO8Ehc7mtcWcb1SMeOiJDheZ2PGXP00nK642S9Rry/yP9IuiYY+kVaztjGQnADw8lA2fSZ9XO
m9B9cgO5wLmMoogWeau7PVKEhfG4XSECG3lCm1YuzfF98nvfd98sIyvp9TTG1X22olDXuh6blBe1
2Frkp9pcJupq4OjQuquYqsh7Cy4JC7v+GHr2bnFWjLm1meXmxpQ/XqcoQkH9mWAabZHvkBvgSWpe
7QVc3i16qau7PbvgDUq2Y/KRNEsClWttmPIr4sWI769AuzMTA4JANiEQt/QFcREAyaTOjZOoYT85
NKOkwhSgY0LkjReiWKt4sBOueclzIPQeOqzkpbBSQUne32M1b3snhul0g6YRNI38aZi5ZkdEEoTF
6N3m16cxwBBCU7CdSHR4d/zrmog8MovCNhJD1ElZdoDGuIQcjZi9vugceEduHmAxQu6RPSNevmul
9eO9DW2hmHJBUk0vBOB3vVSIhuo7HFJtmWuZuZz1GNf8WWBDglR8x05nN6XFQPvUAQDdNAkdXzmc
yaJQ7iX9jbuZd/TxTYcsmsmeIyD56JlpphiJzMdJaVhJhBK2PtMsKPuAFjleS1c/7XhRJr6Dyr5k
hm7uBmLmP1dwfBIn1G3fp5GLyP+jl0/FXX6SRXEwhK4cPI6NRP9PcAD7rDeqRmOuJv4NhnAsu2as
SHlj2pqh4WvR5FwBWXuos/XaGnCvY1w8DGI3MEz4x7b9Ccbz9NxyKt7K8aZm4WzHvQ4BsRkTs+v8
ZEOW54GBn5ELDxwIrb1MprZjunJRLWL58J4ueNzCp5sOHOvx1SdMBdsd9aeiXXPQW05lTvpjgO1V
7suoZrAxwSCnQm64o1V7Xa4MO5hWfzhVX60xRBjDE6YEH/ef7QcavKof7zBU1816GPPx7Sk4d0cq
APi8Uz3tz3slcEm7t4j25GL3Y0h0Kp5b6XvqNGdQc1Ys8yz/oH+Z7FvVpjiTQl05lzAqvJIoBR8O
jHYl08pu795LX1mtFd0+SUPMkP9tGnm4Lkv8rDrUrIhXDZEcsybyb7XE0S+jfoKq7XdxyQgIY02M
lypQguLkCSAAkAT5vy9A2eaB8baG+mNJaURHhBMADLCfPIDfk8FjI1iIW3bbslYIK2/KjWd2HQck
wh8+5WVp5EQQDTqQze3B1vIfuDMGKj73ryd+NeNhCilwB43IdwLujAtKVRfnDYM9YPp1RNX1ZChS
4CsfhBlkpnZeC3JxAV48SARNxZdYGZSedNJVgaCXjDrPEoblh4Y+EsccssbnIi8v2kkeQxqCOpYg
0sLteX/XapqM6WsQaxuZiV3KdMStRuqc6yMS6ws/zoI5e0VvoWHkp7czRJ2HLbLM8oL+paz0/tdV
NT7ECiVT+LMJfxfHGmCl7lCrcs35NzIeTXk2wHTVLGNB2F3n0oqhYMhOp6kgPe0GfuPTCkCYajuH
/75PrTsVOCPltApmIy8/A6g0E+Vq6zYW/U4CMgiqGBIRPvFxx7/+hKpzEAL0I1+mjoDkXLEgwdU3
sLgeU9ZPzJKnO++QbPzoHwfsSCzO6gRoRjWUZ16k3dC8zHpPBG6LkvMADwxkXFrlBRAowIr8np6u
MNHg8CrYOoMQIUe5xxIQa+82wW5lfAL1AIAzG2+KYGqzUTxQCMY4SBICkM9hjgMhLTVphXcIe8UN
P/1v9VxGit7bq/LqJKpmVIGH4gv9WCz+5XV64Zq6B++b5xnRKzJ9drY7dtXNGhhnZOxLS0Ow9rro
VvQVPVB4I2xiMpxe7tKOh795KiPzBQzt81ozZ6MdvYmbVMysCKEvwEcusjEfjN6J8QzZnf5xZCA6
kgNcFIHDusIPd69spVfnlVffKNxJ6i+aBI2GIGzboJ8KIjq1nX5QnXRhRyGE0fQ3sMcFnCZbUofz
BFICIDM14pXytRQnmMFmnDrGeNHqOUc1OuBQzGR5G+E/xPz8GEc/8mFJqM5a1rnxp8rccocLZSSs
NNz/V1PF1vHyaO+PtKetUJD5bP+KTQZy3D9jYsQv9dgSMfPn+JtungDgUbrKvNR4WCM3MNunRADS
s3axbuKzsUsbwk+xmjdUbfzRJU9HPbV0wAIatuFsqLQnhgH26lkfhkm2x9WVYBD3/CVRZHTqLnvl
J0NqwsLFG5HFkTjcq8YwmX4hqMg6u7egAvLOPRe9YMkQ5mA/lqXEZ7opZ2Y7xGpYoIFF8aBcNwuY
BY/7WYgDoFhMFYn2FlZf1k6xDi5znxxN1vIrELnutFLTu0vXKJLN8t5BSgKlQ43OVjNPY5AbV9g7
TfUKeH11v03+LeMvwbJpulFptv6N9w9+k1s5eyLegsigU2Wxmsk9JFr+xR+iWOVC35+clyT9ZGc8
o7fr/oqj0DGtsjpV02WCz4u04h6F5+lhOOYU++VGU6+pr2MVGYNIIOou59vibTRhS9iTK/54Z4w3
m67wZU3KAljm8fTzVgIJVohmyt5/Eekr5fDoxQb2/Bf0RSNfO+NeHWb/irIpDl/roDCtCTpvZrUc
zmoVzGzUswRvMh+cw4eSESc7AkOIYJRbBGr7i9AuH1/Wp80UpZ9U0Pnkq3opFqSw31LsL7YtCe4v
trpU0/xXfF741JxV2y5apMvK3qmdhQsZOvbLGqOPWoptoWVw/hBdV+GtNEf3LYO9k2BzjQcnnO5X
JZYtyRhtnKBW4g/Da2rjpBZ9mKt9EoW4Hlv5+6HorrdEnu0/0+KuotR6yH3LR7pvrwYpBOr91px8
EFpJMpXqrxQ+Tu4WnyPm0RtrM7prkwVWwxAWYZsLzOZXuKBDCUR007qgkXa7XG+iXDQmWMkg8/xa
nDqd/8JsWncFHxKybVgUNnDiLmpzhjTVfLkn+4lpkDEKeCmt7lZcOYpWaTb12xeuDTcJR3t5L/AT
D23p5jjUAVZ8QQAg5UufG/OcTMy0jSQFg23/nIh/ApOWEpCOx4vxp/91BR1dDOoD7++geKEoMxWQ
cStKu8BitV2G1zlGIKdGJA6o8/O1r/65SlV9NL207CYCcBTEwgFoNm2Pa8AQrY3TejkyJWnhnPJX
sFO17X/EozSlziC9OAuaplcV6NeNEITZbH344ojifK6FRwgZFbspL4PPG/SZoX+grp1EFOODal/T
LGUivGzw7IRkhKMDiQMANANRtIk3nb9Fs/ubD2uMjNd8eppPQRMF+lQ4ZvKblIQZiVAsl/L5RhQQ
kMyeGIFxDA+dSLykywYDr4vng9kWrgJpEIrnTU/sMnKo8d7wenSf2RPimf9lnWBKPI+vNmx2OUnH
GNd40uYGKbzerp21EDCNDzERpqPMlLbnIoC/jrw8tYSB/l+HhUABMViR+DdZJnsB4axQK0lsL60r
H+3HiE7KFI1LmFJRugIfi5RRZYPZR3Ik+BGbHW3H/axSFct2y81YaaJnDofTE209w/zcDKU51Fe3
MauUtfcVLFJBHLyKaEqHReM5uqzCd6ZvJ/q4FlxJ4EId/m/X3XHhmcTJfpzpk9uFhyOj0ofinX+T
+We+WWAAXY6J5nryg90DRQL3R84p0Ub+JAGdkNBvXhtKyBPjU/USmTYU400A1GLnSOeqoZjzL4HP
FReSNsK265ihCsgokTsNcYMvZzReP7TGvTpGz1ljFfQzvlXvixotY8050kkx9u6T48lPfx6+4dqz
omcA9sAxAJg1Kwk0oe1Tm+Pncqgwn7WsENXfc3WgMNrCGXgFz008yTtAC7JymSY5q86s6tpBaN7n
sgxkW325JSIBYxPmnY1IruKkZPVPlAq5ZGd021s0l8BwPdWjsVdAXWEV9+byXS6/oEKgqvjpIjzi
Un5JhybkbgQ+7Kzwqb7SMbZrbtLUsOj9AP87O60TslYfhKYKmpOd8LbEOBW4Jtw6PT9t/6HQYbPE
H0Z89I3WQRDhUl/vAV3laVUd7KpTuPIFQkInAldhfYpF+73yNaDGySE9/xfk6U/bsaMH+1X+HM/l
R6yGk16tHqVFlXaDhDfJfpyXdsiA15P5Zu0VGj78R4UeEi5M5cMBbObjFjqUCplbZ1keWrIfChGo
ZuZob6yd8qmujQIaXM8EgDyP8O8PEGClkKafUKU/eQbD5uNuownTsBRxKN2Zz4v+H2qOBshcGXaV
7R/7o8X129WaV1Y2MewB9k+QgE1q4wpHnaPXosd5NVOvaO1sNHDY7AKTOkPopaL3e01km98jAotd
xveYxlhX8VdgFSf9rIPYNwm03diMEYdqiYGWW7LeH7LPGthPeEQTmfCidsulVON8VJ9mJtDTmTaJ
lE5i/WoxhoXhcWisjGEbScpRV+4Lt8f/xb944z3tcpy82znio0Di8qanLOc4lUacQaePrx3acxUx
Tf43dQXF6kp4qjZZMMrJs9e4XLkkUAbdqDHHNQqNIZR66mEFv8NftKd4gWtpbvzUUfHzBVHQOcj3
EtFVpo/tsJ/Bta4vfnBHPEn6nYsq3ovH9c+SL/SrDe68invnywgZZG7ISFbS+omnEiTu+1vl5F9B
S6eD6ktYF0LvMzvIuG04LSzlWshHOi8NlSscCMULA1keydNVqarvtUo1LUP7H6IWMht3yNZDaBn1
areyma66hYkEYOWysM5rh2ZAowL7jTxIG6w8oghFDhDCw9SKeVbV4wVSLmL9nzTn/477os5P1jBg
sv+Chsfo9f3eTMxwopyf5cMPssdx6nA6KlFqSR8Mn+4VDp42sBz9hnqG5bmcLIMrzZVc2H3ggW1H
DIPqWSj5weGHjeZWOpBwmus2glPIAXXYGyrhvmmdvtgSqZerbGhRQ/vBi1nwk44OxoDyIPP6xL+U
QsDAVCRkEzxREM/Eu4wI0B+sha1J+y4YuaegoNl87BXs35E0pBakMX2J/bh7+Gb8UPvS+6cqefOI
8Mipsmoq3kxH3IGcN9bGNkSIzM5KRno9eQmIpXiu+fQU9oYJgPQ6cPz8Diea90x8TA4lCIvoEDYv
MpFTzezt8ok7j2lVoa+coQSa+BYuM7kh6VR4zbQsugEMStCEBHbikIDBz7fOzcMy7ukF1XQZIu6y
ieO/+IEbhCQBj1H+IAe8rbkkXMqxhhr95E+uGPsjdkiJK4COFRuIeHkTEX4NAOWFB9ulZd+XxaBg
kckjClzQmMIPoBT8MIUHwIh0mr6GdAdjPFcEeZo/BIXeLG6yXfEJvM4nnf4lnpPZJsXSqDg3VEUO
zEtxBl2a3Sqsj+m0cLVaqnPXI1HlwQ5XLvvH1GnlW6KwbLFshM1OrDzqsgFmzypFAe+LfC18Kh+m
6WfUYi6CzeRs3mcdNzb7dxn8JHje2dmsQVAAp+CT3cFUQNlyJYZSEaKS3CkQmXzK8Xz6Oyd0+Zjd
ZHv1mGWHAJ60RRwxE6azk6e0hQn/f7RbVqT6qF0/xT9+lDVYz7Rtg8VfTuHqtoJRWmAs6hK6mN8Y
8QR1/1yRGZhUpFVOggTr6RK1yhgGDc6G0ygsP6BLf3RsqrLysingftcbrErL0vERrZcbaHTjELT1
MkgJ5gZt8zlguQ9sOA5MFjTrSjkC+wJw2yrmXUelbDGHI4rO7mcAqD7+dUXo9KBsDoTEtaSs3L1O
V1HWGc0zSDa8GF+8vogiwiva7dPi+S3Y1ZtNe/1QwAX9p6doyNdaEj6y2b5pBJiJPkXHeOrrJyHn
zrQ6wKPtX6WPzqVp/dbSAmtRrpmyT18QwdEhibbKe9Tu4KTB9ocE1bHgrS+JHwNPo7Hj4/UUOiR9
kcSEj5mjEs9SCb6HyGDqu23FeYI1dwaiDQYFUomFFANJMz7adW2fdBnPK9kWR2aFYnZgD+2nTOOM
UzMowQpO8C/B29JP1HkT26dzi3nxrSYR0fP2v1VqvpjkRfwcSiDEgU0N+VWSFBDyGFF0YYwumosm
P4ngMYirNTXzYaFrgl40+vsA+mIxOiwFEIXDM/PyrjKMsUW5YGH+KCiGk9B8nOU+oWkIuNjNVO6X
/qBkqBOL+oFTOwhYDcT0Sp6ilM87jKvBDqunpkkABa5QIJCtLEERa8eMllWuC/jn5ohi7/aQx3RM
u/EAxLzOnAH8nvNn5Pkwa3p5Rc9J2dxNERqX5ZC3FD/NRRGznA3oSu3nsaDoupn8sQ8D7RwrfdRp
6XFFeSB9VkZ6p/6fuzEMpLVYtpUy3WRdssb2LqQo5beS2X0+TUF/Ko/JZK4SZTX59L/n20CVAKkR
tABHs0BK5jE/U+/C7wS5so7dglfKoG1pFQGvJciGgZdByxV0JHqly4KAkyGCB1xuVWMiXybQLgO3
lzuDywk2rH4DTFQHRzjZsgdaE0j9Nm2jsF7RMhiTGMJbl/WAZBRcde0nq20WCqO8y6crAhSVp2K9
PDlHlk9Giq3A3tuYR3EIEsfHWv36Sb/ewpAK3VQubhGN1Hlk1RTeajFzysnsBOBlcnoG64n3A038
6JR363z2TtfA/H+rTtv8+1GHWE+DdzPv/h3FBWZTK/nNkHEs+KmrVOgG3rShaJ7ByFDmy6/vcVyT
qzOvDCCDxiBl+t48R7FGwRfRFFdN2zArCZ/4zsGTt5Rl588FYBGSieEpZPWxD3202m+qPseQGQW2
aWv9kwOI0u54gGSUYTnOYNwWezo/8+i4uv9bjMiOMPKueRVpgKKyvdoZVA8RqSB2xbPy9oztFMdm
e/ieXqpbpOXk94y6tykLyGvXFyXdAlLrb2xmndcaxA4pRSs/YMIiVKsXGvh/NxW6sVbs0gkfPktJ
KhZOV7konjIBH5ZPRZKn9VW+6ffurIzHPDIuFePlHzsZZMLm15ywpcEp2MIsGbJ6PxU694UotwhL
hZKC/2Y669tjsq7MaznqYI8xRKZheQsnGUP22J3O0BjxDMldLh/mfyJAdGaPYc/GO0X7AQMw9OrT
E6mbhJq27UfYuijQplaFWvWfBQ8t4uyNq2vYTq+PI5mH1kJ7iAtrmTepY5BwtmYDLJvj1McBKKL6
ZUuJ+yrWb7n4jeOKRdRHri112mWpvs29q0O7iN3BjlE0A546r0X/f7d0H97vwq9hqbbn21TjBqbd
gLjBFGeII2gleL5XmERnNRyL+8TuLf/IQv9KtJ8Trkx5B/diXL71yUy+/28gj4ldssAw1Z6K7o4c
E1FwoIHAl/MeLfKuDfo4SYluE54nrNVgI2SCkvNbwjPOg7MI54DRdJQewTjaGcktNtQZwUcmebom
NXrQUjw6seo4g8Tf8Dxd18O6a1Tptuy/33yHRrlG1lkVHfOhXFrwrm1rhMjg4FaPBXFBZG5XvJcO
k7sZXMcmklB/13nuismtfx/eCgZHawANRffXLjzKXB9BKa4kFPSwMgAOwhpJZJxLXeIpg0PcNMGF
P68WntDlGlwUfwSqdlNwa3l54DfnFU5DbQahQtlE/tq1fGbMVOwb1PXt2sByh5AmHTNIsqUbM4ue
jaQUgSv7MD6o24epiKge5A7UkwFXnz0qe3XwRGG/1URakdPjL/cI9bR2hOg53VvA4buZBO8ObPRb
kFxEcPrP2s8OhBuJn7vZwqXCE++Acyaqi2tMVwpkmAlh4vJ7q7dRAOeN0bj47WSk76LcVTCDO0Wn
S8VQfgZP0LaQdyOsQAfoEDexlC728mOtoH1rJV/hmoMwB/n1IdeM2YKS/uCxWoxjTkBDb42bPwsV
7WgXnsczsECNO5rYRjMLmCUhxPEhO8ll/ZFGCZDH+Ai847hblMsdqyWnM51QukL6mM7h0iAqitU+
p1X/i/wjyH5GbsmDQY3MkANazPa3wFCOWoi/3/hZ2vbzV1bxDrkyHddPEevpcZ6rGu73zHjzYAoN
HqvtVsG+K8v3Fnnw47Z3yFLJxoLzoA8hD7Kmq01zs21vCd4QM9qEf86SHpvKLyx4nJUal82jkMc9
2ESBguaTOtCpXX/XR1pcbYO7b7xFH/dGhL37dz2SSV4z5LySB8iw5GS/prOYVq4A1veVQuJucLYR
bBd2czsbowVUU4xr/2rrS6Ru2G4hD8JcrhSu2hIAHMuzMR6zwreNeWemh5aqRTi8qt3Yiey1mtV4
EmIo4f2OkocFlvX//+EiahrePSAt9F4YOwnmPtTz8EtYsGb9QBftEiOSh2eBEWN0axOJBWAF5Ps8
mY79Q55T96+KP2LuolsltV2KN+6OrkXRnJp7SKpufVfOU8enJpsomUNepjW/5Jdxyjg3XdEM3rQ+
E6elLPDQtwuQLUt19e8NKinkARm8tUbpLchZbYJdUkRjrN8ECN+tc2sZX2Gpzhq6606AdVrAB4NC
b2YGx5wX8QjmPAQXkJAbPJ11zItlJR6HDHVjvK+exseh8Di0D4DoMuxN/l3olvCpe25667i6ASiA
jlkBHrLDlcoSBzH2yFyjsKEdv1ioNMQ91V/achsdQW3COLpg84i2HJCDJvfeWC7Q8USM18KzX5N5
KjoYSJbttxG+B/DL9xkzVW+vVmcJtX0yfYXMJ0v0mcrTgK0AQR/hWcOo3hOBXaILEkJSlJc9ktF1
hDy+9IOURgCtjzrNxa44D1xjGrgvAOtuXWM7yzD8ih3xse+TAcJIS0QjYMXcBys2bAxRFzbH/mAz
zKGov/j19wxS9hkGhtXyWDpwrFXpoCZB2NioynVBtl9SZuATHB/XVVq6Ox5IRYQTGS+d0jEgSZmj
Jg+bjusFArew0QRaCijcRL1fAbctQzLX7MUEE+P7uES4Scsr63115ytCPvgeKOffypqUDvRzKHiR
SvdyKiyxg0xg/Qz+IWx8BJWFxF9WUn8YjwPgncZ+hyCL+iwJydRkBUuq+UkVvdlmZqMO/dmzXD7B
GT/7xVduwv5gpYpMI0Dmh5RzOmKcxZ7ho/PAkw==
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
C2TuGGK/zp845DpGMieArnZe+Ir6sPFA+lq2ndINnDLwjJNzVBqUthncBVMBhJgb
t2cVGnwKdVvIffraoXvW4T+HwaCrSo96DBhynmxSIS05iUzoObz4jDuMRWOSK2P7
cNCLKlD1gIK1HorZUlaGIIMmF1MEoYWVDHDQzzUzlbw=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 8592 )
`pragma protect data_block
UmRqY/Hz4pzqpYlwWJvaBhq/RFywkJT/brgmdibV6GB7qtUjfOaDwrCLAMrTdmIX
k60yE6Lc+HNvUhQThKi7KUubyFRTvXuu2T/NA2lkBl4ZBThswcUGvcEkr/4ogT19
wRWQLbcFlt7bfR07mKfmj4gKpQdxB0C/JZAl1b5QHw8nGJt5ngLPOX51jv/yxsL0
aO0tLHXxYzcjQdsLg4COIjt+azi8225VNcTEB3Utxyw1WeR9T9VUnanm8mBAYmSE
WYv26kZvL+y2Z+2WBshkV+8XytG+Dulf3r1T53aM6OKCqNpxgHEp2Qitokl8HKel
+Ue+2T5b09IWPzxeh0QKDA0jcSkPnkKxwMFYz1E1BtnIxBL3rTCgI0oDtIqCrLaG
7l14cgXqXfGFmbaYIBfgfy3eyCQbBOAXrdPrbBUWS2NN0hZWaWmYpzEie3nhxq8P
MVFpfmw5DUdeB15hg4mne6JL3qHgPzNSk+TQjpDQixcMSSAfQhryO/zlDy87VlPM
CXTOxBVbkaEI8wKPDltlv3Y2tfRYhFnDkFLzZx+0Tha7pOa5QriBxbvu4WClcllE
Fbvv8BF4R82/vHjU9ekbYZBkLuGIXeqeBjujzushmmpJOCgQy7Z+S5kd+8W7Tu+r
B7a932D6CTHXTFJlOc0+jicBT/vU4hIkyPM6dnj+Yi8rfVJYMPeUImPtYRXH3YNo
w6gCYFXpqHwLpyKcRVb2fx9M9aT0z1+N4CYLXJFLZ2GMaJoq3D86JFS62yTn5rBl
hUf6lkqBpCG4vvU9o/gh5GyUyChi/0XD0ucSoUt68BLylJcThAWSbTBSeHBygxjy
F2tazh3Eu2VOVRRhZ32JpgZiBVRT7lpaELY14fPg1T5+PQcGQ+gU8xHXeM7PCmjD
fKWNOQdkPhNrwGK8zxbGHgxV4SQ574ggFx2PJCIhsiDcX231dIqTrXF6vvH3MPzW
3KoFJqbrgL87WB/j6EW/hw0VcszztElPeiTsx8+JsBsUMhR7Q9ZoCBDwWK6jLsNr
dbRkDo14I2rOMZbZsIaU97rovrnRRvl4s6w4NOcYKVFx+yGtVFxDFqsdwmNDn5j9
PI2t2afnwi5FZ2pM9TnTh+Rz7YKMdXbIGxxwwVcvCeHx/Eqa0WdfkGfvJ2soEe1b
7M5RIVOVyarJ0aQXVeY2cv6hOCIegGQn4KBBsqlmNaMAgvJ5dpFMJ4OYjIXGtgJ7
nm1J/GF4+Vc9YU3Kf9rLkbZK1q6u4Kgee+37dWSmNDS8oGgXArzrJ6gSQx+gqWrg
NqBMpzveDWQHq014L7c21FICKS/tPMDp4DuBEpaNZT6LO+7nDggOALU5iDcUx8FZ
SG/dgx80WGnThQa9aA7P2KFRXz/vtqtTXA3tHyjgs7BIbCrXUMjbYjPHUx3d1hNe
IRa4SUTDjg+BJJPJWZ8C6/NMM701CmuzxYSf8HNZq09ofDc2VHi2mEpViwiGl6mu
cCkyXD+bJyUbW9gJsuvKH+ZkYPTKaLADg2sVa0lERVCfUitrLZAT8MP7xEsuMqIk
Gf86/Yh4KkS/r+m2SyvLpfgh4WcCZVm78QCfIJKj59T28XA8fxgTq+wqNiIXSYZl
1twhX/YQIi8FToVQ97vdyEvAszjD1hZK0ZFe1olkUXVZhVhguDfnRXThTizE7zH3
H5ZZBG4ZS1b7I1FjnE5vK9T7I2KRWMO4w+TVfSjQAYsAxdKWpV+j0mf401bvpnV1
Bob2zVXHrFNnDpDDFHjkq/l1wC/F7YPS+SrHuPuUWS/liHpau2mTSj+EheZ23wIb
gCr0swq12fkoUtOfhfB5oE+jNce3t19jzrFsuhyjpqgOWzVIVwnv1x1/h4025YU+
M18GOM31dYw2JaRTRMMq3FKYjbcb+U7/E4VBzKqEDDONgHrT7UT3TRJUf47v7ELz
PXvbcwJKJW8pfIVSel86bbBGZp9L/XojEMtcncxnodtvpuqivSvYkLccDsuw6kLD
N9QZzs2ubpbkVUn+wa5ydar6O73byfhB/TIvncCwGXv8MxZrHJ7cqCHiORsXiiyB
agL7wvc/NDQhC6ncINI2RhaH4gmuI+AszA51eplvDQngEPabxxG/oTh1m8YJiT1a
gRXKxGJntFSvQZU5+v69W4bUhGEoNgvcA22KqeRhO9iHZZdjVUjgbcbw4jnUCOkf
9CAL2rf/YL369hjiqdsDceSn6wLuHADRzLz2jYbug2TSUsXogPBLxa8T4X429K70
2OGjmg4F34pYV9hf6AGFfCmc7zcSRFuXZPmavn+8th6OByQ4nII34Yq4UjA1HFtX
tGSyY2Z2M+iIJ7mI6Ncc4mF/iyOj873jxAPa61+NYyd18/PT6Lsgr901Z/PVVBpu
wLJCeUY6JMMWnxWEoq4kIA4dq0BUiM7toBF8RnuRFGrVfewc0CvbADgywnq5g+PH
ncbgf08xMrUAmT+yZvJrsi0yjkKPUue0pJOYlaMRWCbgCYUSINslVsBc6o8gl5aa
e1ZO4Am0V7nRm0KzCZeB5au++m1GEpGDagcqff1Y4N7DErSw9bs39vfEzLb/ihIQ
TscxihLKb8hv5bkeV66y1Mh6vJqohBYughh8FX5BhNqrNrP09n5MnrgY/9Xhf3su
pMWmYFpjZBZHcCvAaZiuslCR3dNNy+w2D8DKHzizS1c8YJfpJTlmCYJ728JR4Aod
0+x6qN/+6KXcfvh2e8KsurVfLFdbzAXddJEbiwQ94LiVrlVKWEl0s60N6IFDooUc
ChnRIHeAc3v/HhqzfsHHS1/i+AYvjV0Z+Os1xezi+kLBl/ufw5PWLet/Y86qF23p
QZwEMqj6EcdDNGcmF/6dUSwB4RBOFw8W6yDXj0CjPzwj7lwseqz8jxHbe+jLkfM9
1Ob8yTlaEh1+UAJlnGnX+peHedZUgCdHSRqovpaViXDi22Yo+dhY41dCA4Oagove
uwhnfomXdP+Jr8Uk+XclZ/ZsJtDXMDNo9Q237jRhNFGz7aPCl68dVMqmbToVxxWe
qwBw0ZRZJm0X/kPYcz62J40l5xPrLGF+zqH5JTXVzdVMsJW3Ju4OYhWv1wdAHOpn
MC8qAIm4kBFkTVOMtV1WuGYEQvctYhm/+6jQ0WDA8B9yDbbNEVO+CHzT8BRN931T
CwbWA5wb/zagjA6Dy//xCgc2Wb6Btvk2ewg12ro/de0DN5ieQEWZZukq+HdhOC5B
YGs6HuwbKVsyx5vlqzwQXtsWPaphFdLdrcq5F3XNnj6WimX7QECAaNsaoxC7A+Ar
y2IlOZlItQDF4jKB/2suh+Itq3PxRQNfqNeOInvlN7pzFHjUuj/rEHT4brvq/TqP
eg1Z8mt0ib5KyS4k3HmYT6pTFhUNx8iNtYl4bKEYFWSclOy3f/P5j4MHXX69hvNZ
WQ92hZwi1dyBxHX2ys1LFxLKuFEaCTktUuMYLNblPQriaXXtTNXnhrtg3/FwY83n
sEm2RGPtEaM7CUv5kLQIbQ8MqFjfcMRlYviWThk/Z3nehCZhWVLKISi+wFfUmUdK
lFgy5qxk+OA0pt947zfb/eXdIajTwuntJRnJFObCWDK0fQp1dlEg6i3jsa3Pe07P
cNkEYPbKxI2D1KklGtfS8aW8yOJNDqDiPqXY6vnzrvIXzUezhLKDnSwh0XTEiR8r
V5/psKhwi1nZtJJP+7eRzxTjItjv7gOFEcIs8CkAoWPgdd1xkJ3ZYdabz86p0OXt
LSDS0CRZ1vwQUC7GOO4qkDIwPTp+YazBNtqXz1ktVLbPyp+Jl/JeUGildkAWgoM4
BdKIszhg0snYOk/DM6REWMxulpfoTHle8Ksal2VbA6qW+bYri8J3V3lU+41qFhh7
Cu04lc73WTlQO43JlmgnCb7advD7TYH04JF7UthFm/QWUyAdCUutvunUmn7JBP9B
oLdE59f6Wk3lChCevvIVNC+is2OB9zA43bKCrHocN8Nh/yIiJYPBtmBRHyPtFv0T
VhaoOyf418cbUW+fskZqBBP3VGEBeC+IrXzVi1+Yn/KFmvfuN849BsTaA/rf013Z
Jq84SVGhmDoheXjlyUc9qLEZjK+1XjR96e7KS510erJC9rV6vmNoIo4sJ3B7Ul10
SJ9qyRWqJXrAVU2zncs6AWxdRfpk3SpsZNXOjauhXZPAlAJjb2WLmjodDyb5xK/G
XTc3AAVCibmM91ZmdapqsxZhMvEmv+cAQ0wlEp0caJb8KxdsdHl252XhdZKfe+P3
hIRCtfaWGen7kshKea0jVBcecvj0yvXl5Qt2WJGQmhgmqVtTodtyfs3uSiZChfsW
0HV304a9fGcJUbWqHJU07ZfYYJrnqPvuu/xnOegz2XxGS39fLOogQp/PFN4PT24w
+cJQQh3mF/Ipdk+Wjq8p9IVRNGL/YKGmq7VCD2yDC/iT/mp7SVS1dxyreGpkvFIL
RrA0FUmwkSDYhwvw6EquJ1FmXN2FSms+duYNx6nl4lc4UswuEMcf8Ft6joFImbCm
Mmn23mniRmVMVkwBx1YVcr8BV4/btsQXHPK0DihecJtjm0v/h6CCt+/+PWKwVJUT
o48erS+SR9UDLrNZICDjmRx0YoOWBSkyYJq1Ges0YvnDyvayRNYuXNUI8epL7J6u
f4aQ8ffjES+0sHJjNUGfM/2hU0V76mmVq+Di4RzIccfBf8FETfQAOScoLrp3sR4D
Nvj9OadUM+hqvYu6nPfIXjYZaShMxamYBdeXl4ZrG8/KOhUUgt5K9NucKb98GSI3
8cS14093ItC4x5H32SuoQ2ffP1UHO2I2WOjv2nmy80pa53SuS4Mlh73NXp9F6Cpn
Ym5Kh+ze95SAXibdqwed3HeGlc12b0fiNwHcH/nGcNQeufNpmZV81IODVH0cyl+Z
lkqc9WQyhB/Iy6E4GfrSf1Fs15LY3xJHoBmg6kRIgNHLHTd0MTZml7moB8sTnuvk
0lB2Sd4N31B3oOnyc6vANJIleo/jQW699hEXHFV8pcZG0WXdrnhJDzUpsa8Jf6wI
T8OEE9xIcQdPJSgFxGNvgO0ZczmQbvSLVFXsDaPY+JSiRdmXp4Q7M+8TcJEo9ozx
ewA4iuMrbJQH7yFv6xfoFDemfEgLQuPS+Men4pqJDwbrJyYYxFaaing/366F1WRV
6gquzvAKApBpolUhx4V64AOicc9tu6AugQUszxpmZWZww3Do2ZaQsLk1Gth4LETt
ITywFkZrcPEDhwWc8H4t+g85Aq4kmRRbMGNl7R/lgLDOMfMsg6bT+fxQCw4/l3xL
6F6nj2LHH1S0pr+bOk6l6BnOaGVM/vsLdS3xULY0yeUWJ8To0WAIB/eG8HpB7dsu
xFsIRnBfaEFPZfntfXveiFLKvy+GeAsRXxSXF+0erBp4AgKfHwvtRBDIE/UfZXU7
2Sgrp0hQwkv7D7UENNoiKfZw75BIqGQba2Kf66kZWNA/fUVRmwThRIjms+kMFBfs
zekVrgJnDOl1Xz4HDdPliSzdKwx/nq1D1aUmOCah1bHfqzkGnct2mykfav2dpCq6
A3aMk6W52bkBJphzD4GjA/RndSP6WOUaL+BKG2wftOGtc2fz6ZBP7TeOqATO/Ra1
BAC/ofu6qvLXrFruOIXGtgA/isVpD4MHAORvcezxNNfhztVae+EAoZnYQU35Fzrj
sHLWlSkADY4i7yYu366YBuKqYF3GnbTGHJ/h/ik4bg+j5hAutl+GwZaGsHhJUf+A
4o5oRZRvLZV/pI2ZUdAfyJkxgYnz5qMnBr1XKobEjDpkVQigcwxr4eH7XjAbik2G
+/bfGeoBiRqGQNol0uf/r5R+eVNyXOHEs03/hBkx3xTFauhGea6IyWDlVldELJFE
U/LXwGTPexVzuyhu2wKg05jGY1VlrrmhzzVL+m60DjthW/NdDjgtFF4LKEjYvoAG
50VaC0/+a9eqfunf5j9Cxec2t7vCkhvgOvhk/6vfoMote9zzRDwmWV41In/ScVw6
R6DlabtXyMOZeAfclWicmc/asmfwFEtliisPhrIlU5dWQmYIUcAQjrf+f8ajVbOI
vn1y3h0PSbOw1Cpnu/+80Z4VGHYmEdRvizUcSdxn1hxyL59tgzzlvIBrxCdWTvZe
eD2tqEbhu1AsPCQq5ql6jZyZlO8azZlfbYb1PR++i2ZX2I5u5vysLC+dTrR5ntwj
YyjVipyiS25PiupCQs7qY0BJTZtCReaarLdDeTgn5e2hGB7wayAOOo9bp6HoNFJx
HAqW5OdRnc4f6/NReUl1OTlsJe9ixA2L6yVSTz22bWRp0gMTKlznxdNpuZbR/eSd
FHiN7Jfb6aWlFptQt4ajOYzFUmQSNF6e74F4U3eW0WQBKfjLPLf9i2dAUrFYNP6f
GQXRcZO9Q1ZAKQtYOjSiXT7RIG0AVWCNp21KeDHpaiZBr7p9QDuBsvJ6e5S5k/fJ
SMExM340EYE8pG+B0GfB/z931Rdv4SQkwpnPVzrfKxb1ACRUB6QPzCNLLa6+UHO4
Xf7cevk8azCvjHbwD5xdmDDIIcFrlNu/G9E56uVZzuFQaeCT4ri7VUPYLO3LsTew
sgfMPkGVnF46qbNwfgaw+Hn0cF5YamZEfSsvhaxK9xhZJZog01xUwlLSVHzqo0iI
pZtuOXgtgb2Po7+s25eipIQg8jcg1mXJJYig6nPHCvE8KWrOvTju58V5MRmd1Ksf
J9nYeFB8EC7xep9yPENaDl8O9dSSvJdYxczu8sQzZ6gH7L8WghNaalF/b7xrzv5L
KPLB7QZ6hMHVuCRVgECA/ptkfbFgNX00VwsIdZhODoBVsNdkjcF3azNdMFsF21y3
7GTM0hHd1/A3VtILxcKdU3m4fP1Nju0TjM0zEpT5O8nLbaYJkxKv4Gf5EI/kBWM9
pP8RPqxVvR+bW+Gkmz5olhGFnOlWdKwM5XHvap2E3DKY6rUpQf2XsMQ4C9S1ZId5
onMi7c1vh13Xyti4Q9JWC53wRJtNqgv5UsofkiDkjTr75isIkG70dOf3PFSoz37d
gRcvZ6tGGEDXWs1t3+IQyy7d4aEruZmLZFn+KJmpmjrO0d5nC68TildrK3voQ47y
ryvO3iRuoSE3UtdtdO9TZOAG3w8lTu5w2EW02hWt1KUHB4kjxjSZXdEMJXO8aAGV
xwdVteuhRAu+R/oyGzBDAA7wzxkQcrtRB/hgJpzaZ5Yvni+k96ylzPYgXs3fhD18
FjddI0d/ew86CvZNIfukn5Zu8GWJ867meWV5UUBOJUG5MNjbugjDwJ+WrD7hLj6x
brBXC0KReJJjpeN8Ooa+CHSsSaDCWLP8LSQnkIKC2lgoaljdRURox+qX1BXOO3rO
Lxm04lzJYauOWCBhCCpayJu6TWGw+aPKxidwzHVQCJB3GCE+z/0NgCz06Y/sbhVT
0KSWVkxXQOElTyLd0lxVNeqVTy13RPFbzTZ6lhvXqkMIpYz7h4BthQNw3tSW6oke
I89GJDaVCHsdHok3RC6ddMMGGEf0QRLH9+JfheSZCt8YWsi4ZuMYmzkuA64vYjb7
JwmSH8wjdSBH/rPyYF2GoNXViF6CHGOk3C0r0wCsNIVY5ZBwByTB1/MTqvshWpT1
HYL1LkbSm4DACPhnPBjPmA61fWcDt6S7kI7qfU1tSsiXHXmexaii9f4MqFwVqfbv
SxN4PPiseZeZ05xFiKxrKk/wfwX6U6vW+MeepVsCuQp5LS0tIM5oSQ/RaDvaUQTK
dxR8VXhkS1d21CcYdpId73n4LWdSRJRBn1RlVdLb1DSbvZ4geKuApLsu7gjmS8mi
EVwUmbfyXILe2RDZTeYMxp7LhIo4HAkG7mNIyD6hXCD40CiFMpkjlMV6S747LR3q
tjJqT2LBYLDTTTaZrLue8Xaj4lMqYM4sKwsw5NKwBl2B8X7bohHLS+fEq7AKOvap
rN3tJtJduGzRo6xV5QdNVphW89O1XRnR97qGiVcbGbraV2v3bXw51D+ioGup2LNJ
B7WYImmRs1zz6n1HwoPkpJff2uLWB1UV5gPIonuWoPaS6wZRLgStEW3+dWgIr5/X
Pk/RMNr5Kwu85i8xLDkG3FleO30dGUGxGptO97wyERjliOrk4AQgZ26Ds/0te5sI
TpLwgZRhKLdZNU8ooOIOE4TWc2DTqzBHja9JAVZtbA228LQiRefHMSNrrFtg2yXu
mPWhXGzO68pWhefIIa995z0r1WAVei+eJo6g3K+ssMI1dG+8z8fTg8ir+WxBAbXO
h8yv57GSBqXy3iHzIJiUg8Zlxq1bbBO1MGv8scEr0lPXYqyBNaqlz1C4xh2PyY+E
pJHFkfmA953kgkJ6Rt7kipzLsQTNNa5Iod7+oP//E3Ycx1hGkV/xENbTkl3vSvj+
xUUzWIwTKSkq8os7S9mc4NmQPph2dhXQVGgiM2xyBTMSg91zy+2b+GZ7SHN4/heN
iCc3+A1WDL+mekpZGMcz1xUOpug5vnTrbomfcKbBs0j07FSXmlUtZzWAN2IwcCUI
vjRwU2Dnf1yebWeu/ZIsOP0vSyQ4KTrp2JA+uzZ4I5VcT+tS3EEbo0G7o9Q++7wX
F9hB7l+42q8RKRZaSlpYRqdHNgoNinmDC6SV9HuFrbeQQVwa5vhPR9ZjduZDWnwf
GcDT0p26nWs97nAHortvXiMUizqRDReHOGr07icfYZx4bhH+jLnOySPMokmK5qyt
268h8qxLUzpXZYOoOIKplfxDZnbsABzDFaRIAUiVvxufaGH8IJ3doeE/5LE/3lj8
wxEk849hr+EBYM3Tb4zUX7jRu57dWiTS6BSiiKM+KcXDDfSwZPgC0KmEgklwI66W
rJE0vB47nDLePoG80ofHcG+9L7MhsRIhbOrJzWVEEbCFjjbpYj21oQlP8uzi0ekO
1KPtgccPTjPe8IH9v9vYW09+VzzDhwC8YvHEBvuI7j//LvrGG2fhGj34lCKGUUB/
pxiNp7CJQbxVQiXDPbkTs6uikoXutO81tuISLSQ0n0t7dfa3RdskEZidMVcEatPu
ElCY+q+4XAZJR90P2NgcF3vbNu1rojgPH+1H04sAuA+QwTJsjddn3BzCoSiIfEPO
Q8ruoWicwzoqnS387M8ZaUy+UkwlcwJTXevLD4bNxrXqjNauGKzA2sVu/Dcyn3bd
pa8f62jmrwJkBZmgoIG5TH9rbEu+jTpRQ/B2+4L8SuY/Vyolkfkxs56hdT/jC7RM
GcjRq8gSw91B5tORw6zTzjZntBahuCdGu9slFXTZXtTFbtTWlykPpCctQq8Vz/nX
Jfq3T6Ubnw9JTSKKMYE9T/56qMwGMDfklKe3+ToJ9I24/GLgOHfrnHbP1x/BJ9fM
mWzddCgrkxw2XAqBifahcu3mnEDKmeli6VT3BWLg4EqTmdgbW6SFXr1o59Su8GGy
9mJGPyZUSwvdScvazYDybcHLwDQpcZnXZ4UKTnM/q23P6w5gbG4iWqHjxSYVsTWD
o9fFUPB9YN6lX6ueR1VfxGWMbS+UA72xKgtokGgx+DxG/vV9cAZqr2kMRBsQkReV
wuAM7pCSjfgBRPQYzFNMZimTF+ppMf1OTP+SY7BqdmdObOJz4Uk1fMDgchlBbC4S
JNIkYQrvQ1dNnPvABW77FF/2WUr9n5WHdAzzHqUhy/6UfE/TPBHfoqJoFhRN9+tO
4W4SNbvb8Zz7ppBhyLMAtOPmuCgfClfAk2FN1OeY/HpJ/gquS/+zjQtW9Y3em9aI
DyTumBTjKRtKtg+pKss3PW5toz0Zas2AoQIi4Sk2w5oJhsMuIsOZro/PgpPdVqio
kyzVceX+gIM4z6Gpk0J02io1QkfBlnzqvq7ma0U7Qa4RCIIgNWz9UJ1U3qxbiJyh
cHqbKR/KQ2/BjVIaYNne2tXLnpnXRHRGss3b7lAgbKG5C/4XP/jLB8VVgCDC5jWK
ZUDTQXQkDLlvFpGw5sf/MUn5xwcu4ARyeNdTERbV9TWBt85Uhgi9g2gktqbf5OOO
5Hcrlm2RDxRLqw7cL9kIIcOUCRgpeJxIJ+Ri5F2RONW1gXpiDQlywhhpJFjQCIYJ
8xABSSGcZlV7ZIDjMlTLaj4Xtkj9AdK/dCayHiPEbVxVLgBQgIEYuaMoolkDigjp
6JZx8HWm7RoOjAxT7fu0hnN3O6A3RpIcD9Ax9Cinvwsi4JOcUfzdw0sTXlqC8u7w
cnmY1q+/WGFy9T1/rXA1eYeQSFg+i+lVVYdQxMycHKDGWtMe5ooRcJ08tDsorIah
FWfmflaQLP2QPy6UMwMHTQ+ixeqXCBbo7+KW9BAtRw2EoEloJlZFbE5IwI5/sx+t
9eTCjne8Z2CwqyULIouVeayQgAZ6c17x/LMxmK9YWc1OIwTOvVKHq/+e0i9z3F7Z
YunFilWCDjrmI8YUXDE91cvNiwr/9VVCJ2Ca7q9Now0k+afIkULa9UssM7LOOSuo
QxK1MydSVIct+HMb8C5c9IwCzgUdsO8AhPerJYstG3vOaAP8Kmfkds5A4v+1ASR7
7zYk0nNnHPnVu/UUdwH8CjnUB7ASh6wpBQniVFG5pCmsXSdHruWztd/kfl/ON7DZ
Oy8s4Ce5yBa5cAU7gi7+T2+nIfx2Irv8OCD1zgFwkhf7thGyObcBzqacdVbhnWbC
E1dJKT6CNzjeKc+Ldp46xYGABKfXjzFHpScSR7EiEbgfkPpgNDkWBL0xcEvV1inu
o725NrPUEi+9wYhpct7LRphR6gZHitan9hFUX9l+opRahxtob0rjMu03ZJdDnK1G
82b/zS0F3YRD5VBBRf2E9mLa5l63QjVlkdcksbFyMX8n3x7CLStJ9MIiNXf5MBIG
09WK1PjGnrmAtRlOiay1LnFFUnIFEyYrnsmkX2Wvzsuvpu5gU+aaCOu6Oidt4+N7
ch/15PzTCveO0Y0wE/Yw+GQzEhmN8nNTdZJdrHprwjeD7g21RLMczXxA5oxho6vL
YuaSKz1PLUBygSwXu+7Q1uOaaSopf6iMsFVS+BvClKlQW6c1WOvIm69xz3C2a8F/
5uypRMat7NoXTwxjnqhSd34VYlm2KZZt24pbQSOfM+DIp1JDDb3iHS/75NxDXCxl
uZJdEYx3EASFUx1OILjeg3i+NRrsslcelw729iKOyXfVy2apYmFon/5uoQLJtJGV
zqZeiA9IalDDxEpp/TeJlg1J+vKkEsFkSWv4QgurhbdGAeyXOg5WleBGdqESP825
8odVYk5bKxGC3Bxu64SXn2kmlqpao4ZpuHphkLy3pFxrUq2505OQWpn+wisvFi+K
CYf4ndBe1zWHyOR4EO7SAuOU5YAXOBQKU+QkTYasgLBZDVFsAOVC8DhFbXQmx7Av
hEs67stttBe7d556dPNaEtz/QsFGC8dJhFWrLSid/VtUXIXk3Kwv+pfc9OsBu/8v
o0EzmwP17t9EYNGRcy9NW1kcKDOpkgzArACt335hvrGt11TYfLjGkgKvHz04CewO
8bC+NodVXXglbnQlRUDoXZdrKfXCOtlbi6KdHTXbG0PGfm9q/1cyBb5K+xcNdF9f

`pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
gug/P4JSBXaJmq/mehcO3PX6hyzuF50wCxs+F20wXCS2huYsRc76F61YP+cMMag/
Vv1u9tMMj7mY9TDAGpZ72Aya6Tn8aqtQ2lYvLK5ekN9I0sb6MvnYaGS1JvlF2rDd
sox/R8P21jqdBNqYoEjZ4TPNg076du/0uWWTevtGqKk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5520)
NnKHaN6XGBReEbVuSP1klBhQfhgatGEyN4Tens3NNWjOmp4BED6BW8ek2RU5i2E0
4gzTNa4x4WZBzW2CYJpcsvLWFdpHn0tGY4oKKtQJF7E2KfCLxIGdPM62+1Ww0MGQ
5mqHyaQC99zNazkibgVG9Hf+q7E2u69QYom6AD0ura7abAlKJRfDoFgwVjO+2udz
xUB9AqUFgqqGlCXsZlYFQZvESrSxnlolRBb5tTVCdWIdvkw3la3up8tlQKsWudnp
LYs+99rlPJ/vSQ1/h12aRIMbL3z66Nulva4mFJoFxhrLM7T/ciblzJfGnL7Gwlq7
uhaGF6JtTVP4IB+FqwPlsWx1QhMqCZyQ+vX0HVIUSqdWEMjV268VCE2Y8jqqRzJB
cB2g3GKlOFUzTby59+nwUk57gq4rD9WIZ0rOL6R/h6dkBZ7fL7v+/aSHr8cIvrSK
xV5gSsllaAHGsuGWCf/ERHpqi2b15zeIoDQsxo1MZp/TnJRCyBJDx3fqOgNFdpz0
PUDqIcuUo7A/YTaZhNpGPyfq50jSPR+gGLG6NHnOkUx2MGC2Y9rDtsMh5zbcsHFL
wWsr21c4fz6fcs0X231xSUJZZrcSy41nWFreWl61KyJ6YTs31hezkRzrWp3uUs42
acdeGugYsSk0vdy6Zc3DtHKR5/5n57MZnjereb2sWuq8ntO+qQziYJSwJZbIpfPA
q+cZDtsc7q93yCMxzSflhKXkrFOAkZVtb7Aofio8iXd7M4ePzuzt8STzTjXrRgKf
o2OfxRF61jiSh0XuJ0dqljYGx34wWT3O8xSh0rm6YeReepyfYpXWpJXigKxvocdB
PWDqnRdapD/Y94CTq6uKgIv58//Gaf4Qvl0mjtd7E2KsicwIkXC/SuV1W/JMCiiR
7gi2YsedBqEyfGI4rXunPAJCwYZPk5Kvu0rrnYdmWvdzsuXpVA81tQeuj9B1vTms
Je53Xzvn3JZtl17I+h+OnJqqvDfoDRXatvb/KqkeMSZXbsUcdf8imQ6qqTw1Z18F
Wy6D1T/D4APTHs3gStSPh9gFqdRX2HIrUYWL95jBDoRFmZv8JQs0F8fovk0nNJ+L
mQlH8Fx4huhxvf3V8vPfubd8ihO/9f3347m/8/61uoGTyqZQEWsEQR4omL0VjGK4
6ATyZqeWFwuu/yEDEbBpNFfD9WmQKtg4YrPM7iCPe1FQT0H4otzEaHfVlM7C6H8y
cWVnBOD+hrGJDu29EjTM0Sk5Y7FLEFvZYJb71tww3Qzi3CYMnNwd+ufmKlKNXXHX
0ePBwJCEdXKdaPTX3YdFySOEGQDZwFcN7lQZ1tu5zVFJ5IxnZV848yJxCDbsovXs
40tYhEtf1dxnQMghl6c8EUwExWNgWvFSWXtuolmwZxyQzUGhCSepQWWsc1eY1UBx
2vGJWlnwrRt83TpGzYmVaDAkAPo9W6lpXUss4S+PETkNoE9bGKnVjgfWTWYMiAm9
cIi7YgD7bsG5M67fY7GJC0xd0bNmSEPIIip775qWzMrveXcBG4Ld9vzvqk7NyeYw
zgv2cJLMr2M3VTeaArM6WFpVT2MHjda2RFdXniWL+HI5y9pWn1OJTe+KDwPIQIWE
xpn2RbTiIgCwnhvtqRWYQFma33YxPxX5vOShU8LjQUsz/exQ6qgg8Ll/Q8bLsTps
Du7M0fUI1e+rpTyiTMvzE4TZ0uX1OyB4NUcNt/83b7D2cCGBPc6Tl83knxWha1uq
nCctPYkzFnLDuRJQbHyRiP1YoZZPMIAWb6hCIifNoKnShnpPcwZJAiKajvb3ONAk
MMvPm44zSX8jocPn+8kiCEWx4QRZ8YW2XmPxZShxda+3kstauwpHT2VhdATti6qJ
u0D43ce2ZabgMoQOeAxWSLb2uaufNk9kK7Y7zbJdH+YItK1LC0LF5JLRA2lWzKyK
Sp1Efymom7V6mPiFZcX6N9TfwzNTaBte4uglYYmTiSU5V05JkYqpZnzNGHaQGqj5
Bp5ymRWtNZia6lGrs1DZg3x671hHjPXvyAcrhnk28sTwwF+klHl9ljcmJEqGrMa7
8Nocz00H31pugxUcyPIdrstDKO1Xe01fxWx1ld6coQ3ayMtcmbF0hSCC1odWdrsf
cDcNZrgcZlzwPwTPEjOrki7V4DdT78tzA6WVPxOh/UkNkMTJdi27Qk/NgoVTMnuS
6jii5chUihs1jf/2d1TmoXFGpFHldFVpKQxgkXJFWBJh98AbQx4810XAOgd1hOQD
PFjvg67ny5gOu516Nr4q0fHXKrNeU9ZdD4gO3maM5rXDsH4oAe7lb5tueSZ32dkW
2sH8Sg9Y3AU2I3WbGnIJpbZCABx7g//VKhelkFqzI0dGLx+5N7SNEZABFvOSA9if
HRBUORCBl4zISma6mKIiAGMlqby2xlMrfih613ZTFdS3M5Er/aam3HpPIU1sl9G6
HaRN8CtjD/xkZ+5pEEGv/iQCeBppszVEOyiSJv6Bowj+IwwwZ8YcSYbFQBfrH4ip
59FtgfpSlX/DNRssg1pqSVxjr44TdHHpCeJU6KBUqfRtPln17kXWJh6M6ODihaLK
7QVhNzCvtijmdhLOPh+T0Rd/9Lb7l/KJHaK65PKjgZiTkR7e38gcsG2jhaHak1tn
NSx1a+OPeP26CEx8fLNKbYtJGHergUUwawbrKDdk6G7VDzauTD4ayE/bm7+Y0T77
QY1TKLyBC/hF/UITifRxmitmnVd2Q7VlzVx9TmepL+QW//wF8ZideBuhXHb/E3qM
KnKeBoUQb80dVxti5j8adaNKEFxwQ1dvAqB+VHoSTyhK6Z2gmgcRXr+PuLbuhLPU
Ui4GY1DJ+KKhf/QQopDfeWb0VWhEGjliyEb7G46hggRCOgn485G1zTEYMQD1xkRi
FW/ix+SyFqbogzLtzVC44nXF0nDHu3w2yTtpQEgZyH9bXLuW2SLtwe3xoVbOXQg4
cHSaI4Kvv/nqOBQrr4IklyGMUdNpZjO4ISxD+tE2xPM9jc89qPkWWSPkE15OPNY/
x0nZF/LFcXG4s27WjtCC3dxOB5tQ7MFBMGVXpNUhza1BYwc9CY57+ZciPdYFAFng
O7DQVvmFpKDwUn3XViekqiVt0ciHTsuKKNYwrN0x8eDYYL8qaMxQ16gcyIFXavn6
Nod0hrnpovx2of4CHTBGT0T629K9F9blOZvczWpiGRUNrR7Ov+xwcUPzq1v7A68t
COFu4iXD6Mkbk5aVvjDap3ATyNmSd6eATAR1EH2x5zEvanrfRqf53o7Ymz72PE2+
X7Lp9guWYyVffkj/rTfLFBAGtkgcu+m1iUFoNlpv+UnPbEkIAj/I9Mdr1xtuWmBM
CXruTgUF0gGx6eFBu2oXo7trchu7ZJgi1p4ct9TLW2Fz14LVGkDUa9x7kqelt9Mo
6k3gUEni+xiox74DJeGGxe+vj5Fe0NXxFWMBQuq4KGunm7yVIypRfPvNPlVVGS1B
4rmsdrSRhsDA0xtgzU3EO/VK4lsnuynfMu+x12+15VYhZDgitgtvpA8xeUdHCa9m
ttm6ScNUJ8R+GguR+6RcmxYO8Tl7cUzA3qNXMOtII2baBT+dTjdf0D2JQn34kURA
QI0I+Eg3ESnHDmkGWTe24JdKJTpvwC/D58swfGoiyrHKSxvqhV8pMzI+WHKpCbZB
5jKKhW+BxnHLmJUPKOAPKhP96spwC1Y1lks/r+o0/B0GRsI4ghzU9CMfjWihF+4Q
h+f81JMvNeoA1TLHkKyqoU92hugxAHu/ARNTuNLqA0hmJ/4D7Sz4FaNn5tm48IqW
xVFxw1nWy/xPsBtkI4GDOLVgY0BT7KulmL9KpSUUHiaCxNLq7JFu/bGDEF/3z6jX
7pYdO0Nc3xW/ledemJJ8OfGLVEyGh+RLNaSiaFvVcYHA7T8ySksB2J1kHiBzFMna
mD+DXSFiDOn6epfv52vJjn621PDRab7n3uZX2sS2XX59yvaBr1uHGmigrnuZik50
bbu5NESMRslRBqBcmu01sUm/znDWFn/pKWolw1HPRC7HLJ6KfsOSA3BmzSts4HV/
yO1kqC89bi6GLh/VIejHYTgtPpmjLeMcbHFO4VpEB9VJf3BOS7QJajKhzXXNS5gY
/gp9BrolkoQi1RXyixU/yDUug/t6B23fM1lXiBUxuphd96pIgihXLmWp+E8KUatb
IReK5fWXBTv3G0D8CTVedkHtrQKxWm8iM2TRPamZQ/8Nj+j7Ur2SlG/pWjjh+DoL
sJrKhcMJ2xEzgOiPiIN7q7RqbLNKQkUITYrE8um0CyryKYRHUGwmgybKhR5ZAlRl
MM9V4XcwoUvlXxSwVrYKas8gpsjoNyCsF/dtxv1ChTPysISSPLiklV6z1dnqdct6
CO/iqPrwuYvDuiGVFd8M7bTJLTb4CeXWXCXqtMQ+fIiA123kDR1n20+pSrttA2HQ
SrK+ZYIhM7pDHx5ivWmqArLcjzYwgtMZ/VbVsHu2vujmswgSTr5gfwPjODpCSqjc
4+lqr+pQ9pSNNibqMiIiJsvASoTI+rZ7k3DsCHlf3qXId77GqDGta7RpPPq+4fyZ
KfZ06af64iaY65sYxoiNGKoxLmUOxKJRasjOnAEYnBoh5shjbh4/cxyTduDxEVYM
BMagmBUPQBh1y/6OYy7oDHGaJEF204PkXniaWjoiQ14IBvLgIoJdHogK3VEmpW7l
2K+PpBkZs2qB4A62rQPjvZGyDk0mkHLLP8PmFKZHixiANeRVA+H4N2LzIlIHUeSz
ILEEGQiZuiVZXwfns2nqt3KMRNOGKmT/s2TbuIuaXzJaGyjzZPGWcY0S8rkX0SCx
KiWgw71SqV+7+gzSpc6t0bchX6vI0fpXUy8dlGsDu4vmbtwh4ZHZr1SPvOvDOzg2
nnHJfBj7khEb79ql+SaPxzG+wcnSlFAY/2tLoQWdXk7U8fRuL5Vw6YH/+/n1xm/y
7ADkRonp3XzH1nfGWEMytZT5MAEXvG5S2VRTpSfJ9UcTO6iJWMP6HtUyMP3HYw+g
Vm+sSXMtfJx+9lc0xMCSIl5qPodWi/uhQFXTMDYSrp6HFexE58o4MdionVG/EJ6x
W1HO5FblS7ZWjaiB4gWukcdRCfA/LDsWhVSkhd/7hS8GYmfrmyIhtFt+/3dIjcXf
hTyZkbX7nKQIjf8j6yGfInlj8zoCRSLsrGdBE3Rlb3Ym+KYMov6IqG2ZjKFrL2eL
WItMf8DL4NeDlWYnborInmQ01SYcctZ1knY1ouDHRj2bxzgJL3szLqV/6FIdYSE+
cddyHfD6QPdorcQaSWda8zFETf+kUBR5kyn97r3pFG955XzjF0X6Lr/0sR4zWDki
PFk+kJjje94MTQZ+kl7OjF2iChRcHb9hNYsOoGJrDs9Ml5/ZK62InxTMQwZ7fxKI
48Nn/clwFi7k0yFRTKx/lWXFLGdyUHtk/AGYMjb6suL7wLttY46VqafFdhiHiJ5O
2v29CKYz+lEUUSKfiLUoVitF4Ti4ocvXyALo+NgIrR9P23lBXNCrhmlhJiZlzDeP
igxyysGxO2oaz8zZ4F883O7vRMIrtxOyg1NRQfnwjZLeCexNsKU46eqQLj0ib1NT
cG1wFITa2VZu8d0Eafx6vSZuKaTNt83ovzBOaq2gLdeJsFbQHRhLlioDoeg080nQ
eNa5AamXlfGr8cxW2z3u5BJC/Lb7MedhEvlOWBksYrtpYGNRpNy/lPnWglWtBE18
18SHtEy+9IDYrmd+isDX0NFAr0n1M/WSrzk3XJigHF0/MqteT7dFbsl0xY0ycIbt
oqydXSQxK32Cm8u1v5/7/jW6tDly7ELruezFy/SlgofahvebfnbqNTOY96RO5/VN
aW93bKX4NAbPd0TIWq2+4NrR2GZkIA7pRj8SzBRYqTrHSau/i9FzyQqeXyzKhXGE
5b47nBKRweRT2eqxOqHMwlxpksgzxdYHhPx2Snz55VKnA5Kk9ykgH4QpvWLG/c3/
OnnOUoGgyzy+oMqCcsQd9JJQCNpIQBRdp+pIK1KbM+u5pbnKKKFSoGr5ccgxWSYF
gK31XfzDEMQ3NHKjMd4bx5w7U11aLEkvsTs0Hh6z40jaEv9KydRLE9H8Nh57KC85
VkXdeJ9XvVNzEsHGNba+w4Y/ep0Tfj81qbYmwWto2YVmwI49OfrYwa3ue97DJ4ai
UDSD5OIPlqUUCocosBbRw0UfAFKe68oxoz+QmYLwBkgB5jalHnnqLre9E6Yr+dnT
oTNVR+Jxdfom0zBs+xPqknfAZpXhQJBZDSwh/jO+hyvIIAIQZ2MkQT+rEee15Cw4
1pOy3s5zWlkfgnoz84BS1l6N3nwna4oL6HQp7xBZq7/mAri2xOOK5w4/bBTILbSl
jQWP6RBmC5aerI1YDDr2pNQ3kRE5Jq/616NWgl3JPhSiUVbGFX6JGEHkwts6ahCk
aC0NvyEZkWH1macJ6wVO9qctBuJnTaYyDb0jAsmVYsWZwvuYPnABhK0OkUS2T+Wb
Ldrz68Aupt34BZ/ji3Zl1/jI1ZZk8n0SVfE237aX4eXQqAWqxlNcEAonwJvbtx02
WpHS8NI/xekP2qIp0q7kTFl1AGiDXVZaZPMBaHdKkBeWB5wv+0egb2bRJdswDMyy
oIoWXUvn5si9v7QCnV/lIYi/yJIdF1nu832f/VTqNhy2LZVlvEp50wpugFj+6YSv
Q/PqraysR97znSCaenWjjHGd+kw7rbfZc8hxwkpYh4hNpignH+Diq3Zvbi/cO2Lx
n+42a+7s+1MdRvEDnzMOQmnw347d4OfTJCgWUoCeBP+/NTIltikULIrEekIfZUZZ
VzFSKgtObdOOtdNwB8z1WKrqwAY2s5bgrdXJBJG7w2aLwXjZRVkO9ukk6KON5Z2I
pjYU7TiB9u4dh19EaahvGT24bffqfOwV5aq6YwEm9K+Yfr3XOYoUx8USPDBJpBjb
c5wSebeU+bvce1xLs5lNoslqmGfdHF9UrB4qJuXuEycHOwA7HKyUBVcWPbDysfbc
VjQNoHmpCZKtuMBLpur83j0XajGuXPJUT1RqYszyMYmcXRx5jzh33mJkSpFwXQRi
q8LmQD8IrOxl9lFdP74qnIC91s24xfIlwn9srNvAeSEHsMd9aYB/u0FbRB+sPrAu
mdsIGv8Bltn0EsGTuTx/m50MOjKXp7HWY/CYHC69ptFSOBk8gR/26v/7zEI4WYcB
1Jw0TJuhfqoeOZjardp4FWs47RY+HT+WOW9Pofy6LpyaOAHlaa95pDKDSMmfn5Bk
5AkB2hcqKX8lwTqnFdRCXd9nagiMTdKvU9MArpMPBO3ufnTUlYZtROUHQqas05R1
N4Al/SmQvLm5gkoBoLFv6ggbY+3KrgkvM7t568WAcSKpMofDDi2gQOLFvsTKu9ok
`pragma protect end_protected

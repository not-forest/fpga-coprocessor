// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
SPq3Sg1lFttC16ZSSLGrc9kZoTWW3Rk7d/g0tjSVsbkxthfkE1A6pzHAxFO5zOII
3yhDBLaChXVrQzIOJCTTJNqB57ELLxf33URcXUlMWdTfU7HBnpl82sFeiJJP64An
8ObGqB14baV3Y9EDkIoYuYbZy9e3imvxfmdNZDe6+uM=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 5440 )
`pragma protect data_block
MVns1UXtmp3iDutaUN18RwdvLHNZTBAhoojQ0nrNmUiNCxGvXxItYT6v3ZoqrdyQ
WU/Y4b3JzgY30rc+CQddHW9qm/uxl4kN286rUbIzFOvK1H68sBCu5rq6/VzrflAM
LeSQRMjd1HbSiWazjhTys76QJ5DQFvkypaoL6Q0ewZZbm7WdhW1I+MRuUCyUrTwM
De0DQzr0mOw37t92n8cHgxNeVmT6CS17dPZIuRsDxOjELDb8hg3Nfy9wy6NCRuxz
z/ofV1vHr8+MnhJRIhr1/sVnqKDVNMnlITAo1NYfNqH59p9MD9KhSZXh8duI/rkK
PGnkAiznxGwuVxEQgFtybhBPB8zOtIjedxkG2sNdZ9nkQTx8MHPVFRq0vSPDipy5
2Xd0yzIgXVLflzJA5x6ZLvBYSrO8O+fn5BjQkygSKoYyRxwqwnRzOKTRAxtklyJ5
Usjfy68Cb5f8wiwa511wfQcCblLyCs02/Pj7IrUBWq3tSZG71y15lwHvXb8UjO7T
SCbcrlIF4QGZ29jkjEZmCJ+FVymTjKGH3eBZ/MbgzBUN24+QEMlw8Kf0G4YFZvec
2ahVfbU4qZMYQi6+4FtUoc3rZGf0u+jftdEKEq8EAVi2JnVErNZyaDd3RyiPT1jb
0hKulA750/3ZKJ/SJZAr5vx9XQ5BL04Al/HBXToG1MHjD1nFZyQlmKLbgBvqewEd
0+81HgbMZqBhAE8tC4UCSWEUgYycgcgjJFHQ45/DrJLrmwliztgB3GHpMQkO9q8s
D6M5tq8rflPkbNDBU4THsbhi6n/bLT8wggViOE3FzHqAqvFrWewr9q5mH5g8RxkN
EbEjJRJCvYUVEkEiK8efiXswZLmAV6Tkvt0gTJ/RcobHixjwj3PssDiSCV5Xk5ID
dRfYhwVIFpjH4w+4qEo9ZzRjpW2nkF2QY5dCEpLlu3VkK+usjrqagDS0p1fqtOoa
2laKfWZzMY9u6W8CV+AAOPk3EXJnd7oU9uqZezH+FChJ+Sv4RzlOvsQFJ8AQCWd0
ZxWBOHH85x/k2XMzXtsFENhpAmBcgMx/Thxq+Ui//pQjHIYr64y0TBDuf+zYZegc
ysCzoasbH2XtgeU5eRdulsxGkjgxFQ9VpvAErsQq1v4ESviQAm/1gHqdf7XQsc5p
BiuV/+jmwmgcBGP5wGyFAASbblMA3FIZfRHmrf/2viFae6qZrt40IxvHXwKSNPE2
qMGb0HL1WNbriBPF0REct2GNsY4DnzjCGxwbH064jdWGXY8S/n3/aeq5ko/8ocZW
IRH8v+r+KXvf6AsFNnaSIvnaVPlnBitSRjX3N0q0Sj+wQL9pZs4Ktwr1yiGCzDXP
Qou4bTGw/i8jgv/MI3+eVp87pw6fV9h/2RNma7wvdbTxrr17pOHQ3DkgTt0t7bkK
IQKQwVFV0ZmGnVjAwp5vAmd9T/pIlZfEGOcTUyET3yh9T+YHLeChj+xsm6xc7izn
zAonzi0P1uvpQAjfiFZvc2wWcx8orKvj8e2Lay1+RJO6E7OOe2gq/F/yr2/pSlai
dPwIMuUh84EgqzUGFDhfVWa9exhXDn4LbRgfoMVyozsgmbH8tg3+X0qTHLDMjWef
qofn5oRUYgt5Ec+NSIlwm9OOaIUU4Pa6pLGizRiyg4PVGbE1K35bQPKkoHBUV9Hq
UEZ7eHID24ODL9v/QvumZxtIleZ7OA9m6pQrT7kWixuHQvntK51TcU7RWrAUuOzY
LkkKUK7e7J1H5H4Jd6VbKODKmGaHaQzMyqDM+BJyd6ueXtyRhsJY60iW6UoOOc7/
35q3u4KXtKY3wzo3mGCnUqhZl9aLQebnB92eP8CFHVG02Dh1JczC0Ago3ic4/fIC
qb7hZMOuC1l+w3P+kmF3aTQM4q9XwMbygIHDeaa3IapH7drapVTgb1sksjgXHF09
AnL2GmSpFT1eALjKA5QLGBa1HofGYGnW+EN8ITTgaURr7lvddY4HUB2c/gwhCNvr
4KcLOrsLmGozpMrolHnermvfro9C2bguVs3qWORX93KVBxXUdOre6iDomsdw79fQ
UE7DgWgjH/1sv3ISouAzo2ge8DDYKKfPjuuu8DO7TTHCFwH/nytKA9Kgpku0WIde
VPG00pqH7Bp8GRmhIeKOwT0ue5w3lAKupzK7uf7L9HlUKjlV6GOxucT22yBhk6c9
8drsY/Eh5rmnP5KBmOE4nK96sVPSu6/EFyiWOz8L1fNIIoJarG8o0GWoZYopNU3b
z0O8qSL+OnnzK+gIovHDyKTn8WmkAzoxYj14yA/AxrtDPjJFdiPs/eIcJRRPgqcI
dVMJHf00zAYqdfef4yvQQNlk3ReFh6wZKViWiSqf0f85GIzf27EXcV0h95eTjgue
uNUt8NurEyEpWUv6Rt6Ir7wOsAZ0ucyhjlZOBBYaiuzhl4SdAJZShKq2RkjzFvqr
cYLf0KZHpUmADeb82cVI2yflvBrhW2U+Dpj9kRvdOdtZSuJwbNBMEK9VfeRl8c6U
FMa/avVhxJ1+XVCQGTh6LSCGflDYrabe64taUKCmv/QnVibUtjj7dZ8aOJECQS72
whFSQu0i7m1nVTJTcCTc/qwoCPijHddvaOUphIxga7tXzMSK7jHDgBZdAjUNqMAj
PpakNDVDc6m9aKGa1mro3xzJwLEa3uM2y0khnKcmQD6GENCjK3L2IjyNgYQoxbSy
Z6jI2HFEC/3eOF2NZ8f7o7QRBPqg7OYRN6BhhU3i+jkMOTgCRNtK0knoO053Hb+/
dGkKLPKBkekGz/6EPH0yN8F2b2PkvplcEnzRAxEMpvwF+twzsZOlHJhc5HvcTG2a
F3WeK5/w19qD3+Y38iwJPlVRd1BwWtnnsSZygwHaI1C+dfCoeKh4RFXP3TlQr5G0
BBPDKpPyETdA869x3vJq0ZZIQpKHQVtACBCxiwC7bPRZvEHmPCaKP6DLVvEF+NXs
x4V0S60WK4xM+f7+2k3eyETM5EKK+VDFNOqNeasJvu0y3x1xLt2x1kuejeph58Ss
ihZNnEuB3lbX5pdykMUU/G7MZtxCkQIaJlagccvXn/CznPYP65g++KzqUnjbpoX2
gXee9qlOrxF54gw23nCGQg5ZgbHA8xYXtNu/BzHRPeyJWiHNdZbPbneLRpqfGXFI
RLudh56xL8Aals/9lsLGq4eFuA/Z7nGfrDjpHAsDI2YAkUKBZ3wC03Nhh+MZNmRg
mpiyo2XlEHHoTcwkOe1w1jD2oF0XMRmczs5j4+4vNiBVzmrAqPALGnBF4YqOEa2I
NfCMA6FBH+XR3B9UzuyYRw40krcdmBVn8P4LniIh3oxmrdrm6u7Dtyeoq6MpYtCM
2BA4lpucp5cVYyKbjL+GniXOU17vjn4LXuE16CCuXRTwcuiPNqL2pPk7KkW9cG41
adqAXSRLyLziLItvNHxPzcsNeNsJok6w6E5oQk+cBYBbwdOdfwacTv/oQSjSW9bv
lhqCzANTKFZPBMouJGjgdADTpJhatm9XgsVVf3lFOD/1yXyXqsTUOdAAALjOcwfD
X08nGuFnKy2NoUdvCjK0cik78ztLgH/h+kozS9GPM/M0Kee1D1/n5x7mF4w72GsB
qD4LQqwgmjoFyp+/yujK55Yal3KTH9a0oJzR7WyOX7xKAs/OUPQbQ7HqZBc0F0Ut
flOhDL0bhMJvna6Kg0YLwBoRTu7Km/C5iPxhSXN0TesWuL1TVWgfmdclK9nTsBDu
viAJIo/EEWVnVRHUGQptz1qZIy0Cu8OwD4tydl9q2J26utj/vBbSMr0Sdbg6MacB
LaiIfTK3E2cgSNOjpudVZYE+hnCMVWCLS8KisOHRCVm4i9nwsjXQ8jxq6TeOuNY2
iU/cZqBsDfKXcEoTSPFYo68jxXOzThwZLagPXssfMc1qJJsxSY3/ZjZx/ub/tB9D
C13muv5EXMxliiPGYlrtgGi4d0a0cwjurFRmCugrXiIc1VbQxQjxFcGCJ5pT5YVN
nIxbAo1dLJtebYDBqD9fHmyHpKoygDmUe9jCSZ9uZVFv8AmzkOSbdTMe0T3coNX5
jXGNnyh8kXmoOvbBe8qyHxmNR8Q/RItVnfcn6oCxfmNkoBXO1tc5yf9IFrb0R/UC
wyGID2wfUG2u3l/KxOj8vAorlPe4emYi1924choS0xq1aLfjh13eDUOrMLNOC7rG
2gWKctSQyOtGbmehZoIrsniRNA4BZIGoFiKxgDPYfdSPkrUIH3yrHHOu9muabx2k
KW4hMiajS69F8ga1NXNO7hMjjCirYXjnAvcrzL9DvYXDz5gO+/dXzO/RdWgXWUu8
lygjZWhJMg4bHmT7WIyvE3tu1r0jKJ8amz/U6M+ZMSRsMgPWYq/w1obciIm+oqML
Tu/P7/xGAWWxgeASWdWb+8SNhFMKCuTQc5FvAmXZRGIQ8qV2LsXghDLouriwm0gM
RAkQAReSsTHvC+up+rlkALQIr+q/INfuFt0NwROaH7JcWGQxCTxYMRwAPN6Dwbez
krEUYJFxegtWzcIcxURWE6ep+RrRD3LSFlwLJrQgnzYwh1VdcjSsaHn2PYqjetXn
PaII7qBEv2p5ku260NK21jJTsTrmS44URKGp6HUXBoeIlTNsE/YjSCsgiulEyNhk
cQ+V7JLSgS9bLT/G4bo5xQnnw1kF3zMu5em4RYms9dvL4/V8VmeyVEaaSrxEnoUG
syByGcPQfAYlch4719iZiFnUmp2QGjUs//JKlebEICv8AuXX6wDljKd1RBmF9WYv
2Fz3HrYpslx0Nax7J0OPYKso4ia4PrcnvmVtPC4azyIO+3VG/AP4lt9klyFhBjKt
m3TdolI+rYQqwTFfsMQdM14cGmJT1KnfpOrfSK0WOhwa0HclPF1GdoxP94Vq4tJQ
4ZrvmF1aiJrCB7H/17vaZwctaU/Go5awWUwvxe92ZGrKYtMldCKfGL6w0sl2P99G
rkgxlWILS/XTBXbAVJMsPvr0Yz5cCyYf7vjs0O0j+AA1Iv+4ZlJ9M71hxOZzxu4h
+UYp1dtwbkwNURyGmxLTPnjoOqNp1j/DHPcK4Vv/OG6KJB5moF++XyD/4mITjskV
2y2xdOwgIHuAezKJNDzlMksRUmJG9MNY1AvpN4NNdBkJUubnj2XxsAMJUEVXvQNL
2/7OTUDQX2yyLsjdA2PeEWR5VF2eZdfYZ3TAOujd80Y7jdJsgA3v+OoieP+ZSKyD
cHmDQZ4I8ZbijxDq0pjzDLMrob3ko4J8Gx6PHE2pdJK1BmX/BkC2U/diTrZrSa8B
SGZtHOrDU9lqu1MsPxMpqGZLW8QsDh/jcxbH6CgThTsCTwNU2RrPhaiIsXuOmI+7
hpsfyh6wh2YHFiYz06SYcYV+RBY4qknozJLY20a14NwLIi7ElqIloqL9PiUEssW4
cp2epl7wjKDeTYzLBGH7vsur4XMfnat+38LVzK/ozJqOrd41eK/Q6IteEDssFA2y
N76uK2w1rA7K6iUM1E09LctTFcbfF30OizmKia6Hj7+YW+zTL9jtu+2QmmdzOftv
u910PfWb+bS3UvH8SNI7di/Qkq1Fqe0YlaXVBUEpaTd029GNSVtXa3fqUTpFlhGM
pM/ABopOSmZNOfayXmBQg1qeHsAbG+bO1LIUHYknJH3KbP7ZQwXyzWuWKB5smhk1
GFJC7W0SPKK0jP9dwn1HnN5gQqUnURmGD8wUIboG48ruCLPo7dCibqri774sP+fr
LYbwvcRz5CFOH3DhSo0CFtxh37HDNJOjNBvN8xt1d/trvT6GXc6YcUBrPUmfdzZc
x6ww0pcMxfZ8bSg1DcmsvbNwb+Thg9VxDEnt0KbHbIuaU6+VNM5Up71hKmumrnHZ
L5rpv/P1c/Fjir2OK5E5jRtdcoqaYzdcSABQsm7dPp0qfAUgInQoBA1s/wwYk8AB
iUKNWaocNWZNzjRYUxH4I4bfH/SLwzLLjHxvl4W0U18Qgg/SMrp/ndyYZcPTKHm/
fQdTn3iNyRwHLVgRiTV+zCfQcamZgSs3xB9Y82VAnmVx4LasTYNqz9d1BcRbNr5s
TBodyq965igCz6ZMjVx8CA9YHPGtV1fiskG93WbFRHIfqU2Cw1RBpWYOU1w/KxWp
iuGP2J2JIqiPe6BPaFNfH11O+6WwqbMeDpeGBmTksEd9BKzBrNhRrxyq4PudAzCe
TSr3KkJUrXTFBnlxAolFAxHpLtg1SOVJPb2m9qVyKS/WB4YsJwB6RTDribA6R1hG
/Wu+51aLI+MSdaJ21ebV0Qd2qTaMX7iYRRHRAP/tLsJ7WAp15gjQGzqVT3J9s1Xz
J1uLGTDZbl/Egdie1PybvE5+ktyWQq+bPFLlaqFERciHU7JSCW63AeAa3JepBtCu
+XZ1VVMSItA0l33dalwRJ38m4suZa2BUjTSWZrCyDWq2iqTmWbekGhKYeKCi43Re
CP+ycwM0hznqbswIjwcoiG7t0cU8wCUg/2Bb9CXj+Wf0rLfEe7kn53w2H3Ev5c7F
mTdA0IgOe3lHGRcQBMC/cFSivtO0ekCoC5SHluAV3B55dQHZYhev6bEcMQC5Uz4z
Q5/rWHI1CM+jg0u5LEYsDKAKqm/w7EeG0L1StppyPXVBT66PUUlVlZ5wN8n1Cptg
DQfNUSXllmj83FlrhcO+FkxmF68zrs9er1579GYbYuAof7QA6kdo2uuw/ioQQALK
4CzwChPHFWVkNtH5lYP0u4npoyanzrKpRWT2otcS/3poAl3eSrYfZgjckXlwThBs
uyHjR8Ikcf8EVeJsL5o56WDvzVHWHbeyay4+0Ztwf7wiugpDhlVHuy6DaAyHWYze
uiTqs8S3HMxIqg6qVgDBoCxiuD2x0tIKDMgLjzrhrBuSRutU3egag1gMMm04lrAo
iv8P1nsjcyvbHO6tU1JyceFigXTGBlf1Ji70LUTU9gMjAPj3ANsxrClsw3kfz4g3
vF2VcxBNjS9NmU+pkYZ/7OPb1McuX/I5R4RYk8NNEsexFQFuwQsRZR538zKUEF83
sggiK4zcuN6YOEF/FUI+koQmO3sJjERXX2obCzgE1t9RP0lGBOeTey7cvFIePbb2
HQw8xkWNr9LIeHFkCDc4Br0DjuzV9sqjUFRLs1cxeUf4h0uR9yatc7UeP1yTsMiE
VjXA3TXQ2Vx7Y3uR16jikDAfZzx+PBYEW3UIghXstI2UNarfcjF33M8lV9DnSUwQ
MB8E4Rb9hybKKG99SnSYit711xur/mkXj0BP8f5SwXmiis+h8C1c5T1jY0e3LUFs
MpShR1iGvtBnu5VrUlaIOg==

`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
oowk0D0MwpTXN86TBgeOt8hLi5H8akuARw4U5ATkNjLPDD9pn9jITZQ1yttkXNmh
jRjFwwlEG0pCsPy81WpdRHjv0S9VGPKJF3vGaakf4aiPe/DCOYPB+1MNRNUFkpFF
ZU04ks8OKhFq1UjJ+s7U+zDz2wBtj0O7xc9PEtpK9LgBbw3C6lirlEgXtTlW+q3t
rXJzozfKBR+MN08PGMetrw9ZkXQhAzRNpFiRzCnyRjpUQyqKkhE4eugfgJHaunny
WYHsIrMLzk/A/UKzVtxQJPqlq6MzsQffRBvTpKFE81T18Kn08sQ30+4++GH1qwrL
oBnxF9SVy4iS7/VT96nXZA==
//pragma protect end_key_block
//pragma protect digest_block
GashtlqLH3TX6i5YqApjux5tNQg=
//pragma protect end_digest_block
//pragma protect data_block
1Q21DhHEpPBLfdFM4zc105smTHJMjqhlhjPXMvqrAZcVEyTejMpsjLipC0aBsJ7l
Ti2Kd7VBR497lxvqELRAbnXh0hI/3UvNIWXQgPWlnURjBJ/9NIH8cUHBFOhrcfz3
vQqSSYjbpqoqtehvh8S9MxoaOf4Ukw0oNqOlXh/nO4yZHKGIc0etXIL/o2V5RJFc
BTEjuAjNQFyUG76fvPdM+GvkpplETdfWiUkUlonKElECap53nQtTbjI4EUCsf0ZM
pazB0CqRu7H409us3ShMY61NkSoCvjTD+KZ14mJlWc6cog4XxwjYfH+DO950C2Yc
1ol+H9ihL4Ki7mHf5iN3TzNYhqKIEPRtKrttD542PVJOjyquAwXSEtKSB5M2aqIj
Hos20xiIzIk5IBMF9IOzn+xRMlaquBlwPOktRj4s3EHXDopV8xM3ywXFc2bnllyH
2xODewPD1ABllBlfGH4jSkmLwhDe2ZkSEEdDXDgN5n8tHesXUY9Zd12XYkl3gPij
yvYGE60zRhdOwE9JzH6kMDjZHA4nvUQzq1BSXEZYeHCVGf8lBZijty9EkSTshp/m
vO2HF4ASRzoPdAlFbz3S7xmMSdU1oUekiMXWTHQcDU0SSvaVsADdkOo5P87dql3F
AvKmq8lW+YumPujFMk8g3Uf8/bHvLs0n5IBZEmVeBkLKsq8EKsR774C/ykRR9F3n
uWwyH7T+r0VB/LE4EwK79fnqv/vgF6YS3kLwoe6xAvSJMaVwIE1mGmsQbDIdUeN/
Wt3SqN3K0wbIKcPcZaCSd/3/A1CUweh5KwELCkfv+uIL22vLUqK5GfUa7Mt4UMTY
fxBCs1jRfXjwRDrz7StAtlgpVRW+SkYEgLtLzgRWB6BerVFI1FHJBpZ/vE/leQSR
C5PXFr9OQODFQfDzMSf+O+P0tb2ftfQxLzVbO5HB2kIXiOYwEidDGM5RllZQrrjR
WEQZI1UE9Nm5H15BXi/t1twkoopYvubTW4992I3cD/kswO2ZQFgxQrFqZmC4FYgj
hliDm4GpCyYVAOHcVw5kimoejX0sCvvCMXh0bRfkeL68tSgZQDhGvAiD4Ga2CsT5
HW71eIY6bKi0ugTrwNnOwFVjCLfIfyUO0k4zXilHdsI6Sos7HvqIuKmY7pHvRLOy
g3C+th4plppjv1WXHDAUD7Rl90zd1kc43luCPX8MFo/WiNxHYL5+DhB5lbDonjGY
Z36ZULirQP6tHmete9CA6W3Z6SOGiRzZ3Wgel6PiLmShcKsga36Xo/1W0I8N2xxi
8xaVfTVuGbS7rQFGZoLE9kvbU5v3+Id/h6OIqtrZZsEedvHiK/iuCNxuG4bLStYA
ClHxSCVHN8OJQpIPn3P2XkFG3H9SwWAD0iKG9XHptOtuI6QjGHMZhQg9N0ylZGxn
eAYUwAuNzln0dUdMoV1SB28hIGXlSeag7zdTxqPkSpp9t5PTLJTHLspSYJQD9Cgf
grADed9GI/4zd3Y2czxgcPf/GEXaNigcuDI/7ol78OIh9gWH3jpdgnzthgGDhEsT
vJCRvY38zpyQu6MwsAZ2xp69D60ot9UaFlfnfhR6++v3omVAIN4+OQNCyyoNHasR
skfNZtiuMboUFA7vPMMOSc4re5CKJyb0bM3U1uMX+LcjOvNkojdWRTRQh9JZMQ+c
5/6oqiRkLoJcQZuKZkrk2301WoLupPkICUB4GXe7VeMBcf5SwYrNyiiDl1L3cgfC
eQps2MxWHRbyNwZi06V+ggpIw/FAxpa1Qq86svCvyZGPEXGddHZCCE3Wj/grBSh2
Nu3pmRBvOwrqWC8l0r6BpNG0Lk3cZTGJCumxBXnoZz4kLFAj03xclboSTODFvXdh
9+BzOI0mZJZyv07kVdVcBRGQYHSg+t50U6b4tZjec73eH0+zWJ/FpdAnMRQSp4zB
FBcB6mJun/ZPRDFhNKWZS97xyxFaP2lvxuX2ephZWv6G0TLjsKe3rZbg5JoaQ819
TpIXw2b+Y6W/Zhw4Gaq1n/xVxYh7rUAYR2I+KBKrNFMe07PsCNXl5guhcIcspo+H
zoTT3jpirFcELpqiLtQNyVWDn+x+ut/SQ5lUy310yG6RD/RMHins4gSjsFDFF/hH
KtH7CWsd/HOKdf02wtmy6sG7eXwz2ol6lVo8abSIFlHRR/LbVyEMqZD6SAylakk0
jAs9AdCkT7GfHR7ItB+xvuBEF10EGG/iA+z7CNRGY1fAUqJeTVgPCeTDWonPcQPY
9yD2+c2tR0huZPSxtB3dEPn23kEOq15o0fdLec/N3O26PrhC1cw6xMAJrAW0qMtp
hJicCBrCD7PLuonl+BN+FAQUjFUWQIW08xKUjgg0AC6nYeKKyFexUncSy7dXoGY7
TrX7UIQYy2TA7PqheTsHps1Y2fAWCOukdAKqxJx7gHh0d9eXJG5GFR2awQwGw1Be
ijxLmir9Zy4zSRqWzcRA42vijp/h/lgqrTyQEEXy6BJWCIyYvrBHrXXWXxqEKKKk
Dwnynn1GM2Hedk29Hsc2FwRMeXtw9LQ10Sb7MMIhmt68meVnzma9GBNfsTNYH1n3
IyjepOX7H81qLjgkPsw+8mkeGtVjbSW6HbpQs/vOmDauIq9CEzR0HnkgVRtXVLyg
0L6XjfFS/yQOVzYlGoBNl6SMVJiGkFm1gvMqin06l7jYMwg0z8mpTvDeq3e+TaFH
kIer3QD4LcrcGsimv23WyhsoZ8a1PAekYUrSVs5Qedy6QSGoTeZl0Vh0G7MKHyL2
cwMusgnzlDoLdGbt4hGfhrK+U0lrf9oSeI3Us+W1t95ItMvw1enIxteK0Z41ra17
auDnN8gKJsuXG+rao4C8bwvOgGIGwbMQsEQfOkxTF7ZxD4j8ZAp4xSdIUvPovunc
f0lNJYXahltJ+PDDTaKuIjhSBn3U0YQVDRz5s4sEPd/6cbmD4m86chVf0hUxVMHQ
6y3rNCoUcmOAleU3+wzh2H7btx3k18m1jfbAJJbP0+UIIAUO2rlbfCrlPJ5kbcXY
m+pdIwiUgOXUpRFlzBtv6Qwd6h0XGHZeczppZhdCOPjjkNE1A9x4qxy8X6oHfZd+
9DdWYXN1NlMDIp6QE2QM37H5wVNL6/5jcbXGjpSQDOMx/aYyoGStmcqIeVjQwFEz
mp/6TMSMOnF5yE/v695TY/sdvnJIsYfFa4uCuM+2wG81nGjVxpSpBBw+k1U2mWPh
jNIxkKjpTDdcgpNxbxPU+sWj5PqYFwPYLp56/PPNHRk68/RJLZiQluMcEhmHPFLg
q95W/17/kRBlGHqqs4ByszM5EuDDu+/eiIufwA/5inwPr1RIukUC61MduXgw8kg5
QEN6vclXAHaYJkLvrga3gy24++Ai8eUsOZj1FCg6Sty2ELXRMaqiU2Jr1nv3qgaq
zfiw073RTxC6ADx5XQ4CHcPjfW3M9WwlzFm45LwiPEbNczyGK3TLe2DoD9fPgd2z
Xi7MeNzLV8ObeACKv2y/YZDetJt0AyWfSl+gMmrm90iGmtmnrxoCtgiBNUkCqKrz
EbkQk43rd060jQtzaumrvVQGa4IChrojJeITNW1z0M8KpKxiGW5PMPocQEzLosZq
g/zIFF43hFGXzwwR3vpBWsFX37QFr98Bp/ZVu5eSy+dxd7Xdk7lYvZUaG7HexG/4
VuyfBzmPhatgEgX2r8wQx/2W2oQ24MbjtQITuQJIKJJ+ywtZkceYlo2nTICvVxo/
shyszry9aJXVRDhDsHJ8LcVwyeDTwxzrZHyf+GjbAMrpZYC1MA8o4PvnPhh+oWmf
UIgCc+SgKWLo5aHD6jnsBolNu/YmXd5FDCFK7z3zuK53M6sATsHFA0BnLHfd3KpV
UfnKkS4c2eH/ABKBXDdcgqBc8Q4t488O2j4LpXEZYiqWcFUZRqcZsM/Hrg4u4Ty0
M47FBrtnVcB7bpbOL+wStjhxsxptUUiZjV9LdU2bTcT5PQTLmKqjSP0TMp3iso1C
/Tib7btFWqWp9gk7NTBwOsYfcOU+4Diy5sMK1N/7UVtkNBqY4QBP4uLPlyIbOECy
TDYyLFLQDhxIqaoilFCFaiNw+kFTlMAZyIB18a0m3O4Hoccc8O3c3X3s75fAJ2Mg
MQk82eNY93uXWuNoNok6FaC9LRDSRLrP8kf4PW0szG/GBbfW1j03WeiYRqBSXpei
xlXnMV3FXiBXGVRHmv7AVFxNy6qaB4tHiWDUJCz7l8cDpauUTqY3r6XQ+PDDRIN9
TT66OcjNbgVWBA94bl67AYFj82Yypk50gyqyLUnssnz2zgTM1wwFVoR4ddCd/xHG
zCfRHyPBEWpTqCPP3CArgaTxh1SCfrzICkplHcRM8WC1lX7AWDGa/tGzgysWosqH
DuvOVkGihLIZif+R78XVJ306aHky9nWzCP5S5CAf5pHs/mwEosyD3ZNDfDJyF8op
Y/xL0li6WYKA96kt963X1/xM+OCPTC7djbngbXoLFGpDW7f2ymMvqoYZc7FH2d2T
LBTP21QzV21w9geKc2fWlGMH2SsG4f2ODFcz/pAoB6wZjXoaNVFdmk4+dsPiMRRs
Md3sl83tsq0zy/XfHLF01blgxPzeKvtEt5DAkt2EL8/MlYxidpxMRqqNLvtxUS+6
zqw2nhM7D9UiuE4tsKJkZ3ujXfHE5ag5EydpLVu3ctPK+ToIJzJNmWQJCRw+5cfi
9qcbuiTynZrC+XtuBuWOlfkJeDPP54vnZVj6V9Fbos39F5CZuusuPwtHj9RwPXDd
ySnL1udAHmgFMTmO1A0gz1A7z2+aZi91aPa7pZq7bHIX999DFAq61VW3dC3JTNiF
uBdw+LQ3sK3enCIsXBpjRD17KEmKDk1z3fGJPnmgDM84WaEUxuj64Cc3bLmOgFQv
PpuCmKTa/mMJbllDwnve6Tzly92NR3RgzPEngN1WjEqOVbB11lcgpiwNeBHdwgLp
VapN8PBSmTEI8PjTsKHy4UE0cjND0mJ0UFrLBPHJDG2t9hoWalR1hU7IkpQluN9Y
VPi1Ge0gqooj8MbokoPBkN+BgXcVigInVUzhOcCYRnC+/A2Kx8rVVDehlG0n7Svs
HbuU+6yVLIbSthyi2Br2loz6WjJXvqa7gV6nu6/sy4dK25do8WcQSbar6d+OsAr4
swbieTgh5e7dKQmgrNrzKiODwiw97TTiFgVeuatOdxxMGhLOQsysRJmLwtNg9jvD
MZ+ifG292C8QdKRC1D5MMNUZ7Vha8dSGBZE4jGhh+lKKrqkkEFbdFPmE5Q8ccRWJ
9t9tH+aZq9rxh9x1A+oQFC3sxLdQb5K71/k46B5p/CIB4xXEioYFkkCB5QEeiqvz
V4DX9Wp28KP7xocv2MrJkt4fBRzg8ciZ3Qp1lGAyEqshzOlWzLk3TEXJohMdyFFo
FwZP6TWBTRQzWIHGgAHO0iaLtmtVPICh8EP6Q8Xscr8axNUvUULl18M8gAbrN6Gy
5GrH9XeTCTpHnMcr+JXzOQNCRJcT4cJiZWhmHnhLDPiQMkbbP6F3oDOSCjaLsSet
ztrEcolHQZDRanfY//rVFeY8QLpQRpsWil7EVd12YTs3fXkgdYNzEC0dLOQTCXAF
nzC/+X0ZkY3Qqi9AZjbGyQwPDO/a7SNjkUo3KXsvrFJCliQOHFdqBmD5E1kQhd71
7d2nvOjARfaVpQJLgUe7jqZhkRQy27WebPOJ9lQHsdi/BWgB9Khsc0C+m57/xHAU
MzNkV2SYh1lKhNM/aBy86WiqRjgv0SxOB69W9DYjCas6n3RzLh8ZEYrrv16iespR
ktWNXtK7ACsTe/59nWiw2BdFmn5i0nreKHBpdVptPTwOBfaY2hcl5DIl/6gBNkpY
UqMH2tbG8HSjehQFy8k/DMc/ch9NGpnogbTL7A5JCWk7ogRcvSVyJq+7NDCNDzcP
iGMRleZFNPW1Ht2dmSbrZsCK1rfuVQdNb1YZNJ1tNoW+Scid0NWfDYUCWFeUSWIW
8Oij0DxPBMY3iSDHyGaYowoyeBieJFq+EpD5iuNlXlhVWYuWmS6ABgKQ7TZd9UiG
Fjwlx1NSQ/7oHKl0ddDIvWNjACkNmSoUXypcvf1rB3EYBI+2/p/R832o6U5nK3Aj
iEha5VaHVLoNhsRaWS0u/JEovCWgW22cssnHZVb3WympD+EA8iUsteD0j53NmHSq
DcYrpeiVticLHfM2w3WQqfVKKYIRklDd6Bel9zJ8fHiFQtnWrjTg5QdxE6VcVB/n
giePutQhkczZe+BUuY2h2QwTWimBib0k5maQts+pihZGXIJZSf/AAUwMSM4IZJPB
DHcZmLDIveJ/IvtNRi5uwm8Filq8Qe8FvCyHZyJ3bN+uz27v7RG8iKBF3GT6GUBX
PDO2H9uZ20z/DQV/XB+JYwonqkHY1A4+W1pZSfNOsJCXTw88dOTrYMGPA8K8q+ec
Li+2LkHOJoAKoTiL4rJldDHh+csFi11bxQqLq+9Un9Ha4kQz8s+FlkBeIb3fuckC
HefUkf48HUQO3yCpREdUTn/EnmJgVsRAHb6SJCc/4V6g0JOSAHkR371MlyXFPYAr
5ogBGU5yxvD1dc7okTUdLGnuGi4NnyKB1IYebAJZTEqz/IMxRAS0kid9ydVteYHG
FCaZFupFk40Mrw4N6oIhWzWzjRrx6xjgcKHG+FWzCriU3/w1l3tL00UXAB/bLT3V
qtEbyViVtI42oJfJJI7fDXFk2bqdlga0/JzInJ15dCtapBkgroQwHCByDtDBjYSg
herebWqze7gdtjyJMtS3tUW+kyPRb6SBAhCYIvqOKo8+Q+uTX9IQdKigZuYu9Xiw
lpcS6U2xQ/+e13OgMEFpU+W/vSTRe9imb7HKocVJnIx6SShDVM6CHdXTd7KENGlV
tIon7r9cRVqC7+XJT5hOxDnwt9tZVma4DbSeaF6fOx5oWcCPmO5RPjYEpQCf/M9S
PoBVegcgA8EivVp6QfDTiuAhR4wpfBGn2hZtDuaP+OX5DEPQ/KbCBPy2umFmQwaw
mcONTmErLAHEoh+WfWdKce/vi/a1Krcep/uj25cCyfhrQLBBkmhSS0P/DUBp6WEr
PAFr6p1/oagLFdf5kzhxZI08kRHPpkE3QjHVh7JBdHlCmhgcQsORhkGATc9Jy17B
8HT/pFjY1r58FeUjpKaioksqL854mZb3QAGqyTK/BMTZWvNIkvepT7jOfuGBt8Ac
fA+/Aov/q1oB02DEAXobLm9V4amJTumr+4S2Rc1f84y0VAhi4l/44edMT4OkVnTQ
oY6VrMicUaExZgmXXZDTYXrfa9H4jUP4YRy0lxlvrJYovfF71jtMwk82VXYY0Voy
Yf/aW2AxH2xB3Q9uMFdLBNq+1aeI1At0kdyaHA2wr+eUIPZqkLqMLcGKtWFn9mQx
q3UHyBpr/kaKFDFbWfUojb9ZbNpX65uUUUqCwh3aRH4RxzkTCbf6X5N9vB1jasWU
En1gLmvUVMjCpDq0VK4+tUssCk3Zhweojte4SkSUbe4r5P/4bWXTdV+nfB7oxh6b
R2aT8poZTwVtQSEUhtAgkj2TaeF18WHuNKpfgHvKt82zWA5Vm8swB0qnDsj7ibl2
Un9ltoESSSkqQi92CxQuGBLAgXDQFWTl1QEznNfoPjPoyX/5DP7OC5hXKOGGxIGL
jF3zJ0zX6uE0awo9l26YmT7BQqSLy5B81dYhHthC69cgQS/JmWb69JyGZ19H2YAh
WVi85tjnyY3WiScNIyDS79XrqAAhpb/I/Mvowndd5tC3XuOG6A/RwXQ4WvPjwa+W
fQE4wj+cqpvQAE6rcnhPUU2X3Zw2e3I9jJVcccnMqypkwLbgxOgxLJoG3HpWGEnn
mTGAWs7DuQCrcKjTlt3tV/jzgHZAxjzUofcI4VfggC48pv1qIfJiaBMkfNzKwb/b
sM+ChOcVQGrC71EvlbxIPpU9eifhKqtMO3wM/Dw6I/CsfjF95SH/eGN7AKjcIk4I
NqwmBDDuabLQ6HL3/h6cB+N+c/kwJG96EPaa0cstw+177dyOzWiOukmnOE6ykvb2
v6DDj53g35uB+5LZqP3OnFCjxS0dZ2+NbGkdM2/IV/KjwdmDKhNXq4xIx5m3FHhI
Le2eCV3XjK/ZT+kIj4r2trkjnZtgqeKigieajQ6czw9yCc2fp/yQSyQ0Q5ooIGKH
UHr6wWzyvmTMJCbTZORrh+TdjLHKJAYhDIviNf7U5IwG5PzeFJbA5SwcbqHMJC3S
w5kCuVPJYT6XTNBCJXqmA/87KHadxAd4hv/8/0KAiZPeUKr061ympdflCGj4pN8l
rpLSVf0JkdWnVMHeW8eVvS6D22kyXHEpIcP/AXFzAhHBKdfQV1rcSuRr7yY/oqp9
a+4Bm0A2VsyF35jHWLa58sEsvgOEBbWpxGm5HCu3w8V5XG8St8056UL9tcMfqCt9
YTvxTrBCchqeho4SoqAvuolNdx2dUZlssuG+xPjKAXGFI7qid7UWGZzUCFsw1MNv
tB0fKyG6oItjK+NFCLSY1B1oDfxmkTYuwV5ippj3evDtixGLnRwCWMiC7Q8jWtAs
89bHXkxoomnNpUwoE4E2StkqYjDue2dmurJijwDF8YIQO1N3YCxTJetJqYWBS8ZU
PO+DYE5RnCYvkEuXdolttwhyiMY+YRppyfvnU9tEf0Z6KHPOkWyEYJWk88uX80lY
QZoRgx6FFoBtMTER9W1UJhAvshczQm7Ia4e2hoJvOhyS40HwMxniAUJYomdHLw3l
mmb8EYh1GSfxv4THaxUadrOPhPec9i/SqEtNDKu0TRzoeJEFGkWcQtvQkY1419pL
OSQIASrVEDd3U8nuHvdB1KnG+bBjxZQTyEs7Y0461OJFeXslyfOVmGbxkU91EDpa
c4MPEWx9V/YdTO3y9LQD3gk61dewL4iI90Z0gi1wFPkU9U3XwgCAJ7o3futlCqw7
tK8btm/J0Bi2EtfiqYvCWKxY6vCRMRR/B1gx8HM+Y8ZlObYi4G9i+kxVYSnb4sEv
uWVmTarBua4h2A35XRgUQu2Q28DhuopJKT3+C05IXPl2rajAQvDfIODrq1NPkz9r
bo12oYyDVR9KXsZPfMwEDvjAMsJ9ogprEjyB0EwadgwcBHUFdPUWxaF26qC/qP0L
9Wz+RRouIZwHpb1WYG8LqXg8ONhYkdi0Mdym0W31xGqkRovZ+lyAyXG7EFb5LdWq
HgmOdqPicptNUvrmzke25QekKcZ8Imd53sr4TkcGjrh+joAsDzuiKTnuucTAD6/h
4QfvuAZwi4g3EiFRZaaOvLT7xTrRi4E2OCvg792ZljloruRSMhUAaV17wH+lCA/Q
C1IIw62WRreUvttON6lldL1NalbuD6Z2RfzB4e293kJZRNoJcyycAUzn5Es2cIqP
tcuo3uJ8ChQFgavXuBWK3BPGCCGPu7NrRlOuq2FVEO9XWCFIR+3WJ18OK4JLQxJ9
SWiYIJmUSy8W7OED6akaSRIfAkfSpgkSrKsmOtbh7M8h6uQzRc8TwTgRkWstvjHY
otoxEAgveaU5CFb+v/9xK2bXhQcMsYRgw1JCzm5FBRRtX5cikYAl1UFWGM4+ATCj
McoBGSvxLcVP9G5vLTPoKxrESlLj45M7Lok5idsDGTXLlguSkfQS0Ebr1NxeQ0te
TuKO/1iVGdbNPZMSK4QJ6c6N3FJ8UKGHeEPkJ4aryzjlNl+3hMNwdULBDC9pNNtd
yk21ghP8y2AiolAWRVVgWax6jcLYwOe8e7ZoCh0XiukpbrzkmYR/YXqS3hOfmIDY
iKzEri6LIuC72ysBsOn0RMOufnDWEiJncgys8lR9y6BnRAG59ddk8QWGCTWeKHe/
H6Gd/fOD/MAixOkdu8qig8WtBdslToluUU6UTohsqBoVFml4SAQuyF/0qiuo22KX
yaYKphIwuaHSah6EFBiWW/QEhLE15AK2A7JgWRlTZJ9KgjXhk+aBEI+s+uvzOzEv
cSatZiNxnIluvr1k6EnlqM/5MW/M5kKM4aJGY4u78pS7GF7QV7y1KoRFV03TLIKt
ilQkwpqiCa2tMKrTPCp1JbZplxU4QtDmRYGm75D2uuAG5xkL2Dkgju1hopnJNWIX
Eq6SuvgacG9PmLpHh/AvcigaKFBn5zi1H3inxfO12/VF8LKbJ7WAAELM/1D2TJ41
tOGNY/C+BmHigX3LA0/HQs3eCd4KZpS3XZf/Yc12+WLAGk/yPj9+P5WLoHvGodEc
N8VTEMh5wsvy+SruWikLzsojewdoppx3DxZDgp6ycOnylusJEi/Tv5qLdkr8BRQR
X5c+RFLZmb7KyRmpOTUMWoBSGkdqVe4YCWEOofHwNYWgp7qlkPK0AIKZS9UClIcz
GTVcxXK9NoEhDYamPz/SJNbgYTBRLi7ROJB2D2RdIsKfVLQY/tpibQbkDLJpLxka
IBnnEhVMe65oNl2ZCITP0Lbaa6IRD6sI0RjSTp7JQRvSqdXzqryVl0EyskAx1YbV
VgXo4PYy/EuE2cRO/RMFaPuO7YtuGFinlHgpImtRs31ECV0uswN5pfhsZzeXYwJo
OoSSin7MK66naAIpKvMPOqsHPtvLZfU2z1Xr2y6AyoEClk70f3jNciMQgpQ+hkgl
r0kpLRJW93E5cMfZ1RdhaJOteVzHzrhXOSiJVC3/OBl7jBA6yDxTh/+650+VJLec
50J583ZM+jYqCkyj+Y1X8KFPpWf8Ca5UAENWcty4BCPCBdHyZYDoS3gwzZYDLTtd
MKZO4JzZ4aK2BFB5K7Fx2Y237SFZ6P3ViVcFTTTK59e8nH4jFbBgyMgjltRt91vW
RU5Y/SkqRldDZ4Vm8CFKpEq1ketNktap/7qM8oCaSkDlHISzc0uNAO+sGq+LCLyE
4fGihvmHRK/NWo61kejzEZZOJblzteN74gyoJkphBCwQvsHh6brFfToMxWcmN6kv
kzqULmVhyqYdbF5QgnheHDL5av0RpHr9W1H2lyUHnJFo+CoNiwlfmBsb+I/nEOd9
qrRFr5i4cKNi9iz7sNtcloq4vchSXTM7Prk11JVwaA0nkTjtvLKUAw5ZN3wRaiL0
jO/AbkgPGGzF6yIv692IaSXw0mVrNsBFxqTQNf6phCTFhWHA3xTB1b/CN+8UFcEw
l8TitoRcnjZa6yOsnr632ibYxsSTKVHTAAv7wvKC2PbbfViolqeoh4cSsLauEGuP
PoCGskQGf+p+VXe0xXwVB8qmMv1qdhQR9MbUHKON8pwliAW2/I/alk9++DmpqSfA
2UbMD11RxX1QE4+EXfy1aKDHiDCVbgeObAoa1iCspUth/Pw50/YXGH0AWSaH+qAt
CHE4uYMoxg/c1eRrj1b6yQAFFef48GfMMyEyLCdDRyjXpyP0BGl+dxrhVxSDOWTI
WCtFEvIL6pnpRJDDG2WRLzg8fJtvRuICGMW7c/PCovK+EjqEGgZhz06E0JFv2d47
ezR3T76EJDMNQjrLC2um5MrGv1bYYaa/oZF3n3/rXyh8cPHUUhs5J2tM9A6AW2CO
ap0YN+zqc5E6O2FbFLsheac7LdqAUPT0PvxQUZbLruHpX5GD6ecilpYsNzP0KC3l
ap8AQ394Za/trQHu/N2YaFlKEfT477mr7hQq1qTUW1ZJlsyhowSPXuXGN7f1QGoh
Ip823QVBSOeTDhSafrYe3PNJ0vRzg5TpS15w+8O0PA2/12UPtAcRWL4P2hX8QzH0
arozcYFRceR5Ge4vTQNIfyFLxc1wk5dNK7a9geHi5O8unF+SQaAAj2SHINjBvt43
csDqxtULKZX6/c7dLA3Tliy14/w+x8u/vZ31Z7KPWNXIn6IGUhBczPWjSVU7Gp5C
eJya7/SowuoDsprPJAVB9XAEf9e5CWeKDSiAZJ6nbONnnOEPGxbrREV62Q1SjxDf
sZa3YT13cH/9qSodN0DbNy9Ws/lu/a9zIlGFapPH4GaSLp/i5q+PS7fjR3YERrxF
OxqPlXVhr50SLSwJE/uQipsNS1sihvue59nCRAoJhZRebGIXu/7oEZ3oFsgjzCHu
srp6AEAEEketM+liGkHJ21rxgkupxsd0Klf/mcJ2r62gQJcnA7h9WR3ZyQ7/kmOr
PMjw74kt5K73MRq07aPLwuil0WfmZz5EjRQnNF5Y/KgwUK0YSIki+jd+aTJix830
follmZqAKa3rwNfg+Z7XH8Xxp+0zDLANnu0ZT5eCC1BfA3e7C49XNA3yp6tc6T6I
fwW5kM1ButBs3LbKk6znadSIA4NxVJhsoZ3ydBU/6Y7s5oLwq9PirdCt/Za2dtKt
17vzoWKNa6dnbQZXwnBouE2Ohx+dA4C5HzFlDmpDT9ogARj7YdzBaehpNPvYpYYn
6GKYNum09fIVCOl1zV12x7l+bWPNRC1WQatReUiLbAGwzkDnPlSpApofyISuB7pf
uu9t1NgHix2gmFhOxgAsjdGHcdlzG5yNc+LZSUaafiOb+AJW/7pz8W2NGDDQfEVc
VKC/q7lidw3d7ZcjqMnnoNNzT5KtST0GjquzRHqrEx3eb8RyKSav5+K2c75hIO7C
sBPJPJA6vjutNn7MEobLdC8avaLskF66N4Q30B9mJ+c85CEdAz1cCdsqpkMT1CUo
rpsp3PWvTc3cvGlQqgTPzx0NMrcZ9cpt4kUZ7dpvMwB+iLalp0U/JchQgmJ6i+RS
hulplpZ1NL5TVZx8cxvaFHFKBhesJRAvxpfogWS8FFJR/XXpitkrpZUYasVrxxIa
jVQoo4pm1RwS/nC0+vDTHFhrJVAkeiTm634IX/kI2L6CoBebrIiirFjEH7QFZ8i+
88jooPyp9sSBm68UY97AucgYTOt84/AQh9X3wl2hB6eXt//TyvOPVTLj+tFwqrI8
IeeoTbpk1+HRUkFz+OK5HaZCYnhjtBnbsZLjQ8YOietzRgUl6AK5AbaY2bfWZQ2Q
A1JMts+Ss1Q/VAV8pGXylc+A3SEOkPI7rfr9McQBgSN+W0uc1nbe7hQp0Ki7ADEI
KqYO+B3nbozMFVcUj1OG5UXZ4OAGZCVMlztP022ERBN8REXCFQYRAQDiLUiK9yBl
Sv3J1JFbkMZLTiHzPi0hPsaEh5ZUyGEaJTLzW3aLourCwv7FdmNGFosmqe5qgpZG
Fy6bq0MYKePt1A6VQtCn2BWrtZhsHLqWqXw2BWX3JI2+nxKbHmCSIwwZEg6qvVBi
kODjSPTPHmUeoaaLydTlfKmXynaC10hZONxB6vdOujp/BiWZ3bDEWOG2TJkmvxgi
XGnKFh2GZ+o3GHqnEexIvBnIFVMUSj2xTs4Ru96HNhF8OCLgRrrf8//hdYPNYFBI
Lo8iDK+iF/kaEzoliOaVSsrT4xTVqEUH73kpgPnG7l59zYrjDYKvewkVIdYM8UI1
S34O0cCWIjONkEw5Z4IzjJc/a7/yZgfgpigirpy4fiR7iVXy8GrA0Jocyn7p9qaZ
+1u+6ARUm65rUo4jqZRM/kIbC9uI+rQYs2qa7Bf81Aoj0DpZ890wzHBL3kGqKQx0
pGoxep5b6w638r1IYyLYc6UFZP7hjBRnDCETB+Pi5bPXsnNnheBE2euIx3S2bD7h
l2E3CQ2I8ZUtrcFSn/qYAB9EUesqbgn7RZ+1zLnP7YbOHLCNjJHL98NRrg3oUjGK
Aq96X/7dT145beYipyEqW7yFEhQd8bjKaRzR24DyeXCzreidCcNXLXT2WYMPPyub
jcMYK34pQRGYRi92MslmVp1VXd6/fYeJnKqnhWEqOOz+VavJxoZfVPk0jg8jdG24
T4o7J1uK4wcZGZSBC50HzAQFyqyLFocDoAqvu3YwV/hoYXhcm7Iz+yO6Uik2Kk1/
qxzZNmedQZx5L0na26nqCuaSoKadejB9VcZ/s1xgL2Ih1j7daxm3oNCLi50xx8T0
IgGfbVLNos8utKdIPHRk9ihRFRjyRJaM6JClvajBQs2CyV1NqWg6VGHnm2+8tnty
XR852NgjaL3OJsncF92WnxNO1OL2rX8oOaAu2I56vfb8gNmkP6NY4+kNfRD7eReC
RH2WxkBXpAQSefqYnT2s4wg5G03QOnpQukMPAl2bMu9/CDj/fZvQz4ZiGz+PDh1E
uo+sciS5pYLY3cMHh2nbdxsJiXk9Ht84ecWnJSNbFNq0S8jBG4jCk9/VkuOEl/F+
Nc7EowfcumuAbm9OSLUrcbzrm27OeLXfqiMY5E8MblcZMhGBA1ia9oYeaI8KS6LI
6PGg3GmlRphqm+OUg4ItIFe5oCnCxi/I5CWmoHY7QpLGQytMMbH5m/wyGhSTsfTT
0XsRdIDasIKaAnlpOmWApSdWUTHucOpJmQsoNPXCsCeQI0ogtzN4ubYNO5EOkHdR
7KPNT1Pdu8PQUMVefiL7f1RPPPvc7fltn9KBon9ygPbnY+mUpZjD3qnfr5M4uO3/
s0DWP9ghXGbn1Nj6nHCqTR76tFwnA5n2gUdMH3F/eqM6/ZWwvZzDhzcAGBTyZNhY
R91RmtQu3NjizuCy0p0IBVoqk+PPBljyGAWPIeVj4nRwH9+cV/GJ8rxx16KNdyQT
kw+nIJ6YiD3u3jM+bSFf0S3d9VfzViZa0eEFxYpW+T+s45HiAhVtwZTJ2l1ZQwpI
RY5LeqViuIY+uC0NLeUZ51OBLJ0/SBuZWIaMv2FN0no7VWFWbjKwn3+nmNsLuHcQ
ipGJBq6FeaRM6tVdN5GKSAV1WhbvrygdW0zWZDaYnZTu/PNkpFxcBEdEHO2/sXQB
mxhSIqlaMWmhk16JVAYojXgHXC+PLL4ug8XSvSXt9WoZeRXJYzX69bFJ5Yc9gqDm
Svjx8oduBAdHNHzJVHS0LrS77WuDCpwwEAaH1sJvBFGKrRu0LYEFPvHPEm6R2sdQ
x1C2w6vbMDYU92QPHnpBxH91ZS2E92NTYwjl3yii2qGQ1/OP7/MmV2l5EsSB5KLs
dzd8LO7f+DryzrFcKxuU8CEpgt3PFtYSQObejX6aRAnK2Zgvi7rHJEurniMhMnpD
62z/KOgxvgGh842PE5WvV1EG8uy66t+/UsEJBL4ShP4gNKgdRuyxJZeeQh2uDGi7
TnE+F3Q4aVrAaPleU9UW1OH2uYx0atsZjFL1YOFIxg6Ooh3dIgKvg5ETxlcf7j57
k7/EuC6o+dRc1m4d2zl+Tllm6MyqhDQShxUTt8v7lSNveOfAAgBV79HGXgIiokR7
ZWiNHNZtrdArfH4tr6y9OHGa5R1tyJ5NfayYKNOawYZPK/n62skwIOmv2Z4xsS1K
CJ/rvBepN9kXnmcxxbpbvwYEMT4N6CWEgaY0baDF2uuw7XGPHnM7GJHwgTtSO+Fe
Hk/762vE57fTr8uerVlIq+p29bL1YmITNyhIOuopKQ/vqMUFCFP6IDEjd7I+gYlV
1J7fBfuBchTYpxJIBz2DNu81QHYv3nOi1HPd6ZD8xq/8BH2tjxWXieSuW/OZSvqm
AgXbdX2XJRHAzOdBAow9WL1i7IlXNKdGMsOWCU81kIU7aktbfoXpefKXtMDG4V+a
2XnQ8Jl2JxAJdWGQqrXZVeEYWSDeyu2PgTDjRxHMxuQWBMk5gqQ6aJVUfqRXXBdd
7BgSL4YeXgIzkLXlT3or0H6NMReybJ9jABB6arp6ZZRNnEbMkiq4CdX0y0qLLb0E
ctJ17NtKIB+2eC9RzKK30qPqutclze75B7n8NooNdMP3osVcUxIJMWkVs63xJ6ud
28t4pL1OMVoeIrSrlaMVa7xXlwcUfPSEvahYrmriJFyKyQ1m1/v2POzxuDYTz1SO
a3kDgzmlrZux3dzau/F9UglduBE8N0m6B34oyOmPWRtsKDdk2b0OZn6X5s0LntV7
CMUm+oEuJVXYhiAldOrmdSjzcS9CX8VWXWJSzZZZQK9KnWoYcv7xNvsZ7l1BNRuo
zTu+oO+W4HfsBQPU5HIPnQFGo1NXGRYot3iTGgPhUtfcREpLzQfgrkwOjf048ITE
0+XtEQTPyEeDTEW6u7I+UCVjazLo/GbfErXsjwt373d+A6fuoEUoJl9BnMPALgVb
Kvrl3dtLg7/tJQdZn6XuQsFg50dtaLRKKAtKgwxaPrr+e+T5bf9rMJALt+QobHY1
3uITQQ+0S5lp4FtSESuGgG2zADRs6Rrra3yA1+lj7JzRUp3WZfehaQ3zrQctkmFz
46cDWUd8vx0TAC0JyckbL6655w8i97zAFWTb+hIIsvhuxcAkfaNC2DVsA+k+Zj7l
pwjhZ2Zd1Pqkp9RM7jh140B0WtLfFyclV+HZl3KnQ1PlDndr49NLwg4J+4vX9VTG
P12qnDYfZz87uJf44nCVM0+shTFrDcR0jFajN6AYaoXbSpAUPdMeCwF8w7/Ct1jI
JR2ivni9yQ3s5aWAz47ibM7UrgxcQTJY6ccJGCivGLBGkijjVB0jlAuA7z/z8dVi
0mp6Xe9o633CMjn9R3A0YQT/thUikbnLdPXEvJs4wXw6lcXvTMXXYAFQguvc3AoM
+hVpUUVixSBQB/szNTte/Py6Iug20Kk4B1DCnJTnnU/iGX5KhLEE2rUXqBEVX9V8
kh7hjjb7E2zSNTTVO1ccb2WLuySr5tHKmeK7fIiWx+qxhHTZuk6KR7aXZy162H6l
U/Zg1pALEUhhrheEZw/F3aYJt/VbDWzlw5fhjCOSmdJyfolOE9mhDzbIpo6j7GiV
65ju09QZiEZ6T9uOyl9k+n9OYTjENasW7AyEljduUw6rkhwF28Y+gd4GcVI3dQGX
XWuuDiHrNcMcMSBV/7jcxQvYovLWmLlaEwnt/dxmOz89AVPilzu4oQm2wHjfeFak
dxS1SQRhMoULdUT8n8VC5CjIDuY96zp55J+b9NA2dlG/dUA4UWlme2MMzAbyAFts
iJb1DRuo6ypnfTbPHoL8dLAilT8NIzXN8IE5hm5rAoSztIIVHoUZ9BSz8zmWp9rk
56UplcrxY319GY2tp4Pgzl4wthk94L0Gu9ozgF+4GeDWqty39nxInWF2xD2KELzq
n35he4DGvGj9PSfwsvZzJTfjPZWdqUlGF0gtGnlpgPcqWHMPIrbJQvSudowq2OiB
gMu87dARrVT9Uq4L1QWWMOJFd7KAi5NTqJQToqEm/x6V7UjdnF79XEf+cnZj9c18
r5T/H9Pid92tpjjJqppZTqZK4qxmD87w+wg5jGUytklZXrAi5H9+RtlgV/oVKn2A
/RiFEgkLEQBM94VkGql/j6FBLCIOHB1pYCmu8HcV3ZUj2iBE0Nt4IQ6OTM8go83K
3qkRYIVzWsUV1eE8AYqhEPgh7oWHeoY4FjPXdLuwTS8F3ZQoc75FZRce9ymsUfQc
sTZhss6fF6tjEzGYOMZSjDB1CW6sIznv8ZYdP6a98CWCD9PNO8Cww6hTxHPxJv71
++LvvEmLWml83NjKxQsnQdNIG6RTzkGkMedW72OpAT5ILO3W5mbENhc5iAKmnECc
LM2ebyQnr51ptfr1fhr2kTp05WWSVS13ct7LawzP4g0fgrm5ImXBCcO6s4BKBM3r
ekWPTMWqDzP+t/1QFU+O+qPlOrH5FJ8cK9PcTHlnshw2a5+nY9yacVc7gePVwCDb
ut16GcOtG7gMBheSazuLKomgzQ2SQFX7cJPym6aP/V4M8C7bs5oqP7cT2wrl7js6
V19vxELW2IMD1I52f/YSZqFnsGOT/o9oAGlCELye2mo++J1M4llaUVFVbzvzUyYa
OX2fKxT0VCJ8tzxSn3B57lAJJpVKJDgE02fAi2ygD/ToKk9QU+DHmnxL3LYzIgo+
xkdVa5FlxjAQmB8AVMnttf/Lz8MNtXkZYL2nqhQ2iRgXsHpcD42mlHTkZcX3+3b+
kN/JBE6Mi9APCXNbJz24uMmuU9YZVgmMLgLMLrb3OmABIX973Ws6WQB3UHPjR+Wb
TT7RnSDtmPqwlmbYFPrnOJjGt3/9Dy7CIRHmj+6lrTQla3oqP4ZDoRdqB7XfP5Nk
Sa3uJhOjiQlE2+WCM3HOUb4tHqipgvvuv8ZTlSEvAGcRpUpBDK4OxbUVnl2/j5u5
2yW6n1OL4bkckgMqWnOcfOeIRmUXn0wM7DYUf1xfZSGGDNcUkiqpcw19RMBfrGSy
isYu7hTHNNg04PDjr9mdKmdLoVIDKUsO1FpJpi4gLbTty7FZrxqylxn0hhLtKzCk
XgyCY6QbC/07uKiwBq08iRKvzr3u+/++VjghE/7aHVjKCuSpy4Pq9VBejtuHGSu+
n0YzX0E5iODaojt2x2JjpCB3OVK9R+sGu7eh01MhE01JhAwk7h0G8igcAtDSTFtf
nmZq9cUMYqXhCG2w0Vd6UGs/bQXvQBjMtA3+waNrOuZ3w/Rfe+osPDgYpQWcvsIf
LNAxZM/Oq+NlEy0drR2ErmQhNoa3uqojtEPcwsYXaEQ8Mh1yo/9dtdqVfSoDiH6m
14h6k9ltSb7ktEPuEaea8eEFW/QVkxuu97kL07jFom1ieT6EjwFk/1pmdvOntp/z
nT66zYIQPzoc8mzeuHk07O3HdBPfk8UegMBWB0tbGF5nNs+j8ja8EWkF3UMWNmlr
j23sKkNbatQHXhBALKZmvEEhNbyhoXmIRb46SygkE+JLv1dyu4Twk/T2Hbjp6kZZ
Ewa13QADfdFI0psoEZJD633X5ZPT7VojwfWJk4gb+/faqdjqHRzg7xFnYUg8GGxW
9IP80bj2390LGzidQJ87WXHLEGcOhjmyGzMHw/m75WR6Xgl4klclbcvG62Z6BXLI
nJf8oPEVbkqihMQEboJzrVMMktPU7bsrqMSdD/zjbANORcbDPHWz7mvCfiQ1j8ps
wBHRNYv76w+Ap+O4rgCHRRPxkkGDZrM/tx1mjH6bJRe7LVRU2rvwiNWzCBuGImZB
UyiYXMS61M6WMnXr5xTPEMlgyGXv3bGz/ZgmJYe0XubcLuFOyS6LlIBkG402hxYe
N9BrHvP3zkZtagfEkhR8oWC335ZPRlolStpu79v4vFyx4tGbU0uM5qnVmzRtxHnM
1IS/dflR4PkaZ9OHV7L7kRndYFkQ2SenV/hZkEe1BJqxih6v3qdVoco9+lINIgor
SSBpB1NHYryoCblTVQIl8VF6v0b5OLmoi504txDo5hZoi12f5KUHlGsK5m66X4Jb
O/+pSvKn2fX4R3yOe9UHKZgEs+0rPYuI7WYJojBI8nGwkmOwcaTBaFcatPJ8Z9qH
1QsY1lpy5MqS06asE9To3mMXmfSbZ9EjgC9fs8eNRp7PM1dCFAaP7AiTZNz8+GgI
F1To7tvvSWFZmfgdSekqiNQXZ9acr3vn0AlcB47VS58eHT8Jh4QWwBMpk8b/h37x
3Zes8g3PewcoeK/4GS9haIMygbeUlmu/ioO9bjmfCCgCWrPrPM4imWniIRb4lZgN
SwdtqMuUdUYpykrP33Cb7H+MdIaaXsnI8Ijfnf0XvwmzbjdtjluQ3Be3x9G08rYG
kfGOzvSxHxRqj9beoqWmkqyP9dMQCGu8dmR4ozbNG4k1AoIIsRiaO2iEPjEZ8/aT
+IJNyJir+6j5R6bRQJl5cYyrYl0vLuYEq9UHt7RUvSKCjB86kkyalAqPuhRSOnxY
Ql65JB+O3Hh99u/vXQsQgPg/6aGulowkGkdrNyD2rt6/vEgV2nn0CHzEkGY2EDPe
wEotg/o+bENY1Ma7G6F4h4aLZ2jzqVWWOkBJgpDndWTWuOEl8SF2q96MTH/4l+pz
adygFSAHHRojqu2us5/hx3HFbDuQqRRZ4qQftp5L4sh5/ojS+OtzPJNfoh5gVIzl
jGIAAKbMAdWDqOckUckar+N+7SI5j3hqOnr3EYdViPOfVrVmBSHZ9Q+v4xSXT8c4
gUXoNiLYUopSNwy5ivqQZV/QLkHIFYz9p+Oh9NF3luSCZPcWUk1bYKBx6EiVQfrr
WM8iCiFMAXzFBHiem+dAZarllKskE0L5sM6rN4m64jPTmAyy4nWfW9r7/sv6dhKf
rK9iqlKC+l7XVNz5nt0dfS0oeMEyYFHG+hRmDBn6N1gfXwGoNViXd/xpn8CBwzvi
U/ByvzOaV6p8HaxJxVSJ/YeE7fvSwBQ/vejftKlYu6gVO12lccXRn/7YcESsbzb9
DbEubkKDKCNVqpnuQb1iauohjL1yyJBKPdM73DIw+jeHlWcOi//cItON7w1YbDNg
J0A11Lt+5mYUMUp1Puo0elV3n/t3HsFHieOLrP6iz9VfpcfrcOetm3NFP36OA1iF
Q4cXCVG4YudOt22Xn7xtnKVgtTxKs2PkMtel8WUHU9dhM0TokwapoWWwL8sn6XcV
wSzX7abAufRym8bY4hyzY3V+SumVkIR7xWachwA0f982Dy58Vi3TPxLCnf9xVFZu
fVZnhXvF9/XcUqpA5xsz3LU77nHfb1AzJns2VOrzawlyGx6q+6rAAx7Pwed7L/rY
wcgkf+IL/w896AsQcYgOyVNRpXWClrSQJhezD66aiSu2VzYa50Soblm6elsL4OdS
FpST9509g0uDMu/ryE7ZOz+JcOT5N5sQ9MDBN6Jmjg3QEz69duM/TZn5ruEO1jOz
Pt1AEvLBMUJ4DT5CuxgHYResZ52iOfVHyRoZPK1DDj1V3PoV7K/LQ1vPvlRidqWA
XwPS2y3uFS7E1+Qy2blET30j0+/P/p667Kb3NBcQb+B40uQgon52xABueR2ioXmZ
2+aeyuCXqwnimocx1Am/0ahrce0j8foTDBq9jLvakZhZ6XNJLPDvfQGb1nirTj9f
uj3Zu7c31wxYTBMC9v5Sb+D8klw7Wa8J3ZLBFkru8CQkicLrGX0Ogb3TmtgV8zh4
zCOvkgNff0OmJ28EW12srFESDX4rgzdJnUAglQNSn6mdwcgi3nQSEbI1sjcKWEoc
9Jc2eszyucUT6F3b4sUhubdT5JcrhcUjm3AzqN7nRy8Os6hvGsONhLl8o1NGCHfz
t/98VtBQFxJLvHGK0PNhCPcEK5UX5lQ3mCWIRIYnW3ROUniCQZhld22jBQbak9Hb
xWpFQHotJohHGPbLnwCJatI5nJBf23sVCw/zmP030EGnia25tG9PpPB20R0ClYnT
Ei1c8od3CBuz91/ZHKGwH0H0Yni/0kS/dMJ8OADKXy++J3iYLQIcIgyFA8YZvWz4
MI8V/fmnLC5pZpGbN7zRt3rdkt3nv0PgspVsUrKYNVTp9NRdRLgkBfM0ouIqr6U6
RGra0132LL6ZvF0bRZZ+ZpaqgeJsz+MbWluhVGuI4aepU8y7i/rBEoP2j5eV8q6v
goPVxu1emQmydmer7ZSckVZZP4blMu8mU3fOk9Bhu0Ma0cQ/5wa+K8yNCLutTOCr
T6O1GCc0plZmoiDNkzmhWkwwf7GNhQjFJ3qBdArUob9oMr94TdwvP4MHMeZMsL8D
bj1CwEc9pB/n2cop4dNINHMHA2UXzbXSbZtTFxPiK5n1Bce3XTW3bIaO5GbW+WrQ
ErZ0hC6bYlZ6hhh89d+BEvRfR170BS32HcUbJJb/u3HHTeiGxMlEEC39IYQ4FfeJ
kMdw4n3xitHMD5u/gqNr8OGnpTRAZ+YTZSkG48BitI204/Fio86F903qhlXJkkzP
+Ez4gAqPwkckmTP5sZOlO8mg/WKhL0DXX5SqwTLKky3bSSYLxVphJqKWP6d4nnpg
/+c+LTrq6bRt8Ic+lA7KRVpjgI3CghkvutRwjUSZxM1j+aKez7foVFTccQXD7XWq
AhDgX/VM6AxwfwqP3xHe4YGyoMzsXQKjX1Ryn6ATjF7S8gOloqfyCU913vU7/is1
UGKidsGD46dEp7DwKveIpGkcFC1+sTkr9zb5QDf3VvLtfuEq5RcBwin0RywxSxNu
ZY3XpUrLrnJeugYDV+hIP0yHjej6StH45/TiLJcMuyxYpcoXmiDu6zZycTo88mXd
h/AyMZuncEEvey8WFzFIRE+uwmcepqdSVbktElQPGcVjLLkAJ6itFawb1hf//mto
LQFIxtYtBkSgS2GJHps7pCWhadeJb1/ICMuQkTirmqNsLFfPtEW9RJfcz0J9Srlx
bWsSVhVoRkSxsVkLzVSjD454HlRKiHzS8Tr4aRCWnYbs4Ro96D2yXYM8S58h7h1T
vh77hNTHb3bVdVGQLlULtVU/1tAeAeGyqaMpBTkgf862DfLsHtxhMPLU1E2U5jrg
d9ONvXUtPxqw9V0MCbtcA/Qpha6x0JjAJDw6M7/mmTdukNcN536/FGGvd9v5pc6L
0gzOkIRHIlUc1ukM1AbT73Ko6tFb74eB8/PhYx+mMz7EeaG1Utl6EWGlNGV8k3gZ
dI2qepmXSF4DYlApqT3vyyU9A/H+LHf9OgS15m6jnugzYwUUs5zN906RBJY3Bz7V
fLrTreFTo8ofobNqqFGAxlGNA1FBYdQ0yV2QzWR9aVysdvaAz1MS4BQ8sEIVEEmD
x3V2KgKOonIhvtGgMExLsUmQ20TzlD7W3Ez4zCs2f9KacQrDv8OWZYqrF4eYE8tt
DZ6LCspKq+KNPVLA/3iio/iG03a6EXcZT/QFlZYH2HJeisgUM9DNViNnngf9byht
hO0LD/PWvwkj+gA0L6VMu0vBu4VR5FEfQHM4mnnm6aEqZKlHZAcvPiBSpRgxmGYQ
1Q9YXld+ySP+Co9+z/YR1HNhn+1RZ02Lx10B1BJCYQCXxSwKjCydEJviYpM1mV+S
bYsyuvM4/NOkEIUagaKGMeooJT1qFBqT7LL5WwPNcPQaq3AAXNBbVbRRjr3bVS08
enq/+w2cIKNa/+fMiFj5l8vxZQ3eAFLPoI+COAZ7iTPcElRRRmWWRij3qddm7Mdl
b9kUH73DGkGyTFposALn9IlE6tJsaqDB2i2E6atSBrqhXX1atc1gxsV6f4NlqLQX
HWwLUUkCSdLGWxAWpppiqHjEY4psq4RqMVM56Arooz8JHPCAWQY/WCmDAHRaY0ER
RJj/drJZgsKHrNJz025PvDPiA/b+3HT2gi4kIYNkXg3/zcB18dgVU3C73taFa517
1CxoohJX9vMCZgV8Hl9XFSSM2+tqW9NIMR3eXKZ8icmnbXAjItZtVTuQOOt5Cy8S
7RsBoqSat+8YBoG1gnNeylK7lk49jkVp87kMoEs5KCYMX/wJraVY0/m0lAPK7vLk
jMMvP+IQCz3xYW96R1yEdxv+aYv3iFwmn+GMjfnr7/zK5Ir0JZRAsw4t1vAMbwv3
ivm0T0e2qBfrp9/Wtcm7C9Sl+1SUMcO3uygbCR/lEnwIGsIOK4sqivMLWYgybrJC
dh9398dBPX7JlfRhRlkGPtB7WvY8lCwC26U3g+/fR5Yex6FqqJ6VXcqLZXNIAjOy
luVTTrJ5gZ0HvmhTRpcX97YNW0BNOyZOvAevDSjmlnQEAkS7vUmG3Q4ByjFyRF46
Mq6A87WUwYMWP3rcOrPzAzPbrE8eXuxFw3jGRNGdir3i8ntSbRIc66yTaW09NXow
ElApWJF/guI6YcpxChWNbI7gPCQoPCBGkJp1k4hxEZA6P/GR2aDoqXpoMtLNZ6bO
owmFdErIrplDhPZl+l+Q5g6W8LH344/CCR//NEpuwMGIoGLgP/hrIJzHXRLLHDa8
ohhTy/MNi+VhwEtcl14umYWzQenu6ODdI64iosk4aD0HjHWXhM4GvW4tiMu5k1rG
a8q1VpUqWv0aIXMH0t2vW/S8wUZrhjK78GfcqgLY0Y8er89i9X/3BtqNRYAJIXn4
LEjTa+6+BqV6BQ5Fq5VRMhLZuQYWkwpuGgY2Oq/EqV1YoZAxKuRcQ5cY0XmuIrCr
N2EemAo8sw98jjDrvIrOWcpB+EfnE1dzFr71B1N6JiTz2etd0CYvIIv8i7vvQiAr
jAIvI/DE9SMXONX68cND6K+N7yHknsNnzbTp32BXZPgft5rmuG2I/bu16m4z8whW
/wlpK/9jf5REEWRGTS//jID0xk93QE0zoLn+hK5WSXT3pWlKx4vjQG3lvCARQN/B
YGvp+mIUfLyDHw9KZgm8oQZs/SHZ0x3zQtbsj0FvqBc75K46BfmDhHF4cW19peeo
0KJll4CoItHIyxN1s0U291Os7GuHDUToHB5SagciJAAililnSpFyzVRPIPYpxu7N
R7j3BHHFDHfVwls8nhJfsQAnGB2UlIbiOb0MAapkWgKCp5f4AxDwfun1LH14CrkQ
IG1qzvbyR7QUObWRi76NJyiRAVXBCCn6JDvajq1xWhf24/wRFNm0BfSR+x340ad6
WYuocWkfsnYXWGlk3XFCIPIow9Vw3VIUQvqklBSxn7waNaLcUlKUSHfhjNKfDuEt
8lDJa/bQPHxu0rHpIetVdYt4ur0BxGWF5t9MpJH2+hIsK7u/yB8w1va31/Elo4iZ
ffyHZgUgo+/IDpnbeWsXpuOV7bx9OIlV4U6/0B6tmooq81DjspaUrb/tH506npkU
0NcWkjfzT8Hl46naIoqqUD64PG+hvrxlqAOtXIKuAjza6LdSlcmfmnmuJ3vNi8wk
g0v0eg8K6vbRGNa8ArCR4peRO2GA9YMxoDJTvvuchY52275trGAzW6nz6ltmMnzA
meTN3yzRa1ISDUS6EkuwSlzGPLGVzl5Zjd04Pc7V/vmnMNkI2AeCku4DVw6I8YuR
9ER6YrXoDsHIhVmvO65s/3z1ZcA22UYHWbbDavYTsZOObuhNcWWTg6egyh1S/SNf
VQ87NWqoDcyAI0ga0/hNpwpuPqAVvneQXQzJTXXWZWM5BR3YH7qST7ejTlHEiLgw
y3tkkOJfGMzCZblXz/99aViF0IsXKdVXvwAIldhy4OsOzJBQvfrZYlbVCSvIja8Q
o3+Ig4VHSI5I34MLsYpQIkbmYyOtpBhJ7VGKmrSgoULyN9PJb2a3U1qOpd2zQc2A
V1RhVJeIb97GgJ/qF2DwKSM0wTvQqo7cbSGvqxBpb31RmfoqRDziuc06HwhOHTWV
z+BiFv+ZFabs8q8z9YeyddqCHBlMGk6yxUPF7EsRguft5PK0B6MKqgjflucf8Ylc
po0paH157P2dTLxVxWdsR6u3BYAeqEjH6Lujh2bPqA+zCTeYj4dUc10riNXqIq+k
3c4zvhi2+nn/GyEPmZ3s3iXDYgJ+gmuMzolGQqGsRg9Z/gLQDN8NXHWjcxFQEVgx
9UHkSClC2kn5GoID/WamC+WKeY4gMAQfhiz6eXOw7Ns8AVzmDIKAntjDDYQKrnTc
NR7BUQzcnAmQPscATH8ivyZtT7hzLiKg8j9SfB295ns3VKIcEipUCVY14bojXg/l
L1UCErKSq+2ZFo9kVwgtXSqSgPcr8K/CI/WXuS6BPrEnAKLiJfyD9f9IowKgZr1k
uda6AZ1DVSW3eEVLufqf1EH8CqqnPyH2RpvFjVB+minkGCohKeCuqBUF80Q6zBnN
FAW+9Qbikmp1qPph6vp26XUvOVNUzfk4XDnocWbiJsGvg23s/2cn0/u7v/PQPG6d
zD9fxkJkZegAa4m4Wk5lX+YbjWNX4Z6ycCwt1GM//ZRg9gELSZmBZ9EJbQBRYT91
iZyCSJbdqJr/2OO/DlAjpjR8exNweH1pBo/8b+Ocdybzlo2j9D1RjimofGNEvnY1
ajZ7bvTcxXtIGtptg/pToBB1cAWfIdyJ1jrQ71jq7odlInMtr448/BlDaHJIatBo
2eoWnC9a9mrC50ZUe+56qVOW7qW0sptINbStgbnqrWyyXcIZBeklbwBECX1sErry
qsIEw+y2HU9dsdy7YdmKDXpBLIwEMq02eaXaQFr0aqtlqJZQI32DNLqT4vHydOhH
luhQKNmtY67tHkZy6va6sGZpivsEmatslikywTqCuGHHcb11RXCTYjK4rGFq96mv
gZGmGbC1EHraqYqJlSNxCfbUWyMYnnTcC8DCoSelFWVhgNPhW4Pcn/TpkcOL3Y4H
OwJ7KbdjwgC/5TUphHF6Wl2rhphYG8OaPkuj1tYJ5sX+toPc/IK3MfZLk+W7qq6B
llIRuIlTmNpU7iG5ZpWn1EqcllX/l6aUD621j4+AF1X+jJ+WGAEIetXegHzS6DYb
fPH/ZoAnaDJVb78I6964Dk+L3vgHQoEuCLsGLQTkaTMcOeIdrcT6ASU/n9vNU8Gj
N+nldQGL4lnFFz3GLQh2O9LcTy7neg6gL3MyJJfx92fszhkGmyD7X9D3r9vN9i+0
1bKvIYCHIajU3h3fyuytI3WQSJ9iDkR3ig+OL5v3oL7JxHgTanHtuQmZEjoDf9b7
g9JLcu+8J1hsfuLiFefoIiz+Vu+Fc/eK7Wh5U0V7mU+wyICNPEwV9m0Bwb1Qi22u
uPIrLqFp4S12qQo69FTK50QK9NXQrokP0A9kESwVR87m83rLxutFNJFpooy7PQil
stxuYaxbMlraFLZ7hLLoqe5ALd77eBkcTREsUIWwAJ/X44pHQD/jQ74gpTrUVX4n
hD6pbRuP9sq9o5CVnNB2z/cf1OaKoc3UMxKSosgSvWcX4YuJp32uPbDIruyNj6z8
zVdZ4RbCDfGALA0JkUI3q972kNcav8SN+Z1p9zLLxOqCj365dTuH0HYGh8dzQAxH
HUmlLJ5QecdFMXmufyGIj8kBBE4KmvPDtRdau0knlpQERHcODE9ldofakCQCPdEB
W5h7k0uJ2yrDbanpV1iR/TuLM5bzlmNxzcJjo5aGMnlDZGUQst5BX6YSJoTyxsen
L3yOHlP5rBQgZZiw379HSJRPbbDPdqQ2b2pnYWtIC0EycXmLWektwOyHGijaRONe
Zi5yDKkODlX+tzgLC8Gr1w/xwNsL9WXb9NmfmVp/nvkVGZ/MenZQrwSrS/jKRiZV
Pgdtz/TQiPp+3qLj+R5ZTXkpOo9Qq5rQWNWTumt/GZuFCdp+HsDwl5tfgfgBshHh
XWcEVy8oVOM2UzmjM5w9SipD/Db7+sBVUOhg1O6mWju6ovMJxTTznU13ZdRpUYWh
FwBCZKtBjG2VE1m2z/IvB0OCnb2hrPROQssF+EGSnw3im/Z6lr06AROhOtk8VAv2
iBjIZt3svjLz+O5iYet79v0EyQBNyPbFS2GkLwMkFGmEbiU36PpKRsyoEnNAlzNv
MfDNrQlU1pL4jOLeiswG60VgEmBhmOQXXCrpHUs5eg5FcVpVJLhKxTbr7BlLT+I2
RpknvyYJA6tjfqTRWG+NBC41UDsWpmcEK82/zEcPMUIdj2KpSm1Ihuu+NLN7UZ1E
lzipvVD9JIReEhgwrGFl0+AWkyDiUaYs/w3EIopCtk6YNgHeMydSzB2CpiIvUl04
WDl81s8VcDtpAZzeQyi+PWGiul6EvQKqdAiZ1rxWP0CncHg3S5V0kJp+1djMyChX
ECHIO/J02sd4nCW/R4iAdn9waSqX5OzbJC5HL2WdSYbj37QJrpPhJhUuGDOKH1RJ
OD5hROY7jH/stV+vZil1NyufPUpPqyRe54Q86pagIv2b3VmEm0HyiRraaEU0NjKU
Zgc3onvFrG7+39wsfsKDMzReS7NgDNq5FplVDUaTK1YEvpkPqMzaZLDHGJAZ2kC9
XeKYMVLPwSA4oLVzlxzf8TxQxFEhn4y8nKG1AG8yfe8InkzgppYgSBD6a1OaytGD
mfLUyWXX0tAIRLNjM/Nv6tamSKtuiPOq6HQUyEqfGVzaGUep3TWZk+2lxcIDVeMq
uVp/1+jDHcGSwczBEJzhkvRih0oSYssdNOq88P9Fd3IqHlX4uUh10pxsDGNYL5qK
IIEmHSnHquOIvTf+Hedawv1pCDnwFvyNNALWq7kbsJ5jUU9udKZoRJ8EImn1IVB1
BNnK0/hRnBjgieBZ+vWlsDylB8jxVXxntInbJejyQ6bqOi/jVmWiFXlk9UAMkLIl
25gG5kIbBjSrUVV3lFBQrTcZffGOAn3hRkyUbE7eORDNX29Y8SLyvF0URMOTNxWQ
/T224qmvtaXStY3ylC2Lj5LKUjXZia1/yx9avR64RvzF026CwgV/NobJLrvfmDS0
LPpC8b866nQQdqfY3/hUthXqH4UbImYeWRKuA+J6DCJUO5gjXpINSd9Q2zUn4DYT
+EdbqUTOn0cuh9PgNJqTyQDQlyFkW/MfjhO+cLGM/uWA+0YCoDF6Ql67Dc83uGdL
hGC5imJOov8EsYAOQ2ijVMSSir+HLyRn4YsMv0RehlK1Gd7Aygf6di5o4rCNAayD
u+X4RtjAyDI74E1/nkEl5A/mda507LLGP/qY9/Ir8zr8yNCdFi3anPeDMNt3wISp
phSundcQ+72daalyfdMWBeuUxUO74TxJtS9/sq+a4zMbEyuKaxOJ476KcjwXkXP4
N/8TTMvwbgcI/6GCQrpc67+kKrU4V+lG/78UffIJYU8355c4hXrXxD/dfiXeOnk/
4EBJWzrKpWu7n8b8zkmJ5pKkn2mBKpZXcy4K9Z8NpLbvnx5C8ggI0GfPAm+rLpJZ
/thk04VpCHZmwcOrh+4ams0mt04KxBOuV70d4JJ+wKQsS+dljts3B5QOtIq1hzlv
c5jS6gxJTesJX/Q2vTQpRH7wqFVt6lqPjUhbx0Rcxlfz6lOTGQXowLQbUot7+INN
4sRMfTOfI2C3Dh0Cvcv6UbDBJ8IkQysnt0JDucRErYnamz5PwULWnOuIU8/Y8eLk
wLAWhcFFJL/1efzmIw+rn0jkMK6DGpUTPu9FpUCQH983r8NeLGe46ydS25LNtcoM
sqhxWKdZZcyDPtJRkDPrYb7FMPEnMznx4rPMOA7sztLPD3yvH8iYWt49TMtw/ITs
jgQJHbDVIF/st2u7gXVDKMOLur6Bmra2Z+B53MNEJQplcQCnT/t7j6a9cR+DDR7H
52H3UmJpiviGNjU8fFkNufyVayPx/Ml6eVUvpLfaXvXSOTaQNtpKSkHDmdZCylt6
AwogevWy8aXkmaqIf/r8bEbHHxLtqhSf0ZpqVhhar4MYsCsnSWLKqPAoqRPPennf
r0WEZN/JKmYeNEyqkeGJf3URytgV58A8ACwd+Ik2Uu3HsNDLm9lSacAzCunU5vUc
WeyrNSCUqUFS2RHg0rGJq/pLEfj4L+Zcrullo4NKPYZ9V+2GFIOxojTJKGhD/I+L
yl5Vz9TQ4W84y7frDjffnSAHspgvGpHqPbBFRRqYo6PWOtFv+lKwT8aoZ1sz5pVR
0P/JjDBRTnSaZfOf6+IU3Hkwt506/vxm9Zu5Y/FevjuoonGKZ5R+p7Rtn4vzyXAP
NG+fa885dAkvrgGLoRo7iLiLnfhgaHSZOsxtFOSVSeXLyN6yB1OsB75h5o7GwlAr
c1JMjj4/6Kxp82Kdu+uZdac7ZN88zJYvT+WHSMazB26ILuRloHlHBQVBAlKmOLd7
VuQXd6TJHh1Jdt2JBRb7PWyeQQepDzMNLMabFAtUG+UyNdN7NO09ayLGV8U1NbaE
3Ej4BLTiFdilLo5Xf9eiUNP6vI1ECIxnKHbq3vXTrMZBfUmEj/KL5x7gn43Z0MYM
PqZl8VhOmjCxHegIxg2MUtkKsZe3MfdBCeKTz4687OrdtZMLuKRxEnj4hR9XscoE
33iG9SvxikcjkSeH6TUvZBu82oW6sdBNB/eODxmCQV80DhYgheFmybKxTOT0l78M
Y5Cdq5NXRU95LEOw+lLUeStXaYa9Qt4gZpTg4rU2WwN6ZQFNzKwkBZcJHAmD3atR
zMtqoOvpfMObd1JkQGVzJYOcZ0LF33UV0a0Z3FB2gvaRCuOKUXWKoY0sw+Cs1jtl
34iEc8oNZB0oGgIMJMnTRitnLLapX+AwZlImafu2+OGlNPljTJmGuTgFhuwNocLF
YWT5kVw6fUc39iYKZun7iq8Q5tgCmteEzH1SqKJPRrferATVj9ZiJf44zfEWKkVZ
xp2rIOf3mgI25HOcWORcJD+rtorkNvVLZCbU5A1pvFQ6FbGSHK0p7EQkW83XU7p2
yyVMHyz4yaV5AinEDQXmpFAWjAMl6DB5zMh4uNYdL9NaKa0q3Luf1bZQSiqn80dH
nqpFkugrE5WAfiBb75e1ACIiwvn8dICHAX0O7dsL92CSbWp8zNlPMnkUqHOD5VJu
tYlhVoi00AYMEstNwxiPZeNGq99XYb+VfyRW3uK1LCYQ3P14AN4qaeblmqgvI3db
ap4UHjNc/NIlt5D2Iwy+zApGgzGp+CLse9MG6juMQ3xBdtZkAZAVD3QIwBYZoUhk
be+jM87EeQIpDPzCLdAooeVvrNpVVM3ucOcQfADVut1OJOBAtJENvRHsETbNOZpM
zblI4ve2CjLRJ1N5JEveC7SsQCRKpTNZmAoBGMF04cBoXxLLk7XUZ4x6Rr9WVmAm
wU3z0wWKJSeb1J/nYY+YqwF6oZchgTqSrQVsWiXciwZoBYXuRGRVPsdKKT/pGdDN
5c55xyDslB+E7hqTh2V1IlSgOkkauNEu5mRIR8rv5lXOue1yMm60gTBRwrS050w2
Kz9eQXVxWuvUSgXY6L4b6ZyEyQaQpl2Vu3W/HfgMn3PscjgILzAle9P5ewq1LUAP
dRC/ILxXWx09Kpz2O3bvOolWiAti+i/KVIfqbixxT6EdnDpxkf5hvTMyAl2TdXEl
8TXGWULkfDS3tnqqAd/jL9+GTVdpDT7IjizcVrASfOJMipRR5xzyWAIQgeoPuxMZ
fyZ6MnYPJTsh2qwzCv7XYjg0tMi583lKxoKbhShEAB5IYTZ305CcmaT0Gag1HooL
FQH74vrOaMKpgkgwlMX3KPXKl/fhTC3a6IPKXnml+g0lEOPCUPwABjv1Hb9bqFm2
AMNkk/X5HRJzd1Ld2l8OuyYvQ0OdgZOQjeeK0MGhEAMPJNwiHb5e1TcopxJXyV14
W3Z5TaWOoPsC173gZMByJbObjgvropIZk6JeGo0VCcgzKmeLTfsiJBuedbLaAwzD
5SmLcb1iWqHTdpEoTTeKm3b8YIoqPxxlEjmhDUOzXzvs4mpgobSlxYCn/zIgGpRu
hEeEGvZqk5vT0iIF1be69K9qideqRPEyDdZLKBob9Iiqmb76qFFOcteHkGgn/y5p
5+DoQSKREQWs42AfTbqPscW/GhOQl00hB0uIVNvEUFGkC/oDugdD647ZcecCIwA2
YBe2A3Y6Hb87QKyYstDg0yfe4mGCr9ckosVQqy/xyUQTuNyVmDk3YP7B4KKGqnE2
Ypj9a1PZgjescR9nvh/oS98J79IQEubcVHmN+ZlZV+45bEqY+AAUEgqgBI1nCJU3
d+HCnD067X76g3VWoLw+sU0xww70SkabOW8O1E/TX3RDBbUKX9/JY/DdyKpYlTmn
EKuaC0CGNwJ+tErkoZYPhwTOeUSsIfYDxpni9DmxOE7W7PBNvRh8Of9pmu/ED5o6
fbYJjB1kTq0URexM4b0IeQxgbePrOQ5pXw0zaYSCJdVY0Ud3pUxIWxhPCP3HP3O2
/tTvLj/i5TKnn6QHe1XtkUq1JnLTuUbqlSAXIFTCAmp/cvQaFFhJqLXO3yNzXgl+
xszDljZgUTbr6xIHu6QcnfJKfznkgtCQRx31w3awlCojTvOpc2pW/Yc4BCzm7Wx4
yrzNPLGhRUmOilWjjteESMvFE/s2osf5vmnfpr31bnFMUbFx5raqjoeeHlr45G9u
yQAuKAPLwvNeuss3uXV99qIIukbdVwSLzZVw7baqxhbJ3hjofuXt3X7YSm2EpCvj
H3sdUeP7D3vWjtY49nUf+l5Frto3WPFDg8M82NYRqfzmRuRmluIyESG9EOvy48D8
NvPjL7ePqrLoxHEbaRR08Ff7rxCBbr8QpwvJ48JQIceMQV9n6jLInpHiUzWwXDGn
W/pYVUDnWZC1B4MyeCra7yC7PH0TREVsZ8V+A8dj1Wv3oSyEOjaFFiuI3dTbGJ3c
yQ4ZJxv+kxeQ+zXo9JUGVPlL/qt8e+lunE4C1dRgom5AxPUs32/9BL8vfcJN63Uc
gA2aI4owZ+5mzL3n7wlsUqPQ7sE32PKcqdF92u7Lq4c0QpAbIixRu8wwEgu/6V/W
meKmpHKHBp6uDLBD79fAZBDTlqnX9GNeSY7aMT9ZU320/yXLhFMAnYZWMSEAcmwI
hBeRwOEQxFd+juC8wXS0WekxXA9Iz6r5OB7GDG+8iPFMjjls2XvptsfYzuwjk/XS
nTKbMVzsV2TNgUKbqSRxDpOLLdcWQvVmcKYUltvrg553NANfRilvXfvAPKvoEBfG
mWTfeKsQhwSdE04kQ2ZQsfQ+l7HRYzznveZA3rhatFLxzroeN+CJnfU+R4tIq4n2
5rlB3aVuN4pPB6GY8GI9O5vyWqi60mvUK+34mDqcnk3nGFLgMWc6q61XqyRHTnO7
qHiadqGrD93UgopO7phBttG8pzy9PJrE/OytqMo3X1FMY9aGA3kk80zJVC4HcypB
ZdjpeaCBDSlTYjI9/LSJn1c9NCYhywBy0dKAkHZ3fJhTh/T1v7Q4H1YnmNLEy2dj
kzEJQUyC5yzN6Csjk85dbxFoUgtHWSQR2DFjVn46YuEFn6NgBJh5QfiJg4/wUd0y
oYmXMdHVNnBhsXyK/kd/CEIEmxHvtLZYRpbpPB37BUjD9aWwQZILhEt1a5Qnd5Lj
9KRn1W9zcR5hHfT0mJSwmHRiyuB3RPpEVFR0LFOif6tyLldd6a/K0kusuaX3wl7c
5Eh6EGDPhz+VuVjxYmKM0YjXo/Crei5EOyr/wU9ctsfbqsU3yWzrnzyi1MMa45Cu
G+P50VcFQc7v0mKs87VB7BRH/u/CgWassVcfOIi5Q5TZXGi5Uo3BnwdTCybmjO6G
icTyGQ7IJsy/2lNYDAMgVXo6xGCPvc0oC/tZuws6j8rcZ4tH605lvK7ynu5UbBxp
QoBtv8JSz3SjKcxxBkV03h5aNQKo9TnimkZVLa30HnXWLMOb2fb2IZL7XRuLzAei
w+12XgXo30uLnAi7ajJqLWcXKfv1wNuBFIlDuMuu0byHmvt7vkbxZt3kX3izVoqx
2wTxKoRqJNU8qA3Z+bTSmsJ1CqsCl1Zf70t7JJARKtETyVxk+8sxWe/28943IkET
h29KF9UfW6Q2fogywQkjRCLKY1NZUwNRnXRx+uyBlxwBFiouwzdBgD9ZGNffaGO6
3kj/WINJkdNaCjav/hf24wNISagmWC0SG2IAcb8ieBgg93mFwVGmgazbJ6+OrJ6l
vu/JeWiitTxRZyu0yB1m7Ol63lh55XpKxfWvoBsV3pjz7tPotNxpnj3sacwossHn
N1MgRwq6gDcEnCCt/Mccacvi9C46VZXtxK14LbvSkKW2oZztF136C70lrHTRw/FI
1dWfJ7PL2SS2eDqjrBSSjn0tAjzWW7TFAjjBS99c1xR3nKpyPKk3rcNKvF3gfCDU
756SVp6MhkPdTmAni0pa1+ZNAVKdlxi9LTv3oEOGbO8ScO5rV2U3QN3gpU2t6CGs
vidXx9GVq36n1FrUGClt/WqruHN85ntBTgas/FN5lEmi0wJHg0ibsEgYsbOMScmh
MTM87Kn61NLel1a+pB8oAyn6i+BisqOK6HkN7uHNRu+BM3kVGzHVSEke6Wo5x3t8
/rM003D8IyC6ZHlcYRGXUX2Ve1F0HFYvCPXZrQQwSLtp8xLJmqy/NcraWAP3xrmu
wyPXOpDxPDEmrCLzjlhogV84N6Uj3hGpUS2YJm0GEYIYWka895WdxteyEqmAX6A7
hmo2gcj4YXC3K5VxX7B7iJdCPEw3EPp7ruk8FuCQBH/Ye1F9Q1bk1kQKpkfLwDBF
XSYXQUKk17KEsoRF159N5r9qoBXpE2K3tyoBMXdE16b6iK+IjmkwJ1ewieBQ57I4
zEtZ7cKmV/pA5Ltjfw1uiqEZP/7Qp9P4jqCtuEvSRQwxOUp3zhBbu6BPkoHZ0JBS
BAb/tqzTw4sJioga2fTzIw7AhGX9klokUR9sAT7zkuRzeESO3m0BdHyDL7e1OtaR
UuSrn75zNuNjt7zbXVnuQV7sX9439NEMbBy3JEH1O9x/WJDJoRZTqW1JXM1sG8GP
UdSzE189O7tQJwjDTj+03xjYSVsLymXtldz7j7C1hAsN9el/T2ARDM4vHeIuFF8T
2CVhJ1+wTvDc0bX/faxVyv5EV+WDifvL/Wu3gxH76ylSHsAydCeJQfI+U/yWx2wO
nZBn9c+EiG69LujTDL7ou2xHhpqFbxxEbjMgxMVd1JkfVmXa/ZkkDKpywWfgP1gK
OHLJoLXClNhSUTT4MGBvqGMbvCL9bRAYxGDQ2PdWCNwIC3XQ9332mozsIdycQIiW
F3CCE0W2wCf+ueGZfR0L9DA1Qo0XtvQzwyxa3WnoCEQdbdBFgr0NMZvJFDX7yppB
yvK2gkLHlW+Vme4SFMlQTU0KXP1ubAB44pPL0PxD8E523c6rY9zunb9tODT11Msa
ZqS8IQL7TP6pBzkO2acU3w1jhf0WuEx3wAqzsbpLAHkkTf/nnn1dS2SZnZLCRUh8
r15RJiHMxkInT2i7ltnXBQAg1iXl52GA8TQqgnyivq/B6Adj8HcAkEMW72CIm7qG
Ht6Kr6mdCvS6VNFxvueIYkuQQzSn93keeBMD4SsV7gdQfT5p7ZsVdYBea51Q+Jnx
DCI1eSYcDNmUy3dRa80McMOvjVYhq0bqnvrxPe3QR6sxBbar947IOD+1q1OHuMCB
aEgqujlVAfSqVq0HFYWpOnvczaSDyHIcm3JjffA/seEVB0SC3kE6m9DERO3hRcr+
hawnTyyKR+ubkRMGxH554yf2DhEjc5mYzqHhZWWW1fX4yIFBm7wAc0gRx5/P7gci
B00qSROxUazz2laY0ATWfsVgG7NteQfkI+Rnui95vUtHoWcFiFXeqUJ4Mv3fku8w
IOmVl7W89wd43aiUyut6T6dTXgjWXyuFxMvSCrkbUaA0B2Um1/IVAvEy3T3TUG52
dHg06NyCN/YLIQ7UvRBMs/irqa9p+NLkAHDHOThMzYI4EMdjXrifgwiwnxEV9y10
ILyIBDDCaFoa2w0BJFf+DrNTHVMT40D6/Vc9MFwhr9HATRutDmuihmpZtLqjSjXu
xsDgK+jD1zEfzVDUMX+QQoV+gZdhBgMusvZYQX3wB5Fj6eeNv/l99jDCKcuhxBnL
ViQR3EpS1T3wgEtvaWwUUODLNf0QIgsVovF3qiUUEfGixH5AcCrU0fhzxIpyw2m2
bCv+kNVYXgieb83sxuDUyw2tCRReRX4wCM6c6spBwjGf99saKNzF8B4o9547pVsy
KBrBIeOvPx+PK82ll24XAc/P80rqEAcAYjcdF1/vvcVgzTDC20+ZhUgleyK3ICwH
c2P0YmwN7/kGFa2r6W8P0RnH72cU+uAzHfgxUQ1VinmyerG4L0XPT+GV6+Qa5z31
+sQ+B5kj3grGxzqhDha7zQessimjogLkdschbM06FmOs6Q3HGS6Qap+1jY2dMNqD
i8NbOO0ImUrkGhz2FAcbu3zcT/RC2Cw1RrGdrpt6F5DN8Qj+AglHvbxeDbGyb1ka
MSnUMZVC7Z+Cagcpxj3hyQdeJrshmFJH7oMPOIIY7qUAWqFEIhFjehrhJx82pyhp
pmseKnhInASdzgQmVv/OB3OkBjYkybvIyekjgjTzF3RMw1gKHC5W+rfFOz4B8ndE
7M8s79AU/KvnQrvB9TVwaIMMQDMHZdPXkILmGYsqw0Ht3c0FlN0sTV7TvOCkkqod
/tWOhLO2CTF/86IYEziuQ6m+Nc+bPZ15rZ0RpHHKUXdTASjcPD87kWRtvki9cpJa
H8uxQ+Opzkuwr5klGBi8w8iqSf1X3bvmBU3v3Gt9bpS/5ZlaYz1QwbKVJzk5QCan
khzzBgGQRJyjv6tJU003A35hyIWgEwxLqWy8gpfjD7d0nDtWYfFom+NaLs1MZKE9
q9UlglcILY2S48C73tc/sB6WpGv4e3pMrmrudLTKMhEwSOLaCdtJnQOjPy70f5xj
fp23RvIIHCn7DRpgCRdeNZAGqv/4k9LjA5bqBHPJrukg+A/pWrmYaWPcfSAcve4V
qe+YdKx74ty1ZVQHuCMN+agUopySol27p0va5JnGouR7mYFhmZN8IkwKwWZ2iIqJ
AnfT1gk64Xlj7eA2wj5lYQ7hZmlzKcJJD6I2x2aryXRyPDLsE3tu/MAvrT4WexB8
rNItcR+M0zBaDqJu9AgjJf1RTnM84fdg2WyhHhOICrC0XPNJ4SnOFIq0ei72AwUc
EB/4zG9C5lRblxIJsPTrhE8q2tBVDdQoFpn8MQiS9ULngS3pnaJkXvbfapQgG5uL
kTDg3ogigHRrh9/9lB0adX7RbFnO8zYORronpvI8c7+E1KA8b4ZD+bq9NehZpmWk
t9tKPr5KTM+4aHhFxTriNdJ3xcB/K6+EerGI0F1SqPmmhoPP0ng1cXe7+eUwJ5va
PRYWA4xY2uW5AXiNWj910DaXehLjgzh3UVLGvCebm+uuE44sg+rUMlUvJIAYq/SC
mfWq7eTFhw7P7j602HF45WDPzQkK1QeNxffajwSWuHLspbPw+as/rX9jr6A6mJWq
wgx/+twatVOI7f5CQcssnNjkxNTEwXExFqYm/5Xmwddfu2jCQoAzOay4xF7noKyR
ak/PEYT/mGJGA+Ln/k7OHIWrNAWIxJOKjV4zMmCUSwGyeUfYoeEASe1OWIY5LJnL
9OVpOkx4rgibOfeweSIpXPtqLXNvTFVW7XRiy74U8T8H+E4GPZ73IK06/4dAFlzl
j8DBGKPzazlzo/xfyFyIrywHaQJKoU7gpLMf+LS4ri0stKiujBMRMCIbi5mKvu5P
mo8FpE15e5D98NM970OeCgh4MlAiPMLdKXOQL3xtFZcPRT7bQ10JURSY99nmYHZK
EU3ZNy1DvbhP4JQLRd/CMID500/QYlT+hgJtLSqL5f/t0QEAOorehh0VprPwzLzo
+qnmUkFhC991vkzAPxZ/l1eCSBk94YjkoDg0Yv+xB7KYlG24N7tK7xBGW5Hs3b+W
Ac8R4i2/Pk+3wMAYQ99chZ3OMYLEUysZno6EzsOIT6SDAajpNQCk3ozQb2ZSmcV2
DCwmxENt39NMSfO6SpF+WgKhWZJgx5vEppY1koQSsEP4cAQku1fAaB5YJglvJTW1
JgWAX9RQON4Kb2bYm+CC+UfAZH3PbWVetZiuT8euGQ1yYrB3H0lr/E55YU7NASQe
/5sinpm+s5nc6S4Q6MKHa6yq2rREy17Q5ipwetKcQ1B0tUTHnFJhi9ewIlNxPsiV
+sQM9Y7W+tfHpXbPsY35mWXX1TZ+tibTJhoQ1l/e4wNoia0OQ6h14xr9L9MCMirN
CpvKkic4FxqZuD3y4JtvNn3Ze9V+TROlCDG1cLFS4Tf8xDsmXqGzXmuCD1NWbQFf
YLAIHbU+O6NwQUJOuKB/+PBJzRSn8bHN560mpSLu6Qvsp+noHgUtQG5gymjVY5lk
Sd0CD67PUn2zRHRUMX/9JrRRuhkW9K7z8ZjddmaDGJG/7Y3WtgdJnSRNueABjtxP
LE+iRRVOogDOfyE7wJlWu0gaBBH4gLQTB6lwj2ot5HL4s9Kd/rreNfAPQfkO4M9H
Vo351KF38yHjg5m3e7IiTfJevtB2GBdt4xsMU7Gfmyf6SRWgGmBMDw/SYS05WGx0
OKAY5gKEus8y+DkFcxjVzO8AfNUKyTcSlkQI7YPUVnWMDBbNQ4veNsA1qIY5TBAv
MfQlxL4oW9IbZ1FM8z2Af3fq4CnvzPIu6WRFNjrG4NZwdJO9nMOIwnQKy7Kpoxjn
RFqr9KkR1TIKVTAa8vYN5SssfaFI6MKer0eKb77Hl1lrHeqvigy7QkaHEL2Rrgrz
1hiRWhH47385isOUXXKvil8tmmEAJrOMNaiLybHg04rpfqFThjva1XH00L2Ikf2Q
FHUEZsGfwN0y5t7G8iCqV7U42KcV2ZAARFJKXTSiGRYP3SFacr4YUTcP1JGRPkXv
NsyvURurDJNhM+KNR1jh0XtyLpZQ98S4f57urzF+G2ePMLuH+3hK7t6O1biB+KWr
D/LmTtyQaX3jPQ81o6Ra7jXK1YAGInrO+hBX+aDU32nQbMDQ8eWXK9CR1Uj2LpEv
SyidT1crM8NDydzwPwKGeLWRRQjTI72fpFGgszD9YCIYB9oNRriHq/91A55tHadW
sAIX+AAPdPjMAAroofcx1/69xqM2iLyjvKanSxjinGTKuH9UrPl/R65xvaVzeKNE
uNioxGktYRzGSCOkAgLw0q8/uMy3lohFVrZD7O8J+rkdJoKmJ3t0zxq2Ws1u2ejh
EMouz3gOcxLFPf01mLblz3q4O9F7+Ib8bfhEF/NOjDa3XcDI4Jr1ZJ+WyHlDRKxW
etjp+tH92KeDkSWoV1tifhKwKuzUWPP6xOtRAVp4KcF4gCJk44pRVfdBnJVnrzHi
LbCu82t1bJdXtYOev00ugzkeN8oJ/QYpaCp7SJqN2p+N+MRZFumPlvT1mfaata+t
zqP1wKZ5LoLl/nRTP0KZ4zYiTTk3qyDsEEqRgcnZCwP/2YiaX05RkuyhdxWE7o6C
/f5pSX4roQ7Yk9tfbMJi7K4CU4iVhDLNl1c983Jzz/9G1SPpR3cfDfDwtx+D6CDg
vjWxAAEVmCP6lARDVk7qA7vFfY0jtoGO2jfovq2g/g3X0pxQbd/jUyuCinjZmS/M
GPXXXyQvG6O6MUYxuPpu2xVbKUDsyUcI3chzt2Ob+tAy4o9rNgI3Hzl6J0+DDa93
QasC8K4sne/wjqso3Lg36GyDrq770pFq0UImCnUb+dTmQbaAxObvlX+gz2+v9VKl
k7PUQ0XagjTH0xWn1WtJ+RCpXX+cL50GeEKKTuT34OG5I2HA9WPGYbTAnmhtfROe
Ze8ihoIOkQQL0g0+Mx9XeMlosqp9bpCEtua2UazZg/9u7YY4RyqIGPqgBrH86y0Y
GlhCX33/sw1vq2rKpRYQt/uEamylGJhx/4VS2p1MoU3c9zQpKo1KPsm1nV+inFnl
zqM7csv3awwB8heGgbF93r3lW7FTYVLiZGiTHMO25Ea2P+Ldfl3Mm2MciEwvwnJh
XlY7yso46AkkwO+/VeVx5m0CJcpZxYS8USdQqvB987losFNtBxQxIG8Rno36tpkz
9J/aD60cMb40AFs0KR3tJIwX8B81rYqYGTtlykt9U4HaiWcF/htXzgDQKEcsxy9I
XxjDXyUWwoNXRpw5Yvmr2bqnqj952w1vtXGJ9QpX0dYAAKnXto00Pec+hbotQ2SW
khWVT3Ag1bof4eQIXZPfNSC5IS8tjgJWyqRWj9AaNCGzOsTO1LbYsgdkU+DY+zQ3
zaFNieG5v/zqsoZNfXWWhe6/uGpsuZPz+RUtXneAvQlTXzx0sqiKA2gjjc6nZq5Z
rJgNTmNJBDQkdiiSzjF9+0Rwqcrtx1ZYDpqZdw2bWSZ5AMdZw7OtnMNsDQo2jmaC
iGFGhyBG8SAK6cY/O0MvRJG/sR2FK4hkNd0lJyCUmBkR7Xw3PwjD1Q3wsQU/sWI8
vmtamDXFQ9TRBEm4yAM+gkiK9K4Z1CcM+W1kx47tRfZP34/svfZtWPBxsOdlym02
LwouhbPsLkNJXuWR/HKEC1guZlSF9cNktTUuGrA/zEuiDQX2+jRwFpsejKPqW1dp
x+af+EAA5J0XIxVoEjQaKelhetAZrszGss2Ao7oxoP4OdRS8E2IGhJMBV15Ebr/y
6Ru2lFqINHOm9ZjxCPs3af1HoLNgQpEb0vQSvRVSuo7cd84ZEs/aIsYAATLKRfcL
zaJPu4LbbiCbwEYNQMBK1ZwKiIzOqejwBLVIapIyKpLwj+SsItZDpjPYygQbRv7J
pIukv5Tug/bjdy9PYI1HlmsI+BFVnpXd4C+Kjhv0sCxzMYi7C/kszHobLQ3e9lq7
BVa3Kal3LjqSNKxKGR8ClWM23RvUal6jY2LhAZrcF8CntYpt48MNId5E3qQ7+DWB
RWHeokZpmcm0Fd2ujZSNledoqztsS81dQYcDaP7gCnP3Br4UtLdiKhdSj/VE+PeX
0Xz82aPwzLO1j0Qeliu+useZJJqW+6BfKMkGCaupcHHYx/3afRMBFzeQeF09ADiX
0Nj0cg/y+SoQ4evHyo451HP1KLilgkrLh6Tho7eivSg8uoFXickB7IfCaUA+bDbY
7I4oDaRWPfEbNnxMJrySpGYrTQwfOdYX/3NTjPtuZkcZwhWhyCaWiOpjHF8X8UCE
TD0rCw4S3xaJOlqzBYe2UQL1tVmfxE0cwZNw4+TSSCTSTF6TJG2CPaLBfkHufDKd
MEvQqcKus/QdxBg64FDb0Q9U6Bw6r0iP3x/bToa012lU4/kGHSusFw0nhV4Jrmkg
NZJXJJXi/dqI9uotf6xUS9sAg6kd7AtMJRxlxsjMKbmMFZ+xRW55JM+jFbw/XS60
6cmWa9uSVI/eOS0G8QymnC9YObRoAGh8VHQ/KP8vu1Zt7Omrfz2nwOXnEuawz9Ds
UQclEF8wLZyiaCZObXfBQwgpGxVUHXJpcBdGVAs06/WbX5NWwjskEejfKwESH6xC
Ze0PgnqIZFybQ57c+Z98TRpGz+ta6G8UuM4Gpw7nAzNTerLrmEbDw43SBhGciKoG
DhW10jqvlZww3Wgqut7xQxGqqdYRkcBTQUenOwX2/T3KzB1U3y3pST1casf6aDKR
6GDq3N4+j/hj1NYKsxVN91Xs4u85JyG54r/wM8FOGnLINSHtIYkuWWWkMMnFiSEb
p4hlcCuGkIrWq0J7MqXzl2bVpWbxUrv/jxX7HEY8Sia0tOxweZndirEEmbPQCQOQ
NNwHBXZNUKxzmy7qPGzP1nYujIRYP6r4TMyzFHQ7Zty1uURT1STxAcwHTfxMUb2L
H043o3/mDAlMCk9blQjLGyJkxWr33EngC3972LQeMJ8xA3aRbjAlBg7cg58l/76s
rIEkJHF6tfvxMY/eDQ/iTbSNay+wYUFcx+R0AEb/WX8HWBF14IpXG5wteTemUj2H
31cPbD3/FM0WuwIDszZTmL2DPOT5rB6g7a33lCX1USLfp1QaaxPOy4RMGLIQCYkr
m3M/YUeYGLpHwfWPKPr24aucNOOAqRqkBqKiTsCBP9QJlHJXX0KMuXBhbbSx952F
NULA+os+JzW/UVjEMJnJmm1fLVxRT4lrnJpoKVjnegL8B2D+scVQmiqII3NyGqB+
GOIhVkBQ/3MGPXguIDXFWmPgx76KmG86nBkF4qkl3GiKHYBHhVHhWI3qjMrSl4IU
BWysud9LxPNYWbFFfmipo2Z9bfAU2qzdqzu35CwaRZh2hejS5qtcVqQ3UiJybw7z
ovjujpPO2wytTVSUNJH7ywPMfYbBoMlK/Gq5InN9EUTwpOQEBK5TINdgV24JAZI1
TJIo4IIAXU69HiWFI3WcU0URsj7+dDvxTPh/R9OFCHCJHecspr0xX9zYPZ5hBy5h
7+8XxOsD7gd+7n2C8VHgZ1jYtqZrsLSdETN3vqdXeYYkLfTVoVMbjt/vp0mNhk3T
0QrvA/y9pdQQwn+uB2TpcQx3xHM6kRzp1pTMASxVy1RW8bTH/zcoWcmb1SVR0byR
EVxJ/PUeLp9kkneFi++kntM4jiG0QXpAcIBx6pNExpt1H9ABD00zdAZ+hJBTyER9
wfWKFvMIczr3ogwXizIsSsJ/q/zq6ql+dZpydyBWTy948hFVTqLwJY1vsoppowk3
WesjCKFfd4T1+/L+jdCnT1Fa6n+ZyOEytgQ05HwP07NWS+sONOZUKLae/nL9o/RL
cAPM8yXgscCnZ33Ze15O/YtQAz+VovvUXCVbh2AxCJIo/3GGJ17oZgACsv0nuBg9
XcMYY0ImlOFtAhP9naOYP2zO2NWP8EG2IPKUlKEIlbTYiSkZptk9p7KxdFeXV8RU
nuXzuO5uFbNOEGe32LZWQ1zVJOOf1PoXR3OyHRQI51/uKqb9Z/bZSMRnEbCJ6C1v
sjPbuKSkmebFWxNo4YIcanIPV/to6rHNf2Mu7Mrb+7LDCbDKBrVUCKDm//iN6bGd
W0T1OnpnPUy+R0FunBSW+swg1wlZDLZ3Q44TWzQYgjW7i+J8OnGm8IjyIgtMb/zz
eKpZfLOR+wZSn4WgMbjdjrFdO40hnqywiiN7X6YamV/DdAkW5RMMvWE4SR5uX/AY
3LNmdZevFjLLhdAUwAjOs+QyRNR9uyOc6lDw1smXEaMP0u79FsvEnrm9gBYXClI2
JYeVlnHr2QQeRrwQEhSuYTKUcE/ENVgtlHdNCt54kXKpT49gnB126GaCK7TXjcXp
P+0K44VJTxkxoMieJaNom2qFCus8OBQOcgvyAIxUv8LegrvvlpKyNwp+3fm4sNUm
C4uEZWgB4+t1CB5jiiX47ae/emZHdD8LDFe8Bq3KLYMZWt2SADvHgTDdjRXgEEO/
//pragma protect end_data_block
//pragma protect digest_block
au4zTHcekg/4UTGCCeUEELj1prI=
//pragma protect end_digest_block
//pragma protect end_protected

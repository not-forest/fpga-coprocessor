// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
vODReye7eY99e0dCCSZlaH3kabc//po5yyd6aOg6jbj8xTPAuTeIHK53rAUmSY5OhHVsVho/+xdd
jXFo9KFN6nHxnI8Ctbmx8ZY6fh2PU/Wcl8hciMLPGCKHp8ifg8/hzbRqwsqIDSSgEJQqLyqQsLiK
Tielt6mzySROqLRquFq/pTnHlCrSUuJk31b9ednJbL4cgr9NFtyBX55x0JjMGiCMTdnQdb+2+cAQ
F5fprxQPxMzup5uqI4YUfWJMKxr/sH8B9pW21pPliCEo1jLDIQIqF1pMyCao+GtQ3mQItk3ZkB1n
dT3SRYy1YJ88myFyV/X+D7y2ZPD9DVHVfVVE+w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 15456)
Px7Ce3FhWJr1C3IBdQ1Q8GqDQM3u3mTnL6cVyOAu4h4dGK245rYPb3O+vtqojXT60RFCOAnfpcip
lrDYdRSNBOyoIXYVP1A+W2xHFPB62HiE6GSvFyZ5CCpeMhV/CPQdSH+jLUS5/JVq5Cecw+vPi6pS
XHbvyS8d1lBaNxOeGTUTG2/kKUO08A+qerddn/ubiwLNPKspOkZpU9i9K97ipPmogzIyl9zFpQSm
P4aOxyyCY+ivPI9BgfHoB2whLIL8xzYNptr6KnNbBg7xptlK6CRjikZn/9/7IFA0jDJpvdY+2EtL
xH/PiD4MVD2482yvImPj+EgOg6LnC2eMGrjFw8vjENw94jyBkTERrvaV1PTXjfjB4xGsJEoyt457
9X4iWfST+Gvz0XOHlmGm5s06a3YH7E25rsgYvqEEZZk8t9eITorJ7dzrRLc95AcPk+MzezNS2bA8
b7h/VM7roKP63YUqmLAaG3XKZyYSFg4mthgZo6r74EslgZQgBvFc461kORUWtBwi0qHol7NLGVEQ
SNx29hkHKPj5K2JSstmNcRL/3kojaiGN1YaOABsxZP+yLCr7GpANXoq0MdCXV+qwNijlf+cieAwX
Ceo7iozo2JdntmazYhpQr8zUO79sXvo/oVEXlWIrPDFPZkkv8eUoOGytRKDFRHp/WML1x/9Jxeei
FW41bbJZdUzjFg8mQCEJd15OGH6iqckhCs70jHJeHQ2Wyl+x9paPV1XthKIgGhyecQ3FLsoiat2r
8s4I8nR+1xCiGYLXhGwHoVL93YPZQgsExIzCrzk5lk5s9Frkr1OfVs6toC/9RHJQ1YzW1mC9fy2a
sgedF2C3JQfsQc7RUHZ0QDiUxt3tk/L0ZNkZ+klFzodgUQcoJ99yJw5uE8354pL+nO0Ja6SKwL2I
VsARWj68x3rAcFNfBkSduIHQrgsFhlf/qt+eze2cdeqvAo5nsFmb1LjtB0HIb89WhScxT5sFcH2Y
aGycgbcXQf2pksCw04GiBKhlyuosb+xU+9gm7OuvlEtdAnkHWNvjRkj2XMrSerbrkf7iiWNXG5u3
adlztgCTazXbu1FeZfB9b6sgSoqCiKfCaArNV8QNsSn4M4VXZ1PNi2KnvRJftgazvZZonLqabWh8
Ah2LqnoHIqwLdYbVnXgJuEWEDys1K1QmW4KV01tIkf+JQ2QjNrnR0YanuaEgiiT5bN97yVYNNkri
5Q6YmN3CDDJD2ODBPXUzLvjygozwnJZ7wCup3GODlzIubXTDYzrdynQ+R4Ok2tLaLOE7LhTjklJG
ZwCt1/Hqi8yMucEkZV2y2Zw4wjiLIAK6Rv6QV2TnUXhMDjmLHrUABSPlJn3hBjGXR8htMvj/7v6g
D5jOmO4S4Z9gDcM7DnR9q2hIWsSNH1eNdEInfUGS+OpNpazyw2dKEUP1iPoCM3Y1t/MraX+EEO8O
B2QtDyljckaaqoWzWUi2hhWOJazxmpgy9dmQ18hcwvv7UZLtPsiMhnEK7mz/9LwIhFWrlP+yqwbh
897TX2HPflOwLWXTeeVbdbEEnyQC8Nx4EmstkTMezdy8dyzxY3VbI1xnMb9GXb4H1BM9AuRlqBKz
mkPQa4WxGxrab/SqwfHzTlho04sRomjwre0hSzcb5htb7C1F4/Hf2lbV2PN0AWcPcdWVLF/wlz94
NDTrBJj473g2zy2seQKfKpw645vOprDCXpplIEYgtLzwxn+6oW28LpTGxCnlrzk2Wd1yZFvL14k+
bEf97v+FIQv7LyjuOid3P+wg3icRAfGQHQSJwZJTAKLitOooX4c8M7A67YKMwYVeSqhesQUWplRd
OKgPPa68mPpAZFIsXMP8aeKoezg/x0TFXUk+UCVFvgThPTT0gJrAfLhJEB3jQNCChnxgsZFSArVf
XUaWsBk/ormlqideMEDXEXnuaIwGOxsMOffbPadqyXGjSj5L7zybP1dYO8rP2MqoopTOkTU7wPnh
Vx5Fn622b3sKtdYKUj7DdWLg/nVmbkpqaMRcdezoVw6E+oJWl8WJ/MWHj0i/gYM8hPjxfEsZSwR4
ObZQ/penIHlkqQluKBn28iv64qjq5V70ufAr96jtVhabLpBGRzojEJGaUca9fbRoSe5tCm94coOK
4KKiON+YkMQsqI8vBvFLkU58SMRN2oSmWW/YBM1jBXMYGbcw5vxBJwP6kEGfmNA+yIQl36sf0vqM
9Qdvp4swG3m8hurVCg24XsmtoYG9+iG+g+kvBzVWffeCHMT5hTnKQeCSxwLdVND32sJXUAumyMFu
f001gX6qONFS1jjV/YPef8A0trIUx+xlIYTZAKMAOIfeW0Ah1Zc7Tgpxg3nsKw0/xVZKlt2ORM/w
J9IkaTUc4khT5U1cYBzYezwegAvJF9mLCdQBn9/FQ8HBi/uDtOY2aC/1hD7PI8r+fikMTekZIyWB
as5zRww0FhQ/7Xj/sMCmV7GWtGvxdwar0jy/EMUdoO3AOq29e8FSHd7GMbczi+5A51vFyAF0c83W
qw5/W3EMbNbLVIV+k6iFKKqvUpZDRwNOlXrwUwxKmtiE5EEeIe0a6ZYVcgnyqBydRp1MgNIl3G9I
73wUBarjbPMAeU7IPVyw6TNnE5L5rR8a3NFaeP7W42Aq0g9SAkW9MKDpkiN2gCaoeLQXuRkEjhoQ
8XtT1gY++rBTHWcv0Gp5dYWTGIGXD3h1l09DczqAn6XBOVxM91PdCbot3MgslR6A2cN1LZl8fbUz
WGUN5uO4cHye1s1+AbIQxk3KyqYyuEakc1oEkr4CTAyumjVMV6utJIXdUX0ZEkgow6huDokNARsO
Lg8//NDQ1TKTcgibCmZ6+mTSJ4ky5GOzXpirgNsiq107K9ApuUNW1yg/WqgratJblsHb1zAw6By4
CVtvM5WdeTgFl/EuBda+Eg66wXt+Mu/3V3Qs4PMj3eS173mqmjipxMEe3jRuLdfelQSwo27Bfmjh
BVPDBVpYs0LlWdUFNRnZfqK8q0mC1UsgnG9kLtLm3Q/CTQ7xtZz5l8pd7Hrh6MSLAqqXuukp/BkB
2cKzPp5qgwh4Fz/MU6UE0YAFT5/vXoXty1R3C45R1/txcQw7HUXcNP4y7CL84QjnIFJDQpNq9Irh
X2P8IG0airm0NvLFZ/XDXRBb6wAIoEMR1xHsv9M+m+b+HBx//Qk/6GA3JGaLhEP0IGqos58OV2Ps
yJabP/BaFjJHrRYb6p2Wo9KCN1d61GUqpwZVd8+fv42wRuZFtr50LLggB9bKraxdi+BX7FyeX1Sr
3XsYmDqoYb8F4hUGWHOa50uqbKv/9XomBpoqLWUHiKamM1wu6DPAVcoR66tvl1endTyCLVvGbBeQ
y5SYv7s6zNkVOHr9Uu5saGXhoeXFL7sVAqzHTIEemQvtZFkJhY1cyrej33YqVVc4CxZk6IXFY36O
3CIiz95FJYugll02XAjGkE6GDE0XnDK6Taz79tjB/aRxFvwle8RBcGhEedNoHZDaXhJzzrrPl+D6
2LOudwL24TgbfdN8Pt1vzWq5+mENxuQ6KHzyk9rXy6lJ+ALFdUFeR7Gq8XECCETk6kOx9kW1zq0i
dS4v7ocDnzZq/UJVZk+RHLS22wq5o/e0w/aqAzooX2+b1jkfbEUArivUr5ZqLaVSOrItTsWhOyNC
/qzcFflRI9XDIjhXTQuZuL/LZv3BY+Hi0zBjVj1tBfu3zjjzawlCq6Mr7I6X7KUCfOyWbOy+y5Hq
cBB4cyZTG+t+SPkzwuazT+F00QtgfmnZHj2XaSfunMpr35qYWftLz/cr8UhburojIUf1v+RJMCuw
VhPPcCLTXSujY2qHtcvsUGUrUleXCzA6v3VqyM55/XVfC/c3TpbdKPuJKE/bzJ4cmaxTcd8+/pQi
7el2RPmgjQQ87kvsbKClUlK93lWrYrs+WKI/ObLhm8W/Z58JtcL7zhMYIjyK39D+Vf7pxcP26/z6
JC8OQo/6fneZHHMNg6+hsnPCmZWQFh7SaLn/6c4J6UWHDQ9BEZMsdV9ttDgg7JjLo46PWPl3hSSG
dpBxBPE8Rhh/meBKbePGor6p9NFQXssphciUmrGQL6uYCS2xz2BHbIvBMN4ffQxI2sqjkfrLj1bF
g8/I7HmjCCPm+L0cqw2UmI5FUWA0jbJ6DBJC4d/n7e1iWKxCbkAQNWbPQehfGhyTwVoWj4G7yzlr
SnzUspO11Vmtmf1Svdj8aFTuc6TE9v7DDLbgbaGuzGOQK2egiRswBUM2x4WhRKeLGV6iuu3s2zx8
H0XwWXKdBIzmU51K1dmljv9CNTQ3sv5+cK3637YJADuYAz1uvr6KLZBPHrhPka+FwcEWCbYRR0Ic
O6I2gvE6+JtpzTdBtyevcqCT+8DUSFiKD4pbqx5gbNQSqZ75AL9ZR3cPLwPDdddC90Hykceot6b3
RzoePKoGym22KtvHC/+qjAg+3mQTEAA6WoVH1nLEaX3+sH/piBMFgQOxcM1aLlZQr7OGCLVLM1ud
yV6EVnNWVnoAiv0BwFym5DYIFbvse7mmXvcxr+GZFA4r8EEki0Dk62mMt9v0iHE36tsXVqvF+79u
RBzKkd8EHki5D7X4UFQm49WHppz0rfNNpRfGl/U4TRiBs7YcGjJte0lrLGaxANBwJrlLPF1Z2EtR
Ebd3hxTnAaRNPecge9JdZSbHdvmQXh4riLEctrOCA/h5/otUc6Eu3c+I3tppEd4/3xqth3wwHe4C
Y2A0x4Ao/in4+v3or8D7Ip/EybXNYXDNLn+ykVwlaztrMp7dKvVIVShL9Niv5ndii88qX8VxjIZv
rA1iUuOkxvEckm4V7CRwYVSjhGQJWzSO0z+t1Z5kNhoLCNpu0zyeO+TBJK/d+U8OxhUjFHqhOVrS
7UB1hxEpsXAntJ8EHDLBj9LXyKph08Ma2W6BZrgnkE/OlX0/7eHrsCzUVrz6HSLMRyDycNh8Ycrt
PLxsdlGE2pEr0CiCjiup3XXCvf1T1nSYHx0O9zM7qlfi3kAWCW+hDCscz85zloFGBd782/+veZyz
ktnNFtMta6uTFJIQt3J+ItK4fd4DgVaVAhVeksEgVzWf6TtkX7LF3nm71JUvQ7MmBa8ICbVKU0mq
m8OQrYk/Azem+DrgxRaRkL0L6asmyidCwDNJcQfrzlMDHuNAF70icuiAIiR7rL+sK6HPvRwhQeAe
/Gn+45xfhAP+GsuLMCy89duHKhI/wBKp+3zvYPxlC1nKXuCLuOdrxGhBBbFTyv58/WHtCH4AEmRj
Rt0K33sc8WApjtozOd67tQDgvyCNgLePtoPBH2KnttD1EZa0CAEbFZh9dQ5/sdiAdToU6v3y0NKY
qSwVcgeST+heTOApmjdlp8wlBLDMkyzMGCNCU9/z7PbvgZ7GnJrl43haV3T37H4zyZHJhl2JiiPS
Qb8fIwelDTUFBN4T/Fq9YfjsfJEqZRhCXYOMCAJ27hGxSrZEQlSROSV6EuDUcGJCnPBxyn8nMFHi
jIgxPtdatCg6PixAbnhvRhz+LmRLh8RNhOCeSFDbhVQh2X02namp002YRecgY9EoyR++d1/q5UEG
VRAGEpKXf9nzSLRwSFOuk9TYRmLAnR+wgKn+FhnzZUgaMMaviTkv4o765q4owc7k8PnkU4XMJOii
LHuMhPYV0MPcnxA2DWQRbROgcQdTqeesK7uxa0R2m2nOeBNyOp3vH70SK2e/MKSP4n99jbLPde1A
naIJ0lB2eSlLERiUebXL6msJ8NpIi1UdfW14EvRydOl8Z4fjYAQiXuHaGvf9kHpDbEm0yPGZ5gf4
Xhf5OCj54ZyXh+YKAv36sOja6WGA3umDfyuBP3zCQrVvHEEWu/WMSBOmSJEmarQifyKZ2p+Kv6eA
0iX0m0reRB9i2+YZhUfrkXSOL6DxjI5NQOoRrKfAuJyayXkx25g9+wXTuFIRsH8GvhKivGcX8izZ
gdxZJF2RXNVE7fu00N0qo/d3FTO03MutRUc2KCn4P3o/XNuBwoCS6/0hf0LodxIghx1TjLA4hQY2
KJXDXpsKcb5GJ8El6uJS9tKJTEnzgQqLCUeoztdZ4+Yaqlo/7Ryf7DN9Ua2Zi+blURwfVqkK9vm7
XtNPCfbG/T43mwFD104ivcaQZbxb/DNrYXrTN3PGLgqn5L9kOjo7VJOCvZaZ0OjHEIXOOeSwBwAo
dl8vyYEyBAXSI5VCqcijTKNjOvIgQXgauyFdYxIL6c0tGGctvxLnwTEQL0WNtCq4sKNP+7PY9G7G
LuXBiPylbeHecviAY1IiNTdWe2uLqLrj13VB4o2PuVWNDJ+asnWJ4W028wkma0aACDwXiUhQA3uG
Smrhabf2AUD7QA9BsfveVB4PM+zkL5y7YvegzcJLUeCukrCNOsEYxf6+vf4WyFG7uPa8buj7j54p
qYCSpQ6+O+yFmGmB/Ts3WcGg7fz5JQPuqvZl5D+FjhunhxX1vyO3UK0LtV0r9TdLaZzIpL7Xth2i
jYShO8tFDWUxD6vfB7cKMSLF4LOybVbv8QOja+G4kSyrIpCMgQ+XBwJq15oGAllHyJ/Id/rQqg4J
UkHpPv+kZBx0FCXQotScM9Sn1Fr+9QLm1injQweK+K0ibf4GyTGFjQ8+8Q8EfJnkPVTvTFzMa3N3
ZSbX7bGINFW79r6HqgcH4PCtirQ3PxbcD8yhRKvhPx2qlGEeJPOe8J7Km7bGR62iNRjVws6VVIL9
94xcfvsALnhOapAf8HYh/qWQWEomTNHI5IEATZGDClExGIYRVcCIcJpzAcL7Jg57JqC0Q2fOgDgF
rZtKQLUKkSz1d+fSq/CEQekGilaWHumL9YWH9iDcKFJ3rVJ2tZdrWftT4cpPQ6oJu90EgrQzAgRb
lFbp+N1yL0M5ZNnmOPNv0hNYVY5GHy2zhb7tFog/OeHrRvvRuX3TlWF7/PGnoxUK6Kvwl/CYsvAK
hAfIMnJmbkqXx2rbsEUjUKXIOsmVWwh/lugsghuRdi6zPLyWP+egkDNEPBZrHhjllw9RMYbsVp52
+3YzEj0ru8TZjIXZWf1EMEZMgFiWbC0bt2Wj2lULDqSfnGpB5lX6SfDiWsdlC0eXgZGBzyy5sHcd
YrHn2PqtzCRkUbSCdptkidcIGyfznnmxq5bzp8qIt6FyG8AM78ebQL+D9lnmj2EdS20LTJgTCTbv
CIEzgS//1H15BhJhm6axwSuJee53TOSEepsmLOIl6HnUuUyqZ+lE0KOo/012h4yI8ekKDK9azC/M
6+Cq99B2dcHswARvYR4RSvcITLdxeJV6mnAF5vsZ3S4Rs8Ri3aTyZtpwqhcpqaSXK2v5A+bYctBN
LOYuZbJ6I+MEtB6JljCi2dKOZPjhlGb4f2o2pco22vOHKjzY+c5QYsUtbImKNCstfTKhUtCShrLy
2V0v0dxsF4L09EdI0dW4tS+UFhFfNMhsbivlraI3MnFjVZdq7+/wMId/Sur7BeGwsQ4ns1OTp3GD
8YgLEbZ1AU3Q2twXuw1Vg8VVx7eWnqMGic+/twggk+ztIeqYfxQyaX/sjzq1rlmFJc8AmfyUQYmy
CDoMbWpB2ef8OAtdl6+gNoOLYhmw3xcFXZtGkbo7TQnnHMjDTyDbaU3VF1yMcmJp3ic9sbytQV5A
5hxMO8iVC9DzKbNZ+ZWS7ELE7mmn1hYIa5n1geGivUbLQzggKWbcrqt8yn72mU+XbZqfGVMPs77e
yGZUc+QC/BoPzZQVPQlvmutWOb4ziknNpC3LpVvzuF2NJj6eAnCHpd2rRimctdm0iG9/kkEYHjAY
v5FfGQgv23kfwndgRB662S4DOf8sE8inPBzd2e1Ti5bmLZVKgbkkajoRKjkTMXqXRNDyT4RsiI5r
X0KTd9vIh1Ehw6zxGNaoX2q07tgGqHXczJz7Bm8oYZrBqp/EQQ2pZkzrAMnV5h55ooR0kiL2K6PM
qIaXgayXSedhsjuSaKRvVqxEgObsknz2ebD/MKw7C1vR16cpnXiGq2Nl6McyY16FoV39jnXddj+8
G0ER/T7FhxOOeixV5pqgqIUKols46CF59DVaRkTzcc8wqWJCZZguQdLM5KoxH4dZXqzPuN9BkAyv
4j0adKpSeVw0I8eTZgBxisFeZs1y6T0NVBnhsftev+RQe+HyGIfCZOS6aUtP1cDUMGXdcaVT9ndn
HK7zYqqLgBHT9MrbLr7rDAhYzVMwg29ZqCDJD+LNo8P5gcUG4kj4kuQXI7wnSttES9pIyInHkIZu
3mpQvqJ7X9FsO7uCDiIi/V42Q+K9dq78HivyQVBnd5ksfNV+YmcnAJOUpI1x/jYG5BxYSBMLRyDV
ITfToAlpk93gMaxPP/JA+PITDdrnLctyqQCqC25gHyLFIA+fbH4Ad/I+0N954t3ejmQZw4aEFf6r
/dYNWtnpSxuYyEfVzR1FO+F1XrxlNB8f8WA4Ym23QMFkIcKYjdi4pwNxZ4i+wufIezDsyfG37tI6
EIv6mPlRFQQtyn7zUKpxU1ritbdGtR4dbX+5xAos7gg0eeYlS2lL3+ISLuah+/rHIg2/wZwiKAK8
QibuL+EGrUhafu0SIehLjUY7T3YAEun3toyS7QCu/BlXu8x1x6YIbesBxIISbzFCw4A9nFThwRr1
wOyc40N1tdlpiAso4he9qyY+/BxJhH+RHbKu6wXHbjFRS01TzemsVbGYIxQD030Ci1cjfvn2wh8J
ZMbR0gKoS+dxurh8ApU5csDu1VPtjSI8+tfvgiPB2LAVHZQhAdPBXbSvKpyPG3olZumHA/KJXwG6
q8Ec11GVJyERqEaWdB7gZ58GyZWjUfkMJnlkErWFWoz/EsGDHA6IApwQ3pFainlccOx/VZutpvQ5
ppBrBsZCc9U6TlyV/0gGYHQWMZOqlmiOCHhhSy/RrJSo+9UFdoIUcPdpkkLSBkbj9Xn9hbDR9eNI
Oe4JF5ehigQFv8V6VD8tEaVj/dyVMQxNH2KageqfGGK/jrTTfJ2X880ZkFl3DOdjZAZpKoAFohtj
P+YTuDadrVqHUM8D/fCYE4696T4VfQAiJt9dgRv1ElEtbs8ckkFnexYKAoRztZ9WekNDMdPOYb+8
y73sY671sUPmG4EIQoOlXTqeEsRqpbnez/PlV1c+yy3Do2pKQ2l7aIQ+yHb6wvUTSeIXfVdkQpYj
j0HiHydZuU5VP/Sn8goaoAAKrxTpVa+8uGhhngsKyXeP80WSmd08o1ZEGbkIHaDzuzOpgklviMSr
5UsVzXdboGeMJV7WebvQDQ37lLcZt/T23lQ8NcLSVs6xQv0R5F3x3ZRJqJpGxMK3MBQjmrsypbqu
ImZhOIPlWKaqGQwTBvZKepyDtyxKVVC2watVB40CzpdhOPqa0yo6bGfBuYZvA+/6qhkGiWvT63Bl
ARHur8x2/CCXKBVdaoPgqrZ7rzvTccijNTxsw3b0gL3n7vNi0Ai+ZuQwg8eqNlbVV9EqWbhKJ6DB
a+uRSpqMrqUpgupsncfFNsGgjss3HwzYz8qRHZJBonGVxJVJH2qPc1tPfl5y/HyH4CmL032iGWcC
dqko4OMsv+d48QvO4+JmYx0MkDOnLed8LNrn10QCsmh8PAcoAJQ452xXGRbc3X7MQeh5y1fBfIu4
Zn2Y6kk1h25vca/hPWAJvNvnPbgHZgzad36tiqIKyk3w2Q8zHbiacNfTww0pRHIDjQYT8xKgWnSC
kSXGS+AbHuakhVDxOfaO5j7FnJt0NYrOgHfQ2Jpfcqbe6uBVqnDznNcey9UEfE3MangESbWfKAMY
NlFkPsbrUpDFIvtUYMcMhum0daEddf9CV75PFqcxtyzUcEStwa2g47KvtjbCqfjJh7oKJU93IlHV
MnnL+qTeaVfV/Kh4HBodvptR1hUbZxQyC1Zh3QdgyZ5zNV0JAB9mX/rJhwHr0880L6jBBXWzQynj
1wQlfA0vSrp6KlB5myuoiODoCeZpArUrmPmBnaI5gYV5cIKWzrxbhqyOpr3Hslwl7g6O99oi4DnI
9lRb3uQxJ0xUbjpxOA3aFd6710JXMGHS3vkM59vUICQ68jOlEeM+CUesIBO0ti6qeGopi6g0nTca
6Am5IyVTKHzHeL1eSo/8uWXC8/hwXUVyeQdIxcRYqFBM5oybcirGZmQ3eLmZt6Un1x9xvDT7zWuX
ODN4EtM9Pokkub+b28xyOHL4Zd+3iWhwy3/T09z6PQgXUMPLKvQqQmcWrwiv43BdMSlFo8p0OTPq
CWmFsToiVi2B1F+StsGrLFf0N/LC1f5rxbxBanxqBUOC5+eTZ6wairrW3es6fJSCcDROek88deZf
TJmoVwVm/4FHO9jdayXT3N4qaNjRJ3dRioBzCtbuTDrQtdXKjeKuEU0uNgSUvipwU11ueQG8Yw+q
eU1DUPUW19Ecu49QVhGmlOKLt4mRtWPdhB8b0GwohCjUll5NO4d74Mz7q2Ev4mMfUTbOrwbu4sPC
+4+SSgKUbE8I6VnWXokFm6h0jpygfTGu0FfydYzpQMMnyje1Ss+jgEvWO0X8ySpDPxeLIy8QFLPJ
v1Q0IsYuMqJcQz5+JTDMHP6uAJjKcnlBQ8Hln7rs9RFK6CwF7Pni3VgAHuVID+diSaUeMO+ovNyB
N9P/J2JTXsX4PzoeTC3+oUYU05/fhX7zM1wa9eTw+RyIPFIzm6PtErsOV0aQd5atziIXlz3f3ytY
UTC+rqpENKj9nt1Uw6nVcRhR2yEVTjkvNONI7G+5w9toFGfI3g4uSF0Ft0OiKEOlUS+/swgjN2P6
FLUWxJmCKh+wER4Mk6WaOIyIaYED1hpAIcSFn1MGssbaqGBmlgZkUp0/maegb7j4w+yjLP+vDtqs
+2FrQGkekgGTrqdMHMD32V1N2Nnv7g3ypF4KScJa/Ny7g3vFtFmxnkZhwosHX2lNJAFx+w92tsSP
NLCiBMyPhcijSI4eqC9vPUiOH89mIAfShEwJSBmc/UN0+ajfzPFumegsSbknbJurFcId9imuhjal
6/f1vpTR1zxV7ipzLI6zeY+w898rdex22h8kBikif/k6sd2/OpI5Bkhp3WBnDnP3FfsgLBWhIYU5
82WqwICliOtgxLz2QH8OD1x7H0gJQFi1LHSr9E5FWEPuLa589HoiH0rL+LCtJPaO6KQ39OnGjPzr
ugey6Sf6Fw6qzsktSfSBrKgBzbyD56SkOnmKW/rKxhrIDSiox1916bOI5hNnX4JOBnOJAzaIXCCX
dWFa0OcqV66X6Vpp+qszJKgh3qk5+lHP2IWkzV5EV3bw9IYHA3gDCw3kmfAx1Bw+gzpgzA0ZtaI/
PU2qa7m+3sNkq2LDg0l2SIKZx70cAKDisTFn/jljXcz8B8NCa59iFyoNfubJtLGkRyoHcZWefwDO
XNGBp8zbvwpZrzt5vKVUmyCGxNYcZ37OYudc8U6N6rMpkMyFVocguDCJb/b3IeXdtWLuwqVbb5ms
XYFMWBYluc5pTjsttD+F2FgsaQx3Y5ITwTZmnbBVAnJMv4odsAP/8sOw+kSN2yjk2BYFdtUHN18O
8dPwlXu7O8SrkQXmmGeneH+SwTwzpEgjsESpLVQ4hdpLAAvtkhGdO6oiRJHyJHfG9RHfnhEZVe0H
Q9ntw/0bHuY6pLQ3RkKf+y5v2eAprWELN9hMvWxnMM0fGAnPrS6pO6Wotlu7+WWzGpVzHSG3LKRA
vZKjhvwGD7WiSHmFtgKROgJshioy6OH/gcutachuSaKO2rv4JcfJF+gq56vnZ5S5fWeZU3FFoiEs
NcRAWhtX2ilRkud38LykucT6IK7BfZsNe/kTftelCb0deGe/EwHeKKHQAyUp0Y95xtOJCFE1u4R4
eF1UVk+hxeY7bpjV294bbsRBkh2IIqX2oWmocIP5PBqqbC9KGSphCXi30UgufitAYKonMcX9Z+vj
ceKNg12pyvjFooDrlQL8GVxnXJdvHi2qh/xF9z9Aq0gUUk8EwEYh4y2+qljx2ee+/BxFew3hpG5g
vLhoM+2WWBiVqqEDWue7VLFzN8btLxvP/cbUkQRl1jsnWSXkYXH4xQ6ILuXUdkrNWf5IcZaVWsxP
s10yVueQXCo7QYYXQvWG5XLk0TeWOBDu5TfUMeO9ZeICwCCheJojE549XdC587CqgDw9CCScMRia
F1ajZuqC0XS2kkz1rYnCOVtg/WnPBehWbxTsDOlTItD/vWjEilNp0/4gXkbOILVDVAJBwGeYKf74
VufF3VcV/2EKLEnyo+0vpbpMxyvcQvxaF2unQO2vmpTLZEpBmpA2QSnKkVyzZadL86NPm7KBCZWk
h76TwA2Cs7kwxrYKN8LVTSNm7M1zVoqEEYmbfgHgP4MeqAGTLscgj5Z4HBHCkDolvmHEmvNHKaOI
bbIecLfTndD8CJgVYDVYQHYmZD1B/UOJjdyJiF8OVvDKVonfZX+qNZhT9yHAyAPUjUoz6mUGrgsI
nHgUyBpge6OtVDrhQga5uZn4glk0+v4wSs++t2u943iAFNST0JevDKWbuLWFQcdYdLsuNIxd8Aim
ckvAj9FiHD+5E3GE2rfIiabt+dP/dXFWpVbzHq0Y5EOAOguMHVVC2F9Dpq7WbS5SqSOlJNnznhA3
BwW9Hnz76aJs7bdH9qzwyXXjm+LY/euMZ3ibyMokz1oPgT3lSSJewlOU4MS6taFkXEJjNDhpKTwT
PZ9WUUD1IlVlJCrm6PDmpnp1EnYd6D4Ap0Q/xcVCw7K4Wdj2r3C8eGqesKPfpGMpmhD632qr1rDE
MT7yX5fpg0MoQFRJ0yCoxlyeRAxpOUydApjhTbRoBUiXLB6JApcHyPKUhJrZhe6H7UQbwh1LU4wV
554R1cc6FFMSiHFrH5vMgOjn3Qr7dF4VCjLoFuUmPiKNQsodZarPWQCy2Ze8pUhAw85k4Zi+s9xX
BPLJl5L8eGUHs9ZJF20FKQZKCVPERtGq+lQMwHqorZ2teLmbY4w+QugCYkRTcOfooqfLdwPZPxTN
dYcvRGt+iQGwCKNa4QDryjFwVGAnScSFSrTGhZusDvgw4MTUE0sNRZwy/rNcHxhjh9t9UhR6kqiX
Z/1bGKOX7WjSCPomcYxpOWGbxyAp8t76e3gkTP1BMkXC3LxqMt+E6xtfaMM/EJ9fwkcd6lBz7Gir
rdgOBze0E7XKyy+9DB4N0l2UB3zUU7vM3AhOuZ5AL6OH2kN2/b8sNmKER44NWdJ6LFNWWKbpkYss
HekXoFCUFCRz43rQhWUracF25eECOBHHuBtFmFu1FpwGkdwB3Z8eL1IPLAmFSVUCQiPnJAqOL4QT
QZiLj7ViO6ns52Q03RJQ/XIkDtkY5goPp4uBSJulukQuuHJZFdUOmgbzlmrjd4rIsbqBXnnsnj/4
TXn8oSt2mjy0SIkjZauFUZbD/uW+MlFAUJRjpuovtZ7j81AOJ0X+Q2Hg6I2p+0akb/q2VAgSLkMX
OaXDhaO+NDluWuyDYPJYbnXIShc8bLNaTYvuLUay/UJFl2+Lvjie7+9Kz/cOoJzXP9Hxb3qfaSDI
q5J+PFU5FWZ9MVFV7VC4cTu9R7AI/27p0soOIwg2DRfsPlqTV96CViYpTJrzeGwu1SH7/r+K5MBO
Nrn3EK3e6F5svjE7rLZlrk/Gt1XmJ+flNR+AP6C7I8KmZdU73wDJm32EgGKPViDE+Q7BPlydue8D
VARlwD1QIIhP73HBBnOxygu8RATk4EmwTVEGHtW7nFVAadIISlKWmYCR/8sHK0ViAj6mjSrJiEJr
JQWdPk5KOw6830qywICmJJ0fLeiKKh4SitLtDPrtETtMpgZYbxE7D1TO3EvbtpOEzZXF6hIT7v0B
Zpr7KJ/0jkihLwY1zP18xBaiCRvZRdgIhHE3qXWnVLiEfUgourwfx5SbC8Uu9O8M2VIU4Qb4HIZJ
4K4GrRUudM+blF5Hqfm6+y1/lwLf/3HUZsTkkhi9XNCrR3kGcMSUlsmt2VytVIdROeGLnD/2Q2dp
XDqoR6RX18dDTFQrGX5OxKOye6CpkgD6S0qPR/9UT8moHryNmWGa76mNjsSiAExmGQgHa1xVTpJy
eG/aXKLH36grBnLqD21YNxX58XaTbxx+fCQc62ZpVB5Qxwz/VvwOOeLmF4SSeDJcdCj8L2/4psZ+
txRolk6/TvP9Rf6kKirS8erXv0CGCUDzi1v+bqpCyFZ5BXlsltEIHyKbh4LgUYjYl9PRK9UArMxG
6u9EoqHD0rfgKndQdhvJTKPJPCEzBwyFQsIWj6v19BDVBsgCL8VZCOVglm/ZejnRD8evSAg5GB80
dao/yt6j2DSanXVsra92Kaezij0lcPcB9c8IehzX7SYi3yCunc3r4tPuNFTFqRq2eTK6zU7sWt//
9TNJnQvdXsgK0O2DvD2aZe8nCAW/y49AtqS0AVpTOJ2EblHtZgIQ6XAu9jvDBHQm9GvqwQmarAlU
hdT1mngxD+0Whzzh84618muJqlYl6CpJtv7w+fYmo4eqUFw8k1BIzv9O3Iz0kd/Ba/id0bJ/jep0
3hRY3m1MIk0Ck9yfcTQ41eroaX5m/5+91/eXBjxot/WSdah9NPExZa/PPmM6N8yTrDRrk55SKeT2
yFMwQUnpk+nZJRE6nsvFs14sIrsZaCHHiYzoMxq56Hz6my1tH5xBzTvhfsGn5wYXeQdxZeLvhVG0
CCYrLF2NNgYycn+JNntRb8merqwWLo7pitFt6NtJKVNsP5tQ+oLVEzZZiUZi66Azvtn3VP6auMfi
NYm7HCo/hOF3pclaYTB3WtT9Pf3J5Mr87JELVzs0I/S0s2dFwp5Hn4kf5+BIATe4TofDqAdzJ7P6
L8O7jG9NP1mT5VQnJBJgWPOGKrSJ7QKGhPLdfHO9SCrTWmsOQWfTDxBY+oLEHbS7rjw3hki6HnIN
YWvqgjg1wTZDBwkBop4Cx69xiSQSgQhzRy8ITXDKOEwumXJfyxhQFGVi6tZYRrUJA3Bax5v4hH+R
AxPdUstdzsKEXM7B2Ez+N5KJtDrQb9pDMUo1yMdfHUyHV+E8cgBALd04EcA3hXSsBAA1SabKGgh0
W6h9A8vXh64uzgzxmSUW1cOqpzgkEpnjv4c9LumAWqDeaJEbhktjaesaUPajAvIDnfdpivT3qZjG
fZp9yu+QGeUe7OUbPRqLs6Ur4TVwaWv1ArUA70ye7a3w5qEIohq/37U1pWuDCXQSSAVp02f/eXMc
ZzwmyV12SdHZ4wZGFKZn45GFdxbDFYPYY+1S4MBp5kCCt6mkWAsaP/Ctv2IYQFW+37KXFHq57LD4
WezdLLW5i940ydsDP2KsIuai6VxCnhVNPDm2NCLT3xmO6tvH17Qjd6J54xOM3J27q/7HAE3nmP+y
5s95pTasQfdivtnCVMn7Uo71PaKTcphzosQBvKmV2fmCUW0IuVVpODp5SJmetQEm+R3+W9Np9m33
nQGVfMDZjgoTw7PpnwmmoYogX6qbvOY+htFgJbOR5CC0rsZ7MxgOjY8CFwm2viVtI4EbH1EXKeQo
iELNOPg13opiyzpnt0nDpbia/ZpYSOkb1x/gOrK8kWk/imaP0Cins4/oeRXqeii5vrXlEVQJ6Jf4
9IpgLfjRPbOm8kycZraD5+AMGk2xmdtytvH2UsS4RgIWKCTIyX6lB8k5R3ZITgVC9+lgsPp5VIJe
1OULsICzVqDuMmc6DLVrZh3N513CJaGL+TwOyrC1jNm8JQ/gEChcMsWaDotGvCfjiptM8i6IwXKt
X46itU12/aPjhqr8f+aqL2OWeUvRQogHfEua/LFSxvYXoRkDya+EbUo8T9T1RKCxSV3VUUFCovCb
xXL3Yto9O9DHO2EU5StaHaQXgwyo/AQH75PEAMvRcgxldj8436fpzgbZeN8PzbO9Vo1WkDCLEx2i
cV/nn4u4GTU8IpVBz+JN/NRixhemzQ6gpYs2eTX41UkoROM5znXjqAyRaH1IX+W+yWVK5fvJkc5R
XEzQzM8fuQgO0oImU0nj4Rueh1+O2VFpJmXzPR4DQodBdy5cZRSqJ+fjmRK+Htly6u2sudalIhc6
QP+4/ge6UYxmHEInMXc20u7q02Q04+HdvU8ydcMU0Q+B4Mq35w3wv/ACgndYE16kbXGUKSPrbjlb
ncFLidJfwrCRHqumRcqPTKup7NidlhgxS8g1jle4SHgCZytwFLIZpKdiFRLwsA1xuVjAKlBRD4+h
idxZcvI3FsyqrgNvJaj978g7aaWWmdWFNcIZJ4WpRVwwYZ4oLxDrx5TtUwCBEtGHrjfd8hWaj3Li
Icr1uMVODhjT+kNfrNk74fbW/pZ6qfoPWVnDoWzjP8ZxDHmLjSjAoYS8WVECIWWisLmt3pIJ07DU
Q3jpDpojBVDezZqBkooyFpwm5zq21AHHpmlFvgpKJX4YVeoaGOoxnKZc2BaHLdgNYo1vaTK9LU+q
gnZt7mFGxP+3BLC3OuguQMo8vDGpss6ENRAz48BT7q3SH/ICvce3vtVRnuipR2ubBoO7TEtClpvb
6aaFjllBbMDLw43efSsfsXQC3r8CqvIDqSiru1zrm3IeZxSg7QuU9e+/Tl8bVHMfjiKOUxQYKnFo
JtAAfm/I5GohNe7T+V9/7Sj+0M/AsfpQvA/QZoK6B+V44KHtt3/StrRFrt/lqvrglRKv1PSbOAy3
24HXXnBAQePjsbcQ3XxFxBnue1vI2j1HzPeLBVCKkjY0hVzsBzgMb3SLXzNzx+hMOhHs0Yk/q60M
fwdASspEEQksFOTxbTx8WAJB1YYP4Kk68VrwcJxCCJSFL5/ZWJvk4JvbV93jwLNqBADmw9lfVm+9
0e43pmtuQqmsWMPHj1euffAwZ6RjBfluFnLFoBMNZPyJrLdORn4NiIKR5fpiNgMGPftfnphUzAhy
TqbAj6plQj1iYME7p8Yg1nYIraRsJ4mkJJvrTTnc4+dgdBjlG49XPup95ldgh9Kq72OG1AbDNHKc
p8YusDFjeiYqGGOI3pnnoABZxLUj7pugr1IlwxzhjElUg/DSLrJ9aDePhhkPYciDk1QoMZn00ZDe
rld/r68ZYgJ9UD0UqvqgCLh+qgcQ7NRFjDEMigseB/AKoQ+YiP7Hyc3kUKxcOE2PRgFWtNcQEO0L
gFjvI+tyQOcowH/X9GEkAxovs6LF6uNZKFRtbjg/T5RRiWjDkisygwhcoeORiu2wQp/gVM7TP9oF
mzf1HDmlO4PUCOEKlUzLyoxGY1eCA4mOdWZe3z7pS5jM1uYY0Ip+0uOto1XHKWf/DstaePdZcfZj
sCgPlSp3CB1T+roDaHiXZ7UUjMJs8zbMfLKiJsdjwWAHSL/P2v2reE5Q+UhqMvoo9r5OSk5bgjaI
cwNCF2XIHLIh/Zf+i7pTs81VX1DuOED9/hrc3ye/AUvAbdeLG33RIumRdXw8O6mPzV8xOl/5a79O
6KM7fnRhnQuilNiZducLbDiHUttFVrApTb6TI5BdOPrU5sqmJYbJ6wKLI+8n10qQ11FTk2O7Yn8D
CAW5MjWFUU+2yYsLLENKlKBnmmob2NTpT+QGa6Ukugs9khOFrMm+wFdwzXZXuQ0WYt9Y9fTNLfqV
HPgppKV1hXWk0V6ipu+zMVZ4NawElAqMzxu2DuImlWUEfAa2X84FdxAee+X/oHUhSbSHbDh0hK9j
4lWpmJXMuKe0xJ75Ox9aRBubsOwCvUPiNHOa/XQdjqezWLob/EdV+Hpt03jEEBjBXi16WtajhjLA
MNG50rBHlz7yd0Z/xAhOXhyMuOu+5QvZatpz4d9fPlld+6853IjNjuCLX5Jk9qXnxiG9eae3aEbD
U48HyyaktJSb4qyCW5GFQwoK8BeQU9Acyk9Tq+XKP4L6IgOZ7yiiCQ0CgzJxSq6kkPYPMwL7aBkc
0XHM7Q4cOxBbnl/tplhtxKt91mlma+oacA52jEPJ7Ebp4Gh1eyQL7CaZIf/8Z5ysxk18q23LHqwC
WMKpWh3ur1GiXvrDeAxdYimyAUvZGWc/aF27TOXEIq6g3VPlSOvzEJwJ37DRoBQ4h3cnu4DD4+81
qcKPhX/o7x90cJUgIorCHE4NpV2FbpYd3U4iUP0M8p6oI8AZESjtVMlMB/zKzQc4M8Z/loSfgw4M
G1hKKFWU3uEWWggZrgKOmoMWkz6BOtEfGk0dFonbh+bKgKG2UfB4xrOfLzWLVPtJEt7T/QOfoMIH
+pA9TgKIsjznbao0vrpjgY+BiTdJa0xONTDV8BfC+0cM+QxpLPSy7scZMI3EtNYHaYBpMbdtHGo4
Hn3HYJ5sVP++fNLeLOV3mfK231iuD+N3RwjoE6NC/IDkQAeoQCGMrdYwlYXOngg2RdT0DqMcqRZh
TaCqS5R/S3SIi62PNPxzQiJXF54ULF1CYPR6bDAiKWC5+P9ybns5kH9oHHxBvuXLL8atUAK+F36Z
cbEW/I+MGUY1nqa5frLe9N6YKncW87xvt6LIJP8m7rarK2teVo2QqP7YHaomSuXLKy7ZUotGG9CH
8NDClQNuN5XNYm7T6K0UUNxP6vcWxF4hgAbpbLEYv+xJZ7Zf7nVMhYivCNlvuyTv72d/DbBJ7Yzm
bwQqQgcdRCwPEGKr+iKRLKdzgHVPk3pvaxlBrYA0k1L8WcEC50yCgFly5k6I6Rno3schGuR8MtlG
l9aD5zrImq4ekRZlQUNKB1yI8HEZ8bvnP5Ky0ladE5QpMj7B7TmQEPx2Y2CGZBntby/qymCTmV2K
us8TzGVax5IWcAzGzrhdeVcGWKA3JGhiErdUfZDtaeZADG9OoijZ4XiN8gRhcvmwyLa+N5ewLEGL
A2NpPvJSwiZDuMVXX3zRaXGEUJw0bn6X/kg3AlFYR943xUM+y2J/F3PiFWHiFBDSG4ykGKXUQ42t
qf670diqHHdrKsg5r+XgNGno5BsenuX/bGtXmyptb3B8Ky3h1v8mI0O5yDS6wmY6LGu+t9NQZEe1
LPpx0eeOHBtzYvLK696Gy1V9FbqFXaKYyPeixlv+x6dkwjkkqcegd6Q/4lrt2HahRkqSU3DvE1/J
tgezZOr8GkMefrJGeFLqF5frrgAqf+UXlWE6DCAkZpMDM8A8882AceJhU2IqoiBpnapkK7LVqEog
dCKpBGJ7e5nozBQ7zUGFMYMYTz/fM1fEJOUqRZVwlRfCbQFZZSQbqz4lmbHaf+kZnAhMOnLm3NuS
9QN+GB38wc7PlEHTemWFLT5+nEKjfRMS4eAg0LkMoQqmBiHPREU0EK9BXBPsA9/wY6vMBI49zA8c
xjGpLDxgce+Xi+IqVgClzh6f123laqu18Mf6HS2si0yp5bXgj/YxDrIb73KlMBTwViUf0CZXv8yk
vVLXZQbYg4nYQcorB7S4kQTb8Jj+iuhWuMpN5YvQwZYvowgOZYbCF6hz1zOfW/ssQp9Q2eN6amEu
ZBPrxeJKAYiMKUojQtijHUQMrWWDYNFzE7j+H1c2Osq+NYV5WWjbJzFH0IMXNM7jUWSG7qotkE//
VhmkjoVb6l8JCHL7h0Kcta/9Q5O5+PKT81yUHl8xAdRowXnOvILAWy9MginQSTKwONr+RW91sRfT
2xqk+21lkaqqTCu8jF+sk2xr4lAMY63YvZrnJfu+hLDwXWJ5tt37kC/NxE7XYWaQ3uMclCSlsrU2
U2P+q44gYI8hVv6d8ZDmeba+iCPOJgTaQJmuWCd2/vJGRzLEsygGstQFJY/mpsFBTBte7+XHPPzF
HCEjKsPj3/siIvKB9mBZXF3/TtjxoCCv5Eq8VmMem6ZhtTBeY64GsY3ytvBXEmR+V44eCShGWgcv
2KVg07BGhRs3wvlZ3yPQ2L7XmqkOmfFF+wS46yPEqEBDOV3M+biYFXCSK7UyOTCc1m//L7crFWNl
PSQxIPRQFyRIAUDiSejUGPHFr/wDnXJvWIHN+8l2U9Wl2Tpe0A2hLMzOtc3+hr3ilMYs4o+iSPyG
OhTaI8RjihDYjnIZfVuSNJgOCGf6GzKP7zkQqwEXsjC8truBqzOcAwnbsuw2VVYXA/90w0xpGTnd
L24JBAsbsf/EzvjKTNHC0OD2MqzWnzdaXov6EiHRu8aZBgNx1YwkRS9HsZAruWbfJERMRga+wTbl
zAy3S3vG4R34k9WJINuFw5NAe+vR5D9vWzPfvIjf/wP0GQGHRe0F3qPkQSkCnerYwfuDIIyLC5fz
kNgm8hohUIWlgoHYDrrYxv5ervQ6Gi4H7CnOTs5bn+qDdhZTqX1VndGGqLKPeNUlppUfz+zOw7y1
CwlSLMUmtgxKq9/3R0kzmEudebDLb/jIAVzN6q5gh9E3w5l5YXSmjDeu6Vd5w/yRYH8vAg1mzZbC
Y3vCmZeci2ZrWfokL+n9BECD74/MA2wDovU/z5m7ainZ4LrIEtYsuyNYxxREEGK94h1WGm97JfAo
ce8yVrU5axHUgJ4APpXKPi48hHVY0a7GpW5RG/RgjmoNeU0/3zNPkwUiDW3Hb0MAsas2yFJKpIa3
wLrXrVbTCVZ7cY9tRAkuGD5apbclmFqUn0kki1JIiexXTs/dlWzffBrU6vvGA7SMrKhFzYEl0j5k
5m12ZSKmuz3tMmYua/4eU7mrs7AGTDUc7BfDr+3y4mj7PbPhdSDOBZ5pM1SuG279lMPZRtKlPD9W
EcbFHGeRx/+IHT1tWx+c74EBHQh0ygfWfGel8N7qA+eI9p/ncGLZ/mj8AXInPIn7+LMBWBlwYyXc
CaxXfe0LbGRw
`pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
F5Yi4vJSEQiw1daAhKE90z7abP4jP7DMu8fP61pXJcda7cjDNbYZMmzFyT2gQ9ZE
dSgFM57aJ74IcnqOItH13Ga36+wyvYyoob0IVoJ281+6GlcK/jMpHjS5uLrtbOkA
UICvytKfqWDECIpyZi/jwbJchLXwL6I5SKwWLApp8Ps=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6832)
RLbvAAOfEPsiB+Pgz2142bzm26munoBcftyxfiABT4NEm9d5wFDuvL4qSuHI+RsS
Vu2V2AX6oFvpw93o2ATDY4zK/LJ/UYhqBwsQyK4k03wRUBGFEUpt9qZIT68f4u5/
Q9DJa5RNjwx9akoyvpDogXh/efIzqBxW9S/j0p1Es6RJdLgGtNl2hJ463UY1GnIH
LdG9gCTyJn9tSh1eyEzYZGX/yaYggBSvVFDyO2Yi9sU4pbvk9Pcss65C/anOU2b7
7NqiBhD+9DtjExzWjHa+qAbBFtwTip23h6KU0dTpL96Om5LoVATQ22/AZ9oRMmsU
k9hldxQ1hwf/C9sNFcOBK1DRjaniwVfub33of+R3dqmf7i46s/jiqWT9Zk0rcXiL
dpMFBf6tnlJZwc1ZKPTEl+T+F1mK8ttYK5W5gWxwbSj+5E6A/GyXDg+QgkQTwqZD
Jv+pg0gcdaLrNhznUA4QBBq6R8/5s474BGzvDr6Mw2k8yMS1YST8OuLE9gnZg3bN
HsCdR7+l7cmguMcm7cGghkYQpAjAeH1FhW6/2Px2lbgseRWShqASEYhhdQa1ewUl
eaOkcrULVDbNOufS5syExCIIfXuHIkre9el4bcC+ofMWxoUlnVNqstAqafVAbZJX
cltb0DCX/7sUwMHczzFFc3GBnCmGaJcP61IiF3aj9MDTj20ry/xlYqZ7LXy7dGSs
FmDU4wvrhdjXk6Ft13gLvnm//5PJyZ3yx8omXrpvnxRHN17FYfhs6eMaGUN91aa7
dGP+K4Hft5Bu4LdyL6UDZiIDe7UK2ZP8ErXDIv9icLa8mnFJ4Yd1HwHxi5C33uuw
enonF/iaIHQyVn0CQjYnUMNN7mDuAtiMqOkaBPaX9dtax0YWQE38KZLxvaEAVTiz
8M+yef04/X4fKZULjtktHGdeWE28RRpueXO64hgV68QzQZ8Y5QCCx9baV8z9/OVn
+bqpMg1gvWKgkUM6VEpa6kHNR1d2S5mQu8AoGln7jqCA4U07kP0RfQMj1RDtzWL+
f4RMUnYDrL7bsIESGR6Azh0qFcTiyYx+a5DbVBevhQ+5Xo4q56KuBhEWIdsBHvD7
tLnYgr+8l/COD1p3O1h4sNbmy9tuGSLpgNr78Ek6igzuYD2JVRHAdWh0UR4D8F1s
6wmDw1BPuViSGQ3oW6TlK5cYNHcCnt/OJMEinv2UDHCzRGZ94SgufGLED/una55L
Ot5uSlwUrwf0bFFdwLYLLgPbuOxmTsxodgz4UJXHle3QCyy7WfrMOA/soUO85/+Q
JOCW//xpiGM9ntjoNFTh9tbBXH9J0vBZLXFVr1B7oyS7G7NNt6vQM5WNxb90ulHR
hheLLcZNAQ1jztxy/U7hH9xdhPXaSSySRpg1JR7HjCMwjxazEjWG8QBh7DcD7Qiq
9rdPiPeipSDpnlTuua75/+9bdBzXREjeJ77RL60rGQamCyaInXQQZZTRoZiF/INz
+wvanu34v2jM8lSe8wQlAHScSH+18Rz583lYOnuCmYIXztX36ybbj1V2QsnvmCg5
7AjtCtAgXYNXaxaKLOUZ5Ji9Wu2oB8aCNhA8IZOIuaMSKP+4mZwhUHSCJKV02j7d
a748WxPD7FNyay3qMGnb1bcxESTj/HShUMyp2k4y/9/HazDzusETxxjb/xXhz68A
fkaub4aG4aMij2r/hyScqS8ZoTJVnaJaBBJfRANPJHhsKxeOLks5sk/r5rfiMNEa
wS3GfsVH0MrtHsFzPbrKkrfgBQzIcr1Ga46m8jfKfabQig0K75IfzJBOYdz8Uv2p
bMx3rGMH55v/vnJ2ZFkptLAHSunDgpr+9oiVGzviqmUaprCKJ4OgMa0P4yOolMcM
NnFjWBi6l/OBy60Ye29HpyBFYTYt/9kV9jjnlfGFJbMLi6H10Kx/eT8kfwSNXp+c
juYVvJALqDmPrxIMfII/uT6pDAsMjFnymgDqVM/0elONPHmFshnUVI56rrvIzCTF
eBAHCUZPLA4/2Pl0ZXwlMl2jTmHOurarcueR1Dl49uUeIuQlQiAr7+7xbf24H/aZ
gtrvONnpI8q8D9s0E2OoFmOtZmUSKQi/5Lp3cKbYoL9mgwdZWKb9WTi1xBdVn5S2
ojN+sQK+21IrdNSZoib9KM8iOh9FmaBU+QhTtogtpXXRAOkbj5cIo/zYGcrqET90
GmgdFNaTOlZKtcvheDJtrE5SrVXYUImvMl0IkpATn4cwofYDON+RfmgRBwl6g7m2
xPjwRLE8zjJhXT6wdxV97aKTFN1IP7m2vIV+IdI0xtuY5Bj4UR5Hlzbl2LfBbbBX
B9waTIJklCLcArK/DCKELxUpLEb6YhkYiFFKYQvgo/RL4n1Qnji8+6fPZWqYUD8B
9cc/2qcyHfdyVjlPXdOfyu1dDTMDH2o/1JSRud7XhliU6ocEDBmY7mfvrH3pi/Rd
wu2sXB/F/GNXk95/idafT6H1umQUEasZHpFPg3cMPpXzGLt2EebQjEado48uqgt9
EoZVysUI9nVUag7yCqW36PVvf/gl1ossMoTMF8nHEfqF+Bz06SeVpsXFpEoJZAjy
CU0L7hnZ++Pa4z8eHW4gcmJicK7tueBvR7jVGE5SFRiOwEDcFszxNWH8iEeT0yHl
8yekOFGAODY2RFv+o6FwVgelOm9g2UDcnvOdpy5QADEpRADOezWoAqSgNmAFDy6t
B6ENrgx5qkOzS1gb58btKDMDl9N4yclW0Lb8aIdSWKIGpqwFPqtijpvGcy/7iKLK
6I8kWtvQ5eDkf4eYQXdT96SK9tC7RGDDUf6FMjSOQS5mFD4UrRCNgC6aQlghhX0R
7HfALw+8vyipFohRSg+Vf4hY1s9LdToBCKEUJRGKEhyhQiMpBIRZ0pbUZfo4hWSL
JaHPbYkg7Cmtbm9+XM2Ctq0fs0eh64MjPhkx16sFQ/GCR5tROjTHMUX+mhs0BUIy
TwnNL/alY0IJbL/6UZkwKbeYeRe1uXz97I4B3ngWtjNvXJh3upzgSVxJNpqPvXWC
3bERp5Rzr4/6PYZp0ghdVAEQZX2kGA6lKJDJW71a2vSn8t9ifGa5KHSi4bEqjhoI
PS6xldm7DFL5ZMRGdaf1NVQoD54h2JlF56YsrFSWiMl3Mv5UkFksMNhuGMAJN5Tt
NrmYeLL7jNy2aMOM28P7zJ5bhNflmUccfYcugxYLUjvgBs5BfAIdB9c8vsLMyNT2
TlofL7VVnagiUTbwRmfrpauQ4oQ4kvIvOHUQQKSBNyb5EnBorB4Ui4PM7+2d+nb+
ILnX9IcmJHiVATxqSyhTCnr69eizut/95NveOJ4M+bzZc2BmGr9/hXoFXAmvgxTi
VbGsPHVhh9v5Mpb4bPKIVGXWFboJulT1A92jKAz0ZaplaisTPohDUFMDUjjgfPyS
UXnjmtaQ4H9oyIUTMuZcH+/KFjEEdsXembkbwllkMM2pF7/nEq4YdzCnvUDfZl76
YYmqDmji4+gYK6Od3daidkhMvgebB14jXWFDWy7zS7GxYr07fAstVdkB7fU0o8t/
Q89yUh5MVvCV8WBL3ExKPRhqXPSZR6LiqbYVZMAMiSVtxTQcMU59HMU2ptHA2D6I
Vx2Sq8Oq0VEh/R+FByxfs2gU7oABD5P97e9ytLKKmcL/gGkEdnPjaML1b7/Anmdp
wviz2mcOaF60YzaDnStTGA9RGUJG2lrqDpIp/We5vR3TOgLnw7p5QKa6fPzfO7fg
yzJ4/IDfWT3zTO/RLWSQ4zDPxYBI4DI7pZ1yxEHR3tG4IfDtEa8mD3Th+0LP4yq+
bksYvZvVbyh6GNAtkv4xZ+iX73ONlaRszeXRihCdBKGawylo2sg9LSou9V4M+Lco
oPWwph7/RrS4V2TZ4NxKvzhNZUXQfPxQGg4kPWMQbdXVTs1KuJaOfNNswIlEeYgu
yJgv/JzjTPcxiPNS7DyPkpA9g4bGPrH3xVCUgmYET8Bihat8XxIuybLgEXdCyCUX
4H2+pV8FZ90IF+g1aup7nJ/fam6NBntHUk1a+A/NBGECdNIcEvYwIOOMeF3j3LQd
haaqEh//lWSAmZ7RDgZhmwLYRHSvWv9FbaVU14d2J8jj6r7dt13XjHIODR7lcG6E
FIhsXikwZNA7WvTQ0BTyrVEcmeRlKAPBAKUYQzl1e+/X7q1+xSV61gJnmr6fFEky
eV9ZmD+EGud4SmMBLV8EX+d9iXakPQGl7vJf9mA328EhT9vShmMTjrYxgZ1fHDDT
yZX8xu8mdcfXO7zc9fg0jJp1AXzhZK9tLXx4CflqFafbL2oASg6na+20M2TFDsfc
Y9/Its8Fs1tBQZxmKYNGuMKhXT3WF2e7QWGVrwlNK93hcrIDucyRiY0rG1InDE54
4b/XrE/Cq1ZYmiVdvzF4su1kFckpNPI2snCXn4u0+TuJfpHNsJXBH/QTqWahE7Ux
n1irqtSl6M8v5nqMy8VO5jwK5nRk+D832/V+PPzdyJ5eMVbD36zTTE1swb9q74Da
klOo8ddtSOS7KVoHi2BEhkfAapa2q1FwagsTdpWa02PhhjFDbCjGYluvZvQCnikL
sUJGcM+CHPduCYHLcqLL2ElwqpbVdKzjq4K1Hhnr1YwKZLTMjHj98dELZk39JFpX
YLr4Y4Jw9mOeYoQNuNu2IG3l4dBOEn/Dso5CgNUj+yT252wdowTPRC4NGWfDHW/J
oMjVY5kGwpB11lU4aTQBYbFWPA4sUDb6RbZjyt4lXQbU/eyKyTjqebhJks5o6oGe
YUxX4E8QxtYwMQwkzifC4KnHoqBc4mr2nFQMYJGTG68oDRv/sg+U9tHFbudBtWDf
FQjooehj6FAKpE2HgF4F5U1zba2K0e7gXhfMf2lMUen8fXctM0jIxCWczp4t4TSy
a9nuUT79qhJGDVj9cAN39qQBJ+vk2CNEoLWC3LUFN3EjI799fZXUWA9R0BcszqCK
w+0w4PzQJHZ9LoFw3lp+wYwnj173MAl9TzN5GB6oQ3Wa3ZxFLkcpMSOXSYsborBC
veyY5kuSN0Sz34FUQXubekAe7WTnTrom4epik396gzrmNUyQvrJ2Er/395mBFrbG
L0HrojzwUeJuQeaHDeG3zS48cz/yHh/laYs3gwDYNU0jDMWf10dzZIVhNTMyKUbW
HCnMoTFp2yCqVa1Y+v9LePbdvVKzot504WE21ig/b3l4aZQpiJKxLNCJv0NJk8PI
rjoOtdkvVUpGPPNYV5+/vlCRF6bga08yFVk0sreOZD2SaBOenBj5k0dkaSuvjL+r
cI5QzamQgU3w27TtbPDB96oYmGiKv8Zbanf2/2+Cw09sDD7TvAs/SlULKTcsr032
vkKbJQbA8xFwYyzhO2rDKpVhya6UrvO1N+Fmp9V58xnnnec1WzydQfg+R4KYki5J
in97OdBDIkcdsa2KOveelpMXG1K1GagPPzYF85AIrqG4VFFSDRKHvrPRcLwhgSgt
Mb6A4fmE6Le85aK6x2wKwDhlkd6tVJMs8mlMWqsMGljBTmDAyelmMv0eLOkYtSjo
bqgYauMMb8KdzR7Q31ZmVgGGUCLG6rtAGREUw4sgLe0jui6RaSRsnVHkDjoxEjIL
EZetHVm7ecCm3iPiGmO1QvELE5ZBTcSLlTWvsgZ5rJYMYJ/rXTQctU9xdRPt2iv6
br/klOVX1eVBhWobnyua3eVROahGjTQPzD8IdyvNXYPmg4zaPBmQTUteOjLrYQ50
y6fy015KsdtkJDRUHUTfbBf7/FEh9SZXd/poOlreecVMPEW5IIy0/mmIIxZhwl4J
oQws7ax9NZh2BDK+BIYsz+3jfZKnq8huW3kvp8gmyx0GOZrS1lST5F+Ci1Z5TzXz
hPTsAg6UewdkU2IvJxwRNNEI+Dzx+4q/1TiJViF0QwRupTIfZYiXNLkFPz6qO8IJ
hKEIC6dyJ9gJ4+5RUhpmGJvCoznYaz81jgYu6ecb7ANhp5oCLWsY5eTGQDY2cHVP
ZehQ/h2rpE+wubcnBRVjDP+3F4acch7FcrzwyfN50BQLRz/YhxEpYtowL6wocQ+q
FRqRQno6Y2CnkGV8lMSNWN8Tx1AOVl5zIRoVqjzRaqzR/lsIge779CHQe1IjQWRB
KAfx6zfrc5y7UNUXA7pKndH//V+9JKouacp+EggfHpF5PTlNPhyIEmQH3F4ZRgK+
/7FZuy5pdixHX6wwjl/s1xOFwTJlfkYDAjn7t28XuFQyWQRwr9QTf6E3qm9UJe5x
vOmImQlt+XNZ/+9b/zXPDRQ27MMEQp6H0BgBqntxEuG1jk2JOlPk0SnMMYPCDkb0
Fd/EaAMHT0Lg/EbziFQn3BljY81h6MA8qs/dE9u59Vok7KkoNmwDd+rrzUNBYYQb
+nep2EJlcqdav4wVVQPZEeDRrT/Jz+4G0beImMxjWQiIGeitYXgjtxHjLaU4h4YK
ZKHWGHnVPMiPcHLMiOtIWPB1OfTlhwqmYUHC066R0mBEO2qgrb0BRIVXutksAAwE
p446CR9zzhhF+t/C3Hwx7mOYRxLfSBsYBWYadL/rCu1+fs1/DaXH4sjmGKkqoOxt
sDivROAd/vTC+dIubZvD4pEEcuLBITSkhQAI+qtr4xqgwSbhMY5RFakKXHoO5EAJ
gFIj76ta6AObc0zbg76jmUAwIcL+sifNsUkE42wdf2ARKc0myi4pgoxvC95DHXwc
QVti3MSafloF/GBBGEo5vCDH3wPbVoBIg/um1LoBY9WOwKKlYnx+pLkhG/DPC7LH
cmhgKEKgyf8XmNZgsUzqFwYq2Yh8t9dF3b9SUKHMPQdk8lkk+06dnlu1V/N0DDFG
ffFD3tc23yNFZ4kgAU6tEIQLO6zqwM7NlTRGCgC+rsoGkdYiDPAPFXZcAGDlZOYN
Cw2iSzBAHbd8lGQvrRxEJjtRI4oUjQJnpIs+P/bQ3l6yQyXnbY1oFHLPEXhBdSAI
P8s5PD2XwEFihlK360wRubJf4WMCojWRpn8O0VCGHwmYgJJ3AN0WV/fVQWM0ctzL
DjBobO6Vx66RtuuHwVJ+7mS87qyipcK7UVv3k3F8AeFgOoVtiD4QBERPCt7nwNK8
g7N2L4VNWAaJV8K6HBWo2H7ahVtoOUfyoTwwVYTUHje5/Uaf8YhX32RHRnV2ltkC
+/9o18LvTmmgnwHY46eWqhW1p+nzUCPAUX+anieDLbWGqfws9lUQD+WV4Ktk8+8A
4e60xgiIl81T3emnEbeqVwKi+5zfDgC/Zg/cBFPVpEQVwggA7167U7QINZ7aFRlg
PxDoS6yjykcC1dahrWaXVA8ifcDb5tD6PfhXbnhl2HGYbTIV0tnxTln00w2vGnW6
PzZl49UK+rtXiNaYXX6/mvp2nw6hX74o4LtUp0X4st22L0fGVJDM50QG7Oa9k5Mw
/nTZFpHBmCnDlAxWGJ+Wor9N7JZxqLwFgIB8eylZFgBduRVpDHiQ5sBiX/1h+BSh
Eh+wL1RnTmoblNyUTflM8YD5tTQ/lioP9G3YkiUHC/RO4KTbM46N/S42TAcsMjWb
jencqPTxi24JHMlg/gM7pgU0n0FX4pNUgH9014N3iC3S9sPjoiUw/Eh1tpZ4YmW5
yfqniThqRfb9plxkMjtb4Gi4i71Ibr24P7LMP6eg9yOSVV35ciY4kDA++k5g73mk
d/dY1fvuX2M2H0Df+EWh6zzq7ywIFV89erD6M37v0Dogf3HccMpK6WM+btWMAPkP
mqHFKi3ehtgyhXFC2oRkwLunC7LJJCPtyRT+akSvlXPUJowJWvit8Kf32GTrtZ/E
yVanDNssnSvnmGDZKxzxPMWdVXaFprek/5oS8QQZ3EjxfFW1Uv10rPsBREibsL47
TYdS/j8hdeSNfre5qMGexhMB79xA6raoFTeIBVg/2ALhQU6RobAfjKaEHJkCistl
fkN1sYJ/IfMTNb8G+wynNMrN3J3U0D5/j/5DAg0rnc5oR1YQOGKDl00C/OqSk/Kx
Qt3idTyFY5SlmD0+/DjRCCY3Ck5xi5CItc1iELUfr2nGKIMexjAnKmN9tDxy0IpU
3k0Kx47+oa1H1tV67cys3hfu5uXN2YxBigR8uLxg0wJ7cOW6M7109RpyvJlQ0CIl
Ow2EKsSLMcJmzULIEjw0MvIPjG+oNC0QSmltEQBcKY2kpaizkWKWeD6Rvp4ZayPV
qtRzPlzvQTbxob2MCJ16juG7xwxAcX1BSRxN98ZbfTQ+E64Svd10vIGuN8toIe2c
Vh9aaef44/JTm84+yhQ0HP3rNzvZVGO2MMkq60yMFhWGw8vGZ1Z4EUXwm8FZgIHa
Lpfiy8s/xBJr11xXI3Y9udo6g6h63REdHZ9Dk2WzDJFHI0OQ9OM4+ESv7nIgBADW
ahlaeypg58ZtCJtaDEKZKJ4qv+5+/AxkbefC5WNmELKVx9iybEZvR1b5xVjPAiRF
SFFRXT6wIfdH+/eN94I1v1XQvrEg/4y2I2LuWP86X9KdSSkbTpu9xAEDdYd4zL3I
kg/NgA3fh3q+u5F76dDMHkD7lm9QR/gNEp7v+STnjtTJ3+5rg2fqFAV6fH0+qvud
7Os1+Gk8DmozGqxl3NxOsdHsmlwLL/rdye/0o1ijpBXgiR3ZT0w645pKdSyy+8jY
1Z3L271Nq6fRWvQwkcuZLm8n0GppGzEX4Wd5kSmrJS4c6kS6Vbbo9+XiFGL0pdLy
GFkBM6XcAOEb1/6gA9AokczSwj4cjPTTetZqvij8rzC5TmqKdGSdEXSjkQq97b3f
Vcgdt6n8wAuvicgcjSRzcjad/aoQydyYCsBSbYJrw/20yu2W7LA2HeeDdvOMCFp9
snqQseaZ3KsPXMeTR7ZnT3UlOqUbtdufIwgILtI/dObeZ3bJTxa/FBnkoSIfdu37
q9n/iEi79xl80c0pBBQQDmvuHaaSQu8QoVYgXM0U8kNZkEol34TpyTjQy+/II0kr
Ya76SSM8o/ocVl0Ta+DKj48wnes3EgQIzX6PzO6cRhciWdHv2diVobAnCKTo5RQ8
0+Dr6rWkQOKFqKABVg7WwI35mLCuiGSjmnkwJcEAysnie6NTCILRNPOQJPQ+MEiX
7wGtFzyGJRCEIb+CMomRfk+1Gko7ZhmLvuiYFhMM3mph4NeOOp1XYL7h8Ixqk+ml
rgT9AlLDpcbwmliaMAJ5FA==
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
iO7ra5O5NUZjRG1BOQR8AiatlcrMzjgDW7+2DExFlrRRknlvgzwEkteqDERF6VqL
fpYm4W7dqImTtuGwDnzWXm8xRBt+84S2aWwPHiihBB0pNktTJdmDZ4Dh/a0gpXqa
+8f04ycLdtNtzjqaF7D8LxCeJxfEMrDBOGmtBIclpF7ShnaAohn3KromCZsL0CFL
ehptDBabLsS0q+bVsXVya083RwMEYMUA4YCvUcPZt6aUv4YsGbMJ1rR1jkAQAd66
OzLqUeHRPK8YrGNaaDEWL62ScdZ8Hmg1rY/FNzXs4FaPgeWq8X8/Iesw4ukg+i0g
AdbZXW2UqcgtDdMzqNgHYA==
//pragma protect end_key_block
//pragma protect digest_block
0d8nwCkdqLhw27yx2MmHNpUmeqE=
//pragma protect end_digest_block
//pragma protect data_block
Fmw18u4yRp91Gz63tFmCERUwQ+PIPdiS3FLEZZcYrLD0fGqnpxveGkNxvtzU3VYx
NnMVQJjatXOF555cMQjvGpQnkYyhxp8agbAnz7OefbfQG7QPi0rNUGvY9pIBiWl7
wjc6Gkkzby5iuRA36DA8pcC6eQSZ2spZK3WQKSLiQtMRElro89HfXNxUNswr379/
qjnG0B6sQlEp2r5zi+2BZospDaIliLR3INTVvItpHRkgCvsBzdZ9hcEH9o1QOXaQ
h24unQ59xrXocEkv3/Ym3zfX/Euu36TYCN0IrUKPgDzhZe1zG+8sHaA/MbZpVD6R
5nCRVvVs0HWc6ZGycRNw8f3sovpvXMWlHd47Uy5dtSJjA2SfwvR4YYJ0VZFldO8I
1ysUsuKXexxbn9wHIHId4yr93km163Dkkqx6oAtm9MnEbkz4E5VGHH7jOT0pP+QV
qKGdZesuqc11lpsx77Ie86qzjOVBQqouNNi6DEoshMWGbWuEqQRLvVq/gO1lEh28
+ULrq9SNXHCEZTIBlN4dXKR+mjqfRuPbJIvgf7O9VbsySIGnh0pfrUb8mOe+YARH
/wzK4+5+LMY1xRNkgn6wwWlE42NFraOm3Qeeg+h4X1jTt1H8UOgvKq+VSalDI1OV
mIZaR0Vm9en2CwCYPjw4hQ6hngmz+NQrHLoQEDzctLo/Dq6M+smWlzBLwphhRewB
jLba3nzkmVSdbKafcv8GKQ22HhzS4NF/9Eb4ROgpnFHj2uPA8YCo6ZOvCR2DLzXi
GsFSkneCHAsCvlclYCGS/o3ZSr0W8BkyxakuzX8Sf0UnwNQzWHEdDnnhqDySwYP9
1XY4Tx6SuWCcYdYS64pWIjfPvt+hnGmRqjkZscs4zFSsVdu+T39L3lW6OoydJo0e
kwyAv72d16Qn7WXDUKuoWEUifcX+HRgOkT4amUGeK5nlWIaeirqHobh5POiopiXB
WmsavpfZdFNZNT6Cv8ZJB9bNq3iGMphPckGyI+XSl3LZs/zI2nIi9MakgCSh5kL3
6CMEybQpiIDPdKut/NiItwosUu7qz2ZQo+oQkkn+UndKzf0xxIbJ3xdQgW/Lmbe5
VHFmNbStjq4QfJ65TMDclxjIaKnlnugTa7tIq+epF/uPlMCk4wZ8CpwoMfexvlE5
dHZdOk+II9ZqNOZUDi+uBO4FTkoWvtKqj4u8oJCHBFw8SMYPPGNQu0B4FSJd+Aq/
jJtuM3DxSzALBiLw/QYccHbHurnPnTHjOWRg1jK6nnUtHWCYvb9egmq+PiNmS9dZ
hmByDCWpJtsGDLL5Ss5cPfABy/oUtUFKNMjGnOBRvSXJj1Xu2t1ksYAimlCVXn1r
3kjfGPUNBhDHsxL24tVHaoLeHIrnZmWrWNmNi/xpQ2JcdIsLAIJZz3LFdL8aPw1c
OG4qq76TdOrpaHM3kM92uuQW/jGExsdRKKn+rUYsTWflH4i03qsDs3d0yWHgXPYj
nYmmT7SpQ7vFXv3mjkeQQexuBQ4Wffwi9U/dppo/7689Er02PetUblP/6Fnh9KFP
AakFlAhGVBqDDB0e2Hb6Xiy2Z4rebKDRGimRHbVQDq76GaqFvOjMCFQPfRV+S5IU
p7knoIP9ppJKNdUWlLzSysg9G1RjMN0+0uXGmuiEVNZ9Ir2X6gi8mrx4UueJHQA/
SbLcWGVyaz9M4qFbfF3HAKwSmo+3EhF1JJ8ri0mwM/yLStb877I2CAf1/XdKJH1r
Dy8BhIsD5Ct2g1wrRPao+jh4vEuhhHgmqP1uy4YHXvN/1u1MlPfNI16aMDVeRQAc
lzY0hVjSMiNViqqg/JG6etb9Nn3x2sWc7q5DUitE1SGoq/LI/LgE9gtB9UKTOViu
RGYAj3Xsa6JH4WvT5bCtoe3IK4o9jVU78E/oNSFrN4E031+prxCmD2jxhgy98nKn
9OCPRkIjvvwVG7GDHg8wyOepqmC3O3o99Dlbnv1hgQ5WJDBWml9Ixs50g6LTyzeG
6k8c0rYhAnbecr81hjnmHuobY7ED4xljvEF+s7u65QSXtWkd23Jiouwg03Xl8uyF
gHp0qhpxmxMG+Nt3OyEwspVZsASww3dcdOkoHgJJHA3HRRRsl9obhIm3KMg4aPkb
N3wZOi3SK6cPJPzxtDOFsgqEtflgqvCjBlcGr5sigEozG7lDdP+TJ9fJr8NAfnJu
DruF5lbrhvUl38klyODmKrPpCjOzV0eNf7vO4ZqeiQ3rFRIGjUyFt5ooEfFjbbMD
MPtdNGZ3SDv1v9aq0IMbAXQvdw6wMAuoJPZCiX32yl2sF+b/PDj/A7rPtnK1My4y
i9Z/lE0HQ3ioeF4NEmYkx/Y9WNQToyUGuVrj8IRbYWlCSbt3MG//Nl5+DCFLzO+X
55hKcDfb+w7R+9Vz2ca2aUusWFokw9UkIe/u0mXIBXb5T65W2tvgYr2weN2p0V37
rQXE98JrGd5cKwX5fVz+B36cyXjqJ6fcH1ndWT/Dpvj5kgyY3eT21jAaaXAWz+S5
40WQqBzjNreUKYSgsYIf0GnRx1IDuXp8H1EQdrJMSCZzhjUIVSLqGCYKcWnjYIAu
zGRfIK1pXDcbTZKdy+zXJds+QV+wraPHcDJgM72fx76MF/PIIfCQjYIQ1U91+Gz8
rMzRfJTBSNA+ZVM/bTntOwJfQFalJHVQ3jxNeRkUVmoiS/aMWtHZLskfQVehdxaf
MjCgVsiN16RyIdvpeODKT7rvaOcmCdnoETjbjRInd6ObAE78excFBaPRzmK2Zdmm
Xw3E+LymNVBtch0AKg0oN4sQjqZxyV0rjdUNLNBJMR985GdCMFJzzlnYAHCYjGlz
xf/PpWEHOpXYXQULr1gAjDSN9s81Z346kfguSC3XqokuWoIHZJt4QDjRk5bK1Xa5
92NdVbBT/gpzP7DukUA/IvbJQV+Xnijnm/k8EtNvXgpTg/HcQ9BqylPfleUHV2AF
Bms+365PodzIaSSRAWN2l9gB039jrypyWbcoKFeRAp0Tgw5nQmmg5mjL3UEIIV/j
1dSE2ZRhgTkB0mNYAqtdyhMbCo1HCWJr+kIxZEezgfSfJxJOxD3YlvliX5lgQShy
NBa3gyR0ftuXxShJdjVtBp1ubhkIteHwD+f5iMIL2D/N0GFWjuJMrwS30GnHzgqn
14VYmrQ/gsLQmvcU7KkbqUHIYcRtLAHgvIIXQ/nYthUFzNuV25gGRLKScZw2E+Ct
YdAjel97uUuz0DL8zLZssVTSchlOgj/aOlPfLHSjOBXIpZnJDffQcGpTgcxjMCM9
4tLsX6V9NIgiSJ43U2+o/qoVqldcP7P4rvL5tfJtNi7UguJKwF1Tj8Fntw2nloN1
0H3BGRXObP/gq8fc3aeB3aLO3RiB8Pq2T4/OF4p62J+KFp+TSZxJ7kTzGVuSRi1O
w5R9O5+ODjJ3c2dRhg47QQZ3BGgs/l8f6QsTvAQr8mznRVMyqqgyS9Js2hynJO9w
EpwaE73vC9BDJctOP5jkP9Dvgxze/adrYTWqMXcBVTYEWx1XYhGyegxHADQ1S9Rh
Iwte3tY5xFWBeZvc2at1EBqBPmI+KyeNLUmqKE9E6lGXbqcc7baD98/ecAtM237C
sFY9cjQY+O0AdtUhOm4rGvdAKA4RwjRuowxhlywFM5dTxy4YilpmjR4BJTAJ7OcY
klWtM/niYDA1o+eTVSAPEvsFuOjoP8IM9+BVu2ALNK1dlu9kaFWsnqm1DX8Uc+dy
UlVROBv1w5sMAv+ADU0fmlMuRuAaQMPdGi+ywH1aKibD9ItHlezEZ4JMvgg0AKoC
MUZnWhAXZniXCnvg6jjiLwk5YIopFzbuA3Eg+qPK9cVfmmiLVESzz2+CQ2MWPxrT
e53OnE0RW+zinfBTHoFjR9KRRxvOfwqqvIh8Q8A3Ei3z/K5IT1gPvrvqAWN2waSm
TVUw/K6o9OyhwSitv9n3YkSFmWy+e4tXnjkD3X12/IUlaQL7SGYUcIBmQ8o7Qf5c
hEa246Bx2znrG+jb/Wpt+oQQ7GqabsBKbLvKb3J0gUDwBUIwpu6yaYBdFSrP6bkP
12dHod5rYLYR9auu4gsqy1r4pBUMhcOXfD583fJm6KJxc/sanqFD8/Fb9oE8meFE
Ib7geX27XsaP9+UQknZXklSPXLGA25BFM+hTPtCzci1uuPeURfN4V+DeWso/7yBS
sAo77Y03mfGYIjRUvcInUajZvKJ1VTW6S4rONFS/1xqSIvxHvHamrLPQhuxkM22T
OgCM0ncInCLhn7AHWS78t8U/hEpNh9hy2I4mauuMRf6LXA7P7xgzf2ecjNvmUqkt
5YizSGtSKmFdGNQaYiIg7dLoOdY3Cnq7F6Pw5P7VrG0dO5n9BMegdhZyzhyIosJb
RqcmAKxTmPUqC0IHsYhoyrpi5ZoWXKfd0KQ9+roWyxY7geXDaMSTJzKo8/yS4YEy
lmOAOGrU2VkYq4iFajEa1J3UR77mAOiqPnnfhx+R66UpsAttLhK22vUjOyUp9I9Y
c+M3pn9yZN9ZPeQS2goVXYMyhgVxewbupq1ebaDGiPP7lsiRdsWmctURyOdUljWg
jln3Cd+UG9zeXtUaGhwEEL2LNd4hDmTNznAMR2bgqOorkg0Aqjw7DBWm1e0PZKmE
gN8jaIE9MkV7uPJ/yBwuy9YgxI74NZcuEu2x1e+vrG6rsYldJ4M7/x2DWtpJ7yS7
L5sENI8pOvv9+jlFUeZ3nuItl4nmhXYaY+0lbiFYo8qPN6fPbG3lUnH2T5DqX324
av530aAWfuijVaY2gPSaGAJ8IZLX8wcUcsbCwN1dyIiTNUpNRTSctNYAK1fL0YQ3
eX06b3xT27gG/xWRzuaziu/nTwmpouw485LsQueoblPWFI/3FcFUWditaGhVO/MH
r2Am3t9L7786ytH2dDNvtT+4p4ZX68fHGdc4R69ecGmTB23gOgxwkhdxL9sudaM+
N1AVhS0LW0nkYO7o92yLzL91w/hXGaxocRxJc86K6Gi04LhG2Y3UDl5SBCNTzc3w
kEJpozayrN7RuVOV2Vq7z7nbN7XRpZD7U95mf9lcnJfyqE2Zb7vm5icV02o3f9sz
WydHHs65foBSJcaa6vIEo+AaVko88bZ58waRSCGqMFWeWkCQjElP4bmC3RAziLkU
tKNmhgo8TxtyVBHgCsbEcyDmbphiSEZ8EM9CQU68biv9wR+GVij6MVt225H3VSH6
UmLi+QjgAF5uvgLVQ8yCxMOj1rD1nrL9xusswVDcptEBVo5X1MbAr3mslN9yF989
HbkxQw+ysJFOlVZkDI+CRydmtOgiAQci+YmlsLEfWY0Q/Q/nSZDtfQSsqGofVBba
HXUxGE8b7qNs5q46235SBVzg1O8hxb3z2jb7uRcLQjnB7tqzEbJs/LguLERE8d/W
xK4pWTo6fUZp2u0QfEs4H7UtHnDsKVf9bv92Pw3uY0j6Mz9JslRwhX78AuSqtG0d
68NXG72vPdhRChqjYaUt7u69q+ueQ6MmqvkWgjitvBtYIHKWaw0JFflvfwsgbntn
ezF6knHYZmbHMngA0N2bpgjzqQhxZi0fkWs1BtkOFPzskV8NLBtzLOOFWJvJUICA
sxmv7J0kgxzVzX1xlNW1lpyyEyd8dUPsrTSjdpSBvyxskOLD65A8qeBNY1agVxFe
H07DmRO55shRX2x+SVC4IkslTDl+F259NBZIRC+MCXyZp9Kk+4T1UbJjzLXbEZwb
mrnhcDo39panJVJZGm1KEuGubZx5+qkqfly+Dou3XWDItonGyHKtNQLaRnM77wjj
jofSA+ZrEtRJXKC6ygqW1qe8uqnxt8b2bJsWx9pVx9AC9EdSKhOZQAHwyDiWvM4z
Q1e75Zq3elotVOy7eGTuCFowfxG4odEdc1c3f+QkDfo4ssxlkSL6HfMZlbvg15kJ
JsEg3nATeJp59huy54LHltpA4FRh3voy4fLPu8o1WJVbo7o/OgXlprjinHnXlpTF
fc4L8YVy0MONV0oQggFFeHA1nCXIF723ZAQPs4md3Jx5xyqxY0p+GVnK7H3H+3m1
dxip3niUWGc3tA5AtwlxPUhbtsnblY0o9FV8Kmgs4ygmc/RhgXYCRtNlsT7+jpaK
KNUUlC/RL9jQbdqUxkyE9oaCBJTpTOjru1ln3uJK5t+rbmwuTXgvndc84504FaJC
Qco7CIMy5ZJmCOytEos+F0AwMGpLXLacWiouj0CD2QyszLz3hNliybmuDo7NVX4v
wEgAKnEjtUWJEIFLeS2UTYCjBfLFEAVHz9iVOZ2phnztjPAID+CCHQfwVNBjVTHI
b5dOpVQyaPha7H+cpiXsxgyVMv6KNRzbbVOK/I8r/FLNOHXNNXGCRLw1bLN5p9Dd
sNTyEa1tsDv/hWD6uDNCS9riX38E4fbcTejVsF0qgMa346ChQ5RrwjPsamoYCu+V
Al9N0ZQsWpjB2ZSnD/fQUluP+TmXuAPgVCFrFMAlqjZWnzYbsDaiZY2Vhfv3TYrh
KY03PsM1sFQHPE5kdn5gJSLgHJGD+qHaEF5XgZnv0dyzP32TWdsSb4Q55hVLecIx
+G5K6W5ohTrCayQVjTW1hreAGr7CaKlUlE69DDtk4HeZ2CPnOzRiwgVCFVjn7Yzy
q+GeUrp5SqSKelh1QCNq5LxbX4hcy15MwNGhxijDJCi7mICNPrlu6TP0eCkkBuNO
WIsHhOTOTACBEQtF1LFsuzEjaIKliJkrxpma3cET/9/YqcSus02aEOXv8dELkZjG
yfG/Cutum0cvNBx2GATEZncOMXqcLdJdbhaNv5/Kulkn30KOC4SZ4TNW7CPZuyqo
xykBCTglVm090lvQPzXdeGJMMgZKVMUyvvrMTVvQPJc7wZueRWUSRUWfHHWWmDZ6
+n9Q+0iZfSZ6Q8h1Fh9hhB9OjnDL4e448ysfj4i7ESYLSjraqPeepeb3EpvywJ/8
qmsQNDWdcQslc2btAEXm7z8fA85jPNwDmsHxPcjt7zLw8Gq18p455jpV/eaalzcp
ON7X2KffizazWcP0tgilUnZaq3yBUNdHrg0O3DH2LZntL5TyWmjfN4ui4ZjL1NFy
TG90CvrXoZl5tyxraLgEhnpjtcN0fPuQQB5W/9UbMrSNhJ19St2ZrLo669EMOgqe
dtRSRPgM9ikSFxtFhxsDo2/cs5lvwrS02qFHwEQJoA/+QRQXSkwU5TbvWq4Nyoky
mjeieeyx59U2Oz7Edf3s3zvaB0DeRZjadQAbxjpdfROwb6e62NJ9AGX3Km7gZM2X
jlgPZ4Fy4wWrY8+piE6qzVVek8eTWKLIWZHr0V03vpgntdNWc/3nNyRWFKySLfkk
JPpmGzfotxaWvgFbxPx262c3L0OFjWxSoOfnGQP1rFtI5jWWYw/bNQIKDoGrkEAH
6Qe2/Ue1TsmlSM7wlnGzNk4icFtVGu3UJVQpGj4mWdnWMvD2oTdMe5h62trQFVgK
fJoxIdqKbPGpua4AdG0zsBNpFdk04eQy7s7JFSfEADQZSRbU7XdGAFdjehSeMUDL
on/5IFSowTgosUiiazCrDkigTHQpHAxDeGBwmC1MGYoHFIfcxAxTvIc55MBYZVEx
E6oFnhCVb03JGM1aWXyyAN1MLunoFkUNyCTyfUZgFaS+v0F9QwgHmbauVYuOWekW
KRSo5qUheAWtuTA5DqeXFRbXy0Vbv4+FSx/U4WZXgLFClnONxltiN0nx5WdjsjHE
ehyIquDddvLRoY7rZe/1vclzaykhdQsGQ3fF3RQCCQrQJzcZxIDR5XySdhYQZM66
8fms+DA0NGBJYffyrf4qqCzLemhSaJMJkdAzdMPcyLwGLwcL6OTnw3JwmAKDvGnm
uI596QugdPyA4WRHgHmAlc3XZWjbCpynxUvEgJUhRrpgXQmeoxLS9TacqUQ3wLl2
+cUtbwjoFUbmF6zTbwKcpXVSHbfuXNAKyMQZnjEgEO8jSCs876LgKoDAdm/WVFAF
ZUf/8Cle60bnM4IShfvr6M/ieB6PmYor0TML7CGFl4nSM3iFKgWfodNgn4E1IEOr
ZbtOEBXKLoPpOGn6rd3y5eBHJw+MLbjQMLVJyiP3Tktr5FZZTwJl3MQnDKI/r17x
d1MOaNd+NM/8uPs9RwqLprNEoedNet+35vF/5Hg5RAlMTuDT4dG+tJ38a5vPruX2
KnUDmm5m7Uujfphr37R79XUBlZjD1O3+7QUfZzJv+17C3j+bMuiyMP2+WvpvHFyc
t9Gv6hFY6l1BeBI9QHJvlAhelJeUImqBz6JotyivwWGI0ioW0PLnsfnncVzw4JgW
akg0HFZbjL7oUb6+yiBiw4DqouZ4s5AdbFBCeuYIkoZXTtuRUWJL/wdTOW7ZF+hn
hx9BXFvfMnhZDYpkCASPL+oRj2MDUckiCAoxUG2Ub8UJxBVIfpHBhNFV7Aa9QGt2
IXsL8LceZPuVypIjo1yg2j4VzKxVyexUBN3n6pZnfdfNi/DaWOUiHPzkcUOCK2Mo
mr0PuLghxewHV/QXClNEvAmoP9dp/aI6K6gl0cJUQu1MeU09/MB8m1ztVCeZkoM/
cDHqFCZ6l5FMydVHmHNO9BcEmWGmmfKYVsmNkk82EmQ4PqSBdQP2XKEuOwgu9D8G
KkdFWAf//SOkqMxoKoTim5o1O/yHdEFOaR4jyKKaUQ62fEmLkMYNj5xw7+efFQ4Y
lDBaBxmf4BQAnM3sMDg0uZWZVkYpWHBedXmb2D96dsM2eVyUOXPTOvv91aa51z9J
vGPLYfUnxF9lUb1QryKmdyuFFWZP0VXPGCp8jUo1n6myleNyCPPPc8H56LKYbC/v
hElQZcEffpDMmP5R7lIWzKjsSV4x5vvLGyqy5aRrvUA89JwAz1ch5ndaFIYcBFFA
RVwElNF1KrURjMY0K/penGlHojVmnWFZ3pR12o4VHC1g/Xpe/ad0ptPjm1z8fWdm
lzrkVnT1OrouRAnIlxWsQh2s2J2xyPXA5nkuZb68GDNLqMLYtIpIISWEO/oVJIc/
Usvjv5CXf0kcQfSolCD6BAPgofsvUqgXTmi6RRRlKp48SKq2V+Rt9yRyKtILClGA
4sm4ITk9XbB5hSYutIN8ZZS0VYC1fIi/1Y1oI7mPFumu1CZvhjevBuX7lmlCk/6L
X2IwtffqU+yOF44SHRix00WcTT7By3RL134qhmDugamm88b8sJJReqokjRUJiksH
w+l/uREeraP7gJoynHwAtfY4Ep7edSTiirlWDDQiDzoVjkBbqvVVXmq1e/ziZFLD
j0/rGnG3T6U4lrmQvDlnXEBjge/z3X2HFMJnQs8dVhA0sG6+DjcZSOwKIcW8Zg+V
SMSDRC3wN+ADXFcKU6yGVw/PNBGNjRoXLsGZyAds1oWirwa/cCL5bygIwnPt6z6d
pLEa/Y7vjdCyE28zRJFiQ8E+RIYiGW22Sm3Y/mNSoGBoY2PGVvrzUxGVv12MgmN7
09PrNl6R/2dFq7bLKV06S9qKKhjAwk9XiZCS7oSzbO24n94j7G1QKcMQO9zThJe0
rZiw9z0s0vw/EQB2OkpgMiEFjsztV1h0/KA/xFIcEd94DtAZ5AwurKGvKyRzqY5d
fCSSNl6pUoEJ8gh3dBwITb0ReZQ57otp5pUT7sDbx+pBL8iJ5ZXfLWdTNY0Cz/Px
EIMLxGi5E2p+W8WhcpN+yDsaedWL/V9wiRAtgPexJBWE6wnbS7ibK/ZJzXCqrM6R
ftNajqnRGh5AqpDH4IFzNHLlwikI+dzWwNBTcyz6mVhhT0Orq8UlrHneGeUFskZ/
bSfuEYDm0WKX3z9y6Ei101j9ufk1skvzGJ71f6LM0vsBLjECGzbWR8ESWz3hEvNb
HydN2i8mSJn8ykoyBAiyj8dFmk97gcJeJHhCcUwdmKpU5m4mHkplKqe7fZNFUQOj
KhXSbZqS5maZ03tC0tMqi+BM29Oav4X/XoB3E27BmI0ne6d38u3qOIWEyhpd65qC
4pZByAekuowJ5WQ5B/nOVzOjTxyf6b/iDfriC3bCrDc6JyVvjj02b21u6czxQsCY
K8H8y3OBm5rzDjQgFK8d8okUkA/yo9F/evHUR3mr0QOwg/oCMOh4IHbKBYD7p7Wg
swzOEZNIX1mZzqV9RALW/zPsmUin2ZTITZzuEBZU8qnAM+cC/nrqKUT+gFy7VnQs
Qu92sOHa/DS5r4TFdVQBndDMbsaqEdUxuy0ATl+m3AtqjYHVfcAjNWo7R/198aV5
xUWzFNvOR1x9E6siRXdVLJvX4UIIGyuge9coh8zXKCHXGY47upCdNQgsDcfuNM2V
8mn5UgrZn1WyZL0gfZnr3AWkYSGVbIWeYmqQ3uVY2SnYXLApS09339KBQTGH7fzC
PCPblaBj3ETm3Emf2dsSjroTQtQqAeRJ1ttdx20HlxyGqIm2U0tjE+D1KGbM1z7k
uwApCJq2jqu08vhRoIzCRzSZDqWvJFYATsuuJIyzJkXFE+V4T6JSTW60f+W59frN
Ftz7exB/QMUeyghuf+JsQKVZzlGx1G471/MgrpTbi3FLUxyJp2jdb/WgkpT2oxpS
9xtOfFhac4H+evH64OCXfbPewnANK9ry1d/PghD/wMq2P+ct7gxnST2UK3NP6PLv
Bv3g2U0mIgrhrGh7CaGz6LhBDBViatleGNF31mduWHIjERHG7peoFQR5SIjoYm9g
vAy3dMGuum+K44gHiqcdxsHFUiBCIARszq2f6ldJq/tWKBOXzoN3q/cUidnKYojQ
rD3ZXkKcm5GvSil5blQlN7mRFlEa9J71Y+Mmcqy0aZ0xYKIpy2k2hOJNuVVXkq/0
M78dG5qumqkTeIGUJRi1kxAzVVH8wiPq9eC/vEJ7kFeiuYoC7bO4UYBlvPj92kCB
tUhEZNsZBEO4tV71ZVd9LES8c+0FDRm5vWSq44o4imoxX46GWKa41xuIYHKjhbpd
KOC1HUpKfcfn4TjM+frK7nHgjawagsrNDdjQ3QJTY8fOZKkeoHgpOgG5TiJklFn2
PPLP+zodUnKbgDFDEaJKQ5aNsd+Lsl4bIK6c2i99z3YiUC8h4o4LMKJhM2nmV64U
89dIwIqKXD2rX4eoYDNd2G+gms6AQcocQxKfLFoCcYE78r8dTa0kLjnU/S2qFMez
aIKFyg/Ux8aRUR5S0QAbgCEZkX8MbzOVzGp+deucOqjBfml8uotPmf5ZjUs1wJK3
HsyZ9aNMeqSOogUeJGiDuJ1nIRm9K3cmWGPcEQh1K0JEzpuu6n/QRqlbzE95nPRC
nw7I9iVaa/d2tsSo+UvMDHwuv3EdFublfWKgYzKKd/SJQDdZpDQKUhn2mvgC+Vs8
eGnb/zetGbsmrFMkRKJgsGi5O+BSUBnjLjFjhSXhDhUl3ZoPeq+WkgHp10VwPnQq
UKIATZPsdm02A4Htgn3NhN2yFU4nrE5OQR/GjPqsTNK1tATfn1PqneKUF4BQxAHd
9m8efNbN9SR7aXO45jE4KYaNUclkzNRFLKAB5duMwcLlKyWjJpq5wGbqBjBqUydr
ExpfaDBdvBUJfOOujKTaQ19pPjAZbldzyfWLBw4ZhNSsscHc2eV1L+jDXR22mXpx
7GJPJwc8f1IMaOOp6ZLWsmRyDrcW7n2eg6nyAer8zTszY4vRvUbHTMIqWmZMecER
PhzzXpZ9SYRNWvLMFSsXQDJ1UcV8wdvhVxMuQV3kLDRSj1x2h7zX3txldOeyXNwJ
QQtMjoi8f2l/MPI98QTzADfbzmut8b1H6e6bParRz1Wpwo9/pLwhWRsQHG7aGmEn
XR4wR+ZMNkTZwl28k3+xaIwrbLYalFvJMsEZCCsWM0mAn9OHKkcOqzsY0/PnelAc
3bhS92eQvWF2cSWCpLtWRsYgxsUHZ3mIpB5JPgM8m6YXXo4AvrV/1PO4tOKJUG+v
YlYg5liGYVpxA5Q5F4LPxpvXo6WO7m497KH6I+EWM3Ba6Gsejm2gyhH/2/pnrFHn
NXK9XCP9SlV0SGM0Nql2XCm/5cnH5coI+wvhtAZiT7r/3cuX3WtP4AVWRX/BdP/R
ZPpbRHaaNtahwX2+GgblPgmfXUxVWO0fj+Okj9UCqMXkTFpZ4dgohtkZO8xHpCUI
QQCRmtBAyFH+v1mmZDYQn4ohSvKRk+1GAvwdlrTHuRQSlX/tyX9czh4E6MHCdb1a
+G7nE4F3EjBXVnLsjKD7DWMrOL2UHOLLY2F34n3tT9xqShClxiJHhTRbXGsQygBJ
ETqpp5sOkLHWEeKt9pLCK3CBc0XYcMrxPjgJsxLahRhVSvIMg/ngI2+ZXTiNPoIe
oydcdel+3bZjyDRl/wzXQaFUUHFlV0XWxVCZ6lwgDzpV4lHQscPMDXUbyYGuKJOy
4Hh+Uo1hs+F2Pgy+9xpTxHsdOs6O5e3pfPJCh4t0gV31tS3Zwj+2uoh47X3IIy0r
+XNVgzEcV0BSIqbWx3JBDpsiCjr+hwT36QJ8RtinMFOa3q8cDfi9NssUftIOkZVO
4oTPqjzrJs2KVupi8xqGFx5DeuVQdC6SWcsTBWNyd9xU+MPYkayRx21bTSV9I4SH
VJs9pz87vkRE0oAKVO3tFPY2sc0NyZ63RcC3LCIIZp8qVUiaY5LNhDo/0vNdQR1r
k8YQQs05Nl4UXo+CAwDmE/+JiBugGUzZUy9Zkt1fyO9lZCrzsxIfnuGE1zAFCqia
IqG+CUEo7lF79w7YvnzFtnKdT0w2QMjMRuXNAmTNTc8J0Cyn7ickwBeb/y+eeprd
KfH0oikA4WkhmBKFlx7FcF0b6cBocp0Q4VFgz1v9BDSDCSwEalr/FiCvehjSbZlM
lWE1z88OELpM79tw9whOHZ+VweGdAt/B/Mj7T1wdyclXds4xlQefxeCFhZnbFXtH
YrtNhhn8Ym3+aze/yryMnOir47+xNlfb3NZanuFumPwrjAnOs1SxC97NpMTA+TaV
wTkBT0TL87Xt6hEZcw6+CAzcaWTpBs34g3jGUIs6Hay5TFgFehCDPE9X1LZRQxm+
qnMslZ79wBb8U/nVEghpF3nKZi/+939YAlsXRBBvpQTXt1i2ceEff2Uq8wTPgpA3
2Ysgy/ZwaO8LNDHfV/IHUN6q7xMiFyjGq3C4PDCWUwJs1pYkICmBqL9BrIrHCzrG
Y4zdRML/aM2Fv53WE1hgdzAuutqCkEaInBfdUjQh46Qr7tyofhAz8Pz2BhSGSm1t
PnQszQnTD8wPNXiacK21Ndo0vymYo+pjocAqS3XGVM0XxA3cIJDzLkx0ymTgvPi4
bykJsUvZ+Jmq7KSW9bJ/jLVhY+72sI6N7fk+fCZ9smUDDaaZyM++ITVSVbhef+oj
LOEs811lls0k/0dKQC2DSkFWicG/9hTGHmXRSJP4Wpt/WOF4lgAAqJsznkOaZAjo
/7Gi4YYOFEoop3mBBFf48YQE6LioM93SHfEPduk8c5+byoZGfnsWkdhN77v2VTp6
PEjpPNaVDxmQYJeYMYudEchREdu+6/N5waihX6uVdvZK6dSCY7MakmuIHKIkxJvO
PIqwO1SWZH+JKGV9zzXipDO4oYgRDtNKKEEIUoyDwbAqP3HnMsk1C/L+7S7UFWSm
AmAzeOYBzUlaeG9QpobYBlY+gBPXVgfp3b0jVJrS+mnFvvabTUFi0uhLMz6iJIAj
lxmUm4V41+qZUbz1168PjzI8tzzs8bgdpEAUIyckb3dK+umsXMK0JeHbLqTqYFjd
K4iWfRciSl7I6OJ24TcQ+Ul0e8SXZWZudtlAUTOPed01rIxc1owXLdKyqjfc3WrQ
B8tCRbed1qzAyt0pV17gdlP1KkXUO3ZJmtekHcEnNri64VJD9yrRw1CkeKDesOgt
DkANz0PrUVb3VFP1rynudFOPwAsSTHcusLiDuCTJW773jLXEcb5Ws+bNhrhqOoQf
E1PApLXvWaVUb36vdpWXTbN+cjjYTKsM8Zwd/7YAFL7usKneOj7cStrW7vg2v0Xz
tZVlUjt8bNkan0Sd9oJkyrHOLpe5EjfDeIaeMQ75/QRRiNsQKjQ9zdFAQmpT/N/L
oD1AwwYoUy0Jia8m5LqPlTkdwCnSHB6fL5M3zBvb5jYGNzYV/VJLKkGhPrtmtjM3
Vc7NJrSwcaQ/UYge9z+EenL7yAzcKIDhy8TJk//RowrAH16m3UnE6pY9jXPwePUr
H5yRSdiCpK8hAMC0mhcDyMAflBFoKZNaGxKbp2dGPIdDUzwZSK3aMgLqAr1KAURA
YCz9k6iytT/Css/WdO8zJqRl9urhrWGeY5nM9CqZbBy/40XmR5wZF1pMUEdBNYg+
xey5bWDhNDatmwojlaTkNjCALXjJWXP0bp8k6zarQdyIGhQ3F6WfqlpoGC3mQA7r
yjoWu6UH2ldEdXOTnpM7ohfuPEtR19Cr79El6itG9eNzt1O19ejHTvF6p3v5XuZs
nTYiFaxbyl15IewMTj/vOp7ibsjo+8jd2S5SYAj0tDMICC6ePKAS4KR8WDQbXNSG
+2vKppLxvvGb2jbvV2yWnDoCr7cMN/3FhdTSvv+OpLdCOr6XW4pxrv8YQZzLZknH
kQrUxdMxBoeBycE5gybKj62asotSJeo2Xygck0uBsO2re3h/+zwwWTmlzLYngK5m
w0d+e2YaSPNjpjsbn97h4+ByaheDayfLETRHJA7OUO3f2f7UZeKIf1TNJ0lItsLb
5sqpMrAJHTXGXF6hDWxLjWaG62y3vpz1FNA+AX33MJLG09aY1mBPfDXmUORd5teh
xCDDOk9MY1zmUFJs6QbtKLN2MaCtxVnrD5E96YL5TEAHzln+L2ac6IuvcwImpNzT
HUA3Q0z364Lttc+/DRZWNDfdJFOiBtVFzIC4IU4u0JMdEDOxC0LN2mulfMvW/JsP
zLDIIIhyBtg8w2KlWVzC/mEnxtdacVyTz2BjOvdJZs/C2fszPAujnCHNoDLcFOjD
GpoEH5V/l7foPjbUUn8fpC+MsPjUrLdDtM5nrq8/fsINgO2/+OImBjdLDmfaeRjT
LDki+suBLSJ28VB78Mwur9iRJE+h8kZftpsvgV/zVgkaLA+gVJC7a6eBLjyqm8Sl
yDv6OGJ2vuZ9sAnB3I8pTRMfhoias/6jMxMwhBu9OokhQmsNB7SART8YDO9zNjJI
yxM+RU64keKLi3chVSFG/aFsdBBwlqCd9ahEdyLI42GLzE8XWSbDwxva4Cb/WhSE
9u70DR1HMSrFR0bwg/kUvdKjaI6vBeQZ9bcYeZbHj79Agj6wGzm7+AX00OkAeMx+
G8b4GmLkiiUKQG28HHBGdVU6YP2qZsbKbL8OLeQcyoZviIuufwWnPPKsAna4D9LQ
h1WYetoiGe5zYA382cz2IXV7xtNpcnqcrSrLadEW8hB+M3aJXAQDIkuByGJZeNeo
QNT+KPpnmPDgxAFfFklj1bKQ3VGybQhZ/3nkSpMPgyK600QaQWnnQF5jqMtG3K52
ksSDQVMGiIevErtaK6w7TsG0f+bM5wFssk+7Co/8mH08vqrpJOXhMVDSIQuSxgXo
8Fp8WSi8JrWsdnu+qWEWY5rD/7f8kH35RUs6tR5kWa14kGWLhrkGxoKaarbFjnp1
g9skBn0jt3fbpU8ovyb2os7UWRaiml6OC3k6nLwcV5ZrqkKbWd7nH7DVKSdtxuiW
rXpDw+gNpVI/Ai8MZtUHjOMzCxcvPNc43OAY274h1sJ/rXkVUOQIyHLQc3yl5ZGj
PiPgr3ozeQJsQBE3cYryJH+LBLj4fkckePOf4/l8K3SkQMMV0qmnsxl2cyMPotde
SbU68zsi4KR3IncNYmkN2V9FqUUEP8gWdSD+CiOD3im6Fh3Ar/ttjZz3bwN1NdgI
ttigsIUppNtqYzqyXrHv4XaMAhBKsD1sUO3i8z567JWOeJV0K3ER4z2KSVjzdlph
nmbe7YvHajTBdV3wuSXTsH/MmGUz9IX05WjYdR7EBx6F093sF/yCnfdHSneVpYNc
9KoyMJ+02fPx/X3akp7a42+UtUxemu95bkHqs7hfgcamk1weEbLA1DoR+RMfd6ba
sB9lhNQsf/OGAxf6jF40w1Cz46bkbgvcB4j5LgxgZUdjOycHFRO4+nZMzyRmW5y5
Xyy+TuLsUOtCICF3BSGpHYlxOiatZ9m7mcx7BX3R6iExyfAfi3+PUkPUoPjvnmz6
Lxp6ku1n2qLpFPOxGvYELUnyCl7S4uS2omkARKW6CG5gxyUS0PfKRp73cpfybdlF
C0wtD6v4IaH8vVEbcH5GS4hlBVCcxx7jUHYFwEh5mad/NTjT7f+mLvQBUTjWrrGO
2SWVTA+KGs4hsT5CgSRgD52M8n8F3AYcyhg3RwjR/VvbST8s3u84tGd2ZW7BuQE8
D3M0G9t77wYyLRxv9+KfOLwcBYTqFaxe2YDjjVBjv2iIrnB1ao13XI9fZEYAL/oG
NDifDznGgl4zaPfrTg3JATXQzayA9+1pVj7e1x/oGjB5r7vtGnX8q9t2rwfAKFiK
30TRmSFQwk42/65o12OwkPn/Vcs1QdBSrKqNFlO8X0R5ztPJ/HRNeafBlioA42Mj
tp5lISE63X1rr9bFF2/jRHmxtK63JX0L1+n1e+9Ye2az6NC7LivKxR/wAfzswZym
FsVG5nTzKe6KhjIsfmtAI5j9KMPh8K+UzI6YYNJlou9EIcYN/yd5IoMz9HxsW1nc
Q7f4eQH0kNhQmr8QS5d2sHKpSkspw9usB1BnP7waP/86agHfWEEUC2m6ulPY6oVV
lgbB39JwJ3B9WhHzlfuvrae3epP0eq3qU/yVVIqIR+WcFZb/iioP6tL/77pSgpFd
nUAcx4g4c3+sNBcscAnHNWF2zFwdzcqZGDBKvpAHMyMCfn/Pm6uYq3ChrJCuo6XY
BSGnJlgcn/cmxZxp01R7TetLCosTtA89XXWdcKYu0OGwKxOBSg3l1y4mnsb2z9aP
C8UryKxQdQiJ5nIcnturKgdK69zLNV6ZJc2sa8xW0pV/Uc3+dwyDhGwxOysxoJp4
i+6k0ZIvB2khkZP4/9yix9Txvd5JcDqDylZZSbULCLiBsHN8hHcDopYhFYW3t2to
VzVU2qjL5UFjemp5ttwVz4xgH4ump3LaOrkzmr1oHJuo51V5E18GZGhJG8Kg4xjz
3VU6mrJa8n6HVAaQ5eBVU7ToX9kUJMQWi3gX6JbDSkdjAPITRsViwKBPSaIsYozD
naMWaWb8lOrH/sH0LcmVzzJDyqG/rk4EAVntFFUJTIkVKM3Jk4a0X44pozyqBcqu
ZttlZXBYFonvEwt6zhWdeBr0ce4xc2181amvzYNt1Mz34Si7nbXBMDErVU3VqOif
nCgHo6wtHZMS2BGN9Q6OEDFOOyPsEX069eFoHPmLdr7t7ZIlSWdb+eZx1Y466W5V
KiDUMjC3H3yhvLNthFbXn2arRgqUnTk7AX16qrA+XQb+z4umKDE/QXgoyb4pGgOy
lDjn87GrbNPG4pMsWeWotfft9eUSQQTO7H7cYMokDYZCjTySyWfYG7LhIikxD5Nv
vjTvf2Ch2+GrA6u+7lmhLSO/e3DfqnB7gPBHU4MWXyLdF2QFlJdvYLt0T4YuvTQX
NvllEO7RtddTvyoJj6f+RhG3KEm+SYZeNSATP+ibf45eeXO8cf/YkamEOpy/FJ8m
4Q5hHsrYq/W1/y2AhIZAH1RDtDU7hI0ffH/+cEYiYDsWFkQWTTb4a6Q7O9YXx78g
4O9mjHnY0AT2UzS1w+uYB2M3mGwA8Qk8GuoXb1VyjplGNWTM62jEYM1Yl2TlVxyq
WUfQ1u/orrEVvAlV8BVHKMSPkc837iN4fEaOkZ7gcf0kpaUehZyHOu7TQW2BhYMh
dXeJlQ1c4FZg9n+oofnHIZ+ABcMg9iWE67OnJjh4ddQrMYVvVTEP2PX3kCClrzGB
D+FOH2AfpeGNFqoNCpDjUmzKPzP/cZXjgYPzkpn9LRIhO1vMfzmBXoIXliYAD0Jb
A43tCLV7TBGDlACVNp3oyFG1s4dBTxiFAcgYtB2qcVXaJU0gDPxmQvfdKwbtpnLe
i5WPXhKzYRS03tEfgawaAtfvwmLriUvQGTrcZYirmhaXOOf8ECh6Tvp8Qw7HWiZM
XD0R6TPUykd6Rt17CN8bJ7FIJ9j44SytgcxpbW4tk4CZEqkWeTQvvPE99tCfYBI3
92FAV9LK+vQlbMKzU6+8H9fq98XoCyrFr/1UBB1g+pRBbUVe1yhbEGBfuxn/a3rI
wYzO9UKicwOMK/EgIhB144Ynh9hp0qPkMEsqIB95BacEglIK7zWXL15qR1c+ahRw
V7JYAg4Mt7Lb2AZjTg+oN9y7emqI54F0eSW2LVnwsSWg/f4XOoBAi1nLLKza4WyB
ey9KHJ0F6DLkiNKdaqbOvBwA+8LeruWy895ldQV7esm2Mra39VUTB17B15YUBDsE
Fk4ey5dtxm56piWJUu9d0WmHuCf0yDGxblU9opNJTRmaeSEtB9OTjT+zvR8SZlQr
qwb8CJyfcezyQeHTA4cR5yHXLpWuKol6JIMNhx3UOM5xIilq+Y0ooD0RSRedj/oL
xMP94q2EKkWo3D9b6sBPBxud667lZ42b8EyZ6iqt94QNEpGvlMLuZTkMdyzXYfzA
zSOW8315VIxpzEb3z5RIBvQk+fG7E1sciMpKOIi3X37zFcwgjoSd+Ewt/wIzNGEY
zcwNpdqFzxgKxnXcPO68R9Jk1JgV6P9yi0EdF1c8VK6xDQruENDgvuHRel5MMJSh
FsDgqdTX8hPjLqOSmaFugJPoP2wQmQ5ifdSY3LNRndDlakrEUEbxxB7gP4uRpKNN
koIrR1fmZBrUlHkiEgS5dHW6wpRIwIXBkKmUSkashg0LedL3/x2CcNWdBvw4fM1x
wPwtsojxJPW/GgAFv86kytzBwkrWG7tjIwBFdo1bejI+pQQVHw8MnUjSZFbzh8gq
V/pH/hjrirObUdnkC9yvxoCnbh38ep1TsL6ZCe44cYGTfYs3XAm4La+Uj0mM7QJW
AKrWBMNXXxTvIFW/nKKoPuyGv8AJb2a9/gUgWcMJ6dRlHfS6ktH4sDAlZE/owse3
yaAcifj9xJeoGusnPS8bdeC2xHuLJmwg+V4S/qq1IvB2pdnaLsA4cuMlUND1Up3j
5toz9NCQ9iSh/uNJqx3E4H01LrfRmH1U49mirNxVVyXqmxXYThAMPOzfKOI2ILq5
IXKak+EKDh8LiCo9BoyjLgJV9P3T1lxR8xJvFFhjBlMBWIR/Uz9z2YYs7mo4cIvU
xq1CuL5LBjs3Rt9riclrQPKXjOOB1RBfgOWH8pMQkhduuyk2PYF0OrJmn7oBWG26
rIUCZ35qLKp30MNBcZlcNCv4pd9VMLFeZWt8OvlOpbWzzBJbi8YWOEEusSiVo36U
hr6iJlRu+ya8tCev4g5e5iz2CIP1roiMG/uPlOVSsjm0fkSPVBe5ma+cIJnSfbyw
D4NWQsG6dPMOWvwqm2XC5pjekEPHtZO7jOBjw+it4D2eNxXDfuf8V7lYV8TV3e5w
NxwzuIsduXdvZzAYkc6Nrmj3Z3ZKzVyVvPJM402yyMWHZsN+ra4sETUs7uSK1zfV
nF6daeKSuB0gKYcM5A20/CbbmLeo7IETHow2pm4ukodXdbRUMy6+dwDrmB6QdN91
BOEn6VwFsf4zFdaDeoQWDDS4ylfHAUrFEbxlHiQUfFpj4LrDt1IVvkO6NbhgU7vu
dil+FD25h0+xj0xdyBOOA04tDn951QHXSfpWNNE7Fwu3C+kFA6iCDEWMip43WbNo
OykiT0Xfq2r+W24U+/pMHNs+3gXBRoHQUNFs5Agugzk6Z+u+KLr2GcSrM6rni/zP
N7n39H3ebjoAvRwVhYIkmM8pTEp5V1IJPvA0et7ubSQ2zmH2eRn+ilLoXVk1Cae+
PxItJ003bqpo3z/7fMn7l2gpvyY/o+k0dGnkM3CihXpWiU3SCe+Ptw73MSQC5a3U
zCFeWDM/6EZ3My/DhsjrQ+zfD5dGicTT7JUOhAI3yiIuT1Yf2X254daDsf3kVGos
SpjY2T6drPTlfdVcy116ZeFqk8UE9LX0PYpcZHX3ic6wb0p0CFV4ttEy2zJuXHWT
oVEoA3Hng/h5MNQdm6s0QKLJoN0COX/FoTnqS7VHEVUyHPph3VeEYIoff2TugAor
z3jLmdl5aRgdqK5qZ2QEo8VsCvKa6eV/70lBRSCvttRDLWUI16i6BwKGGJ32ymwu
UlahvtA/zg4S6EVfiYoTq78nAoOYH/oKT2cGewMC56JRBrLP4iUMatXTgnWvdTxr
2VtNCCgf36dXCn7y/sMjxhMATMr84/IQbjRcE6KGwoN9T5mj1POfAz/1AL2wIMML
PbYBAOA7VFeMTf1R+7iXcuiXaGklauBv+DdqsSMB7NPn74ijiiS/1+6HJ6JNOup9
ck6cLLWAaP0db18y4mRzid/y64AsAnT7mjzv/aGqeWO0O03OXmR0TQewVGxsjmoT
wKiidtXTllwe0AdCZ0zFRBCk5rHZfLlA5KySnPHs8rijtUfhzfVp9AvHUMt8dIRT
jALGoy4egk5nUibCoe+yKBZN3mjoosEc3sfE8ESBlPgj3Tb+4+ghcnUtc8vWFtKM
ERfh9ReB4i8iRIYHBvch9wV7SYq/18/kMJM5OG11k605WlC3cSbt3FfHMOEQlxEb
83uwKiXa/ajAumYpnTifeWH30voAUO9AvtWllmoLBju7T0yWx6spxFf0BhS0BZg9
9doKT6jFG3Ow/zjXJfgNDbstfTWZfM6I83LBewn+B2JvO96IDFDdsy1Qwbt91zt2
yj7DsVRDt3MWqvGXPBT7qpi6bFJ7yGm8DXHk21ybPTo5wQigLneFcf4wP9EAPAsm
5vxL93RKbnoS+z3CVkGQp/P9p179Ae92RcPQF6KvNeA5o37h2/GYBbNlMEKur3Rn
q5xDqvkp1RjIWW0nmGsy3Q0stx1p2Snf3sKHwBa7Efgdl/lap0UtE2WF28mNenEE
JGk86IvOHAOzCAOYvrxxK135Mnm/qkbocg1Il7vlRhE4Z8EzSogqxc5jyojyTe4+
voWfNNKkgR5jxg86Oa764k7DvtJV19nF0o2m9Q3jE75Ojd0fnTIvf494SWh9YKu9
O3MjUmL6/tiQzmmHR615G8Gk5y8TiPr2QZ6BVKs+R9LaG82iWEfGw+9Kjn0PCaye
P21GREqiIZ2YmWchDweH82uEOmb8Y80hbyoY9QiZCEYqH5P9nD0o8rfXApY2KXZU
cfUIh2LSyFSQvkWhGFzpq20dMQIlY2dN97fqPMT1EmQfN4D6yA9ysgGxk8WivAxu
tStd+WtOucJ0SDo2XIqxZ/e5VsuhY84vc/qQaanLypiZXFSP+rb3tc5HUfXV6Fhm
W7Ct3ojiiPC4qwTTzyG6jRsxsD3ogUqSIZiVUH6htQEP1DTGC9xzQMIjj1MWFL0g
yc4L6XYbcivSq2myE/thdGqdwCjK/nq+HfYT2tMdlZM7zey8eV8hTP2q7/Fsa5I8
ctN9w1fFp6MOndGBUi5MvVFNk7nXlanHEphQ60EEoeFfhCsAW+hGtKV+bZQvh57U
vv54dFjKrprJ2NgTRR0LOsq4Y6a86q22dnu/1p0RlT6fac1DkS2AN+ljpFds0BD/
8D+GTUWqIgZbnXswSSMEQ++Q5HdJKqJL6f5ohFHNUmwxD9Fwc7l4OhZYLbJWf2cZ
6K8FAT/3Wi3zAci9HgJuZrck28msPSc6GfThv057l9DIder7boMBtt7hSWOStIlr
kvs5oVKRv96701NtepdmJruG8gXBTIbbOgVg4trBEzFPx/MfQHEIh/agYSy5H9Dq
agPGpPHEZo+qdlktZCTMYdzs/OUK/ontblc6r0/XBDZJGKpBXzQyPRQLm5ByAijE
wACo2t4B+Z9NIWPHqfgOR03DHXQjp5wg71jvLKCSu/+Ewx37B2ZwUcPkRAxKasaN
GN60m1qN21wuMOfzmGj/RDbyP8bvwkiWc/CHFIxQn3Or6CsRIO4OXhom65atEq6v
qpmOvVXo+tjKZFsp5I2Zi/dgIJwSbwN2wLah1Shs/2duoYcx0hPQbW3wYD0upzYc
H7Jljq+2ozZyhrS4ATvwvjMr/vIdq2p8r1KZ+4UoVTqeSfpglw1uPgZz7kanFc88
oyZmIqXQg05ZOiLzIIqgpVeHlMWjC5YC+7DhRjI3zpALxZzuSvsw9/UIYCV106z4
wmJhsnwsgfr3DwchFPhise0k8oj9sMnrXAn+FjwtNrf4k9QoIMw3fjcSyNnfL5c6
NZxKCh8gmcTpz6EeD7359iWec+SK8a2KHIuT+PtHE16zfk841NKIWvzLlXioOBrY
Gp1EaG4kVVwBW01hII+hXBxZArdilqVhuPWfWnhDsormh7PAc5yWf1IKRVq/7z+/
4/+hFLdnsF2Abdg/re+Tr4LWbPJNChnzEvhdwk4EW7rYk/9fgKwgxaIcHRlH4Tt1
ujQMgkFlFwnkZv4lu9Qlzu5NosSEPxS19KBLsRKLnqPMrQeN0FImRGF0Fp1LjvSj
F+VYQn5pDD5hFHMJChHc8GfR37CPf2FB9qp7xpFOuvSUP/850EOgcn7asLCRpM8x
R4VVeS7xvsjcz0X2Nqz0KZEHXilaYOBnTZQ6HyxLQIsLpduhnCtHeZ8nVnmIZoAj
JNc9xmJvfCuKGsx95whfRoBRVMNQUERRN+hGFsYCn0o3KvN8w3/o36uT07xPdppB
t9+qEF22fbi4XHfVNVjS568ymMcLotm71cuVtwx0sHpM6c0sRe63eWSfGUDmSR9t
ftMPUTMZS7AIRDXVOqaoeEFFg0KBV0Yzo8joiLQMKdej+I8kjEI36ZEkCCMMRHeu
d7BJgndORBcv6MtJSixl3SZ31eH5dpZdaTDO86zOVb8c9riSBGHBmB+T/VIv+En8
Uc0ird2ztH3wQD+q6UC9s3VHbn5E0alvwIAMW3kHO61sac/iO02d1SeNL49EqaKO
pv5kJHYb93cavKyIW6A+KhUa2PF4Td21z95BTt4G+tBGBsyaTJHm7Edk50iiJb9+
Zj4puN/me948YSWbk2FRcD6GbDvbpaErMqGQAMvhLbG8L/8Fb6Y2ogjKqYIMYBjM
28uAVlBHp+eprQUmq5BjdfADK6AyxYYFOGryhNZaZYQy3ClfnvyC+k7PBS406wek
4ic/Z8pNzwnQmrSX3x28twDnleqkjoQJ5Ty+vsE/4z4fpXPdlGbMhbyzQGuQ5tX5
/tvklFh9ZaNuaYz6ejsGAeyb6ZlulM/74HaanVQtlMpqVkw2fbF7FXs7csa2quve
nC0hkMeCF9R5A9vPSNQX7Fp0dRs/6HC2NVeLeTRipW1FkkBTzGPgOJcBDUMX1/Oa
oPqnxBrE/6AR5F+hCiPqrCHcetSu0QYqAV5HmshOME4QYVtl0CyPnSewgi8R0o8l
lDEBYtZqWl73gzGD3AkmwDLLyHELMbhjCdzH24LVg95mymDGRv3S9mOtp3qaQmMG
44OOgRVLAj0rOrKl7taFPhjQ9CFPXN8ToVP3KHl3PkGFRamJG5B76AtFR2ozTVOH
eNm+tBHk3Pmv15cz40mvQGF7tNBRx8JrU5VPo9GUYWQzkQj5oCWABcFj7X4jppXV
HWUmOe8d/f364nB+keFs6PYla8PQKJp2TgPGpY0XiQL+tB4c59iVuqB+sl0RfHlX
XrKFUmHPR6M4xHA9Ec7f3lljkVSDHVvYkHT8vIuEpNMrf1Wmk6s0gn4l3fz+SvLS
4vnFEaCB3v06pJASiJP8LPkdawxCGjFw67UeGWd7NZWUQJHUYXeOQV53naOTkbYV
GpdYNl8Rp6nDXvI49Z5KniOEEWsAL2gwjEpOAsutSiH1kcHPHmZWEaBSaY2gRLeD
1zP37CPYhA3qSjHWicTkeRi7Wlphx9HMTwt8jrKG7k96rSEe4KuTAGRzxcjCwHmh
h017dRbyipFXOg/00pP86i1f6K6weBnGsCtRDIICFKKsRnWNld8P+M0XuyNcC9wu
sOwf6pZAEIdY4FUh+RMzdu/wOxFAB/ahBobsMx/pT6idvauo7WNUbqNWxjZfHlbq
33x7yZlvvrDMgMUymMZu1AvjDWhG7rxwdjghb8FAKkYOUkRn3EsIw8ku4LPhkLuQ
6PIPqEagqFT+730ueJ7MPLudW6kBEfcV7XSmqSMFAaEE9zLF7g7cAKpb5RGsj/8T
5OxKjOLYWZjapt/DOPD7Q/nljgtninLSLMusN8QH24g8sdgr9IEn3+r/kpkVlsaC
3dTt76vyuomKvGPshAIeLjZvV9en9gLO2m4G+dd8wYFTPJfGxdtQ7NkLjFu23fom
XRr1qS6VmRMEpK57OQoDmKwMaZWpsGhUzRm1iwy23HXf/5X9F9FSjWu2IucODmMF
CFWOyOIGdDjYE9l59qQMnbxT1CH6IQKeOSxm2ipK5GXvGFL8kM9HmsPpwVR5sr6v
jKBoR8htIliOfLeBeZysUu2h1lmD0jnj1yUqKQTgpB7zCrDyo3Qri4W6nfcvHqZU
wmuQNspx5LymD1/2ebVWGtcd8nG85c8GGQc7S5pWUSiR3p70a55gt6uY+uWeNM7d
SvEONaKXc79Sx5o+sxeogjJm5eBdpVlv7tBrr3J5N7irA0ugDnlMCLNBSduVxJzI
JKnQOzJOEBjNBHSkTW+6bB9Y0iyfg5UuYJ3qGe86NvcSGuT2jME6LyiFe40AblEV
VflhY4JNAxG5WFFfkPz/nXH1hnXS/FuVKQtfIm5Tf8zrSkkIHMoGbWAo7kf9OmFT
81DIg09vQc+PJ3N4xEEfHokIUwtJ3szDAXLtn5Cnore742vhtzmXenqNibf8+P8p
qDOv5HPnefYnZkam2/CfCwyk4EHRFgO0iIomFtHIkqO2bfXIu04x5UAORyXBrW5L
EceWzlaYT4mnSwnEe6qXFqJWIPqTDDRJRtFM1OXIfaMC3Ayd4eaQbK/fbMziBqJD
QckN+IfqAkG6k4saDJEtQUWKYhdxuaG/tU6ZNqkY89Znh7HrzSbSUd3vmcvZzIrM
bhZAngmi3mCivvyUzTlTX1XMmXWeVdpISDpmADYKqsg/p2W+NcOWPQ0uqFZEQ1x5
si69PvO5LQhrbsQZOEqSNMM8HPfksZgtfCQqfmYlR9wWqRRzZpOb2VSVlfmG55gv
KSaCabTcCpVhdjgbHbGowbZNn24WRZw9h5ePd8EC4yLFXLKz9ozfj59sUdNt0L+6
YyaGbje8h6Tnpk411z81GCL0SvXi2si7dB/9ffHP7AcUw7q8B48zar3dRhkYQqVz
OyOhjTsuNHhUzNk2dHvXmTm9/9mjjbEvKu5Ai1KFEUbEK5YXjUY2OmN87Vp1bVpi
v4UTxFNAhZgucou2oLuIUiAfloRL69i3kDIymYj+P682jcHyEiZJy7lk7pnlqQ5i
HzWqj+Dbp1tCe8Xm6zLZUrhC9CnV69jm9LcHJy8/myIiqpe2RnEEpYImeAVm2VJe
bjgmJsPpqvE8yy/YoMnlIArA+uBattXEAc7YbVw1RQPmIcYUMh4GUV6YD1rKdYA/
Wn1X8x8DsW1+Fpqi6SrApV4z7oJLZO3tKFEUVsU782DCHDRVFO1LjHoIK9LieNGM
n1k+ZmtfkTmsZyYQdqyXjgbqD2P7bTWo8CeBRDCsFj6tl9tJDYelDip4LtjST9y1
uk1ousYSCJ+gSzmTOwVPmSjmHN+bMy1g8kARFqyButd2k1bOicBg6CJGvVUdovh/
Okhw4CU81Fa+ZxUVSvhqlfs49VqYfQblnOOGVyYo/FNcDEIq/CaXRy7pBNhve7DS
Ipp422f7wO8NJvw4VKkkHkdq0bTef+rH8iqlA9vv2aPWoADEfxdEi1DWERbyRHoX
vpQeiH95qMEMHR31e90iPS7GliqGYeYXRdk94Fof+mbMygBD32eMtrBbpH3jciWI
fpKlrUXw565Bbl6tM+XnyEc5zcXQrVto09eXPWN0ZfC6sC3enyAJjZXjcAc4wLap
bdyCy7ONiNDUl4r7CmbVy7gcWRZkJylRbSONeFO1EcLn1HiLvq/Szj0OGPq7SjkL
85Wx/5k3htXWFa7mDz8Y2HCmDNVaweAP5DrweNoEmnkh2AhaaDE7Zr11en7DwiM3
U5nlNEAB4ZEmZxc5t1WEBaRssaQg2ClHhp1MJaaL4nTy/aPzTNyZSfW0XltRpPSN
EtZmnTH0iQeFMD0UOqq+coqJzJH3qNY9Zze5rOEEp2lg1PvU3z4UBlBAMD2KWJ/O
LneeftBPkC07PlnMZXQjtz87F6xG8slxj33QwTOJ5+b+gFhaKcCKvF19QHMdH926
Gy/h1epRXfETOvuLfrPKD9o4KcC84H8Zf2EhrcIW5M09Vr+ACtYGwv5auhEg4kEc
8WMWOuPNYp9rVvF1/M7VMqfVuPNNn0lSjXsjry0dd0miOz2BKxpMdBXr/vrCJGZY
cLGUTzYPb7KcyXINazDWnmKAZKelOKFH2R9cskXLecvvZBt1dk0za733UyfSMMnB
B2MmJqysroNKiDe6vA0tUdYtPlDYVJPQKJtv5OZQ4iZI4PzLQN3YxDg4BN63i4Oi
7K4cX82Znj2gXRrUqjHcl67DLbPsIeZQvYAApFgkyF5jRCzcPSoEGXjrh2LobmD/
zq1j7udbNf+ZWp9byCuKfXuEDivFafR06cKFB9psVVe264djmK3fFbioQlWpvOVM
z3C0ETOtvRpl/mb8paS54MGOcSuUhsLMOszFf5iTYiAZMhb51YnHpUmat9B2zQQH
2cCZqn5IWeXbHvQVTrdyRiLEitz0/e01WRzAa52z3kMhh2fwMYcsz6aZLcTr2sKQ
HUsrsF8SHcqvpXrw3Or03MI7qxTkcXIvssoGEGQgaDer+VzTeUt7Acd6b28NDBeJ
sdaKxtgLD6wj6sQm20UDqT1bOwc5dPXoiiatu4TgnZrumshOf1wskFgfM1kVu3UM
HGLw4ZJ2zzwDRXFqaax4LkBSW2DGmvG14RpW10CRXtDBA4jU9Tup6KbnkjwMDFex
Po/FtB3zrBIttkEIpqCFq/6xB0pLae4FGei70Q0k8pUxP0psMrSe6r0Zxqgkr+bR
R+zHB6WBrk3wWUItyFbVwrpKY82sDYyKx8WF8qCnBinwpr8WAv0ZS/NscTz1lzEW
JY8enBFklkV7f1d1xf4B+zGqGXnY9+gg/MERqYQfHChTVClVt1GXui66DfV34599
ayDV/WKKoLFoA32UPYoUlmD6xpVZd24X9vnpun1HMAxyJxKqi67RFW1vJLpHRNYp
PgLLOqxWGON939tcKlg5/ebZN/0YPz+Gk7rVfxQ90akJwpCyS8y0tFvrYbP53Y0b
uwICIfts3enJqksW6NbA3q/e7ogqcnQ1xAetubSFv6gnVBNeEbMAe41M++/CKiam
bmN9I8wxuFgTD50yxZEomAIg/3ggYfFJendMXkXnogYSx7D/Y+sT7qyMW2TgoaYs
VjFxOsp2WnGhD+nv3hClt3ft6b2GQLKjYXSxHMxAD02A4xdpXQ3PvCBmRH8GtK3P
tg89MXc7rRbkdY4xWF8IaykkT5EKmyw8h0f/DA7W6OErnUF0JrWbATsrjKTYQgo2
/Cf1vW1vzvfkBoNte8eL96q2CpjutSpGqd/yTMjNgscM/wFjU7f71elPrEOGxFws
Z+W7lytGq22ZzQoYyr1XerJEuCjHlEntTsn8H3+yg/j5NGHwWapEM3WQxDXgPyAq
hUuRQqgvVTfVZN2btR2GQJeWFGkn4HUpgA/SVCA7V9Qfku9wKJ77hRWrzx4ZZBsY
SGifOhz0EKOhQch775Lv9L6nreDB9YFd9jewEoLHlAmeqL21SRMaZRC9a440qsC5
/sWzDT0WEiMSb6QPWWq1/6l4hG+n86zlgr6k20qjO3Ora05G9jxQ33lRQb7NlCNm
7DYePIRSx7Jq8cwiiysfY6jQdZE6GBPtu46KiNuHLQFFDW9LVev6e1UJ/LNMXrBr
q1eNM/mhlbFuTuhoiunNB1cUtvzuKVU3U8O6i0lDlWSm5DkPk0wQ3nC+ZrSM9aaa
cFMKEBNd/YGnrMRZh8diOScoN/qet+RH0XiRo8mTRtMcQL5VSQCxhlvDKI07D5Kk
s3u+K4vYLDtpaZpj6XnkcVqTCdRSM0T6UP0j2dL2oIMeGdONOD87c5kXeiEmh0qv
ObgJPqzlSDLeaxDX9BCncBqY3n3/kAcZNSn8bG2+6ora80PitRtXSyvg1lg6w8HX
d5Y5nf4enf0hCvjEoYoS9z/zDS/87q5BgWqFx2epWDfpyzMbObDYltZLcyMqss8u
ObjoDjcZ1BUijHQP7UOtx00fyzT2xz2f+qmKyFU5HdmkGm6zPvoCIQ9PsUh5ipVV
ET+BhqalZgiUUGfDU3GOi1p1KUKBjvkcdEQxn1bI17aJWqGgY4N025O6wW9BB7zv
IUXHPyBtFtDb26BittD49YxtsVSElKPz/Qct+OUd05zbNsCgFm4e14eV9Ho17aoA
dA/HuhMx+h1aIaeo2WgthhbHOs8ffSD2foxrBIQSO0X9iIJYihlqxC4FJ4XMLOab
zl340G7r9AbzCUzKESThriaDo4Ik+EQhzzzV1kKfXF0x7Mw2X0cx7YrqK2vHr1Ut
c93CzEKhArepVN7ZmBbHcGwte1xSp02cCwMglaizRlqk6HlTu0jwTXklF14X4NHJ
tJmhf8tsC2TwRw3ZWkPyPALHcl44RWOnAYhQVMbYK44ji9EYizB8oZsaA00WoD2v
enUf7Ph3DbL2vZODIrjmbGMh9BYSERc5x9zB+yj9Xv90m8hind+hsba3Wn/fGSum
KvzK/zn4aF0GVmmK/KljEXsg60n/Q2VcQtvzwboY44ykBvIFAA6yws0C4AA3aaOr
WcDdpHm1iuzEp+8s2yBuuP9IDlzWYIXpzucfJFt+ZfkqnTZLOuXQkvM5Pxn1U/El
NU29zyfdW79Y83f1FypFVFpsIJfODKyVIgoppFtHLDruTGkiIvyMRfoGDqYhYrJB
Xq9DXXBOphOf96MA7GA7cxKAI3PGGud+hCdjGVS6P2P8c1oSrr1m1volC1/lp3kS
TKokjw7RZDG4kpPqc2fTd/nXdIe0aLZ/dX4S8p1oIGAlyaQlxI27Uqs/RmVEifPn
U/wYC8FM9fJLQUFA8zSsfmyiE3czYEbq5/KeUIt2w8SyUUrrlfSmWxtYicwMbQJ6
UaB3m4TIZCpBX+sgxNRXZXFtQ/8aEnJgRQl0jVixOA7Y1hRU9NmeX0EM7fKaW94f
Jx8T6NX97woN3ywLI9hAYKN+LirWipLKHN6zpESrsiwEqobOsyXRRvDP+KtSJLor
fLFf2yk5c8myHInjmufJ1XJKQwmgIzGGfewA+H9le8AF9698W3sxYBA70ZgoMSci
Od/5J2Oq29EdsrCGwaKnDvg0HN4hX/Eoa1975qWcgbiZ2EF62wP4RskfDZiSHTEQ
0Mmn96WEbqV4X3mnu6KuMkc53N+Xbc6PvX6bMG8KWtMZAeKn4p7786fFjHRng6t7
+Z1WXn5jJnIu3JBbAaT4gjIdEDJPBDyfgpBAqPThZp9X/9dGJUZx5CeU1VLBdTRZ
H38GzqpSmpVEFCiAl0vclU8/jKjEvb21+B+RQVqQK20AdV1FhDXDjuwYHlH3jLSa
khhLww9k1lYpW4sS8Hk+o8pCvqCHc2OSShXwKKjCs2c5ZeyylESxAONYjdeJ1CaB
nGiXtrWVbum459d3DoODNYcF1GsXYnYwXX6B0IoSbIOEimwFOlgvPKgJCOuRWioK
/dfMulY0xa9YJksE5XnXtxWfQDthWKrSNQWFVISJ4As6RlXtMkTN44zOZzYIeWND
i0UGZ+BLTgpN0bLta4TSjzRDc3BpmkacXai/kInhUTRyf1i0Nm0EI1DdoFTh6aYN
ePPEhpHMtrzlXuVajczHOg/hAH+KfKUvT+O64YekszB32RWvwRkY2WBCSJfBC/uR
2SVRtjIryG2yXoHbZk9lpxkA1yCZUnqPktS1NGN0BEe2EmSWj5ilb2Bcv0LJEEA+
qhh/7zszEnVwjzkxGvdXfH6yCc4JXxRYRqgP+d7qBfp365o7vi5fgqo+gPTRLD3e
2oQHWCUT4y8LkQsuveoFikgGFeKLf0iyQ78e1/wVqoGe+m+gAwYYgOczO680hQ3E
4n8fI3dP73OfXaQhV/fa8jG03/C+k23YUKuREpB+7MOTCvoDZwR1IU2GiiJfkVze
iFW4QOY9wSmERyrhntdp8SPu6WkeTbo3PXvDl6+8oY2ux6rbMspIJXb12Z5VWJOa
l64n8c1rE3Iyq4yhBInRORYutGsOICp7+pQwo8B3UGGkZiRZ7YlNRjhekXQV4qOi
VhEUWkqVp4KuTDFsrjhNdE6droAFr916LGFvZGbobDnYJDHn1F+N2FT3GB5SS3Oj
lStuWyb9oRU2ZBYN2e+oeNWBc0PoRY4y/jACQaK6Jornz0XRX311e/jg8ZLYFoum
eJkKpM5Uh7oBjBLwu6KwBLSEmfjmGs9dTnKGuI5HPUbw2jC0JnxgL/XM0JcNtVla
6Iq8CiRt0CznDM4peAj+GQNjaiKot5iAIZrXdIDMt74tcl5MT9tatUL7WknHnEk0
FCcDgvZtXrM9vx+GnJjOLXy6PZHw470ccbYbJPRETAFkDBdH5kOHzCSAZR8EeII7
Za6dHczwd5N5oAkw5+WsCdiBDQZYqdGnQVFbTlWK3XdpOCaN04FeqVoWBafqUQx5
McdfF+BzcFDigMEYaNRdpi5HrYMBvBHFcOLc7043VT5FG5UuvIobBU7NyU5HVI6E
ZuywrnImqWQBJfiyEr0Kf920lG3MtGnuSibbjhT02tsucao613gIRMSrxuQEEUfA
vOidNH1PAf388KAJZ9CTdbDlC0/MKxcDPpyvU21ypwenenQLhpoJTdi/A6g2J3l8
irq2dhvYIAgvVw4bBFYJVoExauKx4/rNeGWw5pDpC2sqGNIIVy0YRkFPUdYl7kzi
K8FN0W5VaxErW8jYtuEttUR25tX8BXDxJ1I8i6nuuRCROv7ktDzffb6svQW/aegx
G8FuBKyXlAXbnhtmeeCawYVYEB2KmhGuwXi1TRohrxZnorOHPis2C6Nr1r9ATJJk
jLJ5axgGaoN8hevxoA/TmdprqRnrsi+Zbpmq3jotv43troaKiZz/usOtTk7yTRKy
BmXn8Vsl6nUaLiLLqKLqFZG22w3TW91wvsUE7IDeDGhYMoUpUjkYRZ3+tLgDl1Gh
IF6DiRiY9JtbBLtZr4WyLx+ALGPmXImzvrveF6gwQqArlyYLyujl+NUVGiT+UdKW
mJFc2m4faeWrpmfFDEA9GZdwzZAB+wVfGNfMNhVosT5bqWsXpgm1ewTsSow6oKPq
gyUmt/y/mBXVNxHpfBA4pk/oTNoeaUPzBPniwL1Hg39YZcjEpQKEKcqBevr9IgL1
fZ3wqfG9TuX8iE6cfrtVaFvpVbHiU6DxaB6tWEqz4rVWPj4Tn5qZw3QFzcnJF/PX
DaBPC5x3U56TNSo+xQUe+nJD3CO547WRn1yPeKGiPP9giDDmQx7u7hYETgPBCMeF
NBlT1IXAteogs02nj6LV3tbtz2B6ockpuYMO3dz5LheuJA+H3PhXix5E2TsORTvi
oxVOnjhzgEPbp5v/4TSDLYtEM9or2ldz1VXBc0phHcl/ZU4QPmXtyGsXgmi2zW4a
8Om1Y/cXcKVOpzntL7Is0uPKyf0c+hgzOS+9AzLRxE93bBBq9oFyGO2BdV7iIqsE
DGp8/VMFiBPr1PsGsRnzHr6NCl6WQNMlDFwPHUmk0G8URrCjuPNfoUdxF1TYV5vI
B3wUGuZxbd8ldv00GBx+2xnMl12aNOwF9PWQXNyBDvAvCDGH1x2kSJVlKANssimx
1jrPkAhtHuPr+zr0DX6HoPqWQr6BnPq+kD5trgmm9gPt9lEIVj1recEaFT49E3uJ
okvBWWtFNDBumU55hAQT0qJeftgBieDwgNr++8PM8PEnrMp+94pYmLalUS8ScyNN
P/L+Omz2riq4XkNyLg9/pqQd59Gr5pvyjRWGQPI+m2cyzEKSGlCJAJD3sWqJSqMm
Q64mpJjDiWGalGAjSFOuSrwp4YCmFALyJg8qZY4mg1WUMAXUwB17XHKvZ7nmCAGA
BkDzCNerWmA3ebo0O+atdZFa1Z7ByTQ70glOqW6/xdKOV1uiOWIP7B6eufPJKwYM
6bmB9ivaCqCTHOjYutJVUEJMEQQ6yzxPTKeLm2ITRNj3n4r/VO7O7Kwl8853IO0R
zLGCW9sSSuuBvrXss9Qe+7cseJge/UQJXcLCc2jx1ru/2gRHahtEoqhC+kMxYfyl
P6LIc2yYMnEGjD0Cy7R/bvR2ELuO3qTVcriF2fB14JmnXxPO7q/GUrAvYWASDewP
DAE36rgznNJL0a+xAyXD4VVTLVSkOpfGCyfy7YkpASaTazRVtG8Sw5Ekby3FVulD
bxy31rxjwh4ADhrRfitEzpWmsjrxbpP78mJjpq1VYUCjxwvfX9vUbZTjSmlqaspA
CEdKPWc3/DqDtAVVVfFfurbFYSinRRR17dtNRjdceSokEn5Wwx4cv08Kk9z5N4hj
BfH+V5t+5cskaLDI10maf5RNDhPUYmgF2lPORE9MIK+jgzwF/wAwvjdCdzX8pODK
KlniOsYrw6kbNTDTum+GkGNgFLZU6UtrttLNn42NqXoAF9YZL17HWAEzLsjnhc91
ioUZyyxI57Wkgnh92CmtUga+O14fwKbktggqSMXcmaBYYWzGw0V8DkBHhce+/GsZ
orK28tUuqV7dqPJrzEsZIRejZkGG/r/kj1wiP/6msUkRMzbP/p9JqyC8bx1JRAvT
tEFZf/nDA8SZXP1DPxeCD18OcoZ+QULjoNuOw2aoDgM//IEL4+nWfbMJT2MGQDgH
5czBymfJ4PI3Cv/cbBoWiv5H6S0LjFbQs7Nd9G9SRddp7LRlblcAgm/66+qvGSPt
hHnXPzPs2DCF5LNXUgx/96HhHIC4UbJb5bn6zSCrMw/AkM/mVaIgsO3a7ejNg3iE
0yZSc375csI2E8xIqqmkmPVmPumKhoj3MLsdIWfp6qmKfgHZbXJi3pCmssJg9eMx
/SISzRB5MlEoykPPe+PHDUzXMNqgcQlICywNyY13VXrK8oqcco8UrCFP1uhXfVVm
HVUO0Jo/Gnk9tT8WHw5wtvj+np213I25++YSmoDXTednoj1azKRBlY+2irSMe+SC
Kbtlx5wMnctcJlg63K0uL3dvkOPSNyZ6yn4YCDUO3637zhnE5jDy8xaF0DwFZL6a
TUlhOwS8X6nwY5y+2MFU/vrm62CH9p77xtWXkD+AKBi4QbiCiAoj+Sijbs3LH6p7
uzbz+eIPsubTA4RX9VRTi6YMRwttEvQNqntC5cc+zN/bp0MN/zokQaMFvXvqGgeD
fMYgSO32h75AbijDQQYJ8xQlaQ1yi9OdW3zT8c69kzAwGnla4Z/uHjhaN3aq1DHe
dpob8rjbnFFWYdNkR32/BXnUaYoBecwDYk3p60A3BCpwZ91XRTPnwK5WPC7kWauY
K7iS6D14MbLGImvY6GXVf9GlWsVWcEznPvPQ90s3BECCuxeoYrR1/sNn8JKy6wbi
RMNAvOFNCxisnzmi9N75iLvmNgd+sICaN9kbbFIrx+1sydII1OMXJuusaRKrsOMJ
5hH+Y+KQcUIWROs3ewv2GirdNOj0J+RhvyS39waD/ShIGPDnxW6o2h0Vv/cYezTf
mgeRX2I4KA98gP1jVYZEbjTqLJeBwtAZjYaH6pVpdaJZhzZcmqtRPIR2gDKnpb3u
X4wSkJF0LFSfujRObJsMT0qhsZEx4bUZM1irtvC3UMLIzqYyLnuKPH4RQsGS2IXO
qPf2wrMSl0GmnPuqOOFYxydxWlltxE6xWqhES0BHq9vd2m8xnm1SO9wjrGuRjF9k
AVWaviQSWHwI9hnyzbEbcYrnlCsAscWIGiUFkfamldutI7KAiIX4gml0iX+bG7bj
CHex1TiQjJRzJpraLZ/B7RbNt0oCZ0Aa6FdGNY+cpcgqb7/MztTTuZZITTqGo0nl
ysXkp+/YywvAei+md7WtA+ym6Ad9CNSQYb7dOwVb5dHSSHvoXYx87jwY/IHoGis0
pXXQQsc47fUCFPeCjnaGT9LNIqtlKLr013EpLp7jt94GBWCvWE5wUYL5iF29JWTX
gc4VgoFEkWm/jX1gC0sDJJqfv5TcLpdGdJd1/iHd9lTHPJQR+5NQ0X/ISdqRSAi7
FWRMOz2N5hiNUPFwdmbQ4+d4+GJvbhO6b7KmH82ZUSal5hrzWfKVyRzeK9UciZdF
5jxTdHL1A1IJYkZf2DSbTb8enb3fpBij0FhwluXnxjuh4219jnzuIUIgEcj/Lc6d
RqPeHHflq+bG+1kjlr0qjP+RDoYFz/FCVjIwYuyxUCSyxN4kb6Ct6AIGLNyPN4v2
/M3dRk26pa/NNBLNP1Z3ZM0hdvPyhek24WGlDR+2HO6ND5iQi1L4JJz6Um9ROhBe
pzqcp4nRU0QfLjcOfyY5Hm5JQc3g2TLoJv2lX/CCPm54xOzuGZEV1gMuMTEDAQU2
+fJ1+cAh3/8nevheijQWqNE4wTok881ZrJfUoZ/RAOvlAypyPMM7iWpw/eOCagQl
w1G0ydM9mKdH1rgXGPKGpRx5oeXI3JS51b+CNIbWnVdB6naE/zm5wclhkXEWeGhy
aDXFWBeHxFkkHl3ug2FTyj/RxaKeU3yq9hXIeb7fopvh6w6KzsVARyAEjm3j6Lw3
ea3hVpuwd55LyPbAY+RNhmeiV/gcUBdlR7mB3Rq7r8f8c1dhj3wW33uLvmMOkUdX
9TOePbd6RG6iDwWDF0pIJ1HF2+Jf3mqJKbSHs2E3h+duCZTp7SlcNBVoeu0hfIbX
eHJEAswkQmMAMwKmzXLNVl2lvPdEMZoPbNN+nnnvpDCwh4Vi7z/F2S0++ASRERvD
3wwc1+u3DwrL/j7VJd0Br8VYtcsTEDpeCzIAsDyfdq4d9fCmi87r0Js5KxV+nahE
rjqG/aHMhufLmIGPTpRFx+EZVm1IdOfddisQLNjTFR019rbFBHQLsDg2wdpHlHXv
ehFa6yZyWXamXKEvWH3YZidAE06CmEth30jGdb0rHQHUxyHINSQTqjwfWgBa1JQp
UdL6YQSxNzSYve94KTNloK8hJYgxMs3zJ9HCUdqp74J3etMoqBuFlo6eWWZkIp71
YB6SmfuDqCrAjV+4QdxtfIu3uiWL5VCGfHEyXRC0RXFTW7aCVTq+o3Er13oBZ2sV
VGHMergjPD2yb4ZvSesSjXhxuYovKnNxb/ZI9uqUwGK6Bcd/wVq3WldeGVPrIOJc
iSKaH0Y/6+cGUkTNAn17nVSP5GMVMevFAHZI+wKwkJLWcoR+cL2w8LSiSWfbmjsk
aqdSmXNpDOatk82rhSJnsOxFsmZgvMahUtdUS38MwMpj8IZhBIUCVSRh28nQfiLd
pq65Zv2TZVHdsSfTzBxRT+/0VWuUcKiVAUx1YJqBOPWd5tzU8v82N068oYsJqx1g
qQhIFluDYT9RYym/ZmfVrXsp7k4enD9trWuVJSPE1rJZzIzuWhwucQKy1CwpJia9
kOktr/nO4QrVCmyIC1PbxnSDbvhUgwIQFzxFROO2YCrWqOMhX2XddFEk4tGOrP7d
Ace+SW3VcnNeRiQOMSMftav4FkaXswWPdNaysqL4oq0MHic0IFbd/H465/Yq8jou
2tazEGjD+Q+otlbzn6VzFPP1t/QMN9H3nsmZOHh9gZO4NeVMC/SKXiWB0+vM8J38
rLWbzaCdw/JOYEdnT4l9hOe2GkXRoznCpieZQSX75IHHOJlw2Rom74NifvsyJcxK
Gpor9JNtmgi6dEI4Yhy9NXH3AwrffwtJF5SpAcDOMHUIHPEUd8MwoXBsxG5wLFp1
asLprGBGB0j2e9GrpVwTGSSRACehKCUoNmqDCi1cStmpxRFF780qby8F5n572vgO
VVZrE5qDSvEZHhS3qAJ19zaOfu0sWHzBCN8Z5lXAY1eoHAMNaAdN8FHEl/+3oS2C
wMAD44FgN4EQFPQTUrbdsL6V8rNoGPWf0dnV8xXzsluTBYTlGR00gEVxsc191UEy
36xzZF3ZGDmiUNL3/F1eZCE9gBniwJiRjPjr6o7obWc2B7s3mU71SjNfojeLbTLO
6bQa2Uuq5OjadGxdtU+jG3DVOD27vYULWZxiIPf/Iqyf9Htk8aan/VjedAurdtn+
rRpa4nvhZlEig3H6JkOIqhfpsYDfETdDJGttMZBduZcXEUZTAemuvgllGiEqPzJG
4AdVDC/1Ruz4+W5AHEEd8xnrfYLy1tO4gnMumVU7u+XBeyo4Y1rAfUt4qasK2vM+
G3v8/be8cJiM4VX02w/YU6JJknDgueEXG78MPSdQL5ImbbFP8/OgDgDYaSMFt1Op
cRJffqpIDdQZ8+qvV3I+og9mJbtrwlzCxA2VoQXIo73u59Rso5sXFacp4efJEgP+
m51jB6I9a8VNYaBDxARkPcLUbAexmhEOknZC/ev3xvFbCFBqvy8vi7jHhLxXH35W
5jrJ8Na3mQljVuyxwUiK+o1cuDAIpMZlkL3DljKOzxJMcQC0t86vNoFrM/zBBoXK
b5c87GaNXNdicKiEwKiIZf3AHfexAd7eQ+teySuOFVMyUZAmSRcyMtbMQMcKxLlw
yaf1esn6hns6SuR3JPQTp0dkLDbCJu6EzP3Mds7uVTmE7IJgR30dFl6vcQbeh3mL
ft6N5WRJ9AlQ3gHiivpK9o5I4/zRWLi6CBHdOMtXqoDgjPVeD7PNwix7lVJADPp1
lKfv8kWV974DjQaEE7EefcoDd259anGzbyiFlj+a90ZEf0pq0dTnIOCOZBr7tGrd
6xw2lSLFavY41tCFXPZFdd13ZlZkFSHwwQ/ef93R0lhs9MRA8PoeNVQZ1v6GTXMw
n2PKyXwLKgVUImmXtJjQXPGcdyuuN48vcpi6Myd1znAURqkXuQCcPqQEvAlqookV
TFOyZibjHaK/nWlNaB2NJRcUTvVdJq+Nd4EXU4RFxRNWnjP/5EV2f/mDi+lVSp2g
zRwTGPfU0g6otPcNge9ShmAnFhCwy6I/ykz3AR1jt9Ac9paJVyKQeq2wpvdSJuP5
t3GZCTIu5Fp2dVpeOD0xMOWmd90IJRzhYphHlYSsvcnZKnK+mZelXNagrNSYLhUo
aNPmmsdDynZ18N7729X1qLlEXEYGxfdtPVUBPykqf96a9K6eiN9FGmtcE3wKx3Bj
ji7b4YOk0vqsmGWae9QqbewhyNCJL9HLHNuw0+L5VY8G77942LjLbNXN5/2/f0VQ
J6Z/U/3wCNggjb0W+ErGRP+9rZ9/s78DF8zvXUNobOWx50RVls1Vq1yIIaVKDzvX
RsNcMJxB9mHAyrwitv+pqzxMw5PTmd0Y49bKbze0W79iTAJKqNAkTIRGvQTNAdQg
yH6atldlSAybC0zJBL1dxKn00Mv0sY6Ii+7bTqtTUFrdIqGVqRANgsCNCiaPyaz8
C2DKrBk4q0kD2Dydx0wMM26syiad30XN/7ARt+YeiXc/D70OZQoJrC9w0RbdYsKm
y+IMo+3x8GJQa/vIWZJVhNrEFJ3QFOEHI6yJNSMHF7t3GYcK9mYfCMgfMEo2reoA
wF/0fi1XCNbDR+3pAdODXjUWYyp+BwxOSwVTNimaHOZrdzLQTqaw21X4Rsx+iEnw
hP7JQD5C5FrEmhh4ZimuKYbQa3cVEt+Qq4zqTsn6zvDY4W3+ub6Pgow1cc6hYJGb
W+6QKUdjZpq1hBNj8y5G5EDYN3n5ckc1EFIjeleuRMQemBQu9ACtdOgSDjyZFpvN
8J6HZHphC7TY1GTWZa6Yuffv+rIA9KiBjP9wC9tCNjPgtQ/TY89UZtlcC1YkFUIw
6l7lVX4jPM+/1UdTI7uszDDPIW7E4cK1iJ42JLoUUIrxxcmK2Xx4fHMR2F+91HyW
barl7FG1bD0FBOdESmh/MYvhdoLkqlz0bu2P8MpAhxunuV2WQAbaa3SZ7XWKKUrk
elG1lnYxCsu3ZRtnuYyOMt4f1cTBbp9FY0CF337Cd78cUHmcNcLvHO4KUROpyI4h
On/DjHGnbOoax0qmrx8erX1xFPyOTpydoJcoQGQUhXEQUvNCJBCkmp6qvHPNWwwf
kWLF7nR20Umzl0jPvTCU/qTcGuYQObcF46nqDNy2sDpeUC0sF7hw9RN3+13MkfIz
3KHlBCWtUP0Ot29OQMioleLPN/RVmsGyrOzmj5g5xQpuVJWuUJUlNF6r6xUO9LEm
xIkKTGB7BvsAvFGuJ0qf8l+fTNnaAwvEaWc5f3pq1O9MNgltAasuXNdeORMVYZos
KWb91r92+13mqlQi+ILHzPkxQIZIPRL1WHxaWbmW2rKBjc3UMZJXz8OQ9LZ9uQFx
HRP6mwn20mdXMKnTEh+LKVtIAJXisUK1l6KRLcBe0g3Rvzk4FBJ+Oh2LQtKcxjK3
+D7n2Nq2QEalbp/DtBypuMg1H9ywF/ut90q8jFAvGo2iJa8Qdr1Fe2BYa+gGdxD+
X3DZs0T5rLQAIG8rPLRD3a17XA1Q1SFn2gpfwQPAoMKvbryD4npdeVoLWpA+lcPC
mEMMpcVC9iAOpCXfZPLaLIo37PU3C9XfZwHnBfuY5xVdCzILVDrHLdOacuE5BdS+
TupwIiWT7EUxuQB6aofgwEfVT185MNBvoCt2LZ+u6uS7P3QT5k8JkPkx6ERr3Fee
4zECjG0HnGubbKg7Wr1qc+OEQR/o4e2otYweSfyK7P/8XHaumHP1JlIBVpCn8UmH
/daLYRFtMQNfl5GH9dljSmPoN75xKhWXyZhmttAw87Hkd4Fnyqop5NqL+3RgS6zS
drN6zjEBKViw05ipGHGhoGLlqKbGcKT3IK3kxgB2hcM2kfEbYnzXXCW0aOoRkkqR
TJY6aNyfmA/liGy39n0pIXSJ9A3AvDNLtc8jYa2KAr7lUOuoyZqMH3FcQY7A5v2i
uySTwWFdFRekrSJNCAyRKvQ/MmjH0N4+iAx2/Gevwt/v9mzlaYd0r3En4Yd058V/
YvAYNAMCV+GX5sX19XZOj7QMMwmwLkzJ+LUpri35hklI8mcgo5KhG5zKiqXX/3A0
HnORvXuigSHWNvXRhdeHJvdqd6wYphwFqqTF+OMwOMlF0vdcpkWbE6pRz6Y3tWEJ
yW68gVYMcMyqdlbtQmd3s2ezh/70S/xnDDMZwqtf3OIFo0Un7OJmH5+/1ysvqv4x
cjSxnDWVULiMSoofduitejfW8FF3+GCGa3iZvt9hFJeRgk/bfxXVeP3D7aya71OH
OK+lL5pWFx3OdvvI6erDLH7nXzCC+AwEHLeQ7T9FLTCyRwV4w2sEUwAbN8ljDbza
irKUcrqEeKvQUDBfUL+xKIf6VafZtMzPhzP563+Knvhv3pOu4nLwdexQKjsScbrC
1NKxxpwr/jAC11NSjBVIyvWqjrrE7iFFfZBE9xS6r7vtx/Ermh2Avvrbm6ZcAncb
9NAbptZvBKTOL1mi0CDcGwA06DsEJclyYYGNBaWTeHQvcoDORodDr8xtpaFglQgt
xlWOuPedlaQyeD8tA7LydK0+laSIfgQ/uAuwLEEGVG036lPfkvnNOfXrKktMOV0W
6otb1q6aRqWXW9MU+9rKLDmt7lAYzr+T3H8rszims6m1FA8fwHf4E90l8/BXwNV1
gXypF4GiUr/nYnEgIY4TIV6yefxNfbHg0WsWHSTqMX4h01VFT0YqePAlCAg5I3n0
ZWKh4zX/xt18/YUBf9fTi/CC25xLtbJbwMOLbHVoTcBBKGdOlhh1jVLaMsrIvlOA
BoEq8Snr4WB50gy6JyVviufzBDj98UXAZxhFK+dZfehxucgodsVcLWp0yYn80BwW
zjjaz2M54Dv8vGmR9RauaTG7IfhoNVZ4LnOkM+aee09IDQiF0hm7BMqR9s/xVxUJ
izZwP6YbUrSxaBPybvTwdqzFppqd3vFV2Kc+UNno3LOTap9Gv0AP8dUfEPVO8UcW
zFni+S9P9GeCWEkZcX6rlSK4r4j3Z6EGp4gV+csJWKvrS4NuhRaF/1sbEQljzRH1
1gGEgaJcN8bi1NunwPaPSRoFBvrkBL4B41sAlVORaZtRB4p3l5MNrrWJnWhZXSId
cg4Jw3UbiaiZwVw82u7K7/83nutCi/ss4cyavzsmkXlDgb+HNgSAHAtk/8eDDhS5
1UAKJnyzZ7DzC2nCtir2Ou8ughCEFz/zAnwJZ7t90A3Jg1YkUUato9HdyRenJLpP
Qh+imOftnuby7BQx1eigqyzfGr8zH/ktJjZwpyM5Y8Vh3PV3Y2Zvy3hAjOZt0M5X
4QnwRD9xOgsw+S5ocqGUp9OCRrKP1iNYFc76PxXIvR42F0HgZsMvxAkmVuok/amE
xOlsJ+9KLCwashW+KrWljscElp5zy3U0jyivIS20X5lt4zzR1HpVuRylLqcWlxle
+0+nM9R09eECbmCnRstJ+v8SX5p+uAN3vYtVM82XMJmTQJpDDbSDTiG6A8LFaHdA
JwT+XRNfZBSfUcwXlzbW5+eU/Enkl9xRHZ30rY+UL+tiqUHSwRP+ltonA7LZ8BgW
f59+rFg0VKCc/34TPVqlxuBxxKqfOvsImix2OILbnlsBF9ryX/M5kABTZlIuNHQq
e2i/3yrkf171RdEOinMp7Ldzx/5J95u++ajndXQo8tjBjxboBHvCgWPCY6rRa14g
2w995uSQT7O0xC5tKotedd91OqsLkGfnZi/BQCwkUiYv35joWNqG7ifUF3Q/dIue
kuPcMKZ/tFaKNCDmXRgGog/CG3578MyrhBhLqA/bUADlwmpdoPvYdW10u4gDL1A2
0qhW0dEl698FzKEmbsgzFqobCqLtI2P6a9uCtsFoLrS/ZyJ3zpkogs0csvbaeMV7
yXH5Re5IVF9NSzs0hU8eWzn8fX0sRTV1bhefvXEu86p6oPlvaFuo2OAbAZXoeld2
RBuCmCw9mPLgmpfTjHzV/bQBrM1Z40M6l1kbc0GTT+s+8/r/THuMNjDqpmAsIBYv
/QoKvD56yOmZwJYFbqAmpQpqBjtY5BTQECH5Co0n6Fw1fQzn75KXpTXp97u1a1Dm
AFQPcqaAr2x4Md5ef5ktx8yj9jauqUEQtMQyV+TlLWwyRNvs2Gn05Vp+JRdhCt5r
EpGcvM385KU6eTgGF5KYGc3ZwzCzVxoL3GpBmf1NzC0M/pEarZBHI4NbYKn2ZnOD
Spxd088m4XgyueWGpUnM3Iy/ir4K+i+T+1XO5ronzRo2j2jZDDDkqf/ko7+Bn4G2
bSLNJ+AFLwYPy89t8+IjSlSdKnudVczVYv2KSr2M7OdgCopigoETSxJGL6cMyf4D
FEib32TtaLRXwPzQhZ0znDxSVEUZijMwPNIj0+e8afqVTDjUuVGFTUO+/6nCYUvu
LdHB5oUKFChKjnunGxDktUTe+de6PpNolvCLZFrBuOxlqsak072ysL9mhnTo9czA
Tp/ZcGSjuc+z5zb8szbvhU5Dk4vk4LdYjTJchw7uvc/aWaD+DkMOs3ObjBnP9OWI
CtQAFtvpEf0ZspMtVZ0/hkU1g9aA4eGlIcKigF/8DDR6wWSoSgC0xpd2EEBh3K8/
oTZD2sx8CMCBnsDlNCnRWNPo25qpYZpvoEnLTesIW74J+1kawoObx5JfTa9D642Y
jgEOcanaO2Si1aTaevy7HxhDDLwAPEK0SeyB2l2G0LDWHtFnedh65aJkAbLkduuu
eZi5XFewhKOVRPGop6Sy1Ngufd+8SFOGqZ5xk3Ptoim04iJ4tDiRj8ahX7KYoyzy
g+MTq4z4vDHWgHm62AWsKc60npJOyqHY/ms9cNdTNlnApfRdrY6Hiba/NqvoTTFN
Q+FyI200nstcq5ZG8cN5KbQnINjNdGj11aHya1myKK28rLKVrLXnlynI5lCf+0Fu
5cMEJaO30SUul6RZQ50iC30F0uV5zTAjWaQm+aqGekCL3BGwMy2QPaK57OeoCQLO
FK5eEkcDUdsRvyoI7+uQXIlNYUp+rZXUErCRm49CIVJ8B+Jjgb9OOndWH/yLiXCI
lUEIUOCcjJYJ5KNauyWl/ddtCR2piFnN1a9LtEJmzZA5fYTMqg3I2lSwspKQ+644
PUJGhl7Yh/Q+wFoRwOlzEYxi5M9XbqOkAm0NoU3TPzkvgz4rQoq7o8NajjCiGhrm
tV6c3QmhTmaGESAhcml2w4XTXNdZZ6LY7aX8EuQ2TOdtJiu7irYX2X3dZR3Qpksz
mqXkIe1I5MO1em+WUSWFhOOKfZEbUGfm8VQGMhsqagZp2/adRDXGcpzCuhQD9tOE
U1XXIOqEdpb/AyvkI5U7jlJPbkTEtbalc1bf6iiXDOTneoPnIX8VpUAroot7hspx
QgliCQlL4NdVsBT7zvwWFCNsNgcmWza143TEqNnC5b1l8DJYT12aePfuo8Gefw9O
h8vzTtDqIXBf/NYsSfpxxG1hzRfnNrc2bCVhcUXiMYCyoFjtLC0I+44dJ0HpNl3E
+nqZirwNaCZvDOH2o/U+jrOpeZWvht3BHmoueDdgl38Nu9SBhjBQ8wFQaMzvyc+1
cR6HCpCBvO3uEA8hldJC6u5S8W1N8yttO1dAHUai4o/4Q+B0CDJmPJvIjrmHC4KM
EluFkHIzisPzUWS8AL1ldK4i1b/JA/KzRLoevxr1VDaExpa4qe0Ra5kDR3vDy7Qv
vRJGBl4OropAJhKQEAO3+tBSKwzay3ekl2RfnhGc2o1jUlBSQWZl1L7YAB/NIPUD
FfkNC5gjZhd5d5M3FI/UOOkAzq+zEYXAMv+43RCmRp2q7QkQXDVYCZwfHFEw3RmD
Nt4V345NWIeD2leajmxP+N8HJPiY9fqPBFxxYSEoem8TX+A3qicO4knm7Rrnl/+h
jiedAptB2RzIkUr7wFcuwtFRKlaacz0wjxYtGTFJUkunohgImMO25UNufksbjvNP
/YWdSdjWsvp2SLRDI+eXxUeUDlUyJcH1pEmWXT6O84JDmebzw0D+Zfd6V82Q0cC/
Vw/DozLDye3DZlCTUsMf1dTC3PWHkE+lJlqOKjoRjX52RoibHoran+5L0Mcs/xHw
NLyUIxJ00H9+WiNVFS8YUEuG1czNYt6y0KdXPn6qF8d/WUWDzNPC1qgNvvGmAi7r
eClzUEMYIkctt58PUlPEDPm4cNIvr9GO7zYDjN0uNurVjp9N+U6WLCawX8TwhQY4
Uu0aE9AqBVpVcc9VL8MrhqOxCP5a/8Lge1iHtEq3OJ/rO9eBsMeLEeVqPwNy3qnS
QdJhmlmaQ/mzeEkQ40iHEpAfQMTjpNN6i6JidmaYcQqfMVoyagiopLL+YSm5Go+n
SZ5Qh1gXPgDuPWJSbILeWmcGRmrt9ws+9lPP7Rsnfx36tyXqCHhurbb2CIBsSSzJ
GMEnrIEzXed9CpWhdlMYAgJVk/z7wSMb6IBwCQxrwEEM0zuyqNmZVeaarIUqcrdj
g6rg2klHT6SPU7sBQg6xkE7NSbqO9kUpz2tVCS4Ud43cVMali/7iUUVjU9BQJCfB
nVb71cpyIqos2MEYTAI2fzxG2mXuEh2tMf/8G3ZJm7iZ06KrdSSqK9xc3iu5Pg2+
JwGaOJCa5ozwk/UEKIyRPUVA7iWw+HSFVOBGHBdGl6/x7nQ7GnXWBzVNNTy3JJhv
zZAIC9qSYCWMmFv3cxkpaJ7mCADy6TSqoVH3MszqDW391nJndE7XJd3SLx5MqBB8
XkiVF6GN6KJZYgzD65SIfSJgS8giTcOUrZfUznQv6qtAPpkZHl8lHljavkOOlrLw
fg3ez8XF45EYbEk0WvZtAAWglKGF/4wZJXFdiac+guqgRKWDMMw9DaSBl19Gkuaq
RaaNMtGsBs7TlSyGCYCkrnY/+FFY1gBg2xqKPfWxSjsTR1XkdhflLjBVc1nkSJqj
uK8pSRrBQzYU7UD/vtde5wh2Le3eyBq53ESnebFRF0fzlM6jmHmQznesmE8nXUFQ
sLmG8xu+P3QthGceQzf40/IbeSnNG1b3g/AP36ijy8zslaTzAXu7BSp1p1k6V4iL
9V40diPA0TXAbFJ0MNQZs72HpWW1hlyJcLKWjb+ym/tT8tOjJhFdBO22QvgPwU6b
uY5Z4dIcnEd9GioY5zg9HRSPLYPFJp714TpmWlmPsthUf6duAFz5XTcDL8ZpR8cg
jqVwIV4W4EqMzIT0kIoYzlX6jFOknKcjjJYTMQSsO7QEoI2LUuMOvEmtAgluFKaP
5tQ8CIpbg8JgujuOCAcfRPexJk2uTUbsLwTK/SSQ8AaLwiWEn3FBlgHXiJmHXdR1
mmFLu8/IXBBO3URaHrA5Uc8TpXVgl0Zzx4R8CTLiRyJJuPRx3JNLpLWpKLRiqWm5
kqFCHrwYU01x5w35JyqMAob+HSUbvlfcA0FTK/YPOo+iZQvr3UJrAyU5qQLvYewi
DFcyi/J3p+u4j5/K9x9jrQGLLUmU50NrXQglSrBxE1DXQQqblg58s8qDmgW1u7rA
I5zFBXBVYdhRkx8l/mRMOqG3Cs5c4qtb0lUJTICaR2TZuziBPgh0nY7vjAxxt/Z4
/LgQ6w4CQn8TPQXLP7/pRQ6/hM/iX68CKQiGi1MWbNAa/sRlt9URFJ3KIB0BqyDk
/+sM/5hbHC+WcYIKzZYNL0Bf2TDn7Z4VL7k7b5zAKv08aALu+jTuw4KzUsYn8CoH
iCsPKEIOTPa9XBfPYrdQPdlt+unqwOic/ihIaiW9rg20qs3iHnKux4VH4oOV4ysY
pU6bNRh9DnCNBuVvCf93/S6qO0wGHCRy/LNQIAljlF8P6ngmNcL1YIr1olr+Yd6P
DbtfWTaEYVvzJGWev9lwTRDoggVg6ucf6zVoF/bBbIa+/SP4QJ+sGIhsu06+E1nM
5FFNx6lzuPzpHf2bZ0g7l3Gtp9HN10OhqZcGMnTrZCaHyfddrxn+Oi9yevwIFrMj
idj77x8KUajk1m/HP4jS34rai5JDA67f0JYC7p+aaiakYwnkSQCJqJCI8/OsiJbV
SzmtXTR3M8g2ipTjiMXRj2QFG5XJjzg2DX+TcdGgJ+IE+di1vA/Gi3w2cbLU7Ag8
dFlIwR6Vd15lCDIkRmUhL8LgCybOukfElxQGpqPFafE6Swl2TvPqRR5z/NxBOJK6
n1Ep/STPf8N188ZuPZNDGTuZvrcmqIFPukZ45kzg9iMreWqQb0Cf3EGnt//7SRY0
u/eJrcXPD+bKxrdpFTHhpn2vnXvUuGug4VVnXM+PAVqYNEkKJqPHVYsoOSFA8GKY
n2XR6TWzoyqiiKk6hHBqDW20vn1IpSQ7mvJmgoPXfUCJOVdSfQ/+f9d0jQ3cWmcm
rp6YmBGKErk0nWhU3RWiPbjXPpiuNEZeCV17HOK3FuFAiyRWXpain06eLxdVnLQo
zcSBgocqXaVdIEc11rTr5/W/ZEjH9CD8Un04B5KLzNAMKiXWz1wly9NXFKzbQYB3
9z8PR4pEPt77NDHrx++9d+QVI14PVpMttif7HKGHA1LYpkY/z2S7zq1MBfq0zwsc
DrebYTwqflmWW2fjI56iXzA1IYDEBVumJnSEDmzfpkDHxxz7Zv6JgHI86ssWY59P
8436T8OdIHLM+ZKg9i8UUL0qwmHvtiNtWTRcE1g2fzhNzVQZCFkZTlvnZPjEtLFX
e2edtmpsB+fDBDAZEognDS62bgi2KO5nhrDoIfPCM1IHYfIutIynWxxE4Sqpi1k8
EnbSe+a789TbhvxRKUR619d9X+n8nEqu6wE3stZE8GdxIVpqr5g/AOIi148+0CTV
FmHcZThbaZhhT3zyZubkme/saEYhxvtT/hPQFbJt0fHNWiBoAOG61B2OQZhlDtOJ
fiGP6HfE6Fwp01TKpa+Qz+aqCtUFrGGAYPbqSnqgvXDLPZqgPoqUwqnOhzw2DyPz
0JwfcTkQzEC90H0PbQAtlFmzSywuN6AUwHPSV/I62hULlF9/sTkCGNDp8/b2+lCN
la6+WdSbeJdK2Vnnuf/EKro0R6vqi+a3q5IjOsMUWSKnCb5Ca07Hcdl5R7N+HSmZ
U/AJe5zCQSZbLNqAGyL0HqG6gcCPJDNUqoZhuIc5CRxomUjZxOW6mdOXS9GYnkI3
wBTZlQoiHp2dKHYFqsI35AScS7XYsqDPYBpCh2IwIkVYIjoSzI5vjs4XUTemZDb2
6erIjwzTVE9Po60RcLGh2v186Fk3M4Xt7GVzkwJ1AXsJm0qVGwdHLjJhewvZxPHG
ozmMcXXJ/aQF1+XKhCpvOMAS9dqfM6/LHZwdhZeO8NJHPnIgMHexgY1UI1k7sJCb
9to0Kgz4HyFyKpDNLWbpVQD4fH0X9WiKXTA8yY3XSSIx/yQsml5cPE+CmMUqbapF
sRGKW3xI3xBvGEVcNEJ2v0bHxwZ8aJnXDWREFJ4Ab6hvBY1ACmvQSaGaYevkVO4K
4LBXHomfawaZZ2Vwfvd9LNATA0GTi/uC73AG3OYjPq9NZTHZzKJ3d4cGJNEsWzrH
jDqKBmndads4kWzamuIqS8P67wiQ1c432oCE9i0L3HjMFdbdal2Z+zDD08+xnpAJ
Ktdi9Lhsz5r0mnN28YNMftGAy5pczg/rlDRV9Iqb88xPPToLW+SyilStGrSgzvJp
xePagCyV8pVacRRQLHs1xWzCdUsyXdVC851x2snpaoEHeYuZAOmPhQPYN0Re584V
0L3QykyXFlEV8jvIV87wYCDsDB9vHWqOcY/rPlg43Xk/H2xAU2xrDJhD2XqeOrsm
XPF2VBbWDNnx2KwbBXK1/A/B+dLMhkhGw9lEanywhNF1kRwmGgZ9SnLK35LXbEy4
61vsagw9/ikepcQ1c0R5seP+srQ9Yd2Nid5II/wmqauq84xD4zkohH0eNyCnI6sC
hCL2TYBmgZ5t7jhS4gi0HRD5Nb8nGJek0+uZivcZShGkmxbeW5hT+odFlsBR8yc+
7IcF9GD2uSKuWloCHUk+9iibkYcJIipKlzTKuLnLOEH4Kb2Adi3kZossmd4R8Mix
MMWlrent2ax0nHX4uaBJgPqrAu1Onie4UupAo92jDOkAcAEvIKhdtlPmOv+/shHn
mEJZMoUGOh1mRM3dhgvABXcq1qQKQJZIsTXvoefznnsG5mImanOLY31JPa3qUw+S
JbEV5Ghs5+mrp0lj3E0xcQXfesJTt1L0d5874Zv22BNBAhWbtXDI0levHYdHQNlS
GTYbrk3Yzt0MHFfaX7vDNSbEzA8DpqYWdMpfpTL2KLVOjm63TN/VtnmpCoM77F4M
qzgWnX2WBTCuFOjPjvPdElYSALbn3n13IcJdqXu30gsmuo0UmAWWOKII02snKqGP
9uzBBsX/bR+NMKqvbR51X64TrEO0OKaN7EL/X396GIUc87UZHgsj3OJEcBQ3a9eB
ebRs2Pnc/pnc/VpSScvmd5J2TBdSXOI4DMiGLGqg01ROiFXiThv9GGYl42isaCqY
EVpqc3c+/bZtHYioQpnn8AveIH243k7js8cbjBYN+dFIR5CHQatSme3fNvuRHncM
N1b8rtPXM6AKcZRgoj1jcYEN2RUPCBC+Bh3zM+4csZm/TfkxzNhcwngLJ+dSE4tV
g8zJCOxy3wEgR4CmvP7AJTusCuZibay31hMkKcKqgY0hKptnD1pUJr3BFZpCn9NX
TsgJ6dknSd7tTwVXoRH+ySCP2G+0U4/39LqVycWT75hxKEmZ972BDIWyxCnP2yr9
ySWHo0AS8wHQgsZZNbvN1lbG5V1qyBos5M2Sk/ttcww0RBvXO4i4fC98IK/MKPIL
eS/vtD+fdWPIkumS4HrM8t67Dm/+jBOqjumPGSIwJiQ3KyXpvJ0GCTpbBSSfterf
et0sQg988nj4LwPAo6DyMbECZpM9HZkipepPaQlkE1awD8Zi2R7hX+lMo6Ut2bdf
2ZIBmQutRuAYYIkIPdAcmg5ACLIJ/aPlv/5U3Js6x4dDbXIUKUKPZmiIzDkhahUW
1dQ4t26MW//iQ8DOalo1qfINzGXl92ipGxV53p+1UH8g3WyG0VRCs+3m6khSeCWZ
JxjfVGJVADlU1Vt+zmwzz873PGl4O9VOSxi4oWSqgVW5nxdFA9qWA7F5Gch7HMkp
fifZzCxw/Ov8ksKKJRuZKGb8sfZj6aOom6UguDb4OAjniS2WlMR9kw526QfqTIRZ
KFBB+chPkJ1C5zzmYpBCjRIDruUJpj5b+mpuy2szaRE99izUrNrYKAOMxAD+3GSd
ISNVwBxFCce3mWF6Cb0bpf0EsnSpMtb4paEdZxjbbubUZIvlHurbM3+ZUbYXEb1y
29X3Oi0jq3P5CapY/Sv3x9A43tHrWAytgkOCiy5bLoDpr2Ks2weF81+aeuSDJy8F
Z8AM6gY/zI+asPS55+Pql0n8UlHwJZXVDIli5As7p8x3A5v8/W+Yic2bml+VaAfF
Ip8SPfZ6OEGZ6YsrV57zJgDTTRr5WlZGYeg3SGGgivEf49MQWjpGFa6Uz/Jrp1Li
HFzEeGdHSBjlk9LdnZma7Oa+CNeH9Spm9vnmhDqSE+yJexk6lMOsC6xENqpZPllf
urpE1iH6zaCv/uqDaE2kyr5d/jPDlhGvyhCIfIDWmgMe6Pv6A/xsOKHk+CmJ/dkV
gBTS2OlRtjdOdRwFshTmo/h57ZUpI89Ws6y+fpfvayIpzLHrVl17LRHGqpipGgla
rf5rjNp0ISo5HPJcWqnNOcg0nKvWrcTOhP0Fr7Jebi3LsS1RRHkHmQ3LPdMOtuMG
15sbHLeGAFZ45/yH2kjwGRk+yyu6bNI55qDALFXw3kSJ2RtpJqenSjaTzyEEWPMo
pcJSsHzAA6ZrumSo5YNWaqsQTfNq0FKTI/RkNXbid+1VmjQezWYXt29C4uFZAlSY
RhRvwgXaP8pr+xodfszWEjH5WHFDEhyL4ceJtQ4en6BvGm/Bl9kCXycniV+e3D31
alZc9bXRD6cG6XPI1x15JUa97uyrgr1zQeHU/hmuqDua/jxEge3vcByZeQ2jGbPN
CUefOPzjUsRtqZtLyLHd5vKOHJzkg3+gdLxw6/AXS43SQvpOEzRJqZp1OENj7+JG
dpoi3lmFTK+VpkTT+pR5600e97Guw/Bqm81YJIClItJMxNm/2W6bsreek/t0kgmN
AdXNBejw4ykivTDW+2bikAaQTZz8dHR2YtNoYltzY1WLczyMK1SEIIar8+VJt69A
K20c2n9GLT9YTbqh/XO8LqkHtYJMdb39nAVwDl/o/RAiMUbt57hqbcUAcXYZSuWt
zP8u0yYDr6iNB+xNo9jriq39sKFRD3Jomo6+aKsS+OmnB4FRbYxMQSJOnkvp2+eP
214A8MiH7tb4OhArZ3JO/5h+Gyx+Qa9vuJW8jxGwxW7H1y0poYGTryjO3tVPpj+R
C8POWM9eux2EwikPFhYvsU/mFPtoAqJ13PcMjuWcpRlKVQ0DPZP9mZcj9gJbzKrM
r2EZlP7K8xpjgHaGQ0Ni+1dbS9a6GZuQ01ChbhkmXBxKOJBlzb5fPTucGhv26REm
fyOYlR1rG/9owm6S0KC8oByPt2UxGGo7QlL3S1/CCJ163Q+Iuhq9F04lnhUTt0Bu
lkG3mUiEBjr8LCFLxf1Ms7xdrdbMewNNTbXMIM9BQ41IAaf2a3Co2pfjAjTwKaSk
JxZuGq6hUoguA5lmXklA/4CUmSGlr9+75ePVoDcHzsWKHvpem41qPycfRdZ1+YXY
fnEi8ALQLKEyy6xHunbeTIPnX3NcxsilIER+q7lbh0yVpKuoKUB9yQiNfzETIcK9
x36N8QKmdPNXz/6pUVxDBw3jifYctr2Rfq6jChm2LdYULSBOD79mVQCQoX+HmikQ
sgZHbCjICfw9JXuRMwkU2/8h374FWXNJ7tfVXkGibQeOLM6DygiuGR4tnzSBKANl
TnlMBddfWI7kksWIc0lAxZ7zqxF2Y3B7v/VYDHDD1g1zpbABfbAHDVDzK/X9j0vs
YI2H+w5EqcG2CoaYBmKOheBEJaHmsFPhKiVw8Jxn0dXy6SAyt/1OlgXn7kQaBW8A
heJDVctrDX/LcgQjrCzWADwnudo1XWZ4rYCiUA/MTXpVVDhaHcG9atrbOUz0qBsy
BRsCLA6644DMhAo7YA1tY+8zpOz/+jxXjcBt7Gq59AvnTZoWUQC1YzxJvtK5oQHH
s1UWxew12Po29CveRPPaVAFG+cfW1P93xBbe4k6qbub8gkBSuy7BkCeTrBYpGw1l
tdcEltMo3168R4bTeoFf+a0Yf9ghc9ohG/Ssjt6I27s+On5I3fSXmYCz+bbmdp/I
+eU1K+hC0itfo8ajCF2DN2rt0ONbKbkWv8cmWhHqU0USgswamIOaEYcNp1azsh3k
0u9hqW8CxqRh+25RYKCP57wMieOWaDQCxN/TsSUuTLhxTJ7CWoEOiA/Jw+BaqQCv
VbUfEmA14+YTI7GcwKZUkmx5qkZL/p4/DzgX+b1vEdlLY/Riz9QSfwL5JTKRNQNO
7rkEFmm+Gmae4I8+GkTznzi/w6djstwFF9RId5YX2dYUB3xd8uyTqD5VVRmLfikP
BUOsHbTh2a1Xc65NmL5paIgRMP5ByOxWPD7FCbcn5IBBqeWM02smGS4OvJf4TIba
PhIhESEaiw6DYqmiaLQtAarL+S35agX7rN7BIXlTyq80hbwjsUWRP/9k3eghBijk
ACmOkD8+vle1H9mxGpbbCMQrsYO45YdLhWJRUVSQllDWzOb53VRfONCmnIDgX/5W
K8qW9opYdU3hKxIfKMA2BAHGkMTjbnk9o9bgDdMkhoDUVzGxZjvxCyEBA8Q7INdU
PMo+WkaLLrqn5eQv9h9llWl5qK6YqRFRT/IuwBICnTx3p+ZWa1wwxaiFpMh6LeGP
A5Ky/k+cuoM0xAGtZj1ujFL9xaPrRf45YeH5O28Z7+TseRu/oMk/xrIbY+IW0ra7
GnoWvCbAZ5av+5YL63jEPJopL4ehsVUkOW0qBqekE2mtURsm1XpNhPyUKbaQAkEI
hor9Byo1rUWOTm9CpBpueplhGiT+quOWKXAILeKcFXX76Pud58DdZm08PNzfFVNM
U4QFvyQrG120LWjsAdDKlo1k3+nX6jrYyjbQXvKBZACxTnDXMrfXig1HIhWYTNLE
LB1JSw8NUtv7MBOpKifgXIp/eCDq/i2ONq6YP+cIBwIqXVm5WntVcB1SQHxdhLB1
tffqL4di/jl+KR4Gl4KWzpeuV7QsR0h+XCp0x79zRQPElDEo/M+oLPNFOjKtnJk2
IzTt+Pja403UmEb/ik72PQPx9lQ+440/m8stYMqIpV7AuI3nIfAByMXorKYLlYvH
J44K4Xs9OocCd5jn9+0YDcaseETy18fkdebbSSxZ8QIqsVCvZoIp3lHF51SAyUUK
m8OogBSQHF0jkPdIiDJ8nMvQaP2c2kTFQfU2mH20+AJm36vXLYa4Awl4rQ5NhJg7
Bl5Z7TNfkZit4D8s67Jabgon3v8zX1bA6TMHMRzSUJy19G68nntLkIGrtrsWFNTb
v4JSsYOUBEDNlofF+CU36Ilp+E3JUvf8oTeR+PX/dFsvw0uUqwfT90238GBPfZe+
2GvXftJb6dw5KLkl8lx9zZTWhidInTvOcBMtswstHgb2/z7+8rt+gllvScWuPuAq
eVR/nuKwCqo4ZWIAFn6xIMEcuE+Q7uoZmGnN78GPO3/tjGNT87e41Ik+a2G7Bndy
GLYn/KdX3xgI1RYgcjHrixh9GyHbg4jIyVhu7WWBWeij6rtvhqfd2hXI3vAdDLUo
cAA+W45/gi1oX8gAQRWPI4ocorY7DDlEi0/SshHWfUG3GO9QVJx2VU2qrxPc4iZ0
qKiZHKqeKKhaZJnVyu7xOY0bOw8+Gsx3+4RFlCS8a4R0My37osAqr4hfMXl9H9vL
0MeznMSvRrEN5JUkgCn3Ab1izJsDd2yS7YQidn8L6H08a/q2O40p8wTv0pafFZw5
k7zwgl71kOd1XmdMkLTRHmHRBr3uwgpe9TepX2S9Y6Rzs+rhqTPEr8GyQpj+r3e9
EvyWL8PYgkQVlAclYn2Czk/GR0Nd13iGap45FVhaYQYc4ISVnwG+d7SbVtgMSTpp
el8ke3TuFRTOPQ4xuZofx6AJUUNr5QG5lpRz0zivRIZoBPWdbAtV0ZsmA5YXL2pb
kLgqbyJyAQa/3cCnFr7Lj6dn0LJYpYpZYyuIgM8eVnqz5+UtRqnaTxhved5P0lsK
7bAmM4CjMKvmiE4l3U70aIaAKiMLzf9nW2ZKNGSnhdqBMXzUAUqMEZ5dv1d5x/qW
eitIAeT5MCjViHDi4qO8mHNovMSKZ+jy4c5I/8nFkId31HfYlzaKHRd/CC5SqYLh
jH6ypSEWQFZ9ENN1auBCUWGXSQe21g59xfPTAiUKiL6IIWRAmgakzo9+oDbGT5n3
2YE+zO+FG3K4IEuhtPvQQZI+nSB/Rm1Ryl4uhuWyIuUaB2XpJVAilWcT7EN7jYQC
oyvGKLq8VqMknnvOcyd+o2Dob33Ehm44fyzMjXYLUTLi6I0iV/vTxuMkL4k4N0Dp
Ho9ZWF09O9EeY2MOBS973F2BIYOvLKhdq3XvlmbsNtAx9XVC8rJmqtsKJ1VLDxOd
YK8QTT0A3D+OX7g99iXSsRgGYRXBCTtCdteGdMtkJszvuM1dllQ1UjuqatHLq9Tu
ne8Tk0GEM7ROtPD3n2LoAXEiZYiyRTpWbrsorxrM6fz31CfF5s1Z9lhXaeZGrIzD
lvgGul0ZzJ4WO51meYQdYQhqAoA3QNiQMw9E8nEbXNbBo0gQ/FbTmwrIvhnMuXI2
hZ/B3Ep/OBRDSYfP/kFt+SsIazEbx9UhTBq10c1o15+QCfHowf6EcS5+3O7xi3ww
djaW3TbWMRDuNxxcTbudKckWlMaQGFxFzqTCBd80W5BFC1Ro3SvxD4QqsqcrqzSn
M9tcXJX4R/UjzDRv4Vvr2NtRNXZG3GKwZhoE5YbZXrj7uhFfsd63xC3JOMdAvnxX
KmWAgv9e11pXdA1vEDHpzry0+xcXeFJdpqm/YtbovpAUQH4teGb5F0hSM1WL+I5b
OKUhc6ptqmcRSNr7BynHcQ8V2h6IemXQTfukv1XrTi3ht4u9vb0WpqN7Jo2+dxfz
2i45t3LkFBNMwa43kBVK8UxNJcEjmPlWuWe4CT22m7KIbHlJV1HVVrhS0nlPtyBO
NbMvA6ClDZDOBOa9k1xTpwm0A6/sCS1pkHpudYy5rJ18o/d3ICb6Xu76X0p0pahI
UCoFK9dEG4qQN3N0tJsh4c9bqqqdf0Iaeg133XhPQhtkBl5Az6wBgLzDCBTEyatA
OHEXqxYxeNdFwwFPiHji4mVruqIirvnttmEsmzA/Ms/7vm9vqh9yRA/2h9ncedTh
MWWw+G4SfE9Fmer4WlxNVVRvzO+g01HXKewlZOuaqNVCTEl0SGGaoOzMBzE+oVbK
1qQX6wYz9+VcL5e+2KzmSVxtMALBFQ5TQiF4N5H+YqLFPiR5h57p1Kqrkj3BGVwq
4elogba7yx9uNF3Xo0MSiFsIQenprj1nTWcj4mOc3mgXDh2hyan+Gwz/iq6sqKIM
TgTxkDXhOPbWjXgfFssZpue0sWLKxnNxUl6CvGt77p2aVqgldHwV//dCGoGpp9I9
0GDXB5gek2RLAwxrekL04sXdOGfybqPlIv1zTOfbii4+2riFmVkPSkofDhshxEmn
U/N+XjragYSgEnxRIP0oz6fhaus0YQaMK5I9SBTl1hylRe8y8kXpz64vHgUUXKe9
sTUc/C47eirqLwbFZiS5MaOMYFDdRVpg+BOLpMueDE04qMxHCv07zZc4b1WxihEF
eISGBk7NUsKYjxxQ1Keo/XFYXI1dIe0Y1R02xGb0VFjP3JbE+nC2kT3MOOq/Pwtn
R8gPGNlf/KH5H5E5ioIAWwxHrSjJTwzjMiEwVxzbA2N6Hxof4caTShfsXjrIGRwP
uESACiIbNRGM3OAtpGSLOKOrObfAYy3tYUivurIylUrl3Mu4vKcKpTwbqnyDBE/2
Ud3rm8BcFaPr4r1o9yT9JdmzUtoUOSN7FSDDEbyAm/yksd3ulSBwC5jIe3lxNzaE
BZ962TLG5mlDSZ65hSg0skkf4strdKCxRGts7e3J1avS9LWUA9+Io8BOTEPkIrRY
kpB5yO55QMDwTB/Fr4WsspVe0c3dvSbqhdXZEkmR2KAS1vVg2RrlwNQx2lFPBh1k
d+3zlkf9SJUjVitCNW4Dj5FCpbwA0rrsc9LOVUtNbINdxnKGlBqOTHOWxXz7BYuX
8BnExhjfQ74aJWJW8onlnP7sUkx63GX34s0Rdmb56xpHvRQ0W86tLUva0E2POjgS
Y8sHQiVnxKpMRpbKZu4hpsbWr9cMwUBAjRwT8i01zwow/0w9SjvKYwzYStpttejf
9fcdiFjT5D5I/bNgiWGwbdxqWDtrxCQPR3HEE7kL6usA5T+LF8jXqp60wyhhRx5c
nb/nvZdAcz/xJX5fcHmqQXTAd9qqkJfQmxt5RF70LVyOmxBV2dJuYJaj62asdx7B
25nLGlb9SYgp/qfFP8PGJLGPsVvngXViaInwjZVZ5/JS/FTjyjn3Zsh/cC83tjN7
gSwK7AcMUyiKSQDCR9YTmubeouyEfFT1pfCSUd2Kr822oiZGI1YNeB7nATDEmTOp
p2kawGaV37itDplBLLiZUzyRaljy8NXCBm9gL+V1vgNfclR2FVHW6B7n12ibw8AK
P+jGM8FvYKyjU+0s5IU7Kh/KpTJgl/uVzJPk6fiBwobsMB/SI1oOE2xxlyC0N3Yg
333t75aBnCqkV9HM2mgChrhoC7qvVbrXvMpQybF2pX6b8lT4z/aApjs3PqQGWFrc
B5gjTLuPbnx//XzQtCrs56MOY244UNHHyRfdWZx/giWps24DXG3fIYDFnevixAr3
MQ6R2f8Mkl6+YGMAtv/SCa2jfZiKHhsegdA+yBNz4Q/HvT0z7wGOCp+eVJj10xNA
LkYajDXujzxUtThfy5N5DmdTt8BJGHu3UiXgfKQvxv3bi1SaEL5/OcPrOqvoGk5e
uuGfBKoJoyhm2mRcqMiXc2p+yW4ZjSi+wnJ6QtxxEd4mmrhEM5S8V7EDM/dZ33NL
EoBr3Vi1LSx5lKYZ6FenRa+ZYHz0Tc46kFUl7NV1WT6feE2ukp3Pd5JywPDJgH41
CiWdHL1R6GpyzsGKW6yrjaNJK5Wbr09wRs7mVhWRo+0mJyCbCx4DWWSagVEVLkg5
E4MFUeyH3dbn/KRiTMWhM8kiK/q6OIz3H/bbnWjBBWA3dadVg67MTTH5p3MlrCiK
FWtR+90L9x/d0P1/Ain4JYgbm2Q95LL0TIkkFKX8JCKkZCJoGHhxooHJHJ26JMkK
c2dUfHTUJkhptZ1ny5cuqJh3tBFOTUsWp2P40+kTjTL6u3wM0eG9NAk7scYwoqBh
tyjtJqERbniArej7OlUOc+REmEOduikBz2GQ7snb+4q3nPQr0+GM01z3O62+44Dm
F9urhnaTm5o94MtTpVxVYKndlFoRkAxrz+wsMawqn9CsP4UmhsYQhesr9xU5hXbe
YuCoa7jWjC8orz/hybMRrxEv4pDb0xN0h3ldcW2AItNaAC/Wc3c537Y+LEP2K1YA
CwExnHCI20pyqgNrId7aZ7f9ARcUb8fmzxhSpzgFqZIztt5fNKkEBvlDO6pPd+7P
8ErWDW/k9MDljUz6S1E6zlbplWxLUhQzKlPVU/A3dztzmgK6DZjf8K587mnzEI6/
ZnXaBMaqdAkGjObkHSJyvrISHeKcOOz/qhyWgs3ZQASf862w48jSImcr5N37bZ1Z
LYOe4ES+dOq6PCjz8UwkSOogjvxo1d0IKeefGir2aTKwCYVox8E75SZL1hjoZ+FQ
+WteajKn4O6nI5wGxyqHMyJ1BdnVQfSP6oSFBbRQTH2KTVaEzmTV/FI6YR00aJHo
jNTbTuiFGcTwAFspSUcLkvxkZltmtLruZLQ3HHJI74//ykagqOU/A/oGvsxhMQr0
+DDhy4ArUCjNfjm8RMfnhZ52r0xOa9i2R8nRhw3JOuApDwnerMuDWyd4cg6tMBrx
8N7CFN75uiIRtHCW6ixBg9bWpF/3yyBc6fPU5QwUlWWnRYNdHtpch1kWSgKLRxAM
YVSt5XveSOQvBLDYhxpEQs0ktB2nJOkuRYv3xvXLSKyenRizweKXnrU6j+lkJU9T
uggMDkdAYW6Vu9Czg/FlZnljYnXNv+1HGN1xLaDaOL3mReoL2l9LqqSVcNco4LQ4
SAAol31JksSGgZn1LGWHxHKVnoIsTAlqgAr3PSPgywM0tga8JhMNrdmh2Ya7INIw
HR/pCTacYPzQrpeWR7Ff3HCeHTO3TPPjODyuXNNcjW9Z5AbcWNM7oSr9NyLYgf23
BEYosTso+85bJGtteJKcsli1e0fHlBLybzsdtpn0UAWGChJMblDaDZdSr9NRr6TU
OoqjNplQLh148xFbBCAegmq1bl7dlRDpIfzgxnsCBk/JTJPQePS2CXF+ZL8Bm1ZQ
qeEpWHch4xU/f5mJZb1DWGwoL/gnL+fb5pRiDxJtHK29aOcc3yiVclOn2rktm2zD
vbYTBMnZ0/N2eo9eLKNq80NeJZs88EIBerMEt1vpwInBBu5Y1fvdELOSEJsYMQdV
JxjTe59kiAm4w1FigPGVQ6AhiOTklyEsU8gdiyKklJfgqbPWYya32eiK/Cx7OqYl
CN5slpApoaXytPDYoKkNykdBwqXenNRlVp8Ir6Z8hpMUNkMQqAFOwudylW20cL4/
F0yzpMjHlsoHYb2eOoM/mGYI1io+KZG2XkBxCNup9o13HMjZHe3rgjb4qkn6BOgA
bctSuN1yxwJk0lcxe7Bo1LHDelbU6y8xeZSGSQozKCvqt+zFN37NWOIUeVMBfzYk
JTcmD1BnAeoem7VhDIuOnXE/3TdZjdNvE+fJnyJh+du1Etj3p4hapyPA+MJVYDX8
MdKR9pcvR0WjSCdOibZd8gC1ChyXxrdhRpze3q1g8sd88v8F05ULxIXm9uuaKgPO
9fCZJkvBtxJ47T3EduX9FlYmdxdQt1op3pUqhmNTw8xj4xbCSIuKH/W7pOvrpEAJ
48lHf8RI0ZSTHMJ7h3BwlfgFGlcYSL3UjNmXYFiSIjOS9WAGN240wRYjMfbD51E1
8NOQfxhBwi0MMgNIyhID4ecm0zPgIGj9fNU3YA4UWHZICpF7a0omiphYHPklegDB
Lab2QSfcx8iA8H3FkhKOzLgaiiKmOc6htKxWEZcxXD0lN9Haj+PtH+LQ0g6kPHvf
PiA/IEGOFuEyPuYnRjA6kJG8OD1gA4Ct7jWi4cPISNGOdJ1h8tgPmtP1Q9gwhVO0
+NcmdAq/lK0vOCdlkQgg4VsSSCux5mMRmOU1ojZpdNf4TJLgNhCVSziVVTWj3N7I
LCU02r4i6rHZVIYhH83k/MesWyzcf3WqawgtOBLzOFwBY22Sd+V+nGsa4Nc5CP1n
x1CKCqf+TebCjAJjWEy6wJO6/LrvguTezwl9UjaC77sg1SCNBdwJxGPIZlgOoxLq
GPCZkYpV1yEhuOdr1psDCp7QQTq7+REn4eUP9FosmBIqH+1ZxoQK96lD+D5lqtin
WchRa18OyW6rTrx74y5V8aUg7LcdKsgg5aFIHdQhAIYdmn2zWW81kTyeOAnmCwKe
O5BAU1YImQAfybIBmFGgmbsO1tjyiT+W15CV13rP/3c94iQyxYUZQxjwotNXTABC
QwTuekQb7eDa05eVkQXIAwe2S/0VwxcfYLiSN4X48LLxR3VNmiNk6oAW7V4tG+f7
ItAu3DBwhCCiC1oNDqAIc1JpcfZ15RfY/q+FhEn/RKK2tpefQrQtGfo35p4INOPC
eOUiPCC9kvxtC7YW6qY+YIWPlAeXNeHtuWMUbY2nu5/LJWoyc1vDhT9zAethf0Vx
3idowWRE4jCcg9qOxL7IEK7PZQTbTQ7Jwnf/5h3gegjrD1DXcKLoxhTJ5TGhrJvn
4qBCCeaeEjVyLZoBli1xG4K1cE4LKXZOQ8LoV6a9lZlJl/G+I8FkPQhV7hQ1+BaD
h1vPF7Ini9W1KC6icWes8/h5HY0vjaJ5lrCmBReT57ULxaETqnzlhCF/wD79US1U
ZzqARbLOiKzabKYqlqslge2Qb4JId+5wH46i//cEbA++F9ln1VaaStKB5dpyaPPM
JDZX9rb8LEoImPrCKvhllxXFl6IMZnUKTILaGe9B7Od+vpV60xltsgjstZDsPZir
T4nXjvkUjAbDKvWA9r70jKYga0SpH95KDCdlu2Bxlf5A/7nozgmuOiJjx7bflmiQ
YnScfJrnjA34yio03kjnvgIIsfZSyBFcRzz0GF/nPraKjMzqpiMD7J6VV8enwiJW
cWnZYLiqFhihOH+x54wp0RpPorqpk9hfzhHKZKZF6V/32Cj5GLKG5AVj0ZFbeN9s
ImWBvr+alcub2GltkPg31kqGgEo/ng2bDJ1CcUIEwYdvVAfrl0NBLFaIPhkndked
UrEjDqqvF4bsFa2EPwpEcpR8xje1cGaqkd9UoRGmjcylZKpfLprL4h3xWTwfiN36
Phl5RPQo3gV55oVNSw/YpIpHHWpAzjjng3t7txsTSxSq/gk0p9RC6V6Qu4pgjTWl
Yp/zqXAaCZ8Vmm0jdhMsfJoDQic5HK5S7l3qHe3IQWsEFaWPEOzqIPrMBsC0zUQ0
DWwlIhWmQDeq3vlRo0RGV0Sth/hQFusaRYlZWZU7dp69aszwFxThzyKknCOQ2Jse
AtwKt8M22a9gbJQSp58S9CEklG2oF+chIPqApCzBxV8Qs4TNGiQFzeXp+pqBzSy7
JQuU6GKYI7xAa+LxcdwaK7bXi4C7z+umBse/AMX/t2EV2UnvF5ZjvAoFhJfDYL2W
VcPUzFOY7U/XfHII48DvqoIVMU3WUT3pumE9zko3tW/Y+SSZdsVA5qOrwEYU9CRG
3De4pOcwACCOWOeEM8TKOnohTNNIMwUF39js+7G3MxNm7KbXxUIsW/Xdw01voaVE
OOO6xDEcl0Erx9mngGdnsna/vu+tJL0WIJ5cNCdmjL5NNSq9ep3T+KMiGHnSHFf+
OH1m/OuiPXWzB8j53xq33LyZ8Y+W+x3lSrQMi0aYljS4AGrMZhH/Rzs83jKwTIrv
JTdL7JQdjOqDlTrDPhpuBs7ACaZgaoGvm1oEk+l7gRp16CA5Mkv7anhY7JvNq6cf
RsxL+svSSxOfDIxQP9aRxE57WCZ+JuTKLnPbuZpDUD3DXHtJ5tKlFcoSlLNIpNya
qoglN9zuqmfg50UwcACTyO7Sq3iuAnJWfBqFH2fVTVfAGUhz9iEu4KX3iDBvuYEF
CcAe+I56rpn7APT3leH4uXr7DaY+HIRgCUUhtOvKf9clJDeQaS7KC9KSMBv0jnRt
+eJpy7mQwOgHVIlV5BftxcjfPbI6EY5avsWqrgbZh7F4YRsioCIHtWQ8aAjFpmzB
dg418EN7O5xjcfF5/3xbk2Cn3MmCTlIDbsd4YCGL+w6TzUx7/jhQ+AP5Xfqs20ax
jGnyqBBbv1iwEbjl7xtphvt0gU9iUp8QpfuFfpPfxAhom3gkRJQ/JgQ62Vvl8Fsh
YeiCf+tSW2WjW7O3wh+9r5SdPwjg+gDRO5pVTCGbjiV6Cm21QEC+xXqBxNsFiXDT
ozdRSKOxBS4WqX8gtHDR6NkHOzcZ6PdUs+wGqenskeGVJ9jLV5q1bEGWGygQ7hs6
e/YaOJdxNmxotsCguIX6AxyxbeO8XsVuGLX2/Bb7Evr7KgzGiHgvSpT0VbnbCumu
9Mpce6347Dcqpizx6xsSxEz0MB0nsTLEgbBAwb/l0C9319ZEsRmgPh8x1aTkMS18
MhlDBGyMmRVxXnzGC8lfXpX8ZUlPBeNEGmvwaKaLZgUIbmPsAMFozvNozjGbheLc
P3UU/AKSJEfLGoNIhEtQK1XaRVcyGKeSlfjvqxECarUQ0PkrZQnILgAxFk2khxRC
DfAaHA28rE22MK7eBxzUiRafl+TkLL6hgOmIDzhBx3l5RiB5mqA7XB5eUvI/ezVE
+XW5Pd83RmvTHWnr9siu8dZBWKsRcEO25wRa7RBM256BxccZTcxUyLgbBTUNhu26
GiTiBfo2kWefxVm/THMKtiZelRFkKbxDL+qnGwU8ZkWyp2zskLbablXQ+Oymguiu
/dUVOV86ZSC2iZQlqtUNOteQCv4gE6BpIIoigvAVRqASxR9vebN151SVSo2kiQHK
PMHaMb8701U7GHAii9DWA6Mi8nfMyb0Fr4rG0fVj/PvyuNzGv8THvfrH1qO54Jce
VDrbx5d9rSLZQ+oEFW0OayTbLxbDEc6Ug+1QAEtCrbzQhEC0ODg8rBuib8lW4YRo
Em/c4OTLQehpSzXeBawvmANto8t3bgnM7N+q9AI9SobstQ1NJzgWAbaynS1PD4vH
vg8nVWUo+OXUWStFc9cWwtaZalmF1wFBl7wIQDO4+GxxIuL5Ru0XpD9trFPpwkor
lWnwo37yvAmq3/4mYnEwwAfBZkqbvvEtEzCo8FAZ0scB89cH9dr5AnXfpNxoKo3a
qOZnRpC8MNrT5XaBxvbYF78R2GyMk+aY2O84zWDUu0mwCs4KozCfD9x69yk1iwbP
bfcMmCoIjiJcO3F8XuV75CTSsQm7gVTfWTNbQd6fp+60bdB8WfZp65SOGRuUQ7AH
pqRfsTx3jDiRTQNcIzxtPjbgMt1hk7It8e1XLsXK8Da/1HAsy4JleMuqtOT5Ev5Y
kx2Axncf7FyI5SMoBAkP9tBEo/RmOJZIK+NhlhL9EUR2I4niurEpgac2Jhmsz7wj
n8d3ZF/pYCNSmW/nmaHp05HgXAR31SK3m6LPxipPqIrcqY8Ai8n3dpWjluZlKwS0
5T19jOGNHIK05j0Q7/AEJ/2z88PVxhBOn4rarIY8VGSCZsNlCQKmCyXpbhvnqb7U
AY0J3kcMkz34AEzIQZ2QvR4SBErMXklRskmrhcJ1P0GTR7frrCIrHHOSxKfH2SfP
jKs3DptG53ySBZwrKDI/abce97Lq9ZaFqSe2MPMcttfoNJXYQGwHOPFVovKj0iCI
xioTytZjQMkRa8ZuJlat54Y/3msRrvK6/jeblExMZFo6QbeKsnh1wCit2g/NMMFB
yK4tPVH0+rPUQtJdsruVVhxTiS9bbXQlLvHRe+DbgJ7LM+w35bsKkQSyKVi/sIgM
1JZtcDffonK6Mqa0o2yV1zc/A3RZGzqPQSLMtj1g7KLCxmsC78i8hocj3X1uDU8o
L8AQld0LRn+1xb5HGXsTCNtIGzb/Vz9CfFi7sCXpwMuQX2su6YMmJBLn734rDgzB
5k1kp+90J+Rs6yB3sO6+SGTD+llcUqTgCfL0dGM4ARHZuaF3ewXTXckkgHFJlsD8
Elq633DISSqQoCmv862V74qu0emcO/VIvWouHK9JmnI3uzETvyK2ipZlK9IRt4vj
sRQDq7K8SaTWaHRCYtKWcA/p9gp/RAsMV037ZzJo+i6oy2iNcjCRebqc+XuOr1Ze
aXT5bXtFUKF6ADETvtT+K4owdNLnQci/UaLpClL8yCeHbt21YqX/+eeMk0Jyw0d2
otm8ILdGcGkbnOb4KLjzs9qTlFEnyRPqC+GMz86GEoIjesFoSs2KtCO5fspopHTa
j4PveasEtIOJ/ebiEa15d8RMtaTmZRrLR8H7qFCnYbAZqNjiNtEFpwxKm6x3Qwby
fPvB7ygoMRfoIlUdgNsGMlLtmfM5xpjgPjPQ6Cq/nQk5/j6Bvx9gPAr9Zljc656f
hWtqDPhCKQgz51WXjmNTXIAXPFh98B21+of7/ggeevYCpQEVCdQpCW0ic8kJYnFQ
C/j9TrJkATvf6dDi9RzsLyGINQW5ch4zvbhY3ypKB2Q6byLlwJV0x1IpSXaPrz9C
J3IxxoAJl+OqXzMzOWtHcGSmFDA5Kk1ygxfD4XT0OoyooW04dz8yrKMeenNq/2g7
F9D3JNZcktgxvbKbpLlU0xGtvTQhMR796ZmgAnG/ojLBlQy/Dkt/7LW1rsGcDSHg
eH3IO+uDhi00NSvbQ0AvZPxLbKyo1eGEjc4A0Hb6Elhp9GPG1GbiFjOPYijmD8N6
VBKhEIeXl8M/lS7FRvaVMjWPH2ijqys6hMN0qbzP1XLtuNJ+808Qtp9gjjq7FGV5
bhUHDL9kTME5K4ixzLhq8mWSz9mr8oNxqwaoaKhDYhUVVBsILJYomvwn05c7Ji8g
B6jCrq3vF1ECBRGI+L08TjmkOQG+Bdg+PpkbkvOrKkZd4/k2DfbcpY3bLJWqxLtJ
YfSftRDSp/NqqiDfwu+G+CrjS9R+6emDqDNkZhrUBHhM07+C9O7QwfYUNLgjftb2
EyjdxSn2nvYuugyoHTc8VY/Vnm8MHGKNiTy6t/3vNeh65062xu8vaWCHCj/OgBIF
Mmh4lIQ1vB/Y+mqw3ny5RUR0u5COqBElJmCoA9J+rxcTO36noBQEDVRASCVm3E9q
LioWwS6UBjwDk8N6Q9oLkC5gXylciElc+0nub5N41tUW8MEp4R3N+saVuUKr4ye3
DEhHOOGKAqXTet7Z/rISpBL1V5y6e/Yx5I78+5/iscNzpreefvKO/+498PCHeHy4
3tNvyWgjbHEabZ69cM2MpXM2yEw5LKGxgzOLFUWbjFdoTT7IAAsD75UpX3CNPaJf
7utJHOR+YYIvGbUYemEPF+A1XN202oFYYgDWdEYPYfLRhfoWrFl3OaFRBsGwB1UC
iomsEAel38t7LUBl2gTNVAFm6ON51XDoxLxI07NA3zglG9IkozDpFyLE84k8+aFO
gBSPG5u+9dFzcKLhoM28HuajVbHRejy9uiXFbi0rk+msCiVoh4MHn06MIUEaG67E
5NKsztBq/tlnSDwqVYeC88wbX0hnrmdCPchr57wIBsNAWohQ7INRmoyPkvcSgpAZ
rnFqtc5oygl2llTRa8TgCVifrXwPm5TruKF7FQv/Ljk5xulmRbW/Vb4oeh3sCL/V
zaY1KqI8ksqwET/Wx3wSN+O+YWclM2sBlrhtfA1gXBiqEJKSyroLUC6/ZCri94PK
0l7CjWuAcvNriMayEguFjND6FbxEKqyrgYLz/P8RuIwuupLBJNXYdqjBGc1m5atN
jbZyGLaYs1qqxRzK7R1mTRXbtWc0nxujxwuwXdaHAOWkEEpnPBeF8mqZvbhf3KXv
UcszFwZeNpEap+blCl2lmP25KDdiI9T7sKwiqT5Q9njYLS66FgWE4FU7o+wCkCDs
Va9UXe+apmltaUtMAIROLeFTNodku21barpOGKK6TtZjpeb3qTxgf3hfxnQQrIBb
7m/R/+5tTqi2O18ul/27JcrzRqN1/gLtiGKcmjg4cLhCwi1YoyNUuejzR48gdQoa
OWXaPvsLVVM49zXUf1pdXXRWYOtzsPkkTjigqTjwigYzPQwtgcYAz+2xmCk23wkG
NnkDu07ElTS9xC6Hy6iV2C70G6paQGAiLotY4dAnvCgIaI53oKMSOvtNjtW582PF
Z30yXKh6K1Iuk40SpmO1Sa6FrEX/OYyNQoxJc3Ci8qwNsBXX09hIauI2PDpojMJ4
vEdtpgUrn29ujXvz3P+LXF4oQXDO3+W4rQbop1xq5ZYaAUi08TGbvMWxQbcJxvRV
iTu89PeNomBMsKx0bHhQLnJyrWSZZfbhxR1hiMMMqqpxeH32XQa569eyc9mVQso4
9X/h8Ur2Mg3J1Opn5jxNwSIbBUXBGeDEytJQaCtO2730beqiwY6bs3ekDnf3cpkx
TDyQy9SMUm6UP6vmZ91Av3g6mUibdcB0PTPLqHVn24W1YkPZvsChg7z11aXamcKL
UjjRlueLRRUwxoNDsqes7FAastOv/ln+rm0AfSlIWdWwRbsGFgtgq9CFgVr7dLLE
+f3YbBzFdRnCVwkYqn6wFN/PWxbtP7lj2CDG54TKhTxkkhqQddSZ/lvmTWRFgHwF
eCwG/NyEIkAz1876Zrdzh95FcqO3BglLy2gGxUdTtORQvoEKThmyV63My5IZ+Sr5
NwZWeKh8Z1EABygjYbOHXYqc29SzDYa1FWthWzTmpoBfxOpBdK+++hNzNshxuAkh
ClPB88a3tLgPjeXX1a9Pl9egxXz3wYL771lJGEpB9hVtSD4rkc3czz9kuoYsW1u+
pMRWBMPodG+ARY4/6uxIzKjggWnw/UF7asUt/f441r7uFH7mGMvuiICz9eGr9EHk
bpZ3qdAAiGhzcU3JiE2pCpwTIG2s79j7KOLDeoMOA3454cJzWSGlXGVm4xsb0aS0
UlpCtwXSCfNCmTCu5hX1+tHy66l0g+INhTLiUhlH11exFDE8Zuvvb0tGZJ9VVMfL
btg77/DsowkTrl2cJLqhCfW38fiWY83a2JZ1sXjvZsLdZXQzQ4ICEbcaKIyCBzzB
WS/w5oakFnQ0rBEWrC2yr2BXCfFgzuoNMAiaX6OgkRlhURzjuU0NzVT43K9VHQM8
EQD/Do/u6DIP6+1EFqFTCt/KJXHFsFbZMJcOV5Jwq7kc/vh/Bj5SVDJA1/xeItD2
T4oskng0/4ldXCpjq+koKwO4Kp54zcVMw3PIE2HHx2vH/1qEXvtdMLnVwZH+1mN0
PDmYW7bhY+0nsrvWwfl/xblvihNSgMyX+pwRZApvyoP4ksYr0c5/qKaPIEMPTN0D
MlOgoc6ggR4ciahUvofFBeUc+yoIFLhpAA9JOVNBBqYo6XvlxCe5cTnb/Rejtnrt
70w5VOWotxNRH5oNj1GgjCqFviE7lA1yw7QjtMhw+86uS7o2fubJh7RsFbbQuXJb
XcvkvRYK7zhOzV1PIxu1f8iiHNjQ5kWQlHxQ+5tpSwEI+MgJB90qSGlkwH8k9OYG
364f4QXe4wOCy78iu5/H2iihzWsV8KGGvTA+v1Eqfc/e4r2Sr8UzqTBca9Fj80Dc
PKbdUVty2KP52GQE7yWk+88TRkgv+Zg6ubZo4+dEYl7sck8B/WgOr1kyAnGtvOUH
2K/FBBGax/pUj9Cj+U0ylOkkzsYszRiYTeDZRM6zFziRatmmcaNLinKs7NYik3sM
mGrM8WCEjTbicUKxa+QxlvyIoLL1ZhH4ErvuekrHgU4AFTeWbQiLwOczbiZlFlbF
+foqokALWtDNP9XXNi21WJNadYZxPBC1D7abrPO7Q2cZ8HGasPaYDHVSGbH7X4ub
U0pmNmmgr+itJtdyyKX4WLWuI/tKQ/ThEgSUyx+SK1Vnu+NQCLMr/+5UOQuhPy/E
m5TQfqcuDmbQsldWecmRckKtXHlGC0USjUGX2nKxxx1E4KNudQyOayPulnilhEn7
gSMXFn55PQsXovSKESZTu2za4CR3gb3fDchZrCNytvLmMB8h3RhWZDlCGTZu0oiI
Px6rfM/DCEO6M9jCJc9r7seBQpB3Kai0LTAl+801RmJSrfRtwK9qAcRFLD6bhhcx
6aWOdEjbQl1hcACOtTaLdtBkUmgTxGkY9VMbpZm9852N3/xcsvMIoH3C7DnDoQ7z
iW6cbDyZ0K5N2IK2H09CAkzHtw93zAWrdRSIRfff2VcMwJuGYtM6idearoU57dCC
PKxzYnZMUkhJ8hCbXcPE2XVFwhtDop/da3BRAgL08XM620OOO547/pizkQGbYXsg
hXHVatCCbFhiOSYA5JF/kJZfDP9zl/5U1UnGHq/l5sqmZYaGz1ftwUOneyjA+35H
EYBKlXF2+5MmGGqgRcdgACNB3c9t9d2KrX6fa6HTY/YyeLHd065vO0P/dlZn5XHH
uyCHJSTVkmAyofAN9S8mguHKWkblHefinU8gfFYmH0qNaRszYO1VOOVLcBqGstVT
QRG/MlcnrDgqGhIalMsydxUfRwKns6Q0CX31s7PGyjZC8iRx15550ixs2+VoRRBd
vpyteWj+wtKYUjzk/wYZhOjiObL2HsGPtBLTmgeh/l+gDmJO5uxiZQm8RfFUmmDM
O7WCkQsGrgeGIYVGBxXqVkbH6j89lx+rVVfEVx2kAhH7ePOCIRci1e59gfDhkGbw
gQdx2CUvlXd0mIUCThrewIPv/NAD6NazT/pH/t/EzBJ/oA36XfhZ888EQmy4LDGT
9iU9W+MnnuYksNKmhKgAmq3otvNc1YBHBKqH9kFB2eOyaWSsYLlHciD/uEfM8enZ
KYa790mWV+yqj83PK4LbszmWHqnyqa2JG+zV0V7bxy8MzpbqCKCYf5EeqdfxgEpm
GMOcHsCey+PEmG+LdNx2YGO/fz/l6whw5CoFwwWR0KL7GiTBf2cYGjOSmuJ37qjn
RHSa9ko46QxzOO30t7QptgBMKWs6rACh7zRjYC8SYZKuU9QDL8r+9Mzt2/jGqck/
V/zYEhok8YJxXwkBVyzjt8YZk3C7gd0gRcL068cZGXmdUIoPxl+uhFt+ZyJcm8EV
rxs0slCrYkX7nzF8ZnoAocNn1sAD9wmUrOEi7vqJnkp8wVjoaWWevzXq04x17EJW
9jtBi4of7TbDR5Bf9Nz0WQI8Vq1ibrZQhbJoyZjaAVICkEED9eQ2kRFZPLEbQyE6
lhM6xXYFOZcLP1JQLwspuWBmudCXAsADoaWvD8xMpUx8VvFHYmFDNJFoycCaaUhn
l7U6WR4wv9u6/EW3sPYfsm+Q0PYknEYCJO69LvOBievs6HbubUiTfBM+5uE5xIMm
qlNDG+KKpy4OWCYep53Oz2Q0yIFgY+DFeX7OfHSWkiBIENixTRIYjQOAkJGDMdgm
4P24fw6wSLFRFyaUfH/xedKC5HlzViQ20n2TAvLpPECV7RsfW6fsWHL7Lcn3IK6Y
LznEKvq0cO2RIGkzxoEYW46bvQGvl/eg1+KusEooQt/FAB6XkY6JRAifm29fJjv2
dep6R4lBr5BQru/sfsFUrKICWQNNxOMWVOp05cM6nXUPm6qEu3UatJ1e0OG7PE61
NUeXdY76h+V1ZtHrdpuQpEbdcWUSOIYrM6S5q+Y3ZPTVJ8aZpOL+EEj8kNHggSot
MGTDeRkT73vr2dff7jLBddG1aVTciXsiCO6T041vCmsuKR//X1igYg0zvWFRMQKn
3u8CD0O23oY92BEXt5y4vJCysgHNbRNZKq5fBqdhA6rVVbXR8uSBdPI7ZnmY74aU
tGb6AwtT6n4tjfg9/ExBYc0nmVCLt/56QtHa2ObqNjO/AhtbrMxP3v9PjaxbjlAq
kQcD+D5z2wM1nTAM3ZsvL2IUBlQulQo+njmQK6ty1znm6K4ycX5VmiZ5Oo//lJKg
zNJjl3doetAhBkWCSN9kylS7fyxSrSsUk9+uOeOksgjKcIL412nJiCe3qsdRdgLc
geiex9Lc9pBKZhYVGKt95mD0uFi5s6+2KM7YAPGMmmzsvLWk6yz6V7isG1L9uMKo
FJfpKfjc8OpkzlRO+0Q6jK5mM9x0EiJfDb9xIrKV0kbwLAeVYdNUp9aj/XQgA/3d
+sTPqoHRu+65qmhaHKlJdxXFXUtX3A2vDDSg2eBL9h08/N/tnm7tlm9LQkP9k1oI
dMUng+iEhBU6Wxb2vVPrBthJYI7MJjstYulMvHRRO4Z864ptOZ3IkN272xAw5XPW
NlaFfmy3pVfB3QYiyDCEIHsfFKonGyIW8o/v/CFnEZaRTksb8GQaNSZ8xJDN+JyZ
3I03ThVPMv/kzGIp/0Be45+qGygFEdRTJyBSncw3QcLbhKRy1wBzcG/SfBBMP+tK
DGttmTKIaEUj3FJpcLE3nF6GTUOjILw0NzS1vdXzRl/ZzhuI8nj56gkQcTsJ1+sC
l9ZK3tJrWQQMVK/NEAUdPRzXrxUhVrOLRhm30zJqMbS/IYfVRW2ttDvvPPq4WpFz
ehOC/xHYAbDe7bbWxtZbfOIchA1dO5nGIwc+XC3fq1dGMEjcqEe8rBCcljepIPwg
ZCYHZipXrFZfSFG63rdBLPzk+bWBo22CNMNmCEPFcqd7scB0eS9/GGSNUvA62t+j
IHW5zCisr9e1X7z00jT6W/zsLPte3Tx9lm1Nmct/foI9a6+yJOWPR8NhmBPYkhcc
LrgKmnyxbtfk4lQUGaHpmr5hoJBf030DoWlkj85efApvFbmkBFXhuOG7YvJpQ8h+
CJ6/kTxIoDcbsWdYmUmM9p92Hc3Ue9VnX7bwQyMwvjG4lY61ttPqex5dfGUeoOs+
ERAlfUjff69J6uiXZZRnfKcKBYW/BhhQxsvn7RfP0gBeEVI8W0doIpqHV7ue9Pt9
cuasvtpm9MEZLEyewkapyVKSIQjULHGPwsw8PF/PIPE0uDltUgya1bRmiI0hiMEK
keE99GUzMbARG6U+Ucsj59R1vdKN59BNsg/9ejjuws9tE0NfR4ffXSpTMSaGwtk2
w3dR4PJ2zCO/w4j5qkhgJQhJHItUFwWMi6v+oUy+C22kOJY7U7uoHirT7AOi8zVD
rQpiDq14LTWWqXEGa0bRpZVVD3rykX1OHp4qmrtMJBuW/IcdH7YwtU0tzsrGPCbj
M4OE8KS5W6q9KjrhJJclpTq+18vP8EvlyExtaOH9+m28w7DyIRqg3hPat/sqY1n7
u/5Be+p8UV9tGGQRh35LWkMY2TtUGwmay4JWjj618kdZJ/KHbjV75ioLT8S2dSae
P34gGutw7yqp5+5EcN5/A7h/guY6y/Pb68x4JkJI9bkp/i0ZXNmSJdfmeshAxqSK
hzWuvJ6qfD7K46q7T1vyIOqhjVadFCqW3lKBRBblQbRLzRpUnQV02VrlLmieokYr
MHprXhqKliMf1ZBKd8AB9WUJoUTe/OoNfQJw8pqP/UGxwBxFlEYV0hMAWFPUM2fk
+yxFKhA7p80hfnpc8iHYHPrcInKuYrlLAbkqy1UWtcMt+qjdACRakuMCLoldPrLS
gybI+t+UTPLhUmNvJzkxrTSuEXu/VFRujHKuh68XBb2b/L0iSf8EzyjUm9z33ffR
eUIlhthOyzfyl8xptEBrR70CqKLDaF9EvI4trFAE55oYwZZ88aBAL4md2spPE/3r
DxEz2tNMl7Qj54a704f13phtnvu76PhctMiNivbLdDlGyBTkpwOAAzUGpfAIGr6p
GwLPPmtomwFF9trQxtkOErwJdohRLS7XhE3HXAkVkPSJBqHde1NLJccPj6hN9P4c
9xs1QrVMizLt/dIIu6q4FGXkij4T7tpZE00f9VhbK0o9n7CjTUtwqcVC8a3LuoYc
lwW1uSVmUFQpf9pg9b0LR7o1ar2khluRUBfexbGYVQD5aUvmjpF/iyirQPCC2OxB
Y9ISwlEEypL1p8znycuqNg133lOgOnEbmHZzLK8RgR7EO44iusJCO8hqthSN+8rC
TSD0ZbRXoy/6B4zLiW5Qll1YQXnmp1wfh3iVdJOSem1BZhPGE2kt2TPZdS8Tz8xL
2i98RG/cfFPKLpT0v0mqGR4edtKIeIRMHWLiu3gvMSU057+lIs3pQ5TzLt/mzN7Y
tnxuIk+bz9Bsd5HiTnPdYGN4L4qtV9awSQKAe2GZ6CXS6BtPB1D0WcWtSeqLUcLm
Fg6CJbFB6HFdbGfUcnP4iOsqPasFNWFtkP9g8Xv+c/TgSBtLxXhPFoulunfeGUms
pwysaRBofSHt83R1asxVJ45vcrwMZ4vJne13Hhh40fRwotqIC6tiY3fagvPbzinr
vY6XPMLoyPrRX+l1zoL+NkSm0GqyUrER8LEDJLF/IjEzeTo/W1afacFVxqflJoQo
sEwy0+GdRgsKpiKrhaJI2MO/bhI65k19QtOeHlv/fjU8E3SI5UvfifXw2U3bb61H
HVPf5Kb3n8WoVwBOzJMpH7ipZMinKejtu8H+7Ff8FLgfmgwI2/LWRkC6xwV2chF9
fcVWFVGpOmh2/kBX5Yl8BGIr9zeWfb2ns3d9CL3pB8dywxVowMTUj5chwb5VkKxj
Vz8lfvHZFN6VM/9EWZ2k2zl1iGV9uqT/7X9w61ZSZwYUzU6z+WXyXYjkKG0RFf5Q
pq57CCPL4KUXZhXAEndj/61of4hV+sABG0gDNF//RCPzIN/CVl5P1qHkVh9iP63H
U8UI73tRjg5ROeQagl7ITIfhP/ryc1QXYwFsLqn6dex3ouGFEIwxyGnz6aTcZh1P
z4m55c9JenzgeDve+nk++fRGQhNg6CNCEVIDA0S+nxz9d8NqNKj1daAzRXIvcMpp
BQsdbAUj/NGb8wBp1VbGn6Tnn4MfNdnoLwAQWau+IQP/cZ6/1QRaW8c47MnEMA8o
wNosAsheGrEvWbXnd/5MP2lQ/T0ULqfHv2kocrPMALa27uGlvdpKPmTXwxjOsxxC
P1exIsrNyLm33adj5y0Lhv68mlmPV5sE/WwoE086izm0A6twLuPN8yGFMgeqrpjf
eD9smAykQlsxcXSqAIQgxQ==
//pragma protect end_data_block
//pragma protect digest_block
ujwz2z6NlLsNwU4q97/463BGBYQ=
//pragma protect end_digest_block
//pragma protect end_protected

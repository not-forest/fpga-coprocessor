// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
04+2+RZFj5T18xwOmP02CXEbHwNzATIVb7pizr6nF1J4FSrtlNvSVxYQ+pzIW1/N
dLb3dTr9wa+3+Xdtg0c6W6e9od0ZnPmm/O6K9gLWJovlyuSUYHphiH25Si8lWnKB
p++uliaUbfpwYN+LPau1WeeKGxHl0cHsfYviJk8MLnA=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 14368 )
`pragma protect data_block
YVCawzwBct24tE8rMN/EB8m+aFSCgdtAaWTLXqhKh+8arjpErBjYzGOq8oy04OlI
tLRX++zxxL8JBG/v8Tio7uftTAsSYePGDSlFMNU0oaeOe8QlseWYZbFj/qOM71tu
h0yHsTjWi3XTyPachKJRNLFF0DoxtMTWe40Y8/IxhaDjdxJiYana7aEU8yEMkTln
HMz9uGWGoDJuh3UyduloX/RdI3QBgS6D0IF86L7TehGZij0l1aLKhh58a0O1LnXn
tEMR1JO9/pMOQNRDxuhM0u7g9hEDpJxjU4/BvR4lLFR0Xmm4eu0CJJtOywRrfE5Q
e/lKnqBn+qbtROVpFP7IZ9WakJb0CzaclUvJuwNRPedvJDR8prRGyxTQCyic2GO8
M9rk+NjJIJTzsH1kOMT0qvcnt77sgxBDVnBYfGiyCigSkToNmIbVZSJ83rEo8CyP
SRhIu30QWoPqItW109bNpkTuR0cr8G/C8n4UHXAG0XoZ6Na3R5KioVmWJf7atrhx
dhx0vZ7lwhYrENIhcutmX/kDxl0tcICFTvyCVzAm3mVYZ/cbyfnQA5mO0JIRBI2c
TABJbGUNLd2KgV8rRih4GbGankPqMrnj5jxfyJBty6owQQxkKz44Pl4XZ7A1vHRE
6F4HzwKDIZ0l74jpMiIXJA3KFUAMVEFvHuhH5arVrrNI9NQF/FXyvo0Ykf2bZYk5
OWLoNrBDgm/o12KZ8vfqinUOedOpFW+vAUFXA6PQ5rTimKtHxS7jIEThgxP46Ate
GybnqWWCpSZFITYXIBWDeBecreNHkPuVlcTOztFgJgzJDDfORC4PXG/eY+LsX6sy
D1LflQqCWNBD/ofBgEhUk7i0wwgXTfKWLZQkfCDyrcpnWfazrHzoA+nfelsud/8n
Bhc4ZAlIqHU90paIr4Wp6uZbOds2Hua26D0wsLCp4u/yj4SWorswwX18taTu94Ci
Uuz98GlD4a0LTL5jr+7GotbRLRBRFgHviAn/BRoz1mCQj54i11Rd+adXm/JcmW1j
ok85l1QTygIXOirU/7jwqJ7XBUB1udjBVTOqGIbRBqQ5SjuH/KRl/J/4yUlh3wdc
A2YB0Cw0XMBjcMIGGCYpwckwuUyJ4MPzXsRLuaNnf1D06eJguYh2d1f0t/H7W6LP
+rZiqcT/XK5+0glj9Bnt40ceKgRIibP0qYlUN64jldxsRQhADdn11hDhgBBgI/YS
8jKnco9t14bbMfBM4JJv+g2VA/axMLEv5wIBY8zRPOX8jn8GOQZU3VhmracUkfMn
h84VInoYFVN2b+5rFK0UhQPqxB2uQ+Zlwk5pak4oEM+l/pUzHd74GrFS1UBC/vIi
ZE71sx/vTJE2X2GKXtNBKhNqVyQL+DF3du+MrmU1aKLsiq3DMxTqkScJa4caMCr5
cyFtO/JOn3jT4s3f5aQhdbPba0sBnW33VeV0HuTWM91bjhh2oon0jUKKEqJrInbf
1BurLEkCoQtTvjFEGlj6P07UaujaAdc+coQpUJdhUJzkaKz9Krustv0SDgMT/Mr0
XnCQA/dUnBUyImORoHRoJIcoQ1eFa7m+7jwML2ddryklOgDp+ER8ZhuEX3Mf3BM3
qfP/KE4U7vJGxxBCl5hid8sookA68y8PAkJGgfCu3yRSFRmc/TMDTx93IzgWm2Us
Yrc7VqXy4BbK9JsPLW/DfZ8nbybxUZ39BaUbIWFotCIUFniRsJAwxynjQVq8y8+e
47/SelLRmN/azarAcTfpumcG8jFFU0Cjsk502Uv9hOjOO/Z+bKSKbEsUlBR5v0KM
OvU2JmKbaHNGSa0fQMg7rUyLyaZF69vZIbURJ9ALYYieFA+CgPfeLF6Je0sTi3BG
WE/WC2DOX4JXqk4JsYbYn4+B+iMSAi0P+lh225wzvh8O+ho4EDSKXDfZQsOj0GhK
5vM6OaR58ftCHFaQknm5lXu/+2HDnSksAxyDpmxXQ2jnWqmd5lV/q7N/VblSczLi
f/JmXPpUeSxhcbyYFUEHOACZupQh+tgmMLTSsV0MKaefKEFnGbw8nb3jwdT+IOZP
s8dhLzN2u1l2M9SZew1/M+gYLcAoazA62V4ueqmHzqMoPUid9tr6To9JHygYm4qX
A6zSHw/s02TgOApbwSGz9y9SOXXH+VAJ+OutOeAliN8YHMR+tvUF1QLChbdTiCVM
mdnx3cYzr21x8Ujdj3T1ESg4+s0WbH3gelxfz4JvnucB1rN7RxYL8N/t6lAUutXa
/qotXuT/YFnZyDtuT2znVcPkOCjIdeIUGn1DkxLMIr/js6cQ58V6V+UtTz3gNCBN
HHVkp+OoZk7Fp+jYZGaGVqiMQ7uVcrSstlnl1mCH3TCZ9NLZoaDNlPbIQzg+Iadd
aeP+oHg5PdxhNCJk5O7NBuC+P80ua2AwDIjrNpztRT97vK3gLDgCdGLM3nwxzl2B
EC8Xed1rhfgXOOBTrX+/iC87sdSun6m3pLdv+A2EMdldBSGjVEUSk7MAxAdaDogW
PAuVQzKz2kvFMZ3rvn3CvCe8vYK1FkH5GowL1C4xiPVs/99P2QSr7RtRFRZgi2rR
/kw3FB/z8UG1LQXSJMfXJkOgOnPTfovXC0W3spGcEtaPKrnSlIs4a8XaeVsRrbzE
aNsu3x8U1O5bUw9fhq0G22FdmaX+5N5rBKPeOytTa0QPe0dhSco7rk+goxmYojE9
CUH93s1H91YnBMrPpUsyWOZMJAb2x5xIZNIqdHCQXyuRlUOzDIFSrUbjJIomquVC
tmPlVtdxjOt6ZTBFpoCLvldsW2T3+DdNkrtNsOAqnmEkNIZ9O4VR3iFFFaAirzzj
zaXdVmC/3GvQ5XX0mqzPXnp5QF2v55qOuVvHKycQ+JI4cpR9p6eeWTBHRideLf1j
NVdXw+a8mdasp+XkD0cuO+IHC+xEU3/2NOzvF0zovJBgqL27L+g8NvKvhooNFx4r
uufle93ILRFAyfIoK0wYa0LCJH2gx5z4cGwMZtf45CUsQ3XCMrziHyfAX98PPb/F
QDBIKBIUBrb0bWOX4UjbWkqyt9UlJiIkjIOhP42LSDI5iR5j+4z+3TCaLK/56w4M
9GMhdNeQWXnahYTcOrwhxd928a+E23v4MvTiF4rCY7ycd0o9+2DCKXE1j8e0a3d7
o1wckyWt6DqGIN4BZWacumsq/nPIiGR9S3xyD1JuZzkJOjoBVHlgGDUcgotgqWlK
0XL17cRhRTI85LWyKrjfsKYHsf81U/6ZIatMBhSe35d0OzArHphbr8m6fVxaJqs/
P6yFQ+yU/H7+DR/AtPUZ9dhDFPgZY75gXhnuDBXf9+y9PRrzjLWOgjTFf4aJn/4N
8u4WYVOCKwph/NIZ8eEn/DekKy4oZYmjzeV0WKR+bXWthPWs0EOfKFENPUQPIgzn
BAiBxi3NBTYMGXWp0q2i4N3+tBwlfSaIjaeyG3oM0JAChxkfyp+/j3WpO3RCwIyJ
rmYJNlVgWEASfSb1KU3hN1TJPf9AY/iVOhR6EgzbGJQpYvW+GqT4sTBXMhp64rsz
YHKwfVf/qMOab9hTDKgp3+M1QkcjWDEBHmqRhsowl+/JsnBQYxVTn7kmYvjMmeDw
EoQ4lzo8WtCy4qycO3rCl2Xee+JWHCWF2vaCgz04bCMrKIfkUGeV+W/jNw4M5rSz
rAGCPUR17i8oehlpUGHn/horZVwS3I2YzGl5Tt6MXn6B4GJMNOYrzGecEFMpEPRi
vvEIeuKvJ7vwIrjCi8IaAaHgVg60J3AE8dd/lVwHu/MWQa3GKxP4eKHUDqSoxzT5
Ig9NuICp4lYh3+QSlEIPoQ4NSaXboP9JXB11D8LV8bfbqLQ8ZrJO8NS9mOqSSpKS
SFj8Gte5y00N+0gZFlY0kaary7U+DLDUIryzKaZ7kH3vu4pMA/nRvRUMPI2A+vKj
E5VkX6YjcTZvO/yuWno0by4wP7+yVwU7lFAkp/14NEn3bq4sfP50fjo6Nu8OQfhw
BuywQExNf1Y0rkta+BqNoRAkQDO8fAFcIif6zSDor9qarHJyZi2uUgMA98UaWwNd
wlyD/5+QsMsYIW7Kr78HIKVcRIo4yX04tiwB7wt9kV1SI5nbY96mkZCbXPZD8pwp
4m6PjtM8rklNfmtXQ9XseiZW5qbAWZcozMW0yP3/J3pg8372+JCC29upKb1sGX6m
zN8rVxpEZgTK0hYCSUdnC8+pFj6RfjnFYbIAmGoEQW8XSzIVLiuVVI+ja4uPWLiC
WISrEFa9zD4bhQ3VJz1oL30NZiU5q42LbVdBXmiILhyNSIogGfAbMgalBA6Fc5yR
uj7RE1rS2IZ5N5CSX5JSY5ZZHD094cMPnhZMEW4gkWojMwvUR01Ze8YWVW9rU3Bj
SNifyJbn2puPrABdbXoFQR2rsfkfFoSjGiVz8VYb3rt+4KoT2MqYyHCqw0NeKjNK
QkjJfuk9hqlaPWdnCL9bbludXRMHmNfUPjwb4ZTUtA7mahWyV/LZN7zRDfJwbdxQ
ExoD39RpLWFG7jSIb/D821ziZuCY5JiA+Kh8Ns5zQEBOVE46aag8lB7JRsgpHMFu
TbVA5xaEhLDHPGRMswv+V2iGXnbMR8FO/jZQKTuzf6QfcZkEaq24/duysT0Kb9l+
HwnQ8hadUM2WRvoq2654ASB8pGRQUK3fLnw4jkBmpvp7JbEongVEXdctaQBnD56t
+m7VHymyzyAPEZoF+TlC+Hw7FfVQsYQp46/ODT1Urfn7xiUsCswTIwAcl893FjaM
TvW5+IDAbSd4lztVcrzJZRVlr3mH1P0S5FR6nICVCqssurYHWm5pEReXRWybkh4a
hD5BJQNfOkXWFtaJIB3qIwpJtswG8GfT1KxgmoyeB/3M7EqfjrNyCPFrPx+gBEJu
Y+9OAYSZ3pHUVisSvsO/WDv3r829udksd05lAfaZOpHwc4uHpcPTGtwojNvw5xU0
SCj8LA8yAQfhJ/AVqSlaukuPbStCbexCli19nPAF8eIBgaSGbR77jCpoHUHSQv1n
p78tGPcNEWf/k6OakylG4VZh7QnVO3pXcK7BfVAkUrZsfBz7E0BagennbniFb/5w
y7Wvu4AQBHy2UHrv6AmiiHNbG8t5e4SiEtatvgV9i1CAIGSqOdumK9QXd+KbOQ5i
4IPPrbAKHanOJF0qUqs51a26Gh/+dp/mLA+mTxoN0/yc3ERUs/KVi9Zxn0DkF2lt
17IOQgmBD97wemdLk13XImtN7kdHKb8B6coQ0E+ahtLlMi/c56y9rOTrHgGHcjl8
uwYtTiiXhQQV0xrU9oaVxNI2xP8EsfAc1Y7V8wS/P2CTLxexe64WMC06cggKtn2z
FNTYq1I/zpPqa2g72gBFrfFGnT7JUXXZ9yU9XW4I+l1lcxvMQSgxX1So8sS87oEm
UgwaVmQoZJjs+TDGisX78dzaqKb2M/tWv03dxcSpTblNn+pFE5WOUIRNKDb3SEGN
QmdvLcjpKW6rWXdD3r7LryJdKQlXIoEuPk5W4ZAWPHB+I3r1Qe7VJ7NJP9C1SHrN
sfkyIEyklkz8olZeJL6Al6gRfQ5Yf3QZpT1yktINtJl9dZLyzQxOugJY4OVclA4G
df4NJs4fiCv90CP4fwF6tW1DQqKMlKJPV0i2a+sBOR2PsCCqtdPuA8JXTz2QtmHa
BkCvHkrvlapv3/moFBTffw4khbFHpA+3qDQaLccjcn8fhCF9H8Q5LfVtekSsihqP
yPSUwgMuYacRIolf/6WdTZcpCn7INeOb12gFkR8I4g/Mzw2/5qd19uPQ1qPmlpse
A4ylMAna0usDGGJEdFSRYgNqwMCHr/XykerDRahCPXGBid7AG1vilKmI9uJ9COt9
zk1KmPealwfrOg0wZlXGvBbWwW3qzV/nVsQdEIYcjiQujrn8JbY7Uz3YewTClyTp
Sf94jpyGIjbJQduvnw90ADQ4nvolqhDyJ6i4EvxgMGTZBRWCFtALXWH0taEadsdM
Fj30UhXu3It3wfxzIShUa/UkH1QDHzspxsJ3sznFFbvfKaZ7jvb8hVIA7BBAo1rd
6RK5pQgGZ5u1rUrSmyjM1CLF3h/CEWNTEzWyykuEv5SYSmjW0JAso1Xoz0lsG7GT
u77KrUvFTbFjqzgqlJMMwt3Y6kysYyOgVCSlGpAftRpbiWjHNHmw3NlQT+LWJkjb
z2HJDJvdsEfM90fdCWi5iWkCNB4xQGwYczEYj0qMM9y/jqU9ZqJ9Ly5nbA+n9IFP
pjF5Wk65lP70NtnJA5SPvA4aWjDZn82xAXyYNrQWBj1Dg3XbIawM4WraZpiqeoNh
gQszrUB3euu+svl6U55ZTzMSkw5zFklZV02YtP8SV0vJBvgE4rGgrhRQS+WsFF/v
EX9DaioqqCew4KZj1djosdIL5PEbmc3hBj5sVoyTQ3279f97iI+JifaCSrd/ijR/
I89b3f+CPivMSLb9uvI5PM1vfC0DGbcMtvFWKudZ2tG9ItuqiKEhdd17vrXT4LDM
9lnCV9ZZ+7MVZg6CTdHPKkpL7U1ahp6djb+cKrMijxVUq+DBrSJU5IuoUJLib8B0
q+Hk0fjA4fqmJYsUghz3c9flHQ6gDQpnxWXb+g8KnXe7czg9HsVIKtyxuuddprSS
Z3QSHbPZkZEZqIbClr7R1Sj1LKPBiQqwh0YuU5Ncg8B1A0mxpmZq2ggVcdX1t+QP
YMGWN+7tYRcZKEnZ0J+KG7ZZb9Miw9o/INPVFXWIdWbc1vkKk+DBrlO5T5LAT0lE
xfHKhJqozQ+0S7AOGLZ/j6LDLkdjBYAKOYONg9BAYcmTj1x1BGO9wlwBwIytRXSG
uNrpBUTeMvVLaF+hhQ+a1zlqNHfKHdRy4llLK5eLTivR+LHYAS3gHncTvHj3tAji
XKdAd4swm7iRgiSAp8V8kJW4Syz5JaUmASJ7O8m3jCwII20AkJrmu+yqAyzl9ev+
uXl3AFbijE3GkVBuapDBKLyC5y4HgJyhfXGESYVdgIRe0nCIgngpWHWeDdlaDyQF
JDoQYJu89hNNTLjq8A2nh/Bmf9VHQv5DIt3OnLx+rjm8UWH3oR6vSORhnBXeUVCt
UDXG1AuMTwKc+ECQ+9ylPFSjzMOOsK9NZhhEj7ViI3QkZjQQVs7LLketdHaFLoUi
IFGNOHgcAcHGHiPzc55E97fU3XRH5m0ZSQeFdtJ97Rptgi7YZc3rFljvrIB3PyM0
DR/ETX8CqguaQTn5z2rTp+dKnV60QHAvh9+6e1Yf7kzP4kTHKBPCcHjrAQNnsXot
dzH2UrY6grJ6xs+21yVKDd//LURza/zdMBd2//hvTT2r0n9JorZkNKgoc9eyBMoT
bl03u2Yjz9RmryHDFgzoa3NjZxBs9ZeUI+K8OufBbpgATEmeBxz63/kGnMgU98a9
jpFexfywIMm4PXH8T5RDrNTEzGRE7TvREI6+lIdJWmHTPSm4vW7Fk+hy/jYX7BcL
Yyuwf66P0hHUpeUpkCIyjz4nzlfD+xalDtkAmSwR/M3D6QkjZ0gdn2VoUW7WcZYC
TLg6vcvwestycaERTVp2udyDfwOAzoBYKOzPGO9d7IeIzOQRJ+RhoZ3MD0tKaX0M
sKaJyXBaTHnPwK8lbRjfTNnyPH3gHt7VzjAnrrJ/v/0Hr65E72u299j6pixLpq+Q
5PGCW8ytRFVdmb7GCGQ2MolSkWOw+uPdz8Q4BnbOyWxaelupk9Aku3MZRpCo6Rdb
JQ2N+G2eLPsw3FM3njS2NiyT8OeEqqU8WJFGzSc5SZMAtQZWUjRKr/qxe8Eb8WXd
eNfeVGTjgjkBdRuhwu6rVoqkULXqVJYfjo+sOIN/GcMP+J+XFvts7P/mfnUQ5e7p
byaILtD3BJ3Q77bSRPUAZLNNKM8gYYXxNGFR9yV+0zdzM9PmyYvRr00G07Q2uI/j
f9xpC+VY/DeaFCZE5QcKBVxnaXF7RwReHxyKk4Yk3A7PRuwsbtWNrw6FF93pyCGZ
64ssrcnxzdvPaAJ/KLI+YLhBTrcxUZyBRw1TBOSa3MWWalcE2lABF40x/yVHJaE4
BidAg06RNFGbq42nG1B8xR4P1RSyPEWeBtod2AzCPuGg8ul2sD9M1/T7sSz0iiT6
XqYdvqTeccG5l8YrpsrSGMA1Ba9q3WPq/ahnXjhuwUtB7QjkWZkrDYZd/JEyCFk2
oGGHIIgq52nM0Nlc2+Nqy+F10BntbyNrlraJiDgq+fLnU5nS3oEBlAU61LFw5/V5
6iMODNjA5mQl7rbsgr22gfqHYUlPCyM0VvBqbCFFXjv2vZFk6mn0tf/9eiD4z8b0
uPLWe3vDGh9l19Pfb3SQqTiIUPmNMq+VGQPRhZCcLeJEx5GuG7dD4E85eZw8bnH1
t1pEXTO6Wo8FTW8UHIDJxz14TgD4RedxYWOQXXVm6Prt964pL2JcP3t4hfU7zZOd
6Mury9GSxIkAMb/NAOrJbxIdcWBCuOPM/C5Ml6SwpNJE/17Le/hm8bSxhepMO5mz
11myi51C5RWYSCK2T8mVCO4ifWGKlp0iRhF5YTWwYU2D4TXyE7YwDJ8zlvpbo2Ln
FTiVsuQFmei00Uof2C0X4iaPuEktfLY39zUgTU3aRtn/3gOyO7cdIuxtO9LM8duL
Kt/iioIhnAkTAWEHWa7MI0H8Z+3EkEy2PQgFoJW2c/x+22xk7SD/tq5b1BtQ+z5I
tXj+CiUnJn61vCEdt/4JgEaN5hsgKmhspFTgTpU19GsJqJV4/cRX8295qtrmEUMd
m+wBvOyp7kcRDkZYrqd6Ybga2zj4rIjJDKwasyswicOsPhZo22l9cjdlKKwcEk96
o4B9y0PFK4VlgAutqjVZsxMtLya9pkJ57j3oyg3DK5I5PSpZnvGRoG89ujfXvKvm
0gxBnajhA0xdY2YedLvLARKDY+MLHAgVMRmdupOqutDeIcUs4359A2QFL7c9xMzS
cFawXVAxI5/cnj2McUHvFcb7iXCalKS1Tsfhj2N1Tn6OndnDoaRuR9qJyku12EVb
5bjLgGrnLv8Z+kasgIu/rrNnY3oLkq9TIXttXIMxOdja9m3L+CNo17y9o69133M2
2SdNWqwAJhxEPWpjtm5ZBfPIs6FyPuXr05UZm/7/zAdWYAqghAItzo14uAV1iw1/
kuEZdBhnNa6cEiFSvoZUWhg5pxRZw1ssxWRGhCiKWYuqKwrFA3WCLWoBjPV+0cMU
JUQUBTGwH1i+2FBoqpbwu3QMLq9G6My53o9bJ8cqic25rQoZvxHtvr4nZ1lpdXFS
9aAfWskwGvscvp6433xbkMqYlo/GBg6nj037LhJvn/YD3uFpoRjlhwdY7LDQ3wcP
fYR7xCrWjpxC8hNp9KwVKwpeYS7tnGsHqQ5kor5lBWnz+abFmYZeGJlG1FGll59S
2ImHm+ZNfIJZERjDTDtiFSD+BP+JBUstsXcMz0Gd9NWbp1y6cinH89VHIQEk2vjW
kj0K74Vr/ohLwxTmpvnxWDjbWvhIBclLaaQ/7r/DWz6g/AJD47b+Z4JwHoAgCl5T
cBWAe8rrKA6cV2R5h6Q831hZE01p3yEM2K/NLjIB2pr6FwlzgtY0UtBRpdHPvEsM
xWGmbguPpgzPezuB9RKMGftIKHanYuURxwQkQ8+tR+2epLa6DE05RVoDGqPCk+1h
n/1bJIDCAtzFO8sxrT1v00KxiyuLAmsVryMdD1W+drwRfAQ6DYPkiYkHWEK3lyBF
fhINaXpxgMgSRuRblLxCHOFfegfnfbbV519ZizW/JBa4uLV8pywbmkx6p6n7cYzC
shvDTT3zxKVEbPCzYLeaC+dWucATILWA6IXrS8mhsuU1JlKpF7uwfp6XsAYH/rW9
D8VzhCDyyO74zazsCcyInAWiD1ZEOBHujbJmfUYKTWo/0GrVOeU7NvfB1RFnIiNI
rwWCseYTnbFgm6OZ3rv7gPP5chibDLkt+yxh5z+G6wy/BTp4nenxB0XFrIE28kQx
P4e2RB687u5qwEDFQZxdy2CbGGgLUDEuaB0ChnsV5JH6uDquhOtGHD1ZSd6kpBYW
gmCiK+GT4tQCqlmbfKRFxIgiAVOpxwxHkENLSStA06SaznZ6dN1WTr7rDLEwrREe
4XjZZNzUHtvYub0Y5Qarbau88xLubdjUSS9dKsKN0r3Sv89JY8siOOa+EUEle4BL
O6ciNTXgSaOQeoA2gGbYogvqojyxoxU4tfuqTK6hC+E8/ZM9+9jwJjFNl1a8Oc2n
pB8JgWRxyRpXry58CT+chgCk9UAVWFK9VXnx4u2+HZcwxXunBXEct5d7LxcUsoSy
o4MAvaceOyFdE0TpWysVdyhuDSd1QGguhTZeaDh+x/LfV5qPGyV8FxgjL8JOKZ3e
PRU5Jm/+1Toue+Cub7uInAKFvgvjEab1Jvsac9rhbMYMapA5LyrRlqeL4qVFEw4z
DN+LJrAG0FNJ3HEU2WJ6gK3ebMFbmJJpzdD9TetaPaYmKlc6N111L43UuyMryt8q
X4ychi7NAM1GzkJz1UyqZWgxfuNWpGdtaQfBdVGatKXz9YGrxnB/Id8zfUPfORia
5a1/mGwUqRxgr9wIE1M5PtkDIogPUA1TwISrgdno3F9TYAl/v0PH+uqJ9vZpwZna
EfNRmff4TY2tX0jaNywI6Nc20avHr3zXIMdAfaM2AYd6JFsPnXw7a2wvpYMUELNE
SmS77rXD3cwvROMYq0UnpuV2bQ76aODd1cR43toe1F3VBVwrE0P0JNIxKpLjlgjP
l9So1zvB5mF/4jbsrbK5UPpTSV/58WA9Lgnas83miC+QrHT1XBkwQvgdSd17dm2D
Btr0IW/OT74ljq1qbGwpFB0sci1S2O/AdcLyHWO6wcI9b3Iyj0aSEX3x6nQaDlSL
vYjXgGMA9e9Ay/z0NmxWrZTaMUWpyzqE4bOtGqZjMQqXQSgUXpdt+l/RxHyJQcrH
KU2AekAeBSHZYu1QSgI1LGPYZFCPemBRPiYDkt5mtIopLkacBFu+lVEbAQtW0Uw7
fINRI0SCqq0nBZGfXl6wKV36CVtMWhxO5A75+yfFY79Dgk9Fck8Sr5c5N5jLFsD5
sJXDGHvbLj7tBHrqA3V5O6+7ajf6S46adTGRSDMOZaBY6u05heBZu7rpXMp4xFI0
b6EQJI70qBAFFfSthsWE2cgLe4amzD4b0O3qOwP/xuIX4oTOnO97fgxDyHsrF4ka
vPLpBZGUvjPyVe26Sy3gfG/dBfi2BpRuSBUI2m/RhJTCgtLLKkczw9UUr7bKSiYq
OyRYkL5IiosXUhhXCp2j/o1Ebu4dg5EsL//zqktxcLvPcNY5+6ULn9OVmdkIcJVz
/fGhIYcJVUsyrZVTI4wuOcQONB2UjmIACSnYYKwyBu58F+8QyQrmz/4+7g87D+hg
T3PDA82o1Qfoka4k3P+Nq1PyxVRS/6lK9YD215l+FGK4gxzVqVEoo0U6W56XAJrx
W3BoUqevgmjo97J8hbCqAB9CHeIJOW2eejI09FlPtShhb5J0/m//bH7HkAsG2LbO
1wCWntjujbJt4kE5lEkyDsT8DbPOu3KZMYKzcgcL+m3RwI9LxbftjHmomjwq7VAE
NajorKnncGdgYFPzTf5u/Z4UQNGKTKn6rjGlrJRrRO+IDZCfqm3Lco6Ve1xy96Sj
4niV0cFVWZRt4V9L1tLZA0+xOKCkh12r8gbO/6KhhubHeyt9oJZPlqXM+ZRK3g07
MUP86bWUeRxGTLj3uXnIBuy1biPjC41NsEs2k31zcFV9gLNpRc/VmRwImStXT9fS
TZmIt9FHC7VvyA4VPsI3gKDswqX4GNA8qOqr3AbQw2yw+wXuJaV4L2JFi1zO2trs
geYCCV6xvQNs+bhcTHizzS2tg659Ly2eX34QQhYS5aIY2aEU5uSzfDJCyl+d80nh
KlXW2/3f55PhPHV3EKbKqiud+ZJleMUo5mXHB2tdDWqXmGVZQcdeE10Nlbkdmh0M
48R93zP5e/NZciOQgXr4y/2Jd4ibLJnzo+LqlJ1eRpQZ4CX0sI72eacG0+zxzqZi
v6osttz0p/w0cvKIacM3NNExkmWx4GNfJm77i0Z80SrwZeft66ju5gvux5CsBste
Ah9b5ZAaw7D9UXEqy+5YQkJS6RFFTH2wdvCQ6BG5UZ4W6daiLJ6z/qv+7OGqmXBY
05BmPzdsMwS0q5iKXYTY0g16et+g1tn4nPrp5dpnZzNj5EpP2NOQqjS2AQFkaTA/
OA4ROHlEoDzdEPKxtrnm2fiwwMHxHMaoUVPO0Q48VL0s4v8XfFA0Atwjrshmn9P+
9l93t3+8FZx0JnhuwQM1Svxu4o3JQiyusRSbvcXkMFppjoyzkpOQDI3yGdALV7vt
CA4SC+C4IuBa3hj1wSJkJMQI0VJF3VEY0DVCaPdamceMyuAINWL1zIUdoCS9h3TD
tGWpXlt0awkqjqch41HCVlcMwSoQS2Pwv+aIbs4PUUBYlYol9vMSIinRNRoxMs45
SkQtixuIuwT2G4O3pdTitocmsqNAwGVovI8YfyUWpgyaW2xnNElyLVAd+cwsU/6a
34JUxyEnuin0djObGWchIehy/PBltJtLHYFS/NDJWDqGSb5xYoPvsXpqeX4YeHm9
WGH/pxPcXKoNGfuUhnYXP0VRgtEuCM9Ix/bZy8OQOQset1Xo7ApBSaLC3HK+2ED4
OsyLOzq/BwOxPym2WpgNVRdQZa6eZPL+Kv5TefPU5JYGgd3bx7o+ytfjWI3NozPH
yBNqgq5AETWVDYdy/AsgBn8KWGGLqZ/afNxhD5IPbbBiLk1ncpIbSQgYHKCkJdLe
2b0ExohMf2rLpCDGX37Ooe93pYiFY3Mk+hllEIedTPGJ0d5DXD6tRIzKf706CJ/R
DmesrMilwjRlWSiYGcoDP+MP6A4W+tL6X5H9weHm2tarm8y7DcHOUVdswBKnwSQw
/lzRsHUQJwpWEgqPCp7kj6gGQ4bqzNelqzg6N1ZBIVAsrbzoaQsr+NB4PZ883tO5
n3x+PsJ/p9VTaqNuPCCWuW0IhrN1n6/tShj9XzMxhsDCja9hL7TqZccOU8v6rj7D
wqgnXZ59B2+2Khx+SjMk1FUMJ5IDzvIcDmJqyzLkj3/dN+6Z5gTlbqKXvl5O7xG7
rGmLybp2lV8jWfbeqHju2PMoPIUkuXaJoZO2Cl36i1foGDpMKVdpU/xqFW2nvLhX
KeMtYLKMiQC3b/nnXsoX3JFRUzKJKMBWGvGH9j1SspTPFL9vX4xJhpT5TpubfahH
AJkIpPb0t9VRw96Wwf+Cyl3zG7X9w/SsJyoF5wr1zXEoo5Cpw93KagqUikfxasHB
y5GFHgIlXeTci7MinTOdxDNsqF9wMDuA7V9+ZLy1fletapOpQUSZA4zJVmhWnROo
ByVMhwFy0EVT9p2c6oQb1u/oQb0gXJjMZAnHbNasc2VpoFXcVj3dUfTxF+OAV+1p
8TlZyumPgHNfACzjh59pL+RhmkCtrBJc2fXkMD0na5QMhYW/4k6rY3/9/iFG8pd8
RH9BjFZpOqyIl49rUTLAgBVdiurcpUDqj+6vQwh8KYNxj32nuv6PQkX+zag+CtAH
1FLbO7y9ax0bdITjD2EUxLpltbbBatvQBNiUenDD+nTdmE6MQyC6Y0V1RjpdSnae
/SVMIxRoFBYXADAlZsoP2HAq0+ChrsEMfcvgqymMsPnlVSOzGi1xH5ltje37Fwxx
DvovUg8VuBLxEiIC6mLPDoIKr7qh7alDmTzUq3oSIkNTuHml9vxFG/LeUf7HEEMU
ErQgevvUNxFc1oeMkaizHvgA2ZpeOrDWxV8dHY8WZ2yDrs7vqEKHw3t2xMkSitOQ
XuKy93kDEFwU15t6IkLuHlhW8K5V77Wy+Vltia30ppW8n+GXoesHeIiCmPAIbqTv
rK3joLli3+UHroaYYrjNFjBa1FdEVpd4KkK+AN/DUJfLa3+AMEw77FdcBBNu499e
0bar2EfLwrcnciIi71ovllNHVt1epKyhZbJpipvIEmtoN0G9LEikVBRBXE6eXE7+
YeamYnEaBIJKfTiQEjfGM/JtAaOFFVzfFT2GT4vWCu7r9Qwy2IFu0pNIpln6FEPX
GJgbJdg5ixRHOk5HoSfypbH2dM8v2hn4FM0TNzai07JxGW/13khOHD+H/kC1mm38
BjNU1PtVOOUMKmyGud9htBzCDhMq/eEoZm6tbds+Jnybaky4F/g+wmUI9Zdb4L0Q
MPVdEwHgUi2DwPe0kjlxS2lxwJwRS9rQIlcvlOwKgXXQay8U04h6zm8iKYqnV5t9
aCfNjicg0/2u82bRTgj/j56zFlB4i65Lvq5M0OmbJrLLCZC0tzYfZY7raf2Qk6r0
JPe0YrwXXdB2uLgjkRFXCCtrcW7l+l1jqjUu59ccUKW0pz4P+GE9QcVjXVuJ+Bkb
AHvZNANO2HttBXpC9yDFjzma4kATuXw9rUM5ZlKFuu/OAhNb0P/MCj+D7Jbyl2Oc
yN8n8upDg4dX2yPAkGPkHQv5QGz9xn5xfpt+mafHFaUAh7QwkZCB0P3MCL1UKuP2
Xh+HQskXaq66Ww+C52P8Z+f3HllZsSX78BIY2INXDKSABcRQGwaJNggIyZl5WEPq
FRBS5olCXb11e2LE0zmmaKqoc4OaSgmkUjDoTIkgCegH5SCM3AxfPma44qxNhH0M
8yvdyJf8E0otUPeLy5Ll4XMvGC0QHq/ZoQrmfmhoAEjIvck/CkspTZU+qg4xZE8h
wvSl855tKAkIyk0/aqreboiqod+/Yyx2MdWjRI/RRfYfz1Tmfh818bPxzYAJzAKW
nqnZQiabuku0jGxKh4XJQDril1hCRKx86xBUFH5/A4b/1e+E8W2U5FcrN1GuQ21q
gS09B/CK6Gp6MhAOV/4Jaz3hvTM1xGMwBpoHZle2Pyq7ONEa6/jgQIPCZN6xiT6h
0Thp6+jZQWiyTK5UoOmCix3D6Jp4LBHjwfvR+xOFH8uBihUNzbootN26/1wEP5QV
cQWyywFjPmyzgr+ncodxN/84mYhawdtyCOZRt/BZfjOrR9YgqjtzHwxOiR2xPzLY
beRu7FLIdusTVCIt//2AJ6+zDlnwKz7FZyNXvr4W2Z9/jX8TYGYgVHnGaS0ufjvM
t0CT8zn9GqiJiDtLPDB0xoUDwku8oDsHbB8Acn7XX57QmzbrKBlgGIJkXtAjpWpA
Ti/iq98p/Up0wrdCu2J9R8uP297jWe/NQXedKQXqGKu8iriFSwKGL+MgBgt/3Jtm
6k9O5VS7NXjxDyaWRJk/CE+qdG5/QiwWhuWZRgDD9UHhDjdLlTjXjlwk0fQo58bL
xj5jEJokD0iQCJ6J2Hb6rffI8Yzg8w8iMoy/+2aei9Y7ensU6I+ZbRbNOvOILDdC
VWqX3uvAw7VL/Yp+8BlrQugLZAicFB8JOD7VrC0ZUkeGI3nI14JLS4RHa1hvJfvW
iXbiAs9gAnlKR7K1Jq24XZJf7Hh+lNkU/+GD/Bm7JgfOOxcG2cBkylqLjjbYYXf6
L6dyDupup9oJWjTexZA8Lvks3Sy5s3hbn6ZRen8h9rifY4VnDB1JnuC0wBMgMjbo
Ymc11/JJwQKqYllD3bBuJcge9MBK58UqUYra1ovq/dWdnpw8N6xAi66D+M7qUOgb
JcT4xwvfSWVk3jxphFKht+dzKUVCtSUkMuSIvEinpOj+t8EK6F2IK3EzxGlnGbpv
MLZEHLMSxRrRmRxEv2b1HK719Dt9fV3ZYqockbB0WhkYTMvfu4N2uj9sc3MIdsfE
SYUo2MkUuuOrlvIhRMeCJ/f9f8P8tbGwcG5xWIPVY/PbTDAT32UZEcVDUxh0HLPl
7zaQPn4Xx9qIpzHkvpT7eid6ExeCjKzeOz67j5XHqM88/LMTV6XRNXH355pMLx/0
esPiqZxH/xMz46LDcLwr191iUPLBOexrASiO1F1T5zXFydTM7Mz3BDm6Yntsxe4B
YV4Xk/LlFYeKOizOzz8oC9BgJPf3paFeLPW4eMqbMp1i6r6wgU1g6KySWS1TOTQe
TuNuX8XrUMsEd0r/8A9AEeQhPFnjzs0+vW7Qse344j0R71ILqjKEHslRVrIXGCOQ
szuo99jv2xoUoH6Yh0dfZHDEyX/REiK6Fc2yEvbvoPde80ofz50SPcbe1WugRIwn
Zzr5/9EiQRvqX9VM0OoWpyyX+FKKW8b/+4aje7L+oMZaethcvVjXY7fxpnGbBInL
frpYKJdKB37DCrdpJ3gntt+dmb+OtqDsOYtC74RkWQVDXtU7TBkkW36EGC7W7NGT
JlM/4UMW5BH5TuzBxy5eB2f18EcO+NqfjEqMDGFIV1STU2JCKNbIS3juL/vy3EG1
4bu79HodRBop6Ya8ZUb2YWr32QmfzEUiXFUNsWxxv84JOv4yD66YLRdyRnF4IuDU
4JuzE7QZNDxqHtSxVxLILvxBsq95YxXOdpE1MfWDBgetngj52qDQz7XZ3RKQp2Sp
I44GF3Vkw5ch8UzrJdwh8AX/Ht78eRubiVvftehGC8QUQwvKO42eufuMkqj5LLFR
4zD836ru3C2pVrcdUtNlWEzy84n4g/hA/zDSz9SN1AMRGNfD6o8aVpq77CZ6erD2
7Lj42GaslKbbaVE/QP4VzBpFLajQS7MtSbi+ozf3kRzG7NKemHVX1z4l464KC8Ez
6+gXEx4DJkHafbp9V+BqBR9NS62YIkJAIxy/lEAU3S9I6QmSl9I30qfgkdGNhvjT
xkSbvYQUOBwzdRrGIJJaFnfGEZKuGnBt7GyIr5KoZdxwEv+pWEdzHO3+T47ruf1B
HxWsKsGCZiPLqw/sNoPkesL10/5cvd/n47U+daJtuRwSaBML4MTgJE9LdYZmCDqK
o4qWF2jYFQ4D93JwcWNQL4ILsGgGFqOPjFeKJuHi0JGmUQoNHROA0pTkGvUtqw2J
2VwbrCjN1hPKGS8uni3ATHrNknHS83SdkzrYltw/rIK1i44Uy8lHmBVTFsSTNJSL
0jSwXhpRaZX9xGCQDfA9B6I8JazEZ+FRNW1WfCkoS3edWOIEr1QFsRl5iW4e3Dko
v397IoGxvAYeb9o9SQHRuUhXsr4ZnJCwEUi53EVz3KDbJSSpNHdefUdTz64ysYTE
0zrzttrXlGu2pa+ECoep7yIvp8tyqHrJT991VNs5FzAryMDQh6qxiRJo8HrHdtKj
0MbYxHkV/MD+K6Yy5MWW++clseQZlIvR2iU2uMj1JG/eeLG2PnTUZq/erf6tlz8G
cwbZT6Dq87oqdh+RfSV896DCl4wk4cE16aVUvztXP+NIcbLVGD5jOVf4UnVwpKkz
lIjzm2CUD9h86WPf3UmrUOZXizsFtn9oskclc1mz6RXkZv1mXZB1zBPYj+IyjFvb
sffWqnN4eMhouF0vA1YygE5Cpd6kS/e/vtC7a3vxMXVow7v2g25XcseKyuhd06kP
CQkDPdXR3sXe4roLYDUrP4QFvaJg2BeRBmrV8LBfErIsOCXbbhSkZEAYmj1tAFrJ
+zwOwrIWrjcrnOVFRVnD1Uz02hMbq4xUXFt6rk5w7ZmO3h5w6PibsYOzmeiEZcDV
/XK5UQvRwo3WusIn0gjt7DLDpl1szN6veAsTJI2he7EQjIcfdmEz0zuU9iFZL7Xx
bOvjaQ1oz6QIcQg4loxu3kt/RiqJKFUrepoRgB6pFNEWPC3mRb544LEewTQYvy2A
HFDD/S5CaTOD1YG3iQc+1TDA5IVp4Zvu5afkn/ai9lmIY3zvrmQQvJYpNSMO4r9J
5QEj2ZNowMYfbI0Dedf7XMFEV9zpnUDiDLMIWQJMpa8WXAoYx4gLPLA/eDxsYLdH
OmNOQvemgpvqLcO/huEa1S5LRunFDPiIvgEehW7IPzi7akpZx5cRbmhP5+Ge6D7O
+kIm6M4HnqHrG9AVxuqs5L8LkuNLJb+oi3qSQWDN5jXsiW0fxdnx73lxqMPRF8Mu
SEzWqQi4gr110dJJkKH+lu/AmKTesvcnzUp7XvaZwGTIDobrkHOLu0TTVSRa8Rzo
y6ZUeomTH28jqHka1tSR5oJMg8YRiIdHRz75P4r59z75JQJbbslQit6lw1pmMg8t
E5Xst0N6rTSBDZXkkX0hRDCMAai+8SLR21NnSmFF2ZBDN3P7ZDt9b9MRJGZJCpeL
V5jUgfR8IzY2MrUOt7xVB0813bRqiU6Kkvh9SdwxDNdl+05ALB7ae5aeEOAPsvsv
rGE6MnhqQNdk9EOA9OjRD8DKlGQdspujilLfO75fDMm91piYJTUUG0oMJdSkMikY
nttGv6hy45Kz/I17Te4Y3AqJeNIt2ZHML8bsKxt3SuT10pVrvh+hHdgx1QkrDLcK
a3bSYFktqKYc3Ag4rq3bt5S6UGNe6nHNvbSyxe2QXt8fJCoBJHL4NRfCQsKy85jz
h8B6SwlAZTvsvoCF6WLSN8NKOz/ieslgmprEv/IN6duAES1QdSJymi0xwxOLo9BH
XjMyQd3UGhPFoumAwHx2lfP49mept8c09gXuwjAWhq1Xw0b3vamvz5NAAErPizNa
QMKqLVKOABzI3rm6ICCUK3TGhdAH8bIaXUTzpXwpfk7r0j+i1dBAEVkp0q0v+fUa
GsPgmNukB0yoL91oOrX+Fa6nLcBrtwhHE1253jgLjjOep7JQ/cCsyLCwc9ZrvZxY
47nwLYuBaSfddi5a50qKxLCoPu0FQleBvqAktY3yuc06g+19xTScbeqmlyh4tDht
L0xq3ZwEXbDFt0HONJQ4uI+ZtczYuMl5rJiJYXwih0IXQevolV0fTwPY6PO3DVez
4nEghxPfhZeuRsoXcjm9VAwSO1IXRefixGoBjNRMhRJ97B+tPyFxm+vjNkEx9TmP
4qHDwwQ7qiVUPcq4sYqsUywvBprLawY/vJdf3MJ4ZtaynrKP3RvxuOi6ipJsBOaP
N+D3fGnbug1a10csUIWjp7up8lxaLPtny7TsQ/KDkMKFR0EAeL7ILUv3ggdkBYhx
mcTpWmgIvuLbsJex+HGa5ClAWqIS5ChpzTc7OtD01WqMltEGKguXmyMesFKY1pvF
CwjLHiiuti8bHDtrVKnBwUiMCLjXCN+Di6Ycu7Tk/HHIheVs+eaWT+xJ6lsLozfx
TjrwxrphNhtFYPT/geUCHF0ISGC1wKbht121SENmhGkGLOa/7X2CE8njToWANTlZ
RHVFm4zvMjXLYkC8L+GTwpefk7YCaV2qf1WV15LljCnlFfCXIN2zc+mXE+DzWw2E
kKYDJiuc0sKK+aXMFnRBfQ==

`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
B2oafntcZ+fv0MxRD+8sPi7yyiRjFDqiW0cSQrPnFQGPqFrd2XybBGAETOC2WSq5
a8CGiOC2nZWbG2vhxuo8bvmLDAZD/i+DptPqdaJlvITefSXb0DvxcH9rCaNxiL9n
6FY1i+0AMcUJBqMJ+rMJpqTdSTSaX6FyMgGzB3kwffW7bZ+6Dtct9sEx9i05QPJX
eSLnG//90vsDBZbrmJqqCiVptrxFeLwaDE6pCBJeiKseWcefCwtE2JE0gMTXXJbK
gTGiDuJ2+gbYA2PFPzR/6MIS11WulQOhfmztofcUz6QEegx4NOcAMBokh0wqTgBP
VFJmTzyTLJVKEOs7K2Y+2w==
//pragma protect end_key_block
//pragma protect digest_block
/wBcdU+/4JK+wbOadfnRI48Ea+0=
//pragma protect end_digest_block
//pragma protect data_block
bvs8i2+63Chgb1gPSh3f7M9uuna8zJRSoDqPVSP5YVOzpWy2PcK5d3t3JLdwrpKh
owYfnbAtg3mfKqxC1w3quj5nwVxmUdWX2n0K0BwGy6FVqvZrDQfMvqe1QyP8Lo1A
dJniVL6yWXA/rCkJ4KBQj7MA++l+uzwL+FDTXSYw/tyeRC56Rl2mpUhwsD7zgUUl
ImPxPeknzOc5F3InSwAmGzN3/4d75TmmyxMfVj4aYyChdrJj4EKlInerZ7nCld07
xTGdPBOGgpMA49WW8t8QDS4DlBMxUH0EzZNkZFMxGDuqiTwG/M2dhtdxtWaxj+Hs
IU5tPQYIdccSPZTFxmxQ+a+MbTpGhf2bRDUc2fFJ73PLYWjH9uXEf/shrI9pZ4kf
ysFeL5hTUkdXmUkrlbrg4E+DFtew4/66HTV13mPhmq2Wvzm0214ZgIozNK87fVe8
TfQscGZq6mQ2Ny0WiRT9UjHNgKnpPLLzbJf2R4UK4oyrrP1Zo91fYNLszSxlEen2
Tia/DvuL99RXfZnXESXzx9yvzyPlWDGYxLrNythFXPKx5cwBoPGd7JdskivXqQdG
AES854vKk8gVcd4fpn/ykbIXr2IOAzdE6MOox7+mda6BE3ValSsc9wS60oLspcjw
vyB/lC+xK+dPpaTL8s8Omy9JqOrtchF5NeydGBIGCCDW63AG+kK171Ub170yhSuA
jsOcgUMxFtcamiASlH9tuQPoJFCKacRbYU8xL5TxmqMGBawOP1W/IlPXzJsn+eBB
rXGfkacWiPSatdqLgzOQ3CTMCzvE5VpHFI9GBpp5MICBbrH/Tmr7dUPJ7lqooRC/
uFNH2Brk9I7gvtYXoqQnbXt+eVkog7zsaAP1uY1/b6UWeUHEM8O2EA0xZ/m/NCsm
XDLfWWZtOlkFHv5XCCze74d2x4ENz3MNi+Sr83BGBj1gPjJNovlo3HkqNA4iY3zu
JcMKP+eKql3qmVNqVLzRojfCrilnMV/LxITUcsCjd0KB9FmQ/dWNjqBBl35SgLZ/
57G5cgd+BtYiwv+vssJ+900AsgBtnXGfWSPZ9O6KJOTru0sMmEHThpBK1gdxvx23
Yh+40KW+ir41+NaA4rjwRvVdpAN58IlFS5bvLTOmMfd4J5lUOqoFGKAqEhMaWwQS
hR8VxzJLTsjSyza1rpXpprohwGihASIxjkpBcPLJKn41svI9duVCLzWzY04Mee4B
FGKQM651ow6dgCZK4DAThPmQXiL7OVKPU10G0QQq4jU+SGg5N3L3s3pPkxQj1XGh
X78Y4HejD/3yJzGoMfkBxEbZUpIvoyhhcgvaEvbKUlBHlDK5PKXG3wAiz6eMtcXv
JNMD5m/ni6zR9HRhKVKO0U814KtUs8HWtb4+eo1uGlTtcihPpvtM3MBNv/ntClpG
8hZr679zUWBFtnPi41YU4NwtGb8wxdynY1oIu1jjI4qIKUcN2rIUpYbsjwM/Rn9Z
3+2Q8ChjN0VlqDkAS9+YWdsDbb05jsm7+F/Qvpqnq2OxydcNZYPBVhpF515ZvqCa
52ElK6KrgWmZytLZlZ016cyrWtccZ30sju3Pcsi/+k6jlL0/3hPiNIFCRgKWkjmp
ZU5rK7bgrBYIrXT/AJoR0Ub8w35tGBXSgWeRJ52Vm+BAcqxVtAjvD9lrYsrjGd3O
Dr56Yitr3N5eiPo+acjwT+VnD3adBP8PYACGc26SY3JaD0PDltJ4jpNmvCol2uLi
TLrThg21Z52IjaLCOJvYJmXBfOzmZKeHxbTbDxhb6DYeMkWD+w3uJ3WgkMwi+Nvu
Ig+qY0kdosOW3a4WeB/1FW0V1UddLBqVkP1VWJ/jFpiyNc64imYTBmNfydNnNnjg
SGiQzqmg5esMhotO9xnAJ3IANOVavT09vXoohQ3wFjCkIqX7a2A+czevITTE5zMp
QLZmgIIFT7tWzQtEI2HOmlhxE+Mr1vL31y8KH+Xwd115TTjx1F6uTQ9u6t5GiGPt
h2HhugPzkzzX+BRxIJlUbRrz1yzqkvb+XCqkjZQdmWuh2LtacZCumI3gpdlwEE1o
qw3z+UimsRk42RQU5NCdbA4KNk7qHdcXvEOOkt4q7V6q6Fx1uhsSdjsWdPGqf5d5
ybi5C9Pzm5VboBWFhkiiHArqf2aZbkI0VwT+6ozjS0wW3OTnF/ujf+/ph8vSmXE5
WQivx7Twwmws9GaHiRw2SZsgDu9vdauilX2oj1qVvQ83Ug7iiDPCzcZ+DANjWdm9
ywggDFOMGQ3Yy3pUnXW8PzW99v0kqYo4u1q7dR5yePEU5dZNcIsfuMuXc1ktXcSx
Ozq47d7pDjH4vvAxEVL1sPqiM2rFFILzlUTGl7Uo8xwImpQti7X5EIr8DyVRqhoe
JydCD3t+2ucexOsJXe1h2/iAQN/wAQ+Pf6el88iODk0ixoNwQWximDeqLLb7925p
EaeliRkYXvlh5qCc17QDBU1M8QOdHpvY/YT+s1EJl19lXesWgs+A+UMHdF64RKNb
CDsUP8lvidJ+bhSRLMli6i0ABucfE6gZdDfs2sU3i2YDTvxrmf4B9gpnhKkGxc6f
7QrcPgoBVTI7BtwXvtUGwmRh+Tm+RRvVUU2ucGPskfk/E2XqRMXRmxzT9ccWvwVE
psKNm0rKmjPiIwXwaI5cetBK9f4ECmlw+tyCBrmwMUTHYAZSSC3LRStCRdCjIxDQ
NNHk+THgtpYk7C9cAAt7HTejSJ4NMsl9JpoRDIKF0ulHypXLFWjSHJqbA6NbxmWN
KOxu+J1se/5rxC7zO4+m+E8WXmAvuyTbUIKoB/Kxg1d1IT74benqCtf5I8iVfSN9
b4CdFt6MIHzDid2wf1VYBjRQfJtYsIhaqBYUIrw0QVCInomaB8eZkypD/1Vh2tAC
JzOk2D/SwzKNmlvKfF0TRt+zsbSK6QnVGBYwd5YNzNsm+dy6gGriDf3df62NqP05
pXULaPeIwqXO4XBskWPCIkkIWI6bZHS2FHGpamJgkIfLyVT8Yq6g1IfKLCeKLGw8
uTq8IKDCjU7qMrQV4NYHBVF8EWQ1KNA3ozXxrvpZdVI5MGszoWCu05HR6oUdG36Y
RjlhnI1gFjMXAhyR7nFE61vLYilY+gI9ODb6C/7Fxtb0UfeQd3Pi6TFiv/j46uaJ
sHSln/4CNLOiwi5cEYd2pUEWajfkDpvNOBLWxvkJ1REjZMme52HhqqfcN1v6vhqi
sl7q7tRwqnANGmY6xAtRU8bVdj9reKjpUHzfACKiDjEMHgKuLjCdXl7C4A4xTccj
kAizqCqA0mHBI4x+KG0u8CldYC+B1VA8p4w4sfc8s37TyuppJZeQi/mC8gCMjL6D
fxSs3lgOZ2qANdFNyHAV07nzPPSnqmshzTmHpKHDGk3zDv7E24mw85BkT2tOCa7I
nE47TQn3s9pW9tVpanpz28CyJlAsyGnUieXKl43RmBZsSccvHtK9ozFqIaRMVjpp
JgmjmlaMPy8KsB7SzzTiYEqKfrnUtsz3RH42qwuZLfbOjM0LFaawovqyA64KMwy7
+kjFt+N+3FVVZvgITaclg5aA9rRQVbeDBIwXAra8tAh4nnrf/Xf9AvqyvUVtbOCK
00gJhQh9h3bzSblm/iwJMoe9OMIuHc2vgTXk7flRNyAA8IdCaCr6dea6QMXjeywL
htRxGXraBFNJzxsQmOpDujToebqqrue5EmdG3lfppTgRzm6qq3vW9hrGqRk6fvR1
ZP6v3qoC8Txh4u8ibqMCo0yn7zi/t8ID8+fiew5WXptcOWclm1m522hsyd2yXp7c
iRJB8QJHzmOmSLaDVE3DPNJINorSIQvpFDKhSUf2//NWcqiegfBgVLKoH6thmvdp
XAfZTsj7M1DfG7t9fTs6/uvZlIMTrubAkzMdOjAPVPGZr74J6z4eLL5OR04osyOP
AJj2baW/7dD6DixssbQCrA+fkJIcYigTK/pM34dVlJNzNEBGFqqvDgvb74lF6dwT
VfmwX8OruUbVe3crlD07ttpXvAODE1sF6owKC3rVy0nWN2QaWWsJSdhKD0tG14Te
e9/wm9sLrA45LlM/dPbitG0Owbj6myYCNBCGrOQ5eYgHbf4JaaSPHHKCClAzqjVK
LY+4/zujaQC9e8pgdjCba6WutJ62Tr4Navx6Icu6nE8zG9dXh7fWUvhMthJ+yVT3
ilN8gCb7+GKJ5uzaSLVkLaUOIxmwvUD2Xd2NADITW4Md4gEjLFaFsijuKHnf+uay
XHlXHefdNWyC8qyhk8VFXCRqToPIUcepBf2WMhPDPky9deK3R8YY7oLKX2MvhF3W
cAEn72njRXD3O0iPCTu41nULUfG3dJwH46cB0kr+I1TTxf14E+YqBhDxow7Zjg1i
qzB/fZz6x2Y+9LZkU6TcZ2E12S+RyEED2q1rDzWClchcf22NZ+/Uz9A+V+mCHApy
nDYzdqwHuvJmFmD0QqdLOr9r/ni6a50lEcsjGyEWSdm6vXvtwzz5pajwkw8NK/It
f8GNmXtGubLHVpf9rJY918l4rXJioboNnOe4z+kovSfoPiuwfPOA2H/3jHaMuRc9
IfTi7QUJKsiuZxKrhzNEn3M1i809w0Bvg5RGticaIlFWvNERygrGBoAanp4RwsUj
rMhL0sl81Y8D1VSLeiMMNSmuS8A7oiMtcnSFYSWUTg55FGzGBByLamhfX0v8e42w
eNlxm+OyVTvZBQnzYJJYLPkJtRg8NMblzfvAqEmDKewg4lLP8OLvHz2I4VT9PG3X
leKVOjOs0XxWSpSAlRIjW0unWEe2WQqkW5roo84q63HWLRjvmB3ToAYOc4wtgeHR
AdSHaWjWS7xG00lsJ8WNkb9U56Y3sdRszAqf8xPEnsqZ1m8X5eObkw0S5lJENrIQ
ttAlhkBd1S86ZHtRi2RyuVWAc9ylUyueBvB0aZaX1OwNNJOZ/4z8pRB5oPSvGkzv
nDu46w6l3gfOmPK0hjLU1l35+sqSF0zpDICpZ45J3pDqzuxYNJN637WGRjamVB9E
pDq8et0H5/cBDlcVPrrpC0GHdMvvD4+bR83wWFquAq/kLzG1hRXJvYkYokBdpWe5
Ej29qtoUmfWJRKp64/88sdszLO7WJCvs/0I6w9qTNNv7Y48GaWgV/iLPnBzZVoeA
cCYLsAHFiLHrTtYy/NiXRHfvvf8eMMrAMtEw62iXjaxv4FWZODkhQ9Y+JDxgUgTT
kvbTNOyGEaWCbL+6PLpDSqtg08/1FRpBeFfLy68SMi4/ao2eKJWb35BC8+29z0XM
EEDBKAOK1DmkwUBHNkRc57OJJpTWV8D2RDKLl6R2qWPIJA8qKyTpbtfwT3RJrpE1
R3eHAteGnDG4qP9JUUyTC8yn9JkYDvgxxtG3bZ5PeYYEomWWCpLUtjaD7m7zCnWb
yiDezwkC+/rnwyrB35HLEcLY7MiU1vhA1+BWmqbaTeTIpd/KRutwO0hVw7U3kcPW
59NbyOTiyDjn4WN7MxdlvVdCQgM9s1NfhuaXqXd3aNoqdaIZ2PNASN97jogA0Xr4
TOk2BrmXAKV4BnB3YA5IP3kfZr6wuUOPgURxM7V4LB8U2DlBqJbQWQZnkcvSwELO
/4kygx3JKi2H9cHDYwtMVj6sjz2Vuynn6NcllIXWfTFMA0JMZtp/9UivfajdEsHs
bVlYxiY7rCjQgTj1ElDboBwmDOjrN0fFQm+KMszuhVVnFlqLCWOcFvwDxIGjz4g+
s+8PIsUfT2hfYrTCLV+iFAfP9qnA8ax10GlsIrgmq3ux1fcVIREkwAOaftVbAym0
hhVpyRBMZOt4ofNGKjgtIYbv4eZcjujgXWTqYgVVf2DtMqGuQVxlULMIitRqdNYV
ddIkrJcth4pBpSi6hBNY6ECiZMN1DHgKYeRBkSY8euc5mNTJHP9cT4alHW2JDR/c
SLF8I9xxUQd4AjvFEIPOXb5vdtfTtytBGYudl18hmGz/vqR8TBMa6gERoYQdZqKc
B0OU/17LYgNgPcDtr8Bu1uy05NmuRewknYzh0B0FawY10j+htoZO7Wnyz4mp65aZ
MaJuCIpSH4KCmSw0N4pU2PVteXXS8x0Rgm/CVeINX7ROjzDoX+2zs6VJpNEnsSHM
KWCRNfO1FuIG/EK2/lgktoAEaf/er4E4fUo4BM4DgzmRKnbwn2DBZSk2FBX7PJTw
YrEqGfiefBSsN7om1+py/4aZ4lIQLmG+az4Nojwjxa2LuMG0UDl/6YZ+A7sZPuD8
GrNouLuHDOiXDOjjpezMj2BN/C1FaFjOAY8YbJkeTTsB/0BbAUs6uPK3HGnMkbv1
HtpXDcFXgwiuSjXB3nKfUuosr6lGHdtb1A/lWGcvx8cetPvbL7jHW5cNh2GrYZwK
qNcawdOyqKmFQ/zCqvB2If0eFz4l8ImoSYMbA0rNhNbv93IWmBlBdh4+qteeoDfE
uapFlxovgsy5IgtsaYtmFPLpjJc9YmntP4kpVx/2KtMFrOx8xp4WpVhzminrRDsf
lP/dT5GZFVPaB1cNHdtuih3MlBsk0BZndUBQfu/MtUJmJT/5YR2L2xVN1/oOOnCL
5TzAkNYjmXvG/+GVlLBINdnjWoDLAgNSihdiMj37dSz88HXYyxVmXEQq69XRVb/2
COVs/0epjhunRPL/kHBFVhitMPH4fvOthPD6+UNJcWuoW4uZiHTXlOMIP8ShauPa
9QnkHh+/Vu0JsrWeMEtToQFyDprfofotP58eHJoP4OYoFwZ3gEp/1BS4Yix9eoZ2
4DGvMzc7ahsOrYNBA+gM9gIYkOrkVwxt05XNJW5UB86PbpygshBZI84LyceN7GE5
lMKF7Wk8sMLw0vyH2p3EV7xIO49rr0zY2JCFQkHnQTYuBMImqFWR8mkhqIq5M8Nh
JgG90QvH+0n4xCzeh9giUF+g7nh3/TyFCwMHPRlzJSNOPeFiELftfb1VpGDM91lq
0Zw2U0TJrW6LjkmcaXYopmY/YVcttv4W3/nfNKpzJeuYxvQWDtXejN3mbmA8BfxT
+CO+jSfH2AKYrBHSiyK1BlxF3tzSODXq1zIK2ZvoRvwzSI4BLuYabwThDXFqC+X5
ZIB1k2cTqo6NZaZd4ssnR0NLSd8oXYnoI396im4fiSR3Het48Ko6RUn/7WVqhiNJ
opJ9NHAl2Yc2o7FjzDV9mXcnwQsE00XNPuN62XgEKOxs8AktHAkyp9Z7k0sCzLfC
z2PxOO2ln6tynsm4VzryygM1TmS8RHOz+RHCDdE6qV4nJ/UvTv+gLpEoHIgR0wrY
CQr+K2qAljf84C7Iezap//nFUVEEjDIkvQwM43eqwUjr6DhskNthBz4SEr2dTz2l
aHGRp9yrSs0/UKCsRCVuXOWy35999bqcKx0iVf3Y2SqO1ZGRPfWsvXRDuC14b+at
lv2Og8YZPx8/blCidc2FBRcncFtw4lTqVN6Vs8OE/S3PMlGgusvMtCaAh27Z+93t
3hyEMoJx823bhuCmtSecDBBkKMxTSDCg4NFEmU+VHTrUlckIyHZYav8pzecBFqy+
X2N7FttkdW9wpwcrWnqjecC4pqQKRMgaxmIxfhNAJn8RGjSv7upJ6VxugFBpvPE/
3zYMc/NvPoXqg0tT5djHCJ5z0xae6oltXK6vdBjG3WQNG1D8mnB39pBN+bNHoARW
tpXO7rjZRRW7/exwnLDEw4Pf+ZM+Bp1no3iRQxIAwgVIiom686SDClPh7dymzvSN
t0ow79G94Jo2cEbvxG3F6iC0Y3xzNgGh6E79iwM3q+26e/72qJFy2xKQg2ilVsNd
aH6pNb7heFuar6+HFPSTQwQc7FDokurZpV7f42gwzUxQK3JKYIh6JfDFSCAMBgAC
W96BM18Nk5EHbrUrj0kPI961ktXDjfx+buXLqsVG7qxtjiaPAIA4imsSGc5+L4dP
4P8WwKBq2jM61Y4c05mGjQqw6HzQ0KkNsrKusTtpRmJERwuDX3oriyWYwtmoFOue
MRbZwF5yim7CMvrr+thz685/LSE7N7ggiyu5tvaFf4BFRC3ABQkGAAnCuYX2i2dS
mn1PPb4usDVpS98LetIXxRcw8kjB5LyOgnx804cjGiV0HD0a5+BIMa7wtKUR3C6j
9C3VMUCfD7iLpR76gRE2pvh5qbgA2zFsDmK66MSvy2nxEQDPyftKwyvMYzeA8/uB
h2oXltsG+VPLIG3TDx3S20it52U8ZkD2BhdUgkl5S0U0VS4gUYvlUdV3UfX7fkIQ
uAfHQcltTrSLSTgysIph54PIklUOkYF0fgmp8tYJH2iaYeAJrMfN+sdaoKDidW7V
N+jjhT3txlaOko7ZkDH5+MbLrXyqjZwJOnQGjBdVL/EzFpt42CnBAIPbjx4n1D4q
OvA1FYAXhr5qYqiMujuWzlm2GwY5+FdxbyA0H0ycKYSH3zy/NbjXYpuPc4X0nhUI
TluTFlPOpkKyVs5W5MwVIw4db8VyzveFKGt97SK3g5GaKbPo6aIAAiwR55kkiPjW
kQlg4SXo6apVpZy4z8/JoOvv9htVXDH3OuoQ7nU1F3T5P2jv6ssVcmaN2QhqKktK
oap4bIdkRqQog5na0tf0LRswwo98ROOxgyNu1oVOFr2/LPSZvzco2FUGRk72ULO7
gYEHLLziLfgy/wueul4PqEB0/UY4XY76dFr3CHDloUHt3vzBmzd12hmTie8rMOmX
oAVzWtPd4Y644VoXp6/nFC4MDhtG0Tnft72rZ1tq+3bkslwUTbnFGkoWo9hOCRzS
N1LJqRYHwH8vZDEPsCn+RWp8CkbwVgmt4eXNEIzaeIvwO/+9rhnnPLxZL6q0Ew9a
4upqwik+L6m6tNky9o8oqtD/EOna3gNPJ1rWuCaLne8CxYuXvwJmZZaTTQUUo0qo
6TRlC9FI7axWQChppbGxYfX5tC7rlt08xrYpqelmvyjdOvCFgIeKRMucHx1HWp6K
hbysnkNZv7gRooJpdmKZ8fe3O/Cp2rrhy95pj4RAngm2WLwLrlqz5420JwtBFrI5
hElvKJW345MN1IlURZlIR0NQPzbI6PuTssHga2rXicr1qhH8AFdd57Be1nfIqGVA
haSnW1Z4X/AID1xlSINDkM4bzeloLhpTWUXmS8wigpcPCjHRgk4FtICpcxvb1pgc
C/5MlxfPOYbj/trR3C4bmgkjXMst4ruMMTCV9j4TzVRGr50hswc4vkjzFPYWI+1X
D/T4nJR4Oqi4ZvxKto3C66PaCYplw2+ztjq0JjSM4OHsV+t9s8KRV8yiqTszldjp
EGdcUqatYfsYxN57K/4Cam1yf3E5pJFvZJJN6UTTlPWqGhpyVgSgFeiTtzzd2H1H
wkoCnyuANwZd6V+ke3yQzZ/Db5iDbZimLNcIzTVkepoq/7sJB7RzlFGwaWtvqhJi
HwCA5RHKZ0hE0aBhKuephOCvKhSyeds4Wa8oG0+1vYflT7Zi7+mHFuKZq3IIE+rl
okjPMLGrgvIG8tw6vJgyds5E9mgKz5eWdUw9j7JvEMIR5rrirCnXloQLAnF81rm/
d+Nlb743O3mfgNjtYCf7h9UThnKBuzvGOZptiU3jh4LahH0Hc3nk+VGc6GeG3PHa
ELJEfpOn9/+Pku2hXtRucBOpQpxSS62XxVuWGx7VTkEJ3nJlcIA5AFDzwRqJ/5AY
CPM+IeiBxImrlql4F+lNP3qlG4e9ezMQZisZAxMLpWyy53Jk0oZEHiP6vFJ55H6r
mTpbmderLcbcb3Ax6jiYapXSD/3JjxcsA+ghjdqonxu1JNSBKjreze5byyFm2fS5
xYyNR20OGTaV8rMQbp0Cb6pIYXY+89Oge5eGcIrFfpue9RA8cUcPoNpSwsL87ja2
swDzB/72fQQG5J/CEdUBHBDcNR2h6zb2NcH4s2bcQEe0AYr6GF9TVlYbc2zMzeUk
9DFrNvX0Gnjl1BTN7auUDqu7absKiCIDaidAyej1UpYNqiIxsB1i7LCr/SMrGaS6
CE0+lizF0iZ7YmJ/zAuzlsbbnFW4MHJaxN8D2knsd44sGrZ9pb1E4D4y2ay9mxn/
wZ/c/QMSDzsUUodNr6e4/57ssmxUZZemDi4Uvu3Su5lcwmKHX1oQmo2c2eFHiuno
bs/SHx4APzVO5Acna4IKnK09nMA3S+7c4aZlzmHAAVcQBWT0ZZTqSkNqgiszG+Sx
R6zqcZHt57gvmXajD4vARTx6pbfRbJx/KzGtF1t2BXwRWXI8y3H0O3tkvbEp6hvO
5v0pXNa/jjVLMMnaOAywAxoDsr6eT8YGQNdKBFfgAdEUgnTqoBnBWnAKRCn7ZygJ
bks/k28MTCwWji6c1+mrZAd1Saf0E2avIE3/2KzL8+77Kuq8wCxkzqAoUVxcalm3
aLXSwDB4joOBPRLAeFYEW0cl9v7pHXQqK4MIoODq53qUc57J3uVlG5QbuwlzCITH
8fDPMFgSB/Jm0RXlCdMemJXtKzvtMTCRBRvRgUxI5+tYmOiC9LyPLFZ5Gg2IJOwP
0nXfRnYgCoTIZeYXBnMRlkfdRAoSA7X8uza7rNTIrXw9mD73iU6b9nd61cNs4jk2
WxabqWEXQsb/rdHZyluRNXRCdsRWaObzSBL+5mDJN+is7V89yO13u/1YZ/XZKaO5
J20hzsg6REF+P0rU52PLNu4bPK1bQky67WiP2V4nVNpWO8OIylS7VwgKjpOYQsXG
4iRe2zCT1vrvWVJaokbfgL9HVhG+Tzphx0tx5VVixV8sRlAVT4TLTPfgd4Y4FdQl
juBcyHpDeOkDWV+lcX6hY1khD1mz1d7qLuH204fmEkz8ip70YNugeMExk2LZJkbG
pg7T5PEAco42AK9sJRrU5A+tz/f54s7eLkXXGBpVgYSMu080pnb0jVayCGjdIipg
efqApzo4lS91oi9mLFka+ZdteXHNnECn+qqKLghUDnaXhA/FVYqCZy4hm2vgvzUD
niuwh/ZggedzcBiE+yiq7ZTByiYfvrjpmgvaTXIlSj24/q83bdhVI6SbTu+uO0tJ
8cviBLVjOVQoEgtuyN8n0xDVYu8VIw+Kl5BkJcNmqxyoMIfLhjc61MSNR16OpgTm
PZQOx+LP6MajIHfeUO0PZT0YFqZHFIIfjGKRCeoHW2QMrUNMeJc60ys00x27yS97
l0WhLxaL1QJn5+JB8NKDCYBAp91aXTfLqNAyXOh7TSkhalyB9Zn5YvF/018Ea4Xm
fFHJk6FDbu9+V58iVg4Rh8VdH/arbLMccTDihoyPgxRWqJ+yQPfZZptDUP3YrYzV
E8zLmXmfvXao4fMTzjVW12ouoa8fYKTvcck6l78mxG4RYlZ1P1pKHTZD1nXp2TIJ
gYYnhj7ZVMtQSiAQ9rekK+oaQgGzO6rtojrCw6OZ12wlIE9iGl4YLKN24eLHKIhS
kjOcWKpowclZP0Xfiey79uqqMyDfY02pVmo6dP8/BJuQbBmxmt+ChsU4zwi31sTo
+sBBMdOcZrFQlAz8DacPusI2uhE2WYUZYlt95B9kpXfSbA4Xap257TWKCalcYG+v
ZaR38+bjFLyvDMftym4ntXQ+fKdCOhH69mSPUpON6A2ryoL/GEVlTZ/I9LDxRsHV
EBBf5m+FlpswZLGBuzttCmeLaphMtvgadCh6jL8j8YvSr3qpj92vMKfynCUK9d2Q
VbLlHOa1RRx423dSIxVsjIRDMBW6w3v8VZjudv+L7IBpryMcqWEYlkEaNR2BrYcH
5k5vgOcb9aDszZAwZxNe2dv5udV+SglE5X+im3211oQ+pvSLYcb2nGcUVoYX9hiI
nQZKTtJOWHcn1GhZEeRU6UXjWd60s7ThMzUS2d0Edy0YbzDBE2R7rT7NnwlstJeB
yRw6XUbmJXq6oY4f91kxnlmfWEzPyiZjnLEZyVCV4pGFusjT0Hg//adxvgwhmpMX
kEbraKEMoix4+1H4Nda+hC9QGBGBsiy9LOgoNamNhGdrTS46V7AwXs4Qw7YWxfbK
k0xMBRSSgtOunGRmTiMcfXQUWlfxwX60LZyxKVPlTtTDp8LRGyc0Vw9SMnSSEI7a
8eWlcds6RGI5JhRyv1DHnGSRWnkSIRDG6cOBIGH0DO/TGBXjbJkDdDqJqrAar01J
3B0larRG/ntGv+Z6ZtLoqvH0XcL0NGOyZvFjeaz56ytcUi3KD3eMmz1WcLRSjmhx
ddv8LkJRxZO7WkmxeuOAPKpuyVZg/EiFF66Io9KWfJfU+6ujBW4kvRwHqv9xGdKK
uj150cGrJa/iWkCAfusX5GG/C3tb9rfgby/GgXnuoARcfsR8eYqhhcg/l/fcREmA
3eJuxWaVSL8IT0s+ptU6oHuSoIiilbeSs4e1CYiYyNEYTdHxczsAYh3l0H1dek4y
RLBbKFdAbIe9IpNdzon64m+6ku4N6z9RJeh1gokQtkGeyihfEdDIWy9kfVlduGHJ
9hafYoqPfVgSKOXU64ZNm1NVSN47inx1X2fat4nfFRrsOtgyCFMJJ+nu3kWy7B5m
d6KCJHFiqwdQxfT75OQU9t3yn6B3oFACcdWeM7iQZxedvTwHQesYRL7VrdbzgyM3
STMpjxR/ouWHdUVv90gmxxJzymPolzDcRrht6K/b1gMt7e7IyIARYn6AY6epXCt6
SbjDZZb3rgH9QuLumt2pT5PX1MfUPpHKO2VdstyWfP5rHGrE9UflLZzovK16jwVc
bW3CvMmzQAEskNqASTxMYW7GUFm8cWSIfMFldMN8rGMXrZm4ZYJMf8Baz2FUpMPP
b6otOnE5GGg/9R4VYC/SES7QsgXG5OQnDdWMQRSgEWOCl/NXeo58kLW32V8lKE18
t8xgmfYpEmsGMjXtVz90P7fQiVSJZn9TQ8vVZLt1yf7TQyUQv01SthOQCW9wAuEN
SK8l6NboXahxotA51oko8OqJOTKzynwkEZBqXM4RHZdqj3T7i5yH8ZmNy+Fub9Gi
r3EcqRh56ntNdanafxkgPPQNrYoXD6aIAFXw75DIDdQDE0t3y1d29P7prAQl1FMU
Q65ymrWuOH1d5GE1zkqVE7oLexLHoVQT/hzGHkkxWKUUPNO7vyfPSNt01m+9PMM6
SjJ2MNyN+v8ZkKs5KyWU0ziV9/5PxhRzHhCzg10/TUteJl5d/v50TfhkoNckfLr1
iZqkOfsAwmZ3ZHlaPPVdGMRNn15TnNvtOkQCKtUqzD/33+ImTP7oKIfjwN3ZI0sg
jJMm9uc+VRyaUH4lYUdkxejOXXEHnl3QGPQHJnlNINpUWccH5OFqmlnkNKDn/93d
EEVlDIWF50Niiqo7fFz0GJoXeXsnYynOLk9kQF47cxjmFpHPMALhPwFMaCDL0WeF
/vTDSsQMZfXxae7Cehf7E1BjyYFmrYFOY7jWvGyhrs59jFkCIyMETPj0Ts2JE2Yg
8Z+N9jjj80FbI6MZu688ZLlTRM0dTNhUmIOY1n/JPv5RD9ZyOZyBSO7hjZUUZkQZ
WdDD+bbpd1LIUzgsjePF1BhJDdqfgebwEgAUohAh83PV7lWAHpYiYeg+RxzVIYZ3
uTxQxCM/o8ppihI7iCMXGw8AdHL/qpVzodp/9fuZGvYQqnG/poTrgyUdL+FRaBts
v7/E8lKE60ISkBOUddCFJIrjR9vWTYv9/+tckJnMFyujG0vwgvy8UoQG3hfIwOBz
aOn5OoZnhw/X7nFC1R+TUY0rTNNIoVxXEgydxa6hwwUL/ZxJ8KREpoMWdz54tpBn
j8fW2RxpCaaQXs/ZFFFzFuGFb9AYjGEFuQtAvrCibAPrJGJDOLqny5YcIm7NBltz
ni7/Pbi9OZyY7ntfojiCxuXYq2BXgG/QUVLEDxQoR+tKm/GgGvkHGEbPf7l/uDh1
1rZ0nORlM1IhLcMspEh3YUo5VjBHO7mTCa3gW/iLcbakXxHb7rbL0e7ZHgZtFGkV
3JvAPlkpiCyVmULtItGK4axM5uNehQoiH96OpgmrtYkCDffkMPdBB6xyuNRs/iP4
bNmXUwcd8KuiwsEnYvhqmEuDNVYK8ZXwMDSxtGbTcvMzVZ2uHZ4Bh9RvPXbUgPRc
2K+iKNERSYIR4C8vFVCB9cWoh8w5k6E7SQpZxe4m77jqBtYDkXamYqH5xiC1Hkk0
k8olHlmDnRS79vT5zpH+DIBY5lD4oX7+5frPYchHaUgVNP0so9hrz8DmZoQxcd6j
dh7tXXxrIIyeyKU1CGjkI92a94BQRHa2x0BMxvhY8e0OULzgvBfyP+uO/6/UaxZ1
hER1SmJBTWkJnK+rElD550P7XQEXCZn5PG2BU/3NeYmLoyh36iyNh25sHzonVyOr
f139n+/clLecluz5mPjFuN1ApGzSkAbU7ywZrqUQg4OnuLlq2TamYtwXRHOnXjl4
aJF9S4+pjngf8q5gaqTgXuMYFUgSPfQMJJn1vlD+/7PbL1RhU/R6eg5jHyce970D
ck6/qcUadbEnU/dwR5A7YB9nm1oS54CupFsF8A7ykyjv8SCNBF71UWOkQxlLoHqp
8G0H6TUmgq7rix+7CfTiwn43aYe+dXjK4C84pYysiO4P2Yc47i0LQw+EbTIafnQq
1Lr2WsiwzO8aymouroL4eFuIjap5v6zvYRD4RqLRhYOHJ3erMiaNc3945P83vhwX
jmJNk1dirmiEXnK+BFTl5ABIjAyut5sDzyECS3M8niAbI1Py/W4p6XrYuCQAPaCo
DHhKD2DFmQPYMD/EBidt++DVwYFuZ+F0I0WO+Lls9TSUwRi3BZLBfoUiUfqLYlhQ
Kngx92I4M1da2T2/fGkN8crzbcBuobAUpv3vYZsdXfAqDAs2hY3uID73/fK/bvNV
TukfBKp48rSKa0ZqBw/0VwEbWqwrgCiNaiXsG6OB0i/dEejFf+SgB8sXPaWecrm4
LSYHawrPyoE9Gb3QCz6cG74pBx27VvbuX+OlPBts+YLVqN3NeTPCmmupro4kJeNE
ivZ3ow14/7ewr1SEJ21wYGhmCs3csjvhCM+3nDGgr4jZRbQxQRCnq3Ek8Vy5CPlX
MQ0vM9KBBUBPLvIQo26Ezn70zyX/CJMjLptgvG78gsaqjL1UstGMKiCEtp210Jhj
XnxXwxxsdUdpoM4ckut1jlMbVTVXt6YnH/R6sl9hQx8Ng0ZV6bJCoJMmIp39dYfm
Yr/UoeNyWbH1vJx0kv6H4+8CFzJranC18bEfgDQ4iw2uxD48At+exIc8vOc/0gnh
rSoLtvPQ8Ciw9X9c0BBEpMxpqLv163FXwZHN5Rh3NjaD8rvvNMsvlFmavd9ZawzK
OFcl9jUolKpVaxDkQxU/kXWkQyTtIiMftfmTmxU2P03AFRFMpZvP7X9sR5KpVwvr
TxZIF8eBkhAyybtsSR6dVdHF3bo6gPcRateYurdIf12cWHA5/XiriXJU9uSJb7+e
xpLq64FO+qdyU0oqzb0jkmFzrki6s7KxrUoqtA9WtN4V/5icptJDGfcdUUSA9HOl
NigwfktOOpST/AtpwHvc72CcY8Y5LCPyHpf6bFOvYLKnZGDlfxwmXHS74/Gj+S1x
dvzUV8cQLpFodSytcoW1cQBsol9iSK/43mpX7HumaoG6O9jjGrbiT86tUs4fi6vk
yDk9Bwadh48zvKn7pNmEo7DYhNrRRcaqM4Gz01QE5xllSqmXzMcoBtWnzk3gguMS
X5xV0qad1O8zEFN5b/uDQUjqNWyE28lACAgmU3A44luP2APj2tf5TVIbcikiTXev
BffOOtZF8QsfN8ENJnphGZG8/oLN2IiL2jaoVQzWjbynwFeI235BjA2oLBl6yYz9
+MIBOeIZ4ZbSq5HBTy5aYboXqChUNSkOXIR92FywXw675iaAbWJUW+dRJOLRG9CD
MRd+Nk7fs7tBRZDa0lYs7UwlVQcfENTZX8sZXcat/9rfGhwBSkNQ0Aufz66FnBmH
WdAOTDBoCLhrhOA08IW3fA1+3F6Vr3IS+ZDihTpGXg1rwXUitgv4LOPYNtm7tcF4
CBTwHCk9SaUC/K7BkooUnr6M0Y+JSzENd8/+VxEUWO4glm2INEcLK+ff4bUuP5ti
aHq3nxdO4q6FvTyrD5I4I8peKiK/obZ9gkBnrmqgYXCZp2zK6CyO1qGz13OYVNUx
O/lEsdpp8evh/ZfLX3AAWNl6XQIvddXS0gYYmXyC7qGtjVF2LK15W7MJ38WolzBR
KBsS0tRRLZ6aQoqTsyOOT6vR5mDBKqX7v6k0HzSpBVmdXpN0uE+bfZJT1h/plI6O
oREUM+q5MPgxvNGCl8JVSHVMj3C9Bc1C8bZsQdrashDkH+blD/ZlbfzgsvM+Qlrr
VKWaU2N6vSbRzPi9Tx+yVlVgRxsQ8Eg/j67PLwbI4ibVGu7R1rZkKXaBLbns323j
I0QA4qWi2QoajIG8pmkwZ3V6s4czd/chER2zlcZ3yP+Qo1mDWUVDuwpK1xdalty1
4+x8iS4Wj4E25NlGhJNZ5stcX2YOqUcImEwDHLE0LP34GqXWRYeazgN95Dw2jkoV
5CGP2/ND19SzWf/rbRdyVVPNsfY4YdXkIBmaFW4FKlDrU/aXN0Wq9w/TOUKuVE9f
tszVJxUUMgkctr77qKghh0XGR3fYf2/rtTyp2nvlVgO98JpGoExMeeUPF2JWLp+4
Xsp49sH2bx5fA8djiwxmD1ofO9/hUfDoO8ef19yV8iB912/CvmX4Y4/rI/PhB7ak
6W60bmx3MabPMnjtcZa2yUwmAxF73vEo7xmMWsK+iSX0XV/hbh2E0UxsuyYu+zi0
kxOLxJSOcVGRrOZMaOrea+Zh1ceWNvQmn8jndLO1PnUBtTcaCYTN0Zp3jBPPWXGX
QqeNhuPN/Pw32ejU/AXfbRux/otgBjUEusfcQWH5C2Obier6hqI/XJIeBFxjdGVR
qFFg49PNe//xT6xY0zfDR+lOOlq+Qly/c6+cMXoKhiW5s+Cg9WolE3/JcFR+4UsB
4BQfdFHgTqMEmQUkw99Xsww9QvnC5beyU9qRzzOBBIVvv6AW93N/tOfys1ihl11T
nryicunSPLMPfm1s6AqNKA807eRMO5ixEYcpVlX57BFOxyW76zO0qMhcpYuhhqsP
RxLEiOjowyBJDnaGmbGn5Z1QGjGrqFB5DkBfBlIJWD7zQ/2KTarPl5Aff1bImDMY
rQ+V2bzunabM7PPqT6d/esJ8u1Zr5K7Kf9+kAsalIWGroP3u2jAKCZ1A0oj1CYkf
kCtqkiACFv2NBKcKHF9I8JzysGf3dnFkhWJXYXiKG4ylRRId7tWoSvk2vKwPPHvt
spv3aDCRn9LQN2xBfPOz73PxcbonkgeiLh6C9XQAzhOLiypLHdwNICLeicO366gm
kDJlqZNULzrNICRscRTjDA+PHvS9LG0iBDfcfeVbIr6AIfQE4qcitaztIBZtHbA3
9IqhoOPySaZa2h4deW1OCWkYKhq6+IU7NtZCmN4lV/IJA1V48BzKmIzogZ1fN4UH
WeYHkU6hf97ZD8bgxqsESh6ITzd7V9YvE+Cxcf+3xS3gqGwhuDIeTy1hj5ZgMJYX
Q4U+uKr4yuyUnNOZDODJNy8zXUvUiYTfstKUMJ2M43KMJhhvkNJk2QMbwLaQgRPy
5LOlD6dzwPO4fYVj+tZp04BAkkfYl8VtYIKFBS5lQMzQvZNaIatvAFaBAkf3HqVm
e2phs/9fqw4AacawhmS1X82CNi/JaatTMbAOyBqhFVhY/fwXYaaU6uabmrzjrXWq
ty6A2b9kvqKUcYC1Rjw0qXT7hwnJfTpSr8cx1QVkDCN2vdwrhogU8XchdnZ9+lVr
oMcdxLxpK3w3ZxD4IzMAzPdGUqwMYmXuog+k0Q0WEtVp8DBNUwkH404LyIJa2CSl
ooxdfWOVkRPqpfcptjZf7Uuk5gDEpIzRHOAzuukmVhpYYgH8qJKC9PvqWGxEYcI4
eHCEDWU0OYZ4PPtgyetPHzoLdFU8AgLLrHD4RVGDPOKdJiSgff3qizD4bcGGdOoM
vUONoIVNA0zlvPBIrpIv7Ax4njBjoIINRqc+8aMVaMJZkBjgTfU3ydbI1mcHQjEp
azG2r6fMVT5gFFvWZ97RNDwIEsPM5/V8PTAAADhcT5FNm5B+FA3DQHJrfLZuctKv
rJlNi00VrJCqfoU/x8e4Qv54FLok6qiveuLDKX05tU+ZEp3yS09BuvQn50iSM/RF
PyCWKiryyJNb2o5nU/oqI9tQweqlcCP4IJVCFar5NA6IBmnPts75jjfF0BrFQMX7
GO81LCbh1rImSacle7f4SeZHekNB4Mav38ihO2PsYJtrJJ961oExrI5Y1dVswZUy
9xPcps68p8AEZxccHZkvueF/tqmVVDszmplwtR8V45l+e/g1ZpVIQc55FHA1JELg
sO7UasEVzOxQ/Smpffgfuov3THEV7uEi+LlC9lrVTlRkmdwN8aSH41d9HhMGbiCt
jDidN4Fx2lgSnKBTkMZPI94MkS1UfpNGNzzCA3HSCOg8SqGAspT1sSOIiJ9n6NU3
c9cJeDXw5WhGJ0/Zi9/EM05IVSsNi88fxUEbOqkEemkR7nBzkIXquQ3XtsqigRJW
+0jdSCobQOneioghc3F+4Hi1WhB0UtAlMfkQTsg49uhxpRzJFjCYOgK1WqnZwTYY
TOMZznDTd5o5LE/65Hw8xA1gaPAawvxBa7rtPgo8fhqOKbU4ugvQrtuc2ap7dfZ1
j5L9X1VYugtkEEW20Y3voxcXX57aaiDVe/HivJtMI6Fm2z5Uzi6tl/q9n6LjcM2J
G0eTT/knTqWsLM0mrYXlRFVfmxyc7rzP+9pMHb55lnG+mlAw2HMeXplKFFYpIYXM
1kZMty3u7wL34Lvro+JpTKW8GCU6eII+QBbqXSePNwRoIxUBYWLQdftQDjcsEGur
HFp1ttk1FqvrkHlBdrV6HBpajckLhCmZrSMVqs+knpKYFURnby1iICsqDQ4ajuAw
QAPGxDtpfVrmSZTxRa2XMOEcR50JgTVgweNTM6VVZ1WIo25hLwEC0EV3j4Iz5oVF
7dIPLzM8GjLUGcLbevchH6XcRRfgVB1V4z3nIHX8wFFD4fQudW/pxMJUocG6wk4R
giGwE9+6oPeRWmPzB6wSTdlAnUMioB1YUr08jtOPiOEBUh/AhyCW/5+6tMCIEU4a
dzygu3F9Js0SlbjUBUbzaXNQ8LrB+6pOLBC+aEpMlQNekGC+1DXOUzaxn6OchgH9
ZWAmKe/c8Q+wU1d13WmZtFIu0qD8guX5xlDLMovMDxddU8Z6Dop3yqQkGeviGiLu
e4ecPIxA7u/qzEx2ZzdYywhzHX8y4cuMiPlkKj+AeZduJZ6OjQCyNGXqbN84Wcrj
9Rs9I8EQt5p9QDT3FHLCr4VdWBeA98a7l0BknhF1D7/hDqLfxPWqBY7rcWpwGoqO
X3yPNq/dRScBBAZCM2tdg1KAdbbDBnY6p1Llwv5052xxI2driydkvYn1HDycX47F
Ves+p/3+syeZBymgakx6YsTxX3tD7RSZrjWqYqx7+fYmk16dIoTtQNkO9zd/svc9
sAYzApJGS+aEALELG1G9pNhZCkJVCXUX1xzusx/cdKH6TdCrF9pYjwzu4jqVX3mf
D314H6XOGaEAjwpod99DCMd6Y6Jjbuh0UP9GwXmBlBrbxkEQcQz9eXPA/fIjycuw
C/MOxunRFi6dsjZtHBh/TVblvFRpop1r0lNhF2clBZomraBFSNxI7OTso+1n+fMY
cB6z9Nkw+G2mosbT03ftwScQQdL6we8dWvAR/wk0b/NX5Xk4XOJoVnnKJZle7Dh1
UIGmMxICEDiltYUNCPDxAK9uzvTUU7te1pBhZnSQHIWmBgKPhCfOnQ9syp6d5Lor
/Ol8Inoz7LwLkazys4+k93FcYniwBomgCmzZ30ScOkUYxA19CiCYP4GRAz6a+dvr
JA34TWMPdBgIS9hqLMqAp5eR7VQO2cjUn3nWrNergM6W1l5j8JJroi9bx3iqEEf1
Cuo1qHJY1/qPh1csX9vQDLpjSs9I0dZV8+lkllnhK/zILCy2Wv64aSq6LRCNMZKi
+STGDUkhO3XylD0X6DmbpSIxk88omtYg0WcSw6WyZrRdGMk+Mmh9yYFgcU58BZfH
9PaMBN1WBi10rqGNaMHdHVN2C+UB6f9T2ZMdIbB6OwQV0+vkr1uh8IkHB9fe6n9A
ZANgBmEWTZczKiN93Iai1Ms0wFYW27Nn2m1Nnkrnv5G9QiP2GklS3fJEz+xVAzn2
3fPSPT8cTUni5t8V4NkdwuakDGUPz68REwDiZOK61fk5bpTELh5l8wL8nCOhVwZB
RrrNFOhd/Bd7ovBpG2jOF0c1+jW+RZUCcQvj8LhbIJNMc8xNJgkfJplALkjo+qUq
6VeR0iDRLOY65decHdiAUyE7UdeR8yvm1LAB6oay0zuWUp/HRe3ObfIjJzjdXbxA
H62xx2BrIg9BeSiP5s5XOEZZSvxK1pIU2kjhDD73AJRwtyqB3mZy0VqNiMf8JcAk
iHnbIWn1KdV/nrp+2IoS4KPkd4OEVv8Mbs7eMssXn256D91S1vlOvWMHUs1UXjEg
cTiujEsGqaoeVZOlO2HYgVsLzrrn6ZXRn0Ra3ZrbbsoGUKzMsk0kLK5+3xs/VlMU
/WUjt9UOtto9AO18+2Q3ev38z7CPDj+ZkPeadhQaw6U=
//pragma protect end_data_block
//pragma protect digest_block
2MTfRIJ1SLFFYaCYfoZDyGHpydc=
//pragma protect end_digest_block
//pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
VuCHxWNg+Rs8SXj6Gw1FMxVggBQ7vNmKoWUPOuDfzfsHZYdOYHZM/LFgz8x0rXzq
rJas0vFmg1QK9hi1e1cZ3BGQHQoIobLHB3WaOXJk6chrnpZOm4s3fcBAExZvbWrc
UiauSHkpEPYMWAKheOW9wJCIa/Yh3mYnMyNrfILQRMcc3voNy0muww8HMoiBlVVq
9kzGxgsAoOXSPTqo4evCl4Zp/TjvIoTQ+bGGRXqSuMPtTEsbjlEOPB7MwGIjdgDD
tB7coo1LqV86wQcPIGg/rWnaF9Ay6D3QLAMKNYbHh6/diyrW8f6Gtn9uESDFO4EU
JonbeR6gPgDeFik7DPFUUw==
//pragma protect end_key_block
//pragma protect digest_block
V8bzGN+sZHqLTG87Mhv7NWeuzgI=
//pragma protect end_digest_block
//pragma protect data_block
4x/mPKYN1Qt+Tm4MasEPR9GLrOIM7vu4RGfG3243/SWN+mlmL4CmItV/UZfjTvgj
lHZMO9gFm2gk0Tq7yzbyDqPMrPBWvPEvpuQxkVb0KGVnAochD2NpistfrCyQQbtE
cfdNIiAsFV5S9PkTkUZarIoWCBW2brCuHAEyMT99AgRJxRAvUhtj/bnvuKziKrbR
cECH2c1cJZUrYbC3KNYJAWiyXu+JQ9GutxfRLjwpdbFcg9VIyHMwy32CmwUh1KEn
CdKL8EuPBQ4uSG/vEZTBUi51IocQaNzu8F5lAes73Yu4dgu2SYENGbPRKpBz1+7Z
lmBWDK8agozAQu/tkf3YhS3YlI9AaNv6RBZYlaZ8VBrfSW9UyHwEIrhxbm+y2wOR
wRw3CCAeirf1/jnUu2dJ1DmQRGkeL9Z1TuQK1DnWyEmsGEkxusp2dv6xjTMNjlSR
wL80YwM/rb7LMok4Vlrr9+JQxb4jGraWZxvrM3ljucl/gIPTD/vAUFycigTVP4mE
JaqrnLzgyA5d1oTu+wOf3ZFYcbA0JCJi8EDJxnF31uzHEYmvD45G/4KbGnGlLk92
RWgaHRmLYDJj1x/Yl9yx976+eZtpR+GNsHM5vhgXX6ijNhQskwRwDQNibINJZzOi
scJmi+J7sCutXA7dDUPDT4novZb3nNqbEpK9LvJBVGnjYZIRuet+6SqhBwa2q4OB
nwcJlxVj6JurrOM5+KmqhXD4RTXfpLwNi8EWq/ixJB/RoQy0zxBGgW4tD+Glnvo1
7scNR6IuBcAgOUyruD7jn4i06L27fWARQEg3XEpiuNPru2l3bXyYfuxCuqtrnkpI
IImrV2r1dn/gOqulG4tFQTtAxvSzyfv87KOoeTp/IHRdVkzLr4Tvbk9JxEuBkEML
JH7pik10Ib8GYmeBrEnAm2xzaq+N7fVjdYKukXbzNjwxkjvWrudGwRvgKKX+moVu
RXFe8HvF7w5tyaoEkUF/pmkwtr92NCDAUBHNLiFWiezXxZE2+iLhhMmXpfj8ysDR
ZisYDaNr1TErL4ffK255mZn2e1JwawIJay7WrKhQevU9YpBHepR+ZLbgyLtZapUc
5aP48RchbmB7XMy+0QH3AfCSo8OjtqWUWeSi13JQSYaUXhJvoYJ2ivE0HCyQf0je
zcKzGOFZeT68yRB/SRkF0TRyTCpX8/x/eSvPg1Fdqf88KNY4UxmcpUOvbVFf9Z1H
AxoJxcbjj6KEO1l+y1VlKkyuESgq9NbWbYHsUuTgRxLL15/RzaPWkPeQ2ERD9+Vw
iaTL3PYs/rLRBHV2eMo7ybtWV7PFl5bN3PXxwa33vO8Rol+IwFPT1awv03KuKHeZ
qL0EUAZSkw8ABpHNlVqLu2b8c3TMCTNwnBA1uGf7TfIemYOIiul7rry2kjaa57n9
fJY684nMGDSaF8RhzQg87Y3COSzA8cTMh9p5Q8ZUOfVRb9w0gRTzOJRACGv/9A6n
erA49vksnMMX6yo+MSgxjWred1JG3pHwIFQAsaRWUYgWeO2HKsAGtqn8iQpWuIWD
BaJ0vPdpwbvVq0G7gCtKypBXA0liOxo7qVSydme14tvai2JVIDY2Jl1RU6lXne+D
/Zpox4kIgN2CJ5zLXSZBsKK+Id/kCslKVViCXbq7BaEKVp4+FaH83ZXj/p0IFo34
QoWbgnKGTRaxOKoE7sJ/xbbTBmOtys5UvORUqU88vENUrr53urJU1Gauci5s89bG
8Imq6XSV2ma2vkbi0GjzE8vlsUuPe99OhfSCvscQhnWUJBD4lzNpgd4a6wi63wBI
GvDXRYHj9xOpu2wuzODnUe00saqvdBA3tn1dUvXLStps4dFhoau5SgDel+55JbFS
8N1OU7gqWEweLwl61ZwOzaos741qLtXKbrSVZpNdZLrzTPs7FH6tqo/b1obahgZv
IHu4PEJ59dw93JP2CYSLhGAQ5YhvLEWPfzHWHDkZRAVcLN714pQt3M7YogNqoYDB
pduxMYm7k8AJ8KRXf8+C8JWxHm5MRTDgL7gNWChKUM7NMAWtMXKcRBrJhVWbbNm1
w9pMdQNDAJv/EmRxFr4FN4UbcD0llmJZ1wBk8ikIevQb2LDM920/vOGoXYNdNsgV
sK7ow6VRiqq636Fyb6wA7UEaRWy35UCK/+KEqc2kcuNc3MZaZHTAQVFNCEiIHyAy
WcpDDvjKbswurCm5/Jnvzgq3CpEFOjnZNoJxyn8PvBg2zcmLS4br5cYDLn3nyD5j
C/c5Np+AQy8xRKHjXpR8Dl5lki3UHYo/SEAjZLnNG2gjKNl9OyYZ8k5RzkZxa3wr
SuSiG52dG0dEgftcr86vT9DSKhoOx8TKJyVpiF94S6l4B3oxbW/MT/X7NWpcYKOB
8vWpS1s7CcLfsYuX5D84LMNL57jlHyLxT2xcTxYnyDOkDc7/Wd52y7QlhBcAs2/J
dz6APmG8Fdq4ABOiSjitSZ4bhwgrHZ1KxGj+0wyyqMwGQOAsi5kc5e0I1mPtab7J
NbFi+EJJnpGouanPRtRHTDv3RLSGd/WUun+V0W758DzjuAuInPdXaxsEVk9tdpUe
46WqsHP8r7+WOQ/iPK5vmXgSFdiRJA6QFQCfY3RKt1nAmFzJT2YbhJhdPlZI1r1m
0GmWQrqwxb78O07nIAdhciij/V2fIfhZ5C9e1uSEcliRHx+tpmVa5TXjQlusn+dq
9+uMnJtGNOGmL/LcgBjHB2WuIhb0nOE2Ky1puTpxA8CaYvHhgxlxmUv69VqoaxSb
KgbdUsEp9ShvakO45pX7NhhazqT4jamTA9HgLIwLFZq0sbbtVk0EjA6T2HvinXNq
WYaVlDdSSM7JlOi9Zmwk7PJhVt3cjLACzm21VFC9JG+2A/PUOtQP+q4PEqxfx7nA
sSzx92LPA3QpLkZcsY8FeZ2ESzL+9ZZFslVH/W6AaS6+XOfbnxkEPVoXCodN86IN
MTeXwm/JhO8a1Y/jm0MKHmj7g/iRkIp0IpdHsCs6peO4xwg2F9sVJA1nYsUjMYWq
xU5J0WtVMV7v05Oe/UOymGzYvsHEh9YKni0v9fIYYwaRr++kapxTtGuE71pkKKOn
/9cQ6obO7a5gys0HFtyPW8nst3HjbE3S8qESgtILwLW8C408FtRqV16tp/+DeLME
EHoD3ntpHiMBKsvH1SYFuRYe1jPjGNUcgUeINLGnmgk9idwbzMG9HnB/gTQZ9lLO
opvJGtri9oIVXZFu26SIuRvwRs33fqiOAB91yc1qrvLpgXiZ7gin5fFTI/PAHws5
ekBZuNa4b9stLNnACSMaZNbHOQW7APSYS1uU/55nL1ysPVAti2eph9iomi3SlotK
z8PMzF/d40iXa2ErpJ9/neBsvbIL8ESwgC7MYcuQTtausFZV4dL61uDM+wT+Ovre
MdQFMFvMtXT8syYPXN+wAzphIoFNj9gb6fFnkvp902GHe7vOF0CAsnyGSqd6q3Gz
gVy1WJcmTbsaogfmne5WobiMobk3LrrcWOEM3ruEUFoOgSXyZ1iiNoRAEjf2lJIM
Zl62FC13Jt8FW2mBZNd4mWKQ1o5YVf7jRvGSNs3cbgb9WBLacX/NeA51TKs1FE6p
IXjhHumfys9b3VzE6k8P8F/rVmwnrlwLhUG9XD17l/PVJ9rJNfU1600E7lFz/W9N
8NleNUtCdYG1Hh+DBFYP/x3Ff/MgRVpQYDkAZRCFFBHlxz8Rv75+cl2Vm4c9A3h8
y9aE/eKIu43J+IgqNa8m/j+22bEaR4k3WnmXmp67lWtUXgVbtJWNM5Va+BIMb4Tz
iNQElUfEqAR7u3gjUYgApMRHngCMX/xCa57DGuTJqPON3apXKLHL1UfpA5Jt0x1e
wYYTN/sYccE4PK1lEIz4NaZBIX21sHev7n7Rw6Db8vKM+raB3FwqCopU7QojiMVr
mc8/7iABWjzPgNSTP7YpKoBlzO70LFNzGulQO/HmbO8voEkLtua41/2WwIifB+8m
uXadY7xbJCayFiVZsZHHKBe5m6vYXDMY2ZAjOSCFTbbBN9NqRP3UHv2/vA2ftZxo
/WBXNY6l8xO1mCd+TWzuADkJ8VSm/Wqv+k0YvSMgeDUBHus2o/F+bXAeoVJOj1tu
GdUixFXerU5djPJa4uDJYB3C2QUqrj0jbzt15MZEmc2eeNsiRQp+m2ckt8Dx5I9R
KiwBTXFjYkUBRWOL6RjrOePxJJzCRwohCTxJpJjINLS881JpRqufg1P9BpeFFJs1
JBg6UaD0CR0omHZvnAYaSSd0D/jNe65gMsq1z3o7xuDHp6DrYyaBQ3kO1vMpBzV8
kM/ZHPE21ptzRja44VqouTI6te10e4HmTj88J9Ij/Cd5k9bClaiYF4SO+k5iozdC
t6jrxA9XxAwUHVwb6k4XkATfNmylTdSBstdoXcpDC/Ae5APqmfjzpLtTZfk3JZiu
nDCHfT3DDbJrkXqUp6Iu2A6x0Wvbw3hL0obduRVaaoWNlkA8kHrpH14Ckt/l/d2v
MwaSnLzTl5CjiJZDsQmLuuBvVf7zF+8Ab7Kjd6btu1EWwAABqVGJt+eqopKSJtF1
Bweo/uVZPdbk8GmpUIh+RqNvzULo64OPat3FXARPRG9JUv8M/8Y48yzr4zAbXpjB
T6Ps0APoex2a5RIB+C3jUMugztKbvRd8TAQE/MJWrG8+gvDENq9Pw47k0PacXyVC
KZxgPtBDI61AR+mv9b3QzV/7Tr5y0mNM9QtbdXe/DxQO0KuwvqoYFOwHKDOW20Bb
YWiS+c0aImE1+rMKKYKFkv6VbGZYgdy3XemDRsuFD//xD45lm2XkUglLGnPeMA/Q
Kvb4tHz2Ofli2RHH1eTtKtaOrEeM6EewpicNrtgkMY9OLplPMdC5SWNDKKhVtzDi
TyLMZ6Kzdmkb1V4je2K+gef3SAzS/Qbj+1Gxqp4O+RGDN2oIBRaEAI4YZ/J6/XBJ
n33l7o/8P0yqGF/mUXYCX2m5seD1rFvfiapdz6xzlbd1T67OcY4ADvrKc3qazxyn
FqMznXUiMtbHpsMGCKYf0mWFAKGZZQdtvF5HaJ0sQ1V2Z6kkHJXyZUf5YjWBMiAX
5vsCDlRAgdEFm29aTi6AUoWhP2FCCa9lI3/24ZXLiH4Gkh5R8e3mEXmqyAUYpXlQ
ypknCBvbktE14K5+EnFBC5mkidMAbaiNZCAPot5ifhg/MZzSCgASnub4BwWgJXFr
fcD//so9Nn6k+iK6kBywLOla1Wqog2RLxPXKhnFzh8F2OGaCDhsxXQIi9TCuCG/W
7x3GHeBAo/zabea1vJJn/wU6o8IUxDUcmwSqK9y7GT6bt3uE4LzdSYPE+m3vYlJ8
JYGEazfdpo9wkNG1WI5bes6p8Y8nNcHZ5Z6t1ZEBhzpTHV0m6yPnXjGbBayPquhz
JVJUJSGsrMglV1sepBsPtwEVDuK/Tt43iCGkRjtZXsRbQo7lumIsDewOMxJV5jWH
pv7QYYF6KNg0clNgCWmzxRVnkAFcKtJjEYImlypBruq4IKACeYK5I6aYeVobVaiM
5PHdBFbU4bTYJtdQ83Uw1ppbG8Z7o4aPX0q6aWH0NOIonF+FSxq7d7IkGixVm3lG
agOpR/BQQSirdPzX+r+loXuQWFrcuTan6cLNB9gWXpw6GSzr198XyMJ2ahCyfD4G
PGoBHS+HXc39UquJzG7LIwJZBdUulM4IKPYn653Mwe3mc66olxqR+UZV4fXwlnzQ
RiLlTD6lm3DacEoTuR8XRpKvNTORm47UFvroH5CB8DT35O5zOkuJqLCbkz34Aied
Bk+zVAJRneeM4ZfR0/ttJ5dQy4xdnnLeFf4rBamUSmI5DHY2yWQJA4wiLOqs5Rth
rvA8gu46/vYcC1/rICyTn6Dyi3+i39OuXFkrrkt2k2nH+YY+jDIwhhhkogRQmZJX
geUCikiHYgRvdmgvr6BO677vcAJzSICOpsHzAIbqjW3z4Lnj48FXzjBlsKWIrAAl
StXqdTV2E64HtZj8tV3B567cekL/2RnLcHchfKi5s5Ijb61Y7fiBzRRUbcD7m5NP
2qKuvLm+yRUJJC/Mfuo9DdIvS6fesBrUoYMqbSyiijhX20ef3vW7YvwfRrt2Uys1
6nDp1ZNN2n1TqPush6hmpzRwJNRcqmz+o/saEubcpgkhWG41D5NZowyRMxFeXhGf
yXSWb+EB9aHYHPZjxlPzBaF4dUuUhZRfSIUVf5KGKK3aCXrfQ25FWOgPzNsxzcJF
8KQiq0GRUMokJrcyNhbUKEUQkvObYjA33+YLJNflS87uvJiCkkD+TS0BrmJeX8Im
RCOl00bP6/Y8JyMzhgZ7kkTX83460bKpNWlnnVYZGEdPsaR0piCbnMLx71Iro9VE
h0oJ1/G2oZsmYH0Psl7TAakjNdRoLK8Adfm4/x0ET78NQ8t5QgtWXiw9IdLPBUH0
nAtHbRPmvefEgWKVF7C4cqgim36nTjshY/r94vROLrT+t5KO4APnD9kLQK+XKZBh
6Hj7TH07KebeC9CF9A82BjcDdnWIEty8GOOdYgsxLGFxcAYoF8VFuvRpqBI9bp+f
BRUak59T7TYIhaN0PkXUhxItRldFcztSSrgOOEV+UfTSw4kCTFKcKuoBAdJSTVe8
t91Yd0Mca2YFf5F9II+frZRt8tpv/KNz2l/kg7XvnlaTrk8jOdoqGWdYoxVuLMjA
4oplEMKSmgeMySZ9KriUxsPvGJcIJlZWERhIVTMyacQaBC1RciOUqnkId/LaBaw0
Ufe/2wEtAW0hmrMvBkokcUmKxoD6IvAXEruGH0YAz8spkNsZSpepUYYK3yij85xW
gASXzNR11+ebEUI8NfrmDqLHf4AwOb5JzoN4n2BMPTekTzpv0MTeEacSmvbcZYaT
MxbSpAM9+4c9C5JQ/OlUYUTOgIPp4TI07/tkhuwKgxn+xtf6zI00ORWhB0XBCIbf
C/6Z6tJYU/mFY6LxXLhUD9UPcdrLE8ZieaHrf6AcNh4fNvJPZ1uf89U0WWPDYvdB
EkWTg2VgvN1wZx6b+zu+THRD8e9yErWUkloIXghDrXnGQ/K5+s+R7zyxwNhX84+7
g3jp7omdKkvInSHX4C1baLD34s/lm1N5b9gmxooV2H4uDb9LedkbDZVUeV3Auv53
mHeTMKhZctYeQhwK/vb7kcUac0J2xk5BKRt/jZpVkFydmFeU3jAUNg3giVdWg4fq
Nsz9HShbWHt58C4yxoAZLDo9n4qZ2jZixDDxgI1JXsuaVulqHUUAmkieLA7VeISq
dRHPaJy1nZ6sGR+pIm7ukwOlpsv7gCnYRusXPa1aBKIfORT33qffo6LOQndouIN4
DOkoZ9l1/XOmYsmDgY53hsCHAgZz6dQuWe7cWJn8TIWxegj3ZGdrflD9DjEKhxwp
3kXQvAPcVoZ7dJGWTCuxMVFAaiB0vKDg3li8TMbWOVdSzaHmGnqJCwwYHjrPYr1D
sUxFbwbhqiIiG3BQ0fQQjS6TZ1F0d2IJ9LdAptB7aOLtn8IZMp5EZ+k2KiCvR9ua
Cb09PM6f+o30aq7BqLFdOe3S3wSFIYFEFKGa8BkcOtoGieE1gMRE3bP3Iud/41Ls
4LYOvG4J6hYstfBjyEiAQxBOmWs6fguUAPwkq7JTC9ZMIRNldbPtmu2E1DQyTx4z
OwlI4p/fll0JhcmzQg2igvEpcnUTqxT9KdkfyIDw5MmAtTe/CKAkCK6v7E5ptMd5
vI8LSnGTuurAbUfx0bf+znKUi0rV/18QYKf+nSpykRV/fOErtmZTRrvooynphb7Q
bclqVlVCB/GfPxGlT7r+XRw0Xc8N94fCMBGY9UWl4Yw3xqdp9nWCBnd+KLYPUDWo
3EW8gkqT1m4EfrZ1nI5H+MN659eRRs8LGgrxxcRqPgFYGTLTYgn43CQNGLwIkkqV
PU87coYneV7w5XypJdtu4F3tcsB1q4/iRQn8iVsY85VuDzlei1/aHEzpIry3w6nO
JGOetCAUqG6VSXgtBwCx53REwSV0EkEy1zhh5604OKEvnPvO1P7bdK+su5nRGam6
uTSbOenwxJLHnLrDE96wg2nJ/raSYP8FXcGq/M+j4xS9KLeJ2XYZnzdA/62cojgF
4sSEwb76kftaKzWjtxb7/W7R9c0dJ8tWE/7RpLXOtezYhp62v3BfiimC5RMYrK7A
6OP8iC1ul30aCfUfWWE2bX+B2kuYXup5WzZWyTNCs+G/HkmznWfUm4J0+yZ188/H
y9tk91u3Y6RG7GJQ+zmxw2vz54IKyyoDx/eMCW7YHCQLw3TqGDFPMEu8dmsqqlDE
NrHPiPjM9Z3KzyzGBSqqWVv+C4NAsZ5DqvmWi8sL3tgqby99iAr9HneBwimfP5E9
OLzu13Pw6jo6fuQlossLUbEiQGggM2lfp6RHYD+nWq4J6GHQaIAJTnHxHWnqWcpu
qIK37EizWR95ROU0kRNVi1Xmgz1qaA6vrbnclU7FYo261va4ypCFi6KYimD07xzB
xssiFYDjPPjBzfBiE7T0F4SofBzsd+uTnhblSQA/7GYMXDYEpuAcfmmY+BEJYNhA
+B5P4SLH/y/CFNQ6wy1o15GanJlVapbtdYJNIiX5gf0=
//pragma protect end_data_block
//pragma protect digest_block
012mvSYPJ7Sdcw1ejMKOnAJYLl0=
//pragma protect end_digest_block
//pragma protect end_protected

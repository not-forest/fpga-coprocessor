// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
OFm45BnHxA3ORBn4xYF2mHf4ToMNtXr0gkvwW4nct3cUvbT3GYfr2RzlmjSDEVxO
hV+2ifbx+ULnf5+dmsgWvKrCx3KJFCXBA7tJGQMxq8swzzlqbQHEC0IAtZqh9w5z
iQkWBENpK1Jga+DVv7z3RYCein5qOzD9qlXL7GyODxk=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 6128 )
`pragma protect data_block
wd/eIFX8oto8foidZvdiRJMYZFPEHASo7TVrdun52qIjTqszkTyfIMKQW5OHN4Sc
ecWDv7A+FOGq67DIhGQpI0gcPWh5w9ovWZ7bO98+NtvcmTO6aE88STOWVyueEtvs
UCQlNL+mfLwUSpJnvvdKb/fqoTm2yqtjHxeuQVGutvgt1L+UuQDJuTfyl8k4kCQq
+iJT7sGBxmcFAC65vhGdIzndNbkT0/BkhQ4BYru4cDNIlGSD45wmagKltD72Rg2+
/ifRIA4AmLWy5Tuiq1IgI+b3HG+6alym7ohUMhCLehKGjG7qsbXahR93GLhud8wz
aGp94eu60lFF8jFk+pzj5yfwze7gvBxTJdl/V41vvIcERRVpouidusiJtkbR4UMl
QCM4LljCqQXmO0Uv8lRqRg8bigbIBCRnmX5Th2gumQOANf2lzK3ZwWF8EC/hpV7I
VSte3y1B0BB2aFLra9Bbyf+oODmH295HJ1hdsj9rtmqV71CrvTIs/EROUIi5Hm8a
WSUnKJuGYHtrNFEWwso+wblRrTdfEdxoz5UzNqxkyEOMViAT2EHMz9amB2AOF5t2
Ldu+lj9jNyqeUO200C6Da7FNnIjtJVRUZP1ndf+HMBTnIaRh1BanJvmnqyidwMY5
fcP1ZcQkEXngSexSohrXqXtxlDyG05QafbXtfCkfV9yAcBWVtZiA10Nd3jups3Wh
H2QQDJIpktFX55jg0O51XRo06qYhM2q2CcGGQZZ3nWvZwGPIjCCOnylNXCAEKC8U
OEnDTDi0iPHjW/wzqSsuNxIBykHJTd9csVbHPrFWjU89c664YyguPDRyosIdGRJ/
wdEjDYqFjjBo0PI3PPMI6vHMij/FFhe/eXGBSE9yEsPBEVQysbQN14S0y14X/JYn
/jRNMlWR2I+FTHWJQ+WKzKRqonIrG09iBkMaPSb7VTsKmAR3VroMV7JPyZyyF7sx
CMu/AGEoJ2fHP+oLzE4pP97W237ea5ENyXOYYsdmdcvSZuz1eW5+wMEYrVrZN5v0
zxiVX65rwgqvfqY+jxPmZ92GdgN9RBdCKKtHyDvV6D9QnuSGnrPuCiHqiiexcCe/
spnR9eVNLVHrM1VIWf2ndQ1B9GvQv2EtASr6jQotgVU8y5/R5dYp0h0d5x1VAklS
8lfIZ9TQ8tHBLYvCASK6qApbF1uJLuffRjNTBzC3e+1W5HU4Fs3psXzFORG8Zy+C
dLGUKa0ZddIiKhN7eG/6o4CQmxk5zziA+mwE+1pE/jnkg30+oyuK+h6IS15Ju14h
xHyhkqReihYK3uCyn3HAdd/Vr0hc0VoijbqGSxlrIAkwyYY714e8Q5WhxoHz+tX6
nUdi43tmy+PlajoWYZW24siJVcAMskNei5lzb6AP9N4rI+dIrN0eD3mEoPfi65bA
rinURyN7zTFEzGnESaOnoAKcKVlCanW9R/ATLt7gcXx+cXKQSkPzIXDUXtQHkHg0
CmfPzR0ASJ22lDVpHmkRPs0HEakvP0UspwusaohGJtN5X+4KV6ebiTjyWLeD7egm
NsbfTiTezirV/jRZaztXL2UX2RLQmvdSGAtQOKHqzbOqRDbHurk1D/a9BhoId+WI
1MVfy6D+N+OGNFXElKxvHy7C2dOHInaAAva5MGJD9XCDnzbsqqXmuBBBoJ2DR+xD
K2HTkFHR+HX+iKybT13UWsP302gLhSthIYoYLPYKi4SVMagA3ljLvz9JsMw0bs+E
wy92kG7W9iF5MbsL84imX2Dzqko7tuFi9shnY5rCy4+6tG0AUd849AE409uUf4oY
NCsm66e2XuqQ8ziR3XwPKD1t5AJJSbkeWyF7D3JHg4+PuSdfsTK0rqe+VKdwSwo7
FhEotz3BBMWQS1umgvlCFvzLHP4RVK5y4dGKjfWM8j/P3SgO/5n/qxEkHAjjC/HG
hj8DBJk+A5zIsbinqZ7kJ6NMS2gBI7/ZXQEqOQ3TROgqzrIvyoOGzcKqaTY+ylAH
43I8moBdE49f0N1VY0ckAazxErPa1DgTTG++DsRMLxzj6cwRRQpc/FiWQlGmivlB
im/M7MU/tCUFxK6TqShOMXRXu8zdiy8h4B8aCHXaYI+xHRb8KRAzOkBdncSye6gO
kB/G3E6AgjZuysfxB6o/vvAZdhovH6lw2PBRgNK7JMcajjR9aN6ytm957A9iVVBl
G4lusDeCOTQUUx3K1tuPt72dBegVkxYSpSI0zHtW3m3cxNcGFkixqXaJWv9W6lqG
LdQDbc6n0dXgAM77/heEHZvn1E1I9HI0DO8AyguDgT8RuGSM6EZ9glC937rKLgb+
3PGRbcIXutpE61ZeoJ+FnF+sL129aBNwZazjk/gH8VGeyOxb2nFsyTu//fLA1Qxh
//hj0eIB8OCYCQ5X4fmrvZYSWuVr7VbmqKagRfkmD1V4Y2fcqne8F3ixFfByyMkc
BUDCu2ALSFpPWkFQJS3/LPX9Y8ffcGN1Daait1AQlREyieVtmlcLMTK3fthPrx/8
V6NxGeHBhtV5ZLfdVQ2+YAfA2utwMYN92DFl29YKENLI3mcpPNuzIH4jV2Ej7FV/
z6dXXgfTfojtHu0hSJyP+RSNRKA7aAKEtntsqKrL57xtQL6QEixB7H+jnxE7aJXM
rDg5amulTy2vEn+NH2EnW5A3a7kgi9KCCkiOtEubW+WhjM2FaRF69U+0U33u7pew
TH9ErozkmJ1HbjVBtFUEb6lYZ/AT9Fp77/1aFc9xra51O3WgtxXfGF6l/bZrtKeA
ntZ07cZUa+iZxUyCmTjMrmJ4niVDY96ztGiz5zAja/RoiZfid4W50D1yielMk7o3
gI4lUo9nFkcbUMaWMnpQdsLtN8NJAGFoFOXNUrpo0Uk+c1PoSdD7WtlDXOSCZm4x
tucTyYaZh9Wv/Worah2E2JRVQUN89z967sVl/foR4jcnGS5GhRsTKJJPjtHjIzuO
e+KMqGriJtcr5poF20Hc7Pw0aW4BtRHBCQVwnTK6/UnA6/+KLHfMGa+AE1vo25ib
lvytgh+9RiADGC/K2fysxDUT4fBhZIpdS1DufyAEhnaDxtsF1EPxHJiNx86EDya5
wju4/q9D3pkVRU+jmIqfIo0tJmZmaRBylv9iqlZLJPmQdbMfgBaFvnjDZ9qgOVmt
p/fqVybHHaGhtDYZl/RKH7UqMppvwNONzhIco9CVecRfNxXXirMDYYVB2R/SL0TR
9JqxR8/ELsbEeoS9ITur6e7fQrXvDyfhReucrphjoQIgvE9kEPRu5FixVQm/NWay
7MTUTLEzRDGw3kiKT6J7qaiNdSaNXuSgmEkWU2gKh2nysEPEZxU6HbbAJrWRWq5w
91eIGLRzo9FVK1vFmdUBcGjna7DFnVztn/ELibw5aiK2LgTugGz0iHsQ+GmmUNrt
X2aWFHm6XO2pIYPOpnwEJ9kNHnJZtHxHFaTfFRO1MAN8YHhSYqzSP5IzbNPYtkDo
sC/6SXvqSu2qpxfbixVVS3NxVX3YwDPtD7gi8RFwdkIaCnL6EPrXJLvFeNv042ON
kBlvLgA9OWTVT07TtLPnwvfGYa9oH3ROmq9fu8lrOvXW+tlKRuEci0bwAYVKPBgw
kw4nuCP0nQhlx/4wKeG2sYnClPMYXQdEj12DqXeTSNkKX6G1zS5I0AwPqYUrOCL+
tDluB3OTtMtrM5pt+d5kRzAcdShoCgx8vN6AHsMoy+bvQ+9FLMnK2MbGQkKwPxbx
89w2TlLzqUMME+/OgAz2itXUzAmjYKDAd1SjrqoCSwxd7O0zLmOF38VS4C9Fm07q
MmmSBTlm74Qo22V2mc/53HPfP2mhusryFUP+NZQmUtxJS9uKqoR+CUxJv/2Tx6kP
xQHbIOk1segDarJkTZAfNcheDAj8KCW8heXeLYkF6wq3E1VkmBOHjPhhvlj6JfA9
E50kI1no0IGSkKBNYzlYM7JglywOS5B6KZA+hMBPW4fhOvPr0s0lSkWAmKURRmAW
DVKxoBiTZ26bUZP4QeVHlXMgLeGS5JYXGh7RSsXS90vTE685S6XHTUicNorcFV8n
2231pgHffR7zJ5uha1OToBuInvN6HwpKn11d67p2dB4m7BjJwV+VhUvF8p13DOoR
3hYGQ6ssWiEDia8nKBuKdiW37PhDWXObdt6U2J0R0GhLICJJ+8ssx49zW6oRztP3
jhV60sPU3VwWXEKsjAKAjz7QBPeZuJM8d1bRwn6SKpv/b4mOzUEHk5Qnat/OSXsp
omtzA80/hvBfnlL0YyZMjBD3Mr+YiJ8eRwU5zwoxZ0BKRNVf3zlxzGb0LTC4pAvJ
GAcfcJhCJ4uFb1L+eDb3JGmTed40+UH1Ae5XTDRYlKj0j+6rc96ABjHypmaTc6Kw
UNawv94glw0VTAZT5IgLkqkpKCmr2FLkfuH00zakbMGg6Hafmvv5+VRXvFXCaIWY
5HtYgAXhbyzaCk77nbu3Mf+3yqCSKS8CDHTdm9aoXN76QUVEhYtBbb72T2N6kjU7
H1h7/zwquz04Wt/dCLaaQdMxhHXpanhdM6OwlKaPAPPolWe2vaMC/8OCZbIwYQXM
+Efb4c/ghIYQuIAbj574Eg/gUGZ5UphuIpWQz76B+Ib/fxAdIahTN1knB9E2h0uZ
lq1ySUOBknB2xGoMu82Y0NSvoOoGWrz9/aA3DbtCfuC0OXQNdUWUSULoZc4l99GF
2iQfyJGHnV2ZZxDvdhlSbi2w055MQuYeSlhHf6iWzs6H7VYz80yOuRFtWCtCEoRI
DH2Tf0/Kwi30Zbot4pmOjz1lDKJYk8QypcZROIWk68ITMr21CX5e3BMZAbUCR+Cn
C2gokyzTkKSotdyede2tADMOFjTGKNrOqfcoclk636NsRPEOplO/ovUJfy7CxlOg
W2v/d2h9EP7Yd1iRFaTFeEqwzNAaS/6LO5z43aC41NhqXwPrN5eOMkEl8eSy+0GW
DJN67d4msFV7DygpEhaYhd7NtBLbW1YeWP7U4fLtLeY9je82e4gi4g7Gkxs5UNdf
VWdc32UJxsMJk18eUcNQ41Trhsgw6+wW05GzWaeLtwjnHvBqckQE83h0LKaSYgVp
oJbbSysO6BVFWRLXEAczTMGS5IO2xEAUYYNAkp4jEEpzrtTuhy7UHDmkSKSdl3Ks
Yloo5mRdP9/9ZNj7smjoatleVKTn0Ve0UG9Zgx3k1qGo47GiWALR+l3n+43zpmzu
6gA7n5hESCkdIWlV9TSFu+b43qKyXNTD8m2aC7bmhAqv9m5CxvN7CnzsSSVFTsd3
N0pt6McwpT+jvLTcV8vmQqZC7lt+kB7yIVbdy7DrjBanwwTAVa/y+vG0moBOdPJ0
DNsQZNJ1PX4TGcX489iMGRwKSewTRWtbJsmpPX7Kic7gmjrSAEi0ZgRQictwY9FG
HjbmjDX8pv35ZGjdCv+qTP3QlFvDu/NXJnwyuK7zBf43gP1XkR0R+A/Jlwn6M9ua
23022j3NNX6TDw3nl9VI5QXQZlazu/LaIGLEMC8hDEguJvv3yUBJCqONgBrBLyG+
EH2wAcLaHGYu/+23nkdDjaomFm5VfDzMsPY9nvJYgrKjd68FSvEuV8BJ4k1w2OtS
cOzA1QOKBAveL1cKelOqUuTOI/lTvQpUgngqk2+JrWjFfABVgcc04+/SHFjSAtDI
pfr+MF0GZYWxp26szP1t5idas4RrmJsyXYrzqhezYh1xs9fJD2hsSkXf41sfHEF5
a8xMy85DWlOU/UanVeX2SIEthIinl+ZsmLdrWixETecwSh0/+S61GqryWNjwnwlS
j3TBVBwKPz7/xsixOm6auS1jYW8yujP5AGcuNZONI1W2cwKx7KxmRFeM3s6r8zGX
WoS0PX4JkE6ePWwTk0gm1jOXGVKtWZAzmodvoZ89GGjtQUFl8zS8NCy+PHUy3aKf
3Cs+NQZpQBH6xLeIqkxrMQQlI0yDi56Gk6dYEHhrKDtjiP+c33DYE7N/dVGyFL9h
eNrYDiQbYVbgM0YYKq+mGTvaxGWs/7s4TesqgWi95uX2LRQy/erqksBoI8GU80za
TON3gXN2s/txIV13Xkt7bscVdAYChQCRSZGUMvUwVRtcWT/LS8XoF3zFCY7ggovb
T2XbHOPMVIjrZo4W8s9/KYjNEbt92ShgvbW/yg7szjGj+BAIVPuP3LqLtYUT9HxD
La6MhowSFZY1GSfqrS0y+Rs0+IC7rTJDW3ZscfYjIYblaTuw5CvKfveBFD+PgE+j
sJ//xiRRJQputYiWkWaTvpRUxbVPZlcxNmd5CjTqjlfKYk1yZrnsQRDWOtjoSd3b
XyTD1LBDVdQU1uLSz87Mz8mXX+VgkatGmylrCXPS9CMpwLylpbd7UN4umsrwB+05
ZZGxDgz13/nx/PzE3JJwV6FNAvukm69Zoz3OzTsNdFzAvjOMlossZg4H64u1l5oD
y/XCmYrMw0iTnnNNblhygnB8s6GVdooj/S5Lb0NqVwFHL4kFEiiAjYmAjFBAwZ+g
kjUKBE+Da/slIKHZz7bmo6pc+Ixggijl3b77S19k6O0fz11Y7L10ZuLMaJFwK3j2
gQkcTYerUe2TKntbHvTABahd+9cwDtugrEjFZiiCXQ1+8R+H8Uv+zhNhRkEYbNG6
/wTndyV2bax7KOpTxu28NodyOCZ3VLX3/Dj2vScT3TZmIiAi47K57trRSBQLNfSF
Ef9kcHsu7azwgXdmZeacvcGHH5CwJtgU5YDYuTMP4LxbDOj0E7vPq3OOmjh/cNJ1
5+xGns+X6uNWGoS3KnzUuImKdhpoCeNHoy1XFK0v0+EidyP/AVCeaiXcbo5Lx1qD
zYyCsurf87IvRBhUGC+LOsQjR3yPTkqji+Muykr6nf/bDvMzgDVMqIMWhHsO1nqJ
NxpyJP+0c7IFT6ZkleMfhPTKq9g8jV0Q74t6DijIxlSFp1Tuzw7uZ6/JsmmH4yFG
lAmm62Sctz6Skg+dndzkoeMwnqMFQ64qNXc1pr/838ZCjFcijSzgUiGYij/nd1tF
J/zvKaiwI/MC4xb0j28GxQssMx8R9jc0VGNgQiIFq15b3NYO/OK9GFk4bgTVpyKP
uAwE/9s/ROYv/VgMhEYswdHgD8wj0ZCE1z4yaxriztbJHAUVEcvOssitvKrVUxwH
6wUq57n2ChhKeSun//1idEd3HtERpBRR4fNQj2LVjomSOcUIHt+Z8uTyXxny1e3u
LOVo3qJjakHaSvrApgl9QVmNfU0l0Yf1g3ntXmAo7cxMFKNpYW+zRDfGrdGkldv+
itLT5C1DQtnaaAGH0m/D5UmoCheFAfWRr4V1wmKo72pIPZV8EO3Zmpy0QcZp510i
Z+pAQZ1zCH6jOjia0SLj/6ekN5Tn5fscV0B0vVzvH88J2LW4MzvTbvAhlO7CLfKd
lkt/oEoObcym79dZHdfpiJ6DQmV4vyYzD5F5BZ/hzvTUAfvJSm0O3a32JjG3sWj6
nYbbxhXBEEgW2xxZSr0y8sWgzsDVy3QJCtY9naw8/kit2p3H9xGC12H07Y7xJcLD
3OxbXOIrtuquVwZ+QPa16nkHRYbUw8e5bgO8K+2UEuIXmT/xw4LKlnx2Qdtq0PwS
3DCCZIvlkcplf6uQ7rEBBPhMrWaEZ04FVIhtgqrIfTMipq9U4g7n7JLMVEfThSnO
x3RtFhWH1kgzGAspXw4FhWCchQn3MFszkhO8Wnsylrwcz0QjJo/S0vEOd+w9VwbN
GCLevQpCF8QydbIScBhaOajXZQlxGm4/rwblJs3E7m1XfNNRR0vkosZjUAnbtz0H
jr+IIZjWeWJBbGlYIbU9pSNzDkZOj4W85d5qS81Qlm6n2WveSveFd2MRAXZ86wZB
02NwO+MFKtaDEjDcF3CBOfpFrIrR9UlVpomHo9nxfKmFau/4fRswvx75YxSQj+bY
bwdX17qjbrJW3W2FUH6gzbSfVQnMZmDBMk0Da5f2guIAg+/ovzauVOkhryd5Hjhi
TShUH/PcQYQVggCWj7FZyRa6C/B2II5MAzjzfPm2umFjnspLNgTGgT11em+Yga/w
cn0h1BIrTQXazlW6ml5HmTVE86SPUxwF7A8hlxpn/E+MuW1+hwvfkWc53MCmRDrK
ftWqpqBE9XYYegSC9TNKYO+S9m62l+CHldQc2jRxctpO/AhOPX05r9DLkse2jU0U
e9fXe1FQPcqMMSHjzeWyovK4VVs+hi/NhfztyfMtpac=

`pragma protect end_protected

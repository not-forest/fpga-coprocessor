// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
X8cKQbxb3ujgEczWKHX3Vxer0DLhbpANQPIgYHnOIvME68vLFytft9NEsNuizhts
DMnfXKYDpOWHiWH5+vC2Gy3Lk+OKah+n3WVudNWkRJs2ZKkeb++JY+sORHHiJBBx
Wa7f3HTojGmgG3xDbtFvpwwXH7WuQVQfN72XPG3qUKY=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 12048 )
`pragma protect data_block
kutbFnm6o5lhvCDOskB+OQhBI9zkadywYIf4sx6pIoZKP0/D708BslHJ1tE0iFcG
SG1txQzcz9pD+jhaW7Lr0Cik/qdNL+UPunzkWdS8anXnd84XNCi9qM0yYVzYktZ9
t7IORpBANC1nXSMfC2mH8hOkiSNXtNk0EX1tLGHRwYB1bxcghKPBwUOHpzxVFnay
CCM3YRC0PSv6Hv7bJG7Yvr2YJS/VhbKVkUUBgIUhwgQp5WgrmDG1krnhLqrslXA/
ypqqY3/slpUZfEVMzWe5leaxn8K/xXl7HKUfTBn0nqzoMTLitn4xhm7JWbdz5oVB
ZZiK5s+sCLcgaYcHdfnk0oWJraZKafk9blmAdJazIgJ7UtpP94fawlepsANm3pfS
7vCWyEVWYHGrLC1cXz38PIBL5mdBv7nxrblsZjfv9JKV5g1irk4/kn4thQDBjTTy
OpLrm6X6DMxeb89KrmwHqlYeF5R8yIddNHN1xeCc2esuDHcSUvPtI2wJp1PUAWC/
q9EAI2F5j5kMXi1EGG0K3yy6PDrnJ3qImzA+kPCY8C/CBHN0LlBSKmvZl1KUgKZx
uLBtJ9Qf4rE11KGb56FMbR8/IrLRezg2EfSTEOtwyxw0p65o6TPjnpBGrUKKhXMq
qtokTy+sZ8VHlZLc1awHxolRBizbhH2ZjY6Eli2NxNEfUB23IUvfrDXH9Orqft9P
ZgJOg7OTQsUSzT5H02pwlvzknNXQ6+SL0fxguXuHIlbplA0nuVZyR/b4YhqDftrD
MmQ8kGaWh0/YF7S/K+/Kvy1RByILIiM/1BWptsbjkSjrQawZj2gHBm2ePOA6wblu
C/XrQbNmrkir4beh2ybTmTFj0bj9ZE/P7GWZUIveN3QfyMYTj6B6CVBNKPkbf/vZ
/Dj5ntZLsoxekDXGfsVGCsF7ikBbS8KsDMzklrAO3YJnFtYleqWEMaB3nb8swvBE
LmR8DCgSUFUNskvitJNU7bNgby9dT+6BnZJUSIGnOm1hGpRB17cKXaeIvLPAJY13
c2IExcVtYUM8JTlmYFm3bwN/b/Hj1YDK+721YoAkH6Y9ITIpNkMQQfaOniaAGMk8
VUj1Oy0XTGIFMKtzOF99iEz8ERO0aZ+72kYicvhm08EnPhJNAKdUHkLv8vPMOT4E
8B4fkxCuW+S/5glnn1BjYPpYyygVk0lhCilPOJblDngslJp7WlypKw45XvYEp44R
+PjGsodgvfW27jQN+Oe9jDULwcs9hdyTu7be/y4njhsYlL9S++E9G2L8TDr40mCo
FSee7G83wyXc+AC+pPZIOPmMoC6SUL4GqxikS2QEvRiKAzh6X1WJgkTS6HyB2VLL
BnrsHN7zb+vfN2CXAKhd7/iIvTOVyy5Yy0yzjKJ9Mlnk6VWSHeE+0s5q/cU+xhIH
Jss67aqmryNsMse4csw3x1N6V8bIeOca5dvaL1wPNMiuYUi7dTTINkvuIf+WOavD
jAMu+20psdL9XZG1HPPvYJc64kCZW0DGn8D1u0yOxzjDq6vOTm0Bs3KHI4zIgGAk
Mfd7JS4Pdo5o2xVqH6X77bne1lL+dQuD3Hj4Mbvevykjj0D/NLAyC6SQWxJ1/zuK
+XW/eLwxrkDFaQMgFIr7J2Nk6xbdXEoGrijJIagjn4WzujnR06/LQfTXKkMIzWCJ
SoK0paOevz//PFrAJox36syaRyiWcYW6mcf0NLybdGZ1kJ6V0dkXmofrJs5cW6ki
/GkyzamnOKFpfEoOo4/JY6DcIJLDCEl3EGaGvX3dr3zpsVW+yblOUpCNee53R0B/
eav0BkvrcIc8F1IWQcCo0B2cE3vHts5bMBFFF6vj7EBLkrgX1JJTnJTlMpbLY//v
eqSMg3L+9lbIat0DDznaoa3W45Rr3xrmFsAo+lafISmXz/9QNwzmehzXGblV0R9e
Spv6lBEalfxcFjDq2BDmILW7f5eWHviJEo4AL8HYn+OVoVNX6/0vaTnihGUsjsUf
h1+2BKIfFfUc5UPVvGoiPr/nfMVhaTRLlyE+Ct0VEPA4OX2Q1FmkZSprkoxbq8sI
th4W97eIL9OwhspEpgntDzNF/ZOMfdq9V+Z8ZNH6Nf161KK1Gv0s5QsroKnk727N
g6J0Yt7ZW9/u50bLT+tyC22NMJ3zY7vwn3D/CUjBwHKIbAbncR28Ub9qZlLWtkXi
UxXwWQOpHekp0+oMGOV5CZly4VLdgPoC3vIqmb11ui+8p7euwAzrVbe507qoX2/Y
tPNYFuL6eRdBaVdHf50XXSl5rF3PIV0fXsyxdC4D+oiJdV9AhwQTdhC2uIBoYCZU
rtsUzDtH8Af/BV22gtBPp6KiGWa+vq7PBcpsYYmUF11uwbq6Gv21tXgwmj/N1Vjr
BOm00Dlikety9G9NV45li6vywJQjfZSzCACry7CSJr2521izdNRlG77tcSDvQO/H
V6CxRZjMGNW9OotZ95+2eMoYhnPfY6XnlwFSLiwNetCUBmwTSvrBXGem0yAkl7Bf
DYDdsXln430NviIsY280AlzbDpz3f1d7B1OnTt6hXXIxjYewKHGnT/NSHbB7CH/H
dejSucsA8LklhR1EM5XFULbP7ri1xwM/mFafInfo/dxvbB6FejRk2AkucftzPD4Q
Jbi3TLACSKU++1rO3+Vo/dUjuJXeDSlJOl//aMuNBPc5hA2XF8bv9whxPc7W3w/2
EaFe7mAFbZ9eeuLxWHIqsyrvAMwENwb9yQS1T1Laex4IZTueiaB8Z5Xm9h0MG/7I
Y8QS3gEXocBQRLbYXMAo+VJ0+TPAEVyr+ciVjrwZiq+EVS8vfU79o9l1nqME+yH+
R+9R3+8K4kWrskHTAdw/sNgwxYn42LEUJ1r487h806f86sI/y6m85WSFqrLCBhvD
96mWVNYGJVwQ3jcUup2UoPKj+IjKqFl/DKeGD7ikx1ItcGhGFFuSi3qE1G1AAP4m
MaVcP0vgGlwT2u2ZQWwORT9UOYQ/1KTTTPduAiFhQne9eUpa5gofDTANqA9AngM+
aSYVRji65CzN0fUGPcewvowDuhXdOKHXBVXoe7CCPKTkozSDX9x78KuehtNvGrvc
h5PvhEtfB6AK+EwAZNq6iw94jIHOJt0s5UMfy5yo7tyFUSlcIy/HxYH6Cg14LQ64
LyXJee2FX0zVhYMGaxYozI2LPqk8oTONL9yGBgyunrYcdVfLiXZJblOaKrvFnNAW
RYPp0TF1wj0Xel3OS0EzdXS81b26Wjj+3/zZHJDVpF1vrlvEHcHTZkwee/1/qKIL
sgFADzcE4uqRgEVXd6RBfZyd3TZQYInWd22qASF6FktAnDoMHUWzFQCBoSx2OMz3
e6WvCUwtue8LtlFwTkDhB175p/JQNyHemfm4m80FVeLhSUrnaf0kCLPLH93uUPRU
qi0hB6zwhG1T8XSzXJnefoKLieZMhl5127OCNOIf1FhenP9VJOVDgYvQQHUr5M/m
7ZxYk+d85NwW3sdjbvAf3E1bP1pmXGqkuxYMNQwXyTOcYVVXFpqyAluEcQk5fKqV
qc8YnGvhNO4kAU3UvpZ47rX1fBIracDU6ArAUUuqYIaR9iQ7paRAajVZy1WsBN+d
8l6DfebabkKFbVzwcc62lhnkuaxtNnOJPVZjH3dlPfyxxTsTjYa/EJTCnS1SXnZo
GScmQuda9PfJu4ZIKDGPR9AEPGPRgzdP8QDDLSUzQ4H6jFOySHK5EuvUCXGAEYhk
4zkWRczeZ1656hX2DwqzT+t7zy14P6zj+XH2y8dx/mU1CvHVtwOPp2ggy63/sihJ
jWcT4U/j6ZURH3Ersf58rfECv2lgtCPM5RsGTr5/Rdgc9SfgyxarCwn3zny7Po5H
kcsScmSaHVD50QI9l0oVyPriZFlrtxpf6cMEhMQW3pPgNKSUWpslpuD+nsAHeGL/
B6khq9udwXIQ5NE7vU/RGuaQsbnrzkWg5lL+dqwlLLDBb8BGyAc5aRq2rgIarN70
WUTv4GUWFeYKyTwQxFiSp2UqN8Qu7mX4nrhOjs8g+ixLwwWiNDSBbFTYAR6KTmX3
ksu/CtTh6jVnpDTjpKh9zS3IP1B7bIg+iag89Prtqk86ziR61lQITtkBsGgy9MLq
j4J4LYhjAPuHAsh0TdW2jLYWoVEyWtt5W6UgluOrfaue67pLeEZ73ZwyOPPL0Hv/
DvynzXexbU7l6UR/i2oU/DsuetMr3E0Iq01OYzX6M3HqH6fNWPpRq1esn9eN0Qj3
ixX/mGF+2D0l8KF7tG0miTdnRsyLSN9+3i7qeiP/DBfzhw5Z8lFxrSgJA/UeenH+
c5qDdFg+yHOmf/9NWIeAeiMWw0vS16yBiRhmDIFYoMG4OeJsd2KmvFUz+SoGy4CJ
F/AJ1PR6nL6fs9XmeXyrnPYj8BT4lygxp2FhSTv0rnb313PammG07xqvwsTgKX4Z
jRwueIeUkGPRNPc5tYL3L1Hgg7QkL9GOJM1F/8KcGfLnJ7tpuTkOCAGQJ39kLbKT
rKcYdlu+uw7QT1fBNXqGn+s9geLxfRkVarZ/qGCyKjD8Wmv4g3/DYaq1omroS/Ha
u7PQtz8oJ6DRJEbeOACf2sPkE1zQuVBikQs1TRsFcZBQLM21u3D3Y4M5LslNGnuv
QhzPPMJQQYpXU9f1cjMAiACSJWrFVWUUNyTcC/VPxlAt6OVbf/Vff/0SJ3kqxr8X
NTxE/FeyzSI1XA7dagr8tRRQ0/00tSjlXpfi5RlB0q/njDQgSDkNb4eybi4t7c33
09FQKqN8I8GLyf0uBfyRmrnmbukfSUGylwvc3usI83nJpAfELMDiMzwfBMwyZSnE
rJTZpjSYUpUmoz2RIIMnlB61FUGf4xv2kfnOQpJqj+60aRyf84BcVJ6ClMMqE8vM
DNoFR5tQS6ViiGBMNLo4kNe3jhS0EsvZf91DbRcrRa3PTUy5fDR1e1L43aLY+S2C
Hr8x/gMzqxsTsWML3PoUqXkcs6QLHw4BryxP0mP/DhTuytzPia6wRD0M1Lj1ezd9
l6By3I5JLJ2KCC+oFvHQysslF0+ctP0fXxmR26wDPUlTGpTO2enyPVbOaWpkPsuR
KshFRBI35l36SbFPOsX2mav5tVJidnuVnaf2Bk1am4f4BF4P9Xkdg1GtFeFhiwpu
Yoait9yVtyYJN8L83ttkozCkAmPQ9Kyxyq1Y0u6nYh6bu7U2j0xgVZSkItUYjVfS
HiMAGzyQnXCzhY4hcQjQMZrlSfuyhP1H0tAyqBGJ1NzVvHEldKIFVAv0V9s0xReg
yDkU3mnubI8zuu9JFZlLDkZ87DyYQs8jFmIOjnUikZY8Kr+/sVqF5U6QNJPc791X
C6hWGupSlFUgwTe621uOKGdjgvKsnh0Icfx98TW1Rv6ZUAgmFe0+JFDL9D0SHECc
epBezhVX5wPJXwL6qOroNaQ7ASmdz8nOE9L2eNbDBvsKY06sSY7m0OrQhC14xb+z
PUZTNm0l9647l8VEZaeYBLzIvmVV206Mm/5IC2d2e1RSs+dmHYcNUG8onfHIZ42T
Zw5rBMkaLRkfD5KCzF5KkTaI7hbtAAj5b4QAfLh15ktRAjU1T2G17Bs9g5ymrx3O
g5Pw6f1qO6wEcM/ebaiDsrNLTQIzWeev4cPxe9hU4gXfSs8gBkTUPNchxbdjkVuo
+wVtP/QytVbI/yaSkMmJESZRaA0WNfkslBvSx16a2QO4/uqAQ+tYS8vdx1IYWiEb
yw9N4GfSPtqWfgKg5o+3uzSQ7R0+tBJokae9GeLhBcwLhI/ztqdTb4tgmAgFUPld
I29AP+S4bNmECkQTBNj8uElxzvoCbUwAZckaIgwmvY1+ic64LV078OdYzP2Qp7SC
IST0QftfIEvJfxVDkZdsn49NqVaJEyOWUO6u1bX6DFlMysz+X0PVdJP0rTAMzNru
FfotUxYiy8lJl6a4yLVW7C153RFkYFLw6+0Qg0HbNxukee/RCvxjF5/E9E/d7y6i
uh9hsEG9dOXJa8ta2ZPueiaCmpnc8PxsP7A6jCG5IvDsBNyQZUIzTyU1ZxD1qOQg
dzOCV2vNojU4n/UaTcnNnARlNAK/8yPvTfn33u5gcnKWX6cQw7+fPA6b/VVtpWne
+RvWyIUEStJ3kVYh+u/f8MZ638h5TZIVxl+uiQP18DNJHf2wevQfa+cNdCHs3nvx
ncaDT5TamJLma/R+TTgHAkT5itWYG7EFHpikmMTsoiu4zVslWHDs3vsauRO67Xes
67+jP8bF2E9LjmuYxK59WYRTZwTYogDRPEBmlrO7n1SGfto1U+To6i6G30FlmSvg
jDyONTfZzGjX0/Ecy+cyW5EpjxFlzDaWsiyLnkt+qQbcltpO5ADZSoZQPVDrm7ji
jy+RfCj/ftsnYOlnBYi6XzWoy2ht6QRsS6umO6jC9ZejRb7Vh87Arp4qVQEbeb4n
1QLIJO8sF6OIHlYpGw/BFXIMaquDlnwAlOKGJa7w0/USi2+Lt+ANEzEzTpWPyR9i
y7d+Tn0PpZQIP8+RmXCa9D+9XFIQKtodDwghYenH0FoLS7O0a93w/4ZmcTRFeK4Z
cg2Dgy9I8JnsSrx7RWeyg7mUJpjgveT4SRwaRtPhyvWvinEMYecTmip2gKJGUSg9
2iq9FnucgM/3MUWOjrBcZg6Sr0lU4jQ7ksP3cNw3+4IIoFwDusHTiYK2aOLrPdl4
1Vp8vHscGlMrJICo3nWWnnVY+4XsW67MF4Q3MY23LVsxomr9T0LVpMrDRlo+PsTZ
V8gUhZGgcyI6Gw7Lh+m6UTpzqILUaE4bkskp6xZta3DquRvAQe522FM1N7OH7pQy
vbNLL9MpKje34Q9DOVTl1xt/Nfql9JNGW4uRtUC/8lUoJapsrtXFD7z1Z/wpuQVq
PSXVUJge8XUexVJNXyvw0RyfB8BogqJ4QdajmZJMuGjLHwssksjU+L8EO971zasx
MbNs5Q5GENqTQ7+ZTSfOm4Sc+JKLl1Jl5vzVHcunAff+e+BxMni9N3OkiLNOUz1B
FvdSCdS2kY8NaF8talqa+IXksXjpx0bjL+b+KYA219+1MDn+eoFu9cuaC81CgQwq
/t7o8rbdQaoeYRlOtq/eWo4wdgjxmG449pUAVZ1DkMwcWYXsyAIUmiyLBKr4uS/e
q1UGXhWy0J1ogxa7wypMc6z5V9mHCYDzwAHdW8k9/EUmYqCCeceA9+Y3qoJ/jSyn
pk+BODkwQgeXQua/Etvb0/Qtv+MKjo8hHmXk/Y4vND2z01/7u8eAvcyKIS/cdLug
dM17cUkMBR+WxK/oT8Y5fRlj1mB/nRRcrXiqIpSEpQt+c4y6++k3Ce3GlBRfjGVM
LfZXD0OHGLXclESbtA15gmNea3PoemLG9lAbhsTmzB10HhPPfKBOF3nA3s3/hNgI
fbNm574fEtrprvVjB4OZkeC8KM6QHNiZFokgmWlKayyvZ6duu7BOrVDNaQyuNbZP
BLOaZ9vxR0DzvZvGdlVHhlKK7+DujsqueeS8+ba9BkHyFbRt1aD4oc9UULrmzufn
Y8Gbbfoblt1sqiT7++++8G6PseupALLzwosSO1PQj+Fg2EXdxwEKNL+F0K4WK/Tk
FH7w9v4S+oQaQK7Djx+nlKq1nLKupnA4P3j2yp+5g5jgWfdpjVMk3C8jR7+plA+C
Tnfqrp4O6dLjasj5im0FDoGMSZ/4hCdhKUapFW2sKCKPZSP1x6uqAud0pkGMmnAU
NaiHFowh+lh6g03RLyY7/7IJerRnngBueOqke0CN5sQxVTNTuSZHBm4IXHy1NagO
6nREajPA8u2mQXkJHgC4u+DEnq6y6r2s/X4J2KByiJrtyim4Sufmk6N863Fpj0Zl
6DGkk0XM4qyIO8SSf/JtHUzK6RQGeh69DFtuO62eag8GfIItybgGJpH9LNsibPxP
DO8ZbkFN1O5mr3J+xJZsJiXKCytKM+uZzSEcllf/PYZBl5IuMBQChIq1pqI/jslR
atAq26RCvWEuV9hAyyX1IXDBlUVkslIStnlGlYC2x3AUejVdOHalhQp+cQn/X0v9
SrF7H23BZhls337iXqoC/2wPsvJjwx2ySuhgXiIHLaOs1qzw9uxlEsegbzrEWJOQ
xaQuDx0AjKY+BmAW/+t/BkrR659eS3pyNDPTsz4iJ0I0XFNWOkvFqTSz/KX8+xtQ
ytCvr+WzugAfS2hh5IEM7VIshz/btafzFWni9rIdm/bQJtC0ILpi8kYtiI6U0PyD
lwioocLF/HM/bT3HbVX7uMR4WTW5IR2tdO47B4z7KqmRsdvWaMUEp1y4Horvfojn
tzcjiHDKlXG3+rATEtQl3z8klKllMl6vhOwCbWhHQ/nUK77MTA1aFQ4Ojw6nAsml
niI81KVPliVAawgLXJ0YnXsh7Ggn4XXI+x60wNFWQ9yKY+gcV0Cb3YgOn5U1Pkpm
qFwJWpMHrxmDMo7ZmRPEMmNBfTmX/9vTjGOaGY+S0gqHpUZA3rVj/4z4fmWzyf7g
7h4+02UUjwEVXns2dz+SiGdbfEkDy9gzInD/wJSxoVK5kLi5MCQs0Fx149mRxTrf
UutWNUE5KXBiizAUmr+lqKjg8xlB0Yy5j3+RRRYFAThw91Y1l3N1jEdijXF2XMbI
VUtgWkFyc9FUl2rdH1b+XRLwdeP81I76H6nXJ8S8WeXVKE3Rgat6sRYorg3cDtfz
oQEXMHPN6a3SA3+JdLrJcUkaH9N/zTpAmm6eR/qQOfPsE44fUDe2+z2LIYHk8Fae
35NpAKuruSsvWBJ9kUKNx+djChs9jC89SNdbZLeKazTf+dhYlqE7jqnrXOwyeQRf
bjsYbTNcD1CbLO/KPm0srT0688UBZdJd4CTBMgU8xGolRmAaeIcsJ/R7BBGHitpT
5X+bcparnJ+nHEVqEIxVjqkVIC/dJFl7xLIwoKqiKWj6xhMSPaI4Wnu9WQ042a3g
Wdq6+2t1IESXXSergSMUBmCVjSvVY5enUTVsLKFphLYV4JvMR6ihroumecLif+4K
WZGI36eulJG8hZO37KLcZSSEkSy3h4k1o2M91F3xM3ZvRmll/bqvRDEkfyh6yY0E
jo4Y6Z+RG0cFuG22g/n+ZuO7V11GeFhQ8hynaiGR5w3BfKVkjcnJTk7kvX0ZmRPA
3mWVGrHLnRBNbt69QzK6hSPeLVHDx8bTQJSttRIB6jjR244qyK/fEbZ3H0X0A/6s
I+8CfBLgqyTIN7jfNfuPYEABhsyDjRsL2uvCZZiutsrcKCiXq+2syztwwUu8+Q9I
uuHlhwO4K7vqdsELq9p7IZRiJgVgYHbqV531hGIu5dkUx8WS9+jwAUsMIO0+w+wp
aZppuSaYj7USQL/a/I512oBRg10ZFLxtk1fg11gMNQLWDKlqKcYO2XFzrc55OJpN
xtlgAIve/8RQHvFTA/RBUlDAk3N+K9PiwEwSLD4XaILxK7phHz7PDQlf+PinLfJe
YkY2JMOyJfkltyanxFxBaeOpZ0o4fJag707xJ5j8kGiO1lKjyIpTy35yspWyHCju
Z2wp2iZMsimJva3TaaUvIK09lwydQ8jW3XjnjkLoVLlFQZ12FrDW5uPlFlbRJ9LO
mxAviKYYNDjhD2d/Nr0YoqoKXI0MkL54+GdtCxinC2cErMGSIe9zRp20wFCPl7rm
zNv+OB5KWcTKqZtz04dqOoIRIwu6UTxzQu0yAaXtnqbvI+nWlCFeZ+KFm48LQN0P
Dkxfa22gsfL0m/bMKZGtN9htmhnRlNYkAYFLNOSdRWxT8IcFqu++WSl5YHbg56Gp
WpvQX8a/ps3+jqC528UK5UL8av1rsiQsBAwm4KUg2a61WsXNXMmbTRlboj7UtnkQ
GLbXRV2jHo0WqOK9GrXY7NPQibPOiZ5+2D6yieVnXNYsz5hh9wuFaIkBpk5pOk3+
v7Q6VKH9xFrQLLPPUdeuZLb6o0FpjY3vT7i4yjnxbHOX9s+5EK4IYZ6LI6CtOEIL
HdQsJ2j0mrvfDcWJJjQqRhM/ljXypY9zXN0bYltibBYRbLYQchEPkIambojr6QdG
IRQfXDLZ/T83Lu4evjDSBhA5SFKSbvub3vR9Z3a4sGClsdAXovm7RAxOUO+6OwnQ
FoDLO1nSXZ9q276ieHTvlpe/mfy/mWMze8pIksFfRMr1BXxWBKC0dNVv1ZADNCUZ
XLFMEPEa/RP37iW2XBHXBjeaEbk5EVcllo5lmVwIAQRYaSn5LTHfdyNyQhGgiK4M
4eakq7UDmcr9rEuEhTTspZxhbDouamE+EdY+vw9gyD9PHwqBHf+hfRYHCnuYwLkp
WRiw2N54Lmr7itU8iSgpNYg1IUkSt3UVAVbss8r5GA8WUFIErpIBgokvWnXNnZMl
/uiPqsm+emFrOoDiwjAq54mEoTmZuX1AC+qUPjburkvGrUrjsMTjBQPErwLKTRpC
iCSZlue0J7vIeuivubtLLZdAJkU7XKPf8Hgk/dTp9/zmx5RLXEZygykvDOqpNgOQ
UtbEEHCPDLMcvLm5NW5ZDVqZ9+/uQeiIxcvvUtWQgC3fL521SenbOXtBKYDHrQdb
wC516SVZp7m0JM0oNQlxkhJ1aY6DVsDXJRvFpK2/OBqQ79SvJ93MZ/imKiTuQTtl
ZNs/BiCf5kFrUgDbbyZxlFfqFGZFsdi0/a3nl4N2HoKUjT4j3mhSWQPGBhCNNbqt
Ffz63F+650Q2j2/ez6liAL6hRaVun2flkbgYXaR95y1cLCLZnpuM6X3PxWaoPELO
Rw9AKMIvZKK6imwgbIVT9Jqs2cngSzvbL7LUn8raCS1i281VMOkqTI+C6vjoWl3j
DEZKsFrrJOqcKpdiN9c86jLyB9I+vkU/fYoi2AQYCrgwx1LY/95C2bVWtEHO69Wr
IxBqDO+ijnRXzf4igpPuKciKBCM6GnqEwwf0E2Pgvxzi6FNV1raFcJjqYflz6vgh
oh4keIwesClWpZ0F8OAmlaYxEXLlHfC9WW+gKhEF77o4UVtcbjQnu0ISdS55JYHR
hEpJXasv9su1Af53+E3KfCdcuyeUTbuISEN6Ls+SCyqurs//z6WukdO0jPQACEur
5+zAhk/31kltwWbqGqceA97FDC8qv7bZW4H3Ha7oAznC5rlhCqf3q3Ph1pttYNOo
7cAeas2N9LmAzwN8CCcIkFwsozH0LDwn4q9ate3z7AmB2ql5OA4gpJGriJyQ1Tcg
MRLFxI9JCN+G0YsFjXHGQVJk5ThRLQ6nX+W+AtRzMm7FBMGYBtHaK1h3/+455miF
8OKNzOu0b84riYoiIH6UC8dTdHmcRBUa73fXj2kQblJjOUdhkRsZJhse7gBkc8y8
hRuj7OUgN2anCKaaMGhHNW/Gxvm5GyauTXUOd4r8xDLq2MUhY/wUyNpen683dakd
vG8xHonXwbtvyODxpRO/GDJcHnV8Mjj/XZ4ZpArV3kkCUBRZTCdIxGXL3pGcg4E7
Fr0pkEzwouchuovjXsu5F+VPi5ycjOja3kQ19GGRFWNcSb9dAM7uRoQ2HopMy1/F
/7QhvGXJhrXlwh+7w2ETwwU4lPXYp84k1lmaH9X7c64ToWZeJJFzhk3763mifcE2
xTTRI6bS9MVmK0rAT16317SJdsvEfuFlulvC8LXa6Wi1IiG8GNtBW/dzWQ7TL6ct
j0Ej0mTqyKmUZ+icEsOCWxuOTfSMyyCBOVLOBfwIY1lnGe6obU4nVFEmX5+irizi
y4Z1dWBVzOsNEk8gy31yrRG32OwDiw2nDxR+nLAyp8G5mPhxB+wpHCiIeWgtoYGI
he4JCvpf476TzNyDMlT3m3eQvREpcSt676qQv0BIcpXsqc2tAV5Ac+AJdWB1owYU
TWcRqOa0wdwIBczNcN8FPuYavvs/VuxGjeatNdWklfRd9SZWwBFL7ohYwE3Uz2fI
pwgH5p3n0aSltf4DJFeLq2CLg5r5nWQEuQW6/DVRiVSMNNLud7yWS7weRD9BS35B
TeHYfoLxixBJjyBOleTRtT8zGpRt45AyMclABOlPE2q99TERdhf1bUnf0FgaC4Sq
3HgJJjKJnm6v22tBlSgC23s6EdS7qe+itUT0Uy3pKmOGlbL1z8YP2QEoGog5v3By
md3U95j5hRM6E1zjsxs1o3SYBvP02m26opjJtGdBTo8XSKyfFFrKL5r/Pc2AUVlq
laCDpPpZI4cddklyWZvYcREPoNvgT71ePYyW9oTodQXjs2plHiMHQwVEncZToDga
qSk233GKrI7Y7WddRkSuE+EUUaAgW6Io/WQx+3mlvWz+gSBIoNk9VEeh8Qth7Ac3
GSsHwNksegB/oLO0iOcy22vQNSzGsSWKD9PGPYtMG59fvh/+iJoD89JXlnfcbPvx
Pyr/FJR+8/QdvmO8u7WlxjBfYfDVIgJJG2bZ98Z6uHL7rF+gO0OHoq4NJ4d+bHV3
48u+mm1ilZiiOTxNlkIvPE6w6sVskf/tO1qx4upeyiS8tI8i3ZZKby3GcC4MsMed
7tLjSGvc39hbVsSNBPZFkqDHPvIx1xFCS5VfkGet2BcjHpsHKiIZ6SKfMsDkOmcC
zxsOCYWnTo1YiSaYfDU4VHo9xcQmirP8jsOG+bAisRFiLr5RgqHFAtC9hc7bJ3bc
Eo6M8aDoObVsp2pLuVg+FXpjDZ+e3hp8FSE6LVbNJPc+XhwWTiv6Sx3/sd7NXh0y
B0GUKdRNdwdx9nalbHEWuxPn90+4VznSqNt0Q3PPxhZ0jHVnCGtGmVPbPah0Z7n4
jyGYA9hKtEUv3fJbtvearMAC1v89F/MXXoPPlgrqoJVVUci6Z0DH65TYZK2eAvv0
ytLwsolz8mk4LspOdjK1mTATlvmQshJg3GsfGtU/1Qzso1w+CbQblSvXrY4R+J9s
ar3fy49pUSuDPiyqkHj2oW0Qf+JSCibGzWgeNNMujXq1ij+Om4FdNlIVXlqRhLMp
e+9V0fjy2ZZO2W5moAx+20jAPP3+Y2Ka19a9DfKSUlPlWyE6ymRm+QUgyWXS9/Gw
1jW7SX1hlU0xiFdSFEf4XvXnpjr3Qe58gm/cZ3dJ23o3p9Ulvv+SePh4TQ5twsMH
EcqlE3e982ebe0Bg8hgo5X+ifd/36S940I9useQf55ta6iVm8LFmq7TqhjRfs6OQ
r6l0RfxlwxoZHy6BP/haodVfyLjxAlLFHzxhPvTkqtglD3qV3bARgu2uxIXAEYDu
islG5f2h5mtvqtqlkgTWfuVSKxVJRMgFDMfpVpisjwRheoNMsZwwPlMuqNqVESBZ
Q+BlrlxIRRzx22IG0SQot4QPAD5mCVc3qVPzz5WB+fbTwn1kkeZ7TF8BWl3vB2Iq
JEpvDrP1tUIvGbCZf+gGFpa5lTO9MA+s1viE6CMCoSkQ+zPWXFVtuRQquzn1HWE7
xJiuCB8U56o9heGwIkSvZljeCrd5oMlt2TQn145nJ3OvW5IJ+fGI3aPb5YQRMJcZ
ftW7OoYp3WB4139faFju6LneOwbFj1fwWiV/O8kdwu5u1jH0ol16CqxMfcbeduja
FDzhaUFwCqvYwGH+KzxGofkA97KctWDAqsIVlLpZf7po4rxS4+7f4wtC8zwTCjl1
u+FY0fZcpG4DFb8i1c57XOACktOqqBYRRAFmQDMbRiNdiIXV0duM397vtROpFpH+
wnNMm70Dq6IPEgcb40cvSHOZJCYZGX2wq++Mo2fOuAOXVhy6odV4xgYgZnzyOo4C
w9KT3zoMqd7uw42i7uioYd86DuawR/8xrgg6ro7nBYiVfVHsxRud0BAfc6q+nkza
o2QrOFlUZDEjulcYJiI3eHCgWrXuXw6as616oHxt3Y7gA3xC8Y1Wql/dI8D1Fy4I
YW4TyMifU+SAXczbn5mM+U0hbmtACmMU32y+1/4JUF7XvFH625oAZ9h6XpxJr97G
iwiPoZGJl21WYfsAgsAQ6qNSXcu3JvJqlvQdj9GK5LVgOuJrg/vRg5kjv0bYbNEg
QikkqGmPWNhBmO9eO0AetHKk8Kj7/L2amW0MWkx6uuap10wfwo17HY3LlO2cuIg7
hncYHcQZzDrbSO0NPYcOP2b7GwB+I+GIfchhtFgp9gTguEJ7VUb1bt4yQ/w++EYs
B+/ZOr8FRsdeooZCWf0KuYHV1zj3Q5H88ZHtUplDSpSEfSaOhe8gfZdACAjCbCLr
ufJXBIHDTm2kFXQ1/4iLyz84hxBD2JzaIYyOuxFI0E2L4j5snVTYo4J0Hw4oeWQm
hawrqU4MiQ3c1BpnAyetJGN8rvjk8A2EIOwRVGf/GY752QjNbT+V15G04I6dm2z2
cW5ULMbNjUBd5c5f7CCwE90UdVYIpvpfdBqlY+qvgaelbTYMA1wKFGq94IpD66Yl
yewxgXXnzsMvucwEwU7wXzmByUBO5AATUoyJrDH7JCzjkLzXvzpzhACCayECckAt
nORKmF8U97gaz1M58RfsbdBmK+ZhY2Sx1mXrqmFOpQmeOy3Npvr9G/KgSyXiVvXU
PK9TnFzypGrAwrpTxKJaD140Lt0V5Sh+KN7UZNWC8eRM4pTfvjKuZycxQa/gc1QN
ip1Mq8HEOsbGmoe/GZGu1arjrBPYWNq1VmV5mN7Q4SQHGBVI8Ikiua4TricAWrxN
zZQxzXsl8VSr5qGaGhFg9JBdJ28yiBJPYiji8zZa6j4k9r0/NWkpT3aHZt50DKA+
T+1LJNMzHHbsWBzCDPgDpeBVEGgXyxBFxsOCL7pbYrT6i7ncmMPF3+075IZ/FqRb
7AoBH8lt8TvIYx4yjhIui7wtdkBY+Z0ebFplmkh6tRRFt2EeJ+GKS2jurRtyN8mn
b/t2AF6M5HtqraKP4wA/ecPx2okQjy3e/AJshO54+dRfZAvOQ4J80mRXT4Q4hfsx
RK1ifr4WRcxHemVHBTrrFH643xtiq1Bt4WwIQsfw77yOg+HYcgZbqHBxw1kDfGcF
ZkLuICvjy7hUBrfvN2Y/i2R+kE9BobWi4/1mlNrUuIIoCN1nobnGDCAYk+O2Qx1U
BLF0y2r6ee4SLtIOT/dAlpRiCQSAPAbZQT4WzZozuDdC/UR6WlkO0XruImEV+Q23
uevpgE7yK2ngtWHpclSfmtko6Op0LEoJ8Buc5u717hak0qgoXH7MWiVNwrtyrgzA
XE2kYYCHH6C6qgv/ABc+qIHCAxmyI//KCuoMl4utXZJhZCHS8JvT9lrBOqzd9Fej
oYae0rA28RTxcOydo5J/9SxPxvszm7daSLfJ5+1MVGjNMHYDv3yZB8NFimps2+Po
IRxdyBsNlk158KyjIoQzpu8h5n96lfN65F9P/bqs5kQYNgzHZnz1yDsl8mZCHUWL
h4pSGbHcqv42CiGDvY3aqIaKjKwaAieGI0hsE5XOYVGpXHMlPENc1hq6yTf+8vO5
HksXQIa7aDK96aRrlY2UMHoDV6+ApyL/4Q3z4f6NOprKk0NFBI90fBpNm+m8ncmF
nD48HCWbvxU+s42Qwi5D+tMwmmCXos5agWlJZW9R41FBXxtpAX52ELk/yoobT4Bm
YynV14MB9Cx9Wfv7Ef6pUx6faeeoAU9eodRMlXHdn7DKBU0zKieP4A9m8mOOZgUQ
emyjnweo+dYliPbJxPTop6Mo4MzKFQdfoQD/JNxXzZJo5uuv/O/R3NBqnx1F576d
c9xQ0Pdn9RNkfyEA1txnWhZxwCPEj17XXMj7i+pPv8xDOLeA0g5E3xPkURauucyG
OsFNCxT1m/AfvvB31UtteknaNUeONSWTZ47sbWMzrwhzHk/dY40X2UzquwI/jPIv
xHukHbVQhNfUj2fBR3yI5sYOe49ep8fWr6I7u07kMtTpxWsOmZHUbyu8AaFZPR2/
Fmcv4z3zPw6BANDELk5XNTdpIUeqmlXchMhFQEZhEmpo2wudlwRr8B1XVgcXRZBU
UKyUzZVdZQIlHwBCc7UwTYt8TFX4oWkzEgpOtQBVkmlMsIJ/mHKJurUn6GeY0/Tr
HLU3jkghkTW9MJQEgXgl45orCWXM4B1bXc2eKbSu10rCuRk9zGLnLA2VyzRdDEsD
NRI384Ge8THvfILa0faElbM4VPiSexUJzqFdBAvWoVkZrmuO7UTFzr7hgZnsQ5gY
SwkFt+GvWPYAEF82eksBE6X7wLfuicy8umu8n2KI/J8V8zq1aNSqWVDlpVvbuYZQ

`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
ZC3aCsYaUkBbkrvzbKjUjVuNhY1KjTlFuzddXxzXroZjV4taXK4W4MQbQWFm8v6ziaq1fV8dF0yB
SPSpAm7hN9EBhrg2PZobwRfeeM1ujgBY4OweUuHMe8ZMF/B4fzGAdhXS+jGjmU49w8U3rZNRoLoP
H4oIiSfYH+B/GsJvnjLAeSjYPxWzhE1k5IA+DDdE2GHZSgffRe71KSa+chz1iRMEa2Gslw9+fx5f
BevaZ0zhAbBIWK3dJz0tJqYIUqpIMuB+9nlVnu9C9TEaH8sLSJMWIHiyRsfwjx0LkN1PXXyYpoXV
j185F5pguEUWFbZcT7zmhngOdDSg2C/GT54HLQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 36736)
cSsuP5s52QTAWJhtDlgzkhn/iZFIby17MI5kfj0qne/FkqoClW45XxO98w3i1WbsRrYlf6WeiDyh
7XSIlN/s1G0J71pLDMUgkPx69RUjgFT29djffIiCjSLenTRWrEImZ+6a+vm4OXnkP0TgvlpadE8n
U0Isnr/mUeXnRNWUSB+69dGn7zznLsuaHjayAG7hmLmVsIiOthm/LuQOl375SuHU2aRzV+9hy/fi
Gty8NRZcdI1xcSAMXfUu+4vtxA9qUKFJt8O7f6jauEyzP81YUcCk+wXUPHkfUUy4R4WpkTZr5lq2
36h2t6wY5Jkeq2sW8tVEj8pRDdpz2TXO/AUWKrz2nG6RDNsbti4OyYaNOEflB4cobwJFHyYBbhYp
uuTz/IRguZ6rj8At9qFrztABGMygs7GclG3f/7X/ZSSOKddmBxe8TpvC+EbGaFBrOIR7IK/rQtO4
yz9mnJWYy473SZa98PhSP0iib9DEdniZu4PCK3BBqTm/ppfX/rPUtVbqvi2ot/F9i4+rsE8UAJNt
ZHLr3ffg/vPNsbdAyOhYKZdNFEwsrbEZVhsTbvT8y0iYH8BRdecCsW1ubBXEBbu1in/zy6mp1ZjU
DVnG+l8R7wQoW9HAh/wMBCt868b9VdBoSMhkxQFsMDhI/XuqpqqTbi3Nfqku/+tbUkc5i4zUUq3B
94761U+sXhE9JLXvOIYx+U8EXiCoaORf1gJ3FQ6Y3VsmPIzxfMbCK1sepSDdSyuu6o3tP8sa+FuM
9vZH0walnbfp6ifFE6O5g7A/8XpxAsI8B3HwdDgKzjiTXbQkuF/KmQMLnQgRPQRMbBLzy3joRoN9
gYj3Ui24Kmxd9vQCtbR6+p05S99vyIq+BoZ7E5Y6t7TX9clNtiyLPhy6vd7w77YCdWBusUV+3k7I
VYb1X5qnLpKDgDkMjmV3j+/MTTv/v3azkGkLr3OmltlVwT+zYG1X3GwTHLupJXYGEcLTOTnItsFp
u8X63AMS00/EC9wXLreUG+/k60w5vZartyuTF66mGkW4E0CztqVCjLd/8Ix3QCHkigkavO9etVbP
zB0dskB9/ARmCXG6xxfaPa7QrahEg2LatGXsRcq8Cmgo5h7NT2dddob21usqV1UJLnhi+mb8RK4+
yvEiagyPpBUQf5XU3oEBWTi1EWrxqc6C1Ki9BlmG5/4ezwoIyHGUZnnOaOPn37BQMYN0kz7IylQA
YPIXXNo/CapFZYTc+qsyiV2nVz7dJQkcL7rMXVShzICO+nWFBpR1BYkJceGEogJdubiH5kNxTsrk
nC5cO9JS9RiHic1oVJuDO+dIkuIyTfDcRvy3eH7gUFBkOPwEJ4uTIoBTKkUqchPr+CtOKgC4JZ7E
59pFzJHz1doDe+CcOgovE4n1hANlOrVyKxkmf6fhfoo+s1yBwN3O4/WDmKBIA6QwcD89H3QiUnDQ
COhB/6GrdPJB9Z8kk/7oMbWYb94qEzEtTrVKHOLDqQEJkTY3DJx+ncuSccnKl3Yf4JmvYOgUx0gz
aR+W/NwlXkVnaKbTaF5Pf+PRx8q3GH/8NLoXYq/Wl4Jv9dCGIKttSFKgLBr46oHOGq/mvq+H0j7C
CVnW5RHuLDslC/gs1XqNuuEPa6/Ot+inGuXM8kCXWc/ZBb1Cff/rBGNs8AmsSsuQTcwgo4+YEWsq
G67gk2OVFQAnkxHErPJoFcMqTf271aATIK8nPGEkV0BUUj7AF0pY13RUDKLxaJb8llqENjiX68PR
3T2bH6u9Mmr2psUF02tiC2alPj1I2XqeXi6xWU0K4DkGi8Ez3T979Y2OJ5cYtd9tF0TwwkRy4sZS
rIK+7SdoINVmzR6U1Wh7OEiCS0MO9O+W2bHq60UP7Ozy/Ms/fwaxC15R2NVENLpt9b5q9VgiAd0x
5D4m+AttVPX+zHCK11uCb7QwMCISXE8uVptoZQnrVa7elEeGV3ISg4I12HFXrhuvNnEtQvhyXfAG
CH7X7ZNJDDrsug7sSYPWxtKlAgPVnqZt1Ym3JDZFcUm+NPU4NLxVIYfMsUj6RzXJuXnCCEEC1wlo
PneNquhgz8O/CNMtFTZO8Q0GJ7vNTO2spIUWALX4X/gGQB7QP8NrmCQnhDCrRFgBVea6ht4TLqhW
M613E8RU/E20w6hXXI8Ea9qmOQTYwg2onmNBz6varwkHIXtRMaZ8ooWTxTacqqBRChU05dU7Oysv
SJnQUIaiydWSlcbI8OhrSayVQffI39jkZSSBvVybyRSxbP8Vf75VERGl1kKVtCIw2JhSwrZqL6eL
uQvvOB48PdPTBo5da9Fo0Vb3iD7GEzyTk8RAB1XGzR39FjAXy3JvYTwnYImSNPsIGL3mIKW89saY
X876kUygjvoJsGa+ubI7dE1sxeK0H83L1jIb8gQkKUCHdrIjiYPHspfBgw6500SBf19SVrOoQM7E
3q9EdB5RFp3xClAI9TzGn5LM8TB0C9jk28pq3s3P85zjN0ILy24M6JxqO7ukZYrHEGj2glvZ9NBb
mNsvHst+B49pT0d7qrDuJZgTuJJJd+RnxEYDRAiGtdm3getTUt7YnV8k0AMGmasfyJBoM3KX7b4z
/SN8P12Ss6Cjs0s3/WXMsvkGRMoihCLpXqkA4NDOffTR4i12eBdUFfBpQhdwpWYnT+6wV/gtN9y1
7TsfNbJgUGqwBPT+6pVJ7MUJqSli/M5Hf0eE/u8BWH0QUN+WJbtnKvbW1VLAaa7+dKgxWUrujm7+
BiW5eAI5w+R8tAhvSbDgvcoZKWR8GOr3bgnxI0MymJj4vticEtXwlDfmb+z4K3mMyWTkXEcAy6DF
Y1hphQ7yozuLbiDsAr7FIgbaJzGJTvC0tN1Jo76wx/P9Luz0Y+yvFPf1hhrrG2pFa7OsOnO3wpXi
xF4coFR1rwORzFjaJWHrY0q2Uq/zfYZ/HV8THT0OTUJi2LgJGAbZOzmhnMkK9mJhNp6uJg6tywe3
CofiuNO945kzEt2ZwBue8ttpAix5z7JVEeGzOGQY0MjIveui1dJlF8zBwKOXTXS6bqoW7qIbxpFW
T1df6g5v28ebl57FB/MYziWuhi6auJRp4zUguDlKJ3D618wiAHT2ds6dQErrEiE/JcdZyex/0ybq
pQu+O9j7wjpfOUWcPoTD1T+uw4nJBdl5NEE+QF1cwkD1qXMFkN3wWTUOfWTLKboRut1/sOHF4F/b
gV+WirNu4ZAJswUoa4e4P+6kPawWABRleUnK+VsCH/G3HXEPNVuj7KzeVyuipJdc9aaGJLMVM8RE
+Wx7MxNo7SQ3TR+3VrKaBCOYbUWuFFJX3T3yT6O5JtCCo2ukp9AjnaBZBJLVk0S+uSUsKxQVEl4h
fAARyDMWnWi22pBcvFCRkeUEFD2JeRbgV/his9MdeUpKSy+H5jU/d3TcT5ktgT/d4dmxl4Yt5IM5
40xLVxwhVVJgvlXvpFbniz12ADFqd1haS8ozSepfqZJMimiLqengIl6x96mFmUQv+0tC06lHfJi5
TW0emFNimht4f4uCHwPQgM1DZkJEsdHrju8gTLdggniPbqvuZRLdEa2suGHAjvudaifcECK17yo3
A8vzx4StjFIi+g0cEt73PufVju2SUfadNud33cfRi8TNYL0m0d5e4Dhq7068Kq04nMrE8/ovCeve
pOlYFB9nAJfHFcsfrzyf+tsJPp80fjfRCguLqjKekTGIoN8vtQAJumRUx12Z2jZQH85deGz/2mrt
xlrl/ZHlgzit6HffIn4AhDLwUqkjwLbkae4UYYdLfwPwDeE7/J9zbFYNy++2zOluRZg9Dxyy+ZzN
UeibNOBLvBRpe0FtTTjx1s9BewMYF6ozelmcHLR8Wz1coGeNcZ+U61f6tfnRKl6qUjmUqdrFS1ZU
WAH0hS5DnQZ8HG/9CJ3y885qmp4HqXN2opws+m7CAb1o+Z3EaNY+5Ju6avnGXAIHMwNynYJ5VWRZ
sdlLNG4//VyEbB7Bt5OI/uGIx6dDiPe9wcaAZrZOkeV+otth0cIitll6GDjx0WVOAHFoVFSGncvs
/yionLCINXVOJwj2fGyRbnJz+21abmxpwSOfX0efVPYT8Ir8MjqO372sM8jhKQKDk0ZwpaHfOINd
1sB2qow4fLBrQf98lbvoDFPFSrKvBW1USfmI5Aqf4QrYPukwN4AfhmX11Rpohr40bb0kNFce0h4F
27IOrz5K+NjGG3npDa0fYMgxsRu3+bPrDrevY5PovyPtutgPLocjeo0QHCFWbKGq1WIvDgdmC3Xv
4XlvN03ZsrVXNOPYZ9wfCeYgxKB5cHjwqmC5NF//VcECGQY0SZ1OpfzvrR62oNxeYqvhXhhxjid8
U1cdCmCXD+x63YcHYAzQ6c8FG8n1RfEfUe8f7r21wXLTpKJRgyMG8sPiuzoIo2TVWxcpD9VMaOIO
YinKO4+NXo3uEL3De/m5l6JU+IFOO+7wlVvkbm2C84hssfR7c4ENA5GXDWoPxb6PWLTz1sAeM8j4
OUShFApJL2X/YGwItW0DBLz8BB66JPleMrfBhMMiyZwxG8RCejEWUlACK7iUOx/nFSquhHl/Zxnq
gYJOBcP0QT3wdwcd2jwdhMfrBm14lLl0hbev1Y1uAN3ak/BHdQgA2GhuWnv2GchgxfuCmtvsuoqW
DhqZKATzvmP3ZgVLqkzj0LuqlSdtHqotdBHfL0iSG/oT5RlBVdpEyzDa+LkAxDpb//40PBRGPMyz
phizLEmZesJ1JC00wZVBaad9itULMQgM9Ufnh2VTwnls3g0QlvB9AJNlh5xrCNESNMm55dLLxoe5
UH8O/vp+RB5mBic9Sc4knFseXpqdIj4Ki9rOp43QsS4U4YFWfWePs2fq+CCpx8Y+ahx6aqzXyv/m
6S6o34nTEec6l2N4b/zq7QdrOFnrpvrbDhNZhRA5CXxBzq5r33bJxbazzZM630g6R8QCO6C+u+9F
SmzhzKCWxoHKW0w6mlFgoO98FsS2auOoIZ6ZcelRfPAYp9E2CC1wW0hndFhm3vJn0UkBWrFbzPny
lUq0zCrVDGRf+FKDfee8zkgoStHxFB+OQqXj9c9vl2uy95Q5RGXH0BttZlblfRFt9wfpvLnuDGxi
dz+QvYoLe76Bf9hVu7v5z9OnaUAtbVl4gG5SiaJCe5L8Ue5olMds4saizIdFd4HIcatCnMYa3xtg
wDXyk/+sxniCsWbgXFd4BFl/DTMtgJF/62vDlLjs0/AW3Swq2+HYMgKBJW0zsg53vSbxHCwWQCJH
m0IWTJWDBoU6+V5RTZ5hKnRPO2c8i1HeV0ThbT+SRyA4/WcP5tk37gzgYSN5gqydmcUMfqZXzHV8
/Z98WxBy93SB5D7b4EIggqzICZvTq7sIDRy9p0SqPeGp1nbE4+icOr6jYru/r8cZV3e/qdWbi9tP
RfIgQZ14JHpfnLz9+wqXU4PmG1lVOL6hGSmjqBpY4lLaV9mV/Ro1Negt3nt15y226nMHDp5wFFDM
BnGoYp1EhnL2GQbsjwu34k7qXihw8+KVu9cVOyncRm+hSkImTFrzXMyGkTnChRaGb//sjpBNHmSu
lBsjRnFrtqLAZS8S9EE6JurPIKSoMXUSSuKw3RXCXjMLwZbHhX4LNxSvkEWGsZnz/tBycZXFkd8W
LO/ezm0JAkXUoG+k1r+un/QWlHXn4Wb9zz++6doNvSza45lQytTWpQ+h/rrHYyJyE1n5wmbzY8Jb
ihbB3Blc/jHI1XH21ThBuNCEIFDGHGtHsnTB9pydvsL8rf57VIe9KbozsKG6yMCPIp7X3Av7umPh
0TAMzVTFBwUpkudUMhV8az+NXbd/T6ETOlAvpcffaR8zcTbbnj4U+HCuHwuqYVyjWgl5HSpGVfjx
ixhJKgcnFE2sPyaYcQ9Zaazs4qf0mWB/M4smnBQZwRgS3ORXZefOlRdCxDQvwCBtnfWtjmCNmmxD
EeKb8MJV+I3i+m1RvdYEW7E5U7Zh8a1Yftmh3gkF0LWG3V0WD+PgXShH1M2h5MhAiHenqdB2PgpD
Bj4xhXLN2ScdmvKaydhvzhzv6quGpugJNiY1JEatSppqkVrsyMDWjhikN1K/4S2+QiuuHv1YEMvl
7jZZnt0KwQ9OtV8YNx7erbwF54d398fRvRUuz6pOaW+DErSIyl5mGKHbs8LltsazR6Ilds5SACFW
dJA8+5LJFMscOSS2awq04ZjEtuLtwnIf8aDCuFRFJYmtIBs5GgvUWGuKrjQqUMIWPwoSWvV9r9/K
CLM+PVBPEyD+CmQ7RLM7l4qAFejhoHbcqoK7knuvxqBx7fZhq8fQdVoAMW1T7t+/xR7hocdzp3dc
W+JFJD5C1xrpS30pjDMhRbe4sSwVRb/SG45+oe0ZAeCYMAFkdOyfTUYJ3WsEVIUpOqjXZ4eONCTW
m9INTQkbS8ra/G49E2ZoYqP4M12t2intiplcVpoDJbW5j56y2OfqT1zCemrWm91VSzNE4WYVQGbV
6eVPdcpKB1ZK/VLVMg8yZiG6/GXKHsIYNSmYV6ydNrdUPXdU2hIpX08iqNmtUaWpMEfM74AN1N/j
LjQjvQYOC9Arf1sqeO3jFKyJP8OQVSNA/INV9fhOTq4SrArV2kCeDhfK7a+vDyiMyy6CyY0uQbj6
TI6E5qbkNlxbEikpoJfE7Tio5OeNiwwsjVl+fL6fsoupCSqKKOPynDVF70f13ELy4l+CjjrpnLbR
9oNeSPb4A2QjvYXInvKH14eLeJ4A3V86h02HWhIkWyOLmytf1CrSvd8dzdSYVdc8F8v1bVwy6Bvq
WgnUrRy35BDh1pTf9h5lFR7wrnOZDf3oLrUf0q10bSe6WamXqQrBjCjAKy4m4OkKelB2/TBYlRM0
jonRaAU/3f1XoOoL3i8g9FQNYVbEf2QZFsFWxa6/g5aWxOXf4dCJ58cvKKIJRo5SA+16VW7B/ZL3
/EJfv35wC/6kHS8FZA21fJbGoHUeiMTzvIlY7OllWQ1/dsvrBPfqC61uJZGWkYTd/qpzlkA0xCdW
IFzOQt4enucIEd6qROwIpAFic4u/aW/hBeteWj9STN08RcA153bvmhAGchdHPt/inVJpHsj3utb2
V4Ncaoo8O8X5vCmJMQygsnXf7tneFqU9QPkVxMGkLk22jQNtgNJUEeO1kkXQDr9SDXe1Z73VxCN1
EZo9AKFEzYxDKk+INowmeKUFqWR4DPWphPDUjrOWvTIfTns2ZL/UfyfIPWQE/EQEteXj28u8eZMr
qDNh4IYse/7WcvvfizxHO1aKVDia7xIrk+kX6r0uTa7IgajLgJJpjI7gNCDSivfiurtcW4AupuQJ
P9A51ZcNzpHzTQsb3AuMtVhm8mvcjB2Y1lA7ItaYlP/tsITGFqxx5LN6y1y3XNJ6cB1HkHd7ZpE4
jE/WPsXDbs7IvuVozkT01Tl0ussFdd1/cILA30A35zG48Vi7ff2531DpPGErxNYVHccaJ/57VIdX
1b7eVP3EakBUBm3rB4ZlJezDAkq3u+LOcki+8Yq16FWsAnP/kd19SXWFia/pZz/H8xLD6hQvlBi7
0DUYnRm899u4lUVhdRoqBH15BMW6M3rpQfFKB3rhtZF1eflcSwenUg8+WOUx81iXC31jjPPtVOKy
alTJ8sL5sXjVpmLHc99cLXPCwRYPlmiUXbWLPDzf/7RA9P3wRxS174J3GyJ7FGw9caaG0xMUviNW
GRW+bz0xU3r6ZiJjmlixdkhctiK0mA429rJAgUoKVGOmwSqpI7ZvLitFFywjCpqkURdSa+89t4rw
1sk164efKGbhNeqSqsFN/G5L/tulp1F6ijvlMEB80dc6qELO5VZbQJciAAbp+Jdn3wmq4/1vFMNL
tyrRNDUo6OhPHMI+baF25Kl6uCTCgwdzwBdmFpmpD/sfM8Om327rtRGjE1c6Jfz+U8i0tsMDefqW
gFsOQ21fQgH3dg/nezCwhnLkPsmlN7O7AzJ/gKMMbXZI6L7zBz2Xlnm4aY6/WdIsmACbK2pxiBM8
oGphnPU2xUbB/zou9R/Fh/52/vJMZj0pyoHuJCF4GKkSaaUojA4To8OWKpn0jKYrK5XuoBN1tLUQ
KuK6u/PzIO1T0idulLcqFmpbjUphGnsWJ6Us11u4MnfXT0rlPACjp3jG0Zl3NBMByJceVzCYOFMY
xNPvkwimw+dDZg/HDuScwAMYu7eFFQ1rOThwadM8KphVMLTWkVuh3cAkyZQX+/UOmo1oxxd6GAzA
5xH3sLSH1hwTH3UES3BQfN5U81w9Ao4VILLccHCnC/VwhKsan70X0aN/kRzIyCQkheAU6VI36DpL
htqVGQ88PI4LL3HTWQ/dEx9tcd/65xdkvnk5jXstwmjRMIqllr8GhUJCVJuYb7I4WHfwIuK6LJi2
ieEG3TW8UMdVxDu8BOFBXkcuSn9Pu7A8RjZcUqjK1LQNp50z/ZXG7G3GOs5VuUVx9GPBYJJbLV9W
4nf0bPyEWWMfBMiCcAE+jVFYO2Hpk6PZlHGOnmGXNLAp+Nb/CSpXUJniXqpor5t4SA0Af/6ts4Im
x8EeYNCIOxxpNJ4JpS3DK9vPspi8CeOeB8/4mcKK+qtplaY3vZyx75wYD9kMnq7OyMa1rQJwmTb9
1JVW2VusQjYSGfMAtmR8QGlMKsjn/x/sjyIdgffhQ0D9B8S/jKKKv6r7GeJ3l0rGDScf2OMBFPT/
i5kvGITX/bByAqucENTIFMoSt5ne9U1D2erfcN+zV3SPxNDjaUeYSalqhfR88LLwNtpKPmDTxmqE
iBbG3sWqQTUIOt2xVGK4PpzJquXuMmt6q2ODck8Bn1inTrmU4FQswXHgIeY8n4jycYc7OIorUAQJ
iIkaylkSvkkpeWq7tuTUMQJ4+vRVEttK6aZJvXuq6Nuxps32DWoXOT9YM55KwXWJtZNKr5jeUvSe
iGzMj5sCJBvOG7CqcLLNAKbZ9G8uyksNepvFC7i2IYIIS5iKnkxHSFBdEzG1mQHBAc38I3VZZCqf
vuNQjhbOGergo3768b4G/y8TU3/dIg85PflTJwklfVpaelPB4BteHj2MjnbMAAGoUn7x7RTIk0kX
ud5G9A74v/ROEHKxBJ9gFUGnbscWzQ36BJ+d7dAsWnBOG2Txq69jNd0PyD3ePQl9LJgzWNhaJ/E1
Mbb9ukdc+UpU2PMYT2tbDAi0JaJQ9k89zZGMfXffj+ijSYyUYTF8rLIDEjsg0jWsGVA7S0pd6cA9
YvXjDmuGH18YEHNgp61Q+nRBNU9NVSuHnGYu7P/oIYlW68zWefzKJT+JF5KIelMtvh+fU2wpNjk+
8A+RdN+Ftc361MtBMxxobN7astAqkDS+ItsgJmk6t+r7vzDCLACETtspUIv3GWTb1l+ifwG2KKBh
SSV9dBHqKaHcsEKBNKzB9ggrfIctCCiSRLXJRbP6IET0YwcmFeIjWa9dXJ45YGUUNPWKjc59hGBH
wJD/ga8cjh5KtePdZTLgs7ydOgYkjqUMytQftGWq4DrOETIBXrkCdNoDYShP1Jpw8bziG1q3zUgF
IqNYKDRDtFkzMjj0jCOA9cKTvUJu6NeCQsVWDxvxjTicB+IZHNOMAzNBOSf0wtsCFBYgE9ezI7ic
KypbZp8RpTQUtNx92RMpBBECb3SRYpnk+SAu/DhUAa3kJEGX6qF+iSUetxS2ZInipklmhT9cRtr3
7wDuL+Cd0GcV8nc045QRH24siJ0SVQhSuk16IAL64hcqHbPTAngBwxJkSdyCVRTKbD3P0o+yDQ3k
XLCT012jQnwNGzDnpM1OoIi2dFEIb2GqqMpgazxR8z04kHknC3KWBkAdvCyHnHpv+Fo4js3XcVV7
jp+RoIK5AiPp/Qp9juelO/FLeXfqe/Q1icVNJFyrF0tLZSuqiAJebF77dbVR4YEtVmCPj0bXA7z2
IwfXPSZ4iBX/sszuFwGCvTWdqFvD2mrErDlpZ4Uchu50QezL/0pJ5uyveDmZL6/B/Jn1wDbiPD+i
a7uiEcnGTwfKxDNFuhk3aA0UZIrkNmh+wwKWJLC6K90obw8i6f3aJMDBxD+NSpgWoVWGdrj93F1l
/XpqlnHLeYiAPS66D00KcR6LE2TuFa3AhsP6Qrr6WOB2ILH4leVZ3WplahedMkHPubyf6OnWFZgP
/XNBZO3rBkxyjIzDqAqTIulOpEKpW+qy4eGtoVtiGqxln7ZW/U5MbaHlkO8IXBT/HYb6vRTQtWCo
o44Nr2Xx4UlM9aYJClbivhAPCG9/wKz4axKhSEmpyZTZuZDqFXHHjKiBoActurXbtOKHDDO4dv2/
ztejJTscUppRy+Ux7qP1+cIEYWOMEIYUERJUO07esipGx4jWA5LpSHPhOJaZPDL/T3WbxWtgevoZ
UowqQiIOwgS2Ru6t+zPpl1Qi0SzDLCrq+L+WF60V2PsJecKrMfH5jKEDdJ8hlemEoCZbN0ESJmvx
G0yXdokU1EXM1mjNx+D8FPkVjAktvDpfUDWJxtiVdxRyuSLF5aSO+hWBQawdEt0Lv+ZeyKMftaKZ
HF9HWbEoaAqxJJpuXHr8m17Vj/5KT12knTXVhaSAKMLDH1IqAqbIfBr0GmlsZKOzM+4ZI/tdr/8S
PGLFa9QxsJdINhJ1m0bJzA67lxiitoDsc0+kt5VZ0z+OZX56KLrQwYrciowqwypfd0G9KAtQg5w1
RXzmbAxcEDBu7u2jBDo2G4WjV9s+6cl8IuJqIQotJEFOVttRhFb2rX4N7vX73LisL2m13dwUvfhj
Qgj3qaa6/7ZcXX+wgEKXXSnIPK1aYyWrvSKEvAJauX/M3oL76iM/686bgeW5h3Y0Ny5Xy4V8QKh9
o4UxxV/BLSu91/v/JOIhfBVRSGFLiYbo4Byui4ElmbDGyA9IUPn5s3+w31OI7D1w+f+W73Ssn4sK
2KWanNWH/IWK4M/Ev9hCAiap65kkvYolpX0Pz+H0Dlz+pVBOVUMtKdvESfkqqYA9cAQBc32rStw+
BlyRftKpCvAN8Z5buqwm1BFfzUyuTWRQGGdR+800aClCt5xlU/xTdg6EMdvn5Zs2egK7P8twuHP+
lLguP+PoF1iWILuqeHXajp5b0Y6WcWiD4J76gGe8bAkaDJY00bYRgLy/9H5m6LccQ/VsVmCkBO6i
rXaOQcWXZXXFj1/oCRSbgDJTdj+Y0p+aqffY/FXd1oZh7SV+BKBDwm8LzsJzmwGjfZLepZQbR6Z+
gM4/bfmgJ8FxUAgNPcry6RCOTbUqkXBvy1tU1jpwnmVcs6E//AEaPQJ/2mqkLjgMBMb0asV4vyoO
wYA0bEwqVCSq0EMLl9zWOtkuuxKc3aUAky8yg8b84SIfYZNJqPEqOxVVqeV6JyIu1aPOZdcAXU9l
mVSV0qS0QmRf9hnn7LwXJm6g+d8YXwG7k2yHHU/50P6mhkuiy+uKqIlO1kk9SYGJqZezrCSxzHtv
HVXduKxmTeQ8z9v7pWrLPomn3pLg8BToPBT1uwIvdq3NClRdsjsKODJyfrzW7uMvn5KAaXlaB42M
4QRUIu/qVwBX99GHA7Au6puW85x3RbemC8q6Oe0il8vt/wDSgOkWo33zEUnlpIea9sJ53G70ZlhA
H3X+8idrAZrhTeJg+mNHd1EUmUPmrGwEyPIVm+Cv9s2JnIk9xEvyD3PsQf9Gp2ZagG4jjJOJ6h6x
k65o+5n6GCL8Nxp6tQatbbSxU2MPkKME0bErdpZzC2TsnoY5Zrtc56d/B/byWdrBq9YwVemtyCg3
w8ja5fVn86T5/2mZmFQSO50U8QphTwvHElYVOMA+vwsdIwo6k2Hh0gJsFIM2uaTpGu7Rz1kZU6AF
IKyOaXxNFRE6xrkwk2om/1dV4mouzXbmN1empZFReTfWS0q6v1kEsrMGAdFMy3d7Y7umgw+/alMJ
say1D8CtU9DfPwewwNCQemZc/sdWVFVugf/VlY4jSkrwbIx3nHUKD1DoNC0v5XhzjrsbSlJ3X4/g
VLIr8YdRP/ZnDYXFgEz+D80Q9KD7WORnFP9LJc2sZdiVwGICCC4vCvTlkDnWLiE9Y/nRqwt8Wo/l
O1vyPHSmYXNEN8sa6IaOoIu3rRX0hTrLM9tYnavw11Ggr29cPnPPcZexnFCkAAaL6B6ho+SA5bKD
xQre06Ks99j5jMN0GjuKgzrJVXFn2OgQFi9BDiDSkIqZmkGqB0mM0hFR4coLNn7FJSamzGg5O4jg
aXg7WgiUIORGAEY7bABRZbqNNtuRdiLDvrvO2MQ/C/nxX9Wd+FdB8MCfI+smwgvnAskdc/iQzdEg
xVn7NAN+SgyeOS57CGzM1gp3fuJFNWemxaWgtk2/ejqv6cHN+9KDKegKH7+QoTDzD8W9DLIwUx8h
evJM1cWM/3TNEDwkYEE1rNGFiBEoSC4Uys8K/B8+zjYfLyeYQUvOjLFkUbFrtAPn4VYnWDnnXOkS
nyWyXub7ZjhvbLx7fTq023Yu6Kx2yQD45rMiQEFGVxqcmLgP3V1Sg6AXn9BOb7MLLu1ebUbmbpQs
0OO06bHa1vrqIfPdso2E/hAL2xzaQeXubbUUfAhJx6GnmjmCl+VQb29o0f3yriI2JacsqDSeonTo
jRN1aCazcy/q9+DmT9rz53GQ886UX34h7ZaaEXW3fiaey/9y9+bMV2O6dmPe4ROz1SnBb03pL82n
3AJGW9tASvSHIXpCoTa6f5JjwFDC20FYkSbMz5ERp3IjjnzJn3YeWGPEBHBenlpqOtsWl/p4Pwoy
5bUsWg7jJHQrl7iw9+Ip0fmkcoJLH6k94UzWJWULk4jfuddXHU1eHzAKeVNwkrgPza7tZQ6dNTko
NsTJKeMHhxvZNIG/vtuTNjGMVXYyK/bT7WaEgrwRA7yC4kOwe1egTO384BaQxC+/HzYKRYTlF8qd
MTzn8lPiCXfE1dNPBbykRpjj0/+OsnBuSga5kfiEidTJfe22abf1KgyI2KwgIk6dlQYSSOFcO6A+
k9rzgpfGV+oddXvPjEu/qH572nzCLcwG99e1A8FxNiof0qbnb52LBI/DsOsr+Z9UXpdPK3TW38zA
y2Nk1LHHOLnXK+HZWGPF7JJwriIvIcau6E6jMUnJ/rSdoMZBKRFL/l//t4WSQnPafbXbGucij7tY
2qH5/IzSGP2+u3iZSrPKIuOQjQ+dY60SzlxzqTy7JzukynhLnnolDjbr7EQwdUk8hCYDCdDA8hve
TfN+ejIdlvIrVTrQmjmFvEbKES9aBk9Yi/0ORcju9E7zhnwQ+ro+ZBKCywRNFl8p7jF6bAtqOYP+
J0nIYAF0aREoigBAwxN6otLhztltZmZ7O/8q02BDbOeD/7My6GAgFLrRUqVGfN5PrMq061wKWMQc
Q+eKqLCOPcDtn4QNGGD8GT0iC/08Y3mW0xRmq/PxoaM4He8p1f/b4s0SrwCR79Q0nMWm+JYyf/PQ
HxuQjAIe2S79axFDejn+xDranQlSpcw2TlOlGBeOZlSHDTtTHUQ0sNJmpVdt0zzj8dNZO4qW4DiH
Yq/xtr7je6FxA/s2tP9XSF6WJ1dEDD7p3e/RDeYp1sgo0xaKCk5vqWZK0O3rTm47wjKPeij7e6xN
oM0icXQrAXDfsVi/wGB6hCWJKWl9VsZpQdbVrrcyLNQDahn5OriYq/AeXyglWkrIukzxW27EEUi0
3YmoOAfWClidup3qlWIi3c/lwCGyMotyhbxInCCM7FyIWtTxfk3x689aB9U32Gu+LLa2AuvaNq3V
a2CavKnyatj/C676O3mu5NOZr2wgEITuMpy3CnP9C0GwKFnrtAMusrEd3qIdo3SYxM0mGdCzPsgt
f5/WEAngV7rR8m5hsEG2pg79migU5JKLufdq1MBoiq0oXavGoWYybjkMk3JBdk1kD203GGBCLp6S
22JTMeek1MQpCSvTImW4JLIrGIlK5Lbx8tpkeBq2uTkrYd+5aUX7wj3tufGQ50+/Dsy26v4JnHbB
cQ27r9eRjT/76hcWh50SmRoOJXR8xj2uzgVc4kPonyWRJ4BcPf18M8n85OtcOOPpeePdhXF/PJMO
o5u+zOBnbC2HHu5YQreJUN6mL0g64HEGh2124VfL+USMsz9jYnz9CWgE8eRjriFwg9bRaNOLJubZ
MM37aYEwOkJC8i5LF0FDK6hDNdYFbK4Rs4LGxlNFEPH2NULZ9mbUUcQhjhmH42mkGlwR1/Id9fFI
nnLpqG4cQpkmGCM/2fFRtNoo6yzaUvLr5B57VmQXy8GMocppfqLMT30TDpqVpZqHomFQ8wlO5Hhc
S3QGl7GZC96qL/oEVnT0GVIRWPsgL8lggQeGOwBXhMkmzsuUumS3t9kMEmSLYlw8U9UObZLR5DR1
hRPAa/e5gxMh8wDYMYsn/B8aiBhUwlaaYdNfhTCdyz+3Sglju2DDLxwcwiot60F1/r9RHmNjeiwP
sSjiUvv1b39IdMPJKRaj1WJKhJzXWOcPb+lhbrD4M2UIrNTf+dJiTx+chKzbXrcC+VzZsZo3YYt5
hhhaJUMZbKEYfmLx3RCUfr3JV1e+EcGioriUtEH1yKO6t7v0KARk9BUtk48Px+OKDuZplksRPli2
BS6dB/dFLE1tIMg+cV5u3Z2yE8Axb0PK86yTda0nJYzUGezYKqpzUMC6YJAYdLcJiqTIk5/eb577
pW+X6cJE6ruQCK8kjIJEWqu0WOVrDWdUgZ6LeAAggQ0gmpq3dHI3t25P2OPDrE8+V/XGkmRG6x7d
wIy38Yjxz5jYKVITHV39XnqBm61NHKE6EdnOEgJOaKymS2M0SekSI9Bu38yyjPVldkP3U0/HjmAs
2TK+b8dK2E9fYPG7JvJbGy7RJ4H/ga9/23vWJq2ODiu5EJ4ogyKPr0vZAeoEppIdYDRDJsne18J+
4OaKCmoc5o+vY+DxuJ2/TrLrj+/h/RGbC9Cek1w+9d92Mo02Lx56AkGP5yaUUixerFkag7gx4xiU
Te1i3Ew8CP8flvreUPGb11T94rVA+Sn4zKdMlLBwv3oT8xV+Ymhzdp5XUedP3fiqOcZMhM9K/TaU
TaeaV5mfrlfBEyeXn4TjO5fFXe4aDqhp3cZghb/Qk+bLys0WBcYqUaGbsBOUtclW5o+XNeMtfwMZ
ye83LUqcykpc7YRi15RuObhZkuGj1RZ3DnynQMLlACYZhY6jEYc347DcxzpjtI5U8N7FeP4DTrP/
3r5mjRVJTGnTNYn2MqqgM9TnhLjaDZcOqBNWZcKTiJRxjjyFPeWnJytnI2TmzG3GSO6NPk9wgfa+
THMXwTkLPFkCNCeS+3QYtns++U3KJHC9n6T9pytWofKgbnHFSbR37EAMGRLQ6scdh8CEo/skevLe
H7vLZqCUBdCVeE+L92TpaPCfz8h9QsWGd5i271n6OPNaKlJAne4POCL25oJUy0iTJOr/p/gYJEW9
2cmyD7QUS2R40fB2uqEuNqB6lxTdXplcQuG5C4dZChzgZjwe3Pw+xdLa/8layznt3npOncAPtud/
q1szQ5l3BGn3SSVUgC52OqLx9deYhKbRsn0xZI49OE9cyRH3NYHq/yw7kcPl8Ns/uPvqKsdGW9sh
3Xj9fSH+sq78/AzRDXNfqLxu8hYTPEAnddotCFNt7oDlD72twHHhzIcGVXS87fqAe2RaV/BsUMo+
siYJenDEhtInfgQsY0S88y8OoD4+wQ2T49n/tSFg6qXmItQOY85JLLkRKkmwVEs5p+F5gwMIOxxi
YmT002CN/iGW1/nQ18U7nE4vzanEZE6sDwIHdGVA3dpYDhBtzfojHg+XZ/Ntwnw8A6X7Tlhuzc4X
XIa2qfnNYLPwLye23dY/C4QSXh6bTi2sEIKpwHvZz7BdtpehFsLoSiC8gHeDb/OUrnEcVz0mUFIX
Ko8ZaGoEbP2VEs6t8MX9sF06+A6AMPbaToSsg5SKCGuwnUpZCQzxylwisw89PRgFJYw38OVHVIl5
r+bQmGrANLgoM9pgEx2vxBbcux8kHhGsaJ1XiZ1qsyEa7WnoCDNk2vWLyJZaLW1cB1MSPWeoEt38
DrbXKkmdE+YKWIUAhLlyW02SQiSzF2wBQ+FIpfQ/yiDkQA92t4NSgNdXSBQqiO2LGm0OXWQGx1xe
/XhbIxowOBb2gKT/eU58kbHYX9DpabZuGvp4wyLFidL2X2wZGEo/9FD15KZZbwYMHsaKeOKamPJd
XvjQdh5RSQQ7UCmjJ2ogm1Rw21SR81FZEOkfF8e3TGw94wG/BQIgOm09FeEsBExntd+RzoEhrxMO
1BFfpvBVwJmsRzQVtGIzvALJS655Alpm0JwCfROvJqK/x+xwi7DxYjDr+6mL3yjtgdKmNDYAavPv
pSQD7fFeRyvV0toDDH/kAbFKsgMl2cA51+ASwH+tGHG42OTivlOdP9qUhNf448+th1NngZB+rTi/
Mh4Nflp+zAnOKhGXn493aiKIT1VAiLJRfpCxj2aejPoFG84zveHBV0n6vCRFNZFFfWQA0dnJ5MqA
vfu+Ct4yjnyNL8HEleFqKsFQe0zylyaQ3cLDC2kyoR0BQIDHelae/f61Qq9lKqbRn72qRX+5mgWD
vc8BMQiNtch814i1PiQenNV7hrZWKbFCVOp3OdQNff3fkWTeL/J/2CIYqjfddtjrMcOMRiXpmbs4
b7A2GMrEP4J2EkdTSRnyU8FsDRjqHwjRJyU0VM5XlnNPbQNDQqXR/TRjOydcUwaA+UeoKDPZNqNz
wnfYRsBRxjOzh4GQZpKi/0QgtOo4c6ot0CGIsxSdR8/0FvtrOEQp+nQo8r8ANp2JIqAgQO8DKI2+
c/U263SZ7ozrR/f2THW4NEjjsfXi9qaLR5BcgmZG5mY+RIV1GRUqS1HedxdKwbGKWjJTAjutni74
7JtxcXJjLqR1AZzEjxkafJsjZSsT9O81FaWP0/7xVeCWoZ1maMKzo+/KOH6sTYC3NavBvzIKmlb0
ZGjTjvo0lshdyE2cVChxjvqdhSNmP1Hj+XplRFhQASjQ/47o7g2qGBXJDqr3NCdaLk2YLTSuV91e
GWJXhEgNKB659sbAZTc/IpgrzTfE6le4yZoF9HKWfU9ZBd8hiwq+F2DuhNLRri0MpKXny66XZehx
OeMTsjyOp2Eqytuq+eX2ZbLe65pr0F8DSmgMrEliCgsdaKFl89u8Nbg4c8k7ltHvrRohjEwhPDUj
/NyCl/BRIqGMtMvS5cVnMRImV0f2d/IEX9IQPiUH/fA7v5QSvGtSxucG845JWRvex2mdyUTiHose
5aF9ctqWOUrzAzLrAgC/ABnwBa2ukGJkmsWmmAF84N0nZ4w1L6THPLC5yi78HRoZw9LWuzYXI8Eu
k9o9sx1pHwX4xoEQvzV9kbQsJgACtvza+0rkTsXOLqzdLMpTZktJatko4+5orv5ifYCiQxNBRs6k
7hKAynxgs68nPTB+Dq1ULG8Evzv5LGccU+2t9wLEjynck8Jrg3hos33kewGU9k3uEa5d/nZm7EeC
kFyslOEFaQlkMR9OPQ/TFxlYsK+LnbOUO+YLggM2nCm3FLlwZN9INxC/PG4Ec6WsZ6IcNRrJuzXg
kjRFxjdPb1FNoxu+oOtRrzOTDj4Chj7AILfDBzVT1Yd99mox6tcyF2RkobG+f21ZnWfK92IUMWl9
ERxvKMMRYwjNizZoGe32RV8N8Oz1KvP/kVQ0YMJs1X8EUrap1TfsiI2tDtMl4mD7dZYFoCYuDypz
c85luEM/ZVYYOS3yFgIu7Z4hQN8+fW2cbdmRCX2BM8bd8k7a88L4vSHYbl/4PPRKUdUXOfU1ioky
jUzuAugwIttKTYjAA33tTj2OS2x43XZ2d6b5YsWjpH6LbmGU3tR9E/qZWSYy5QUaWBgrIo6wn8QY
vpLN9Jp7ORwpMzgpkp/R6HkbWA+7DXRypja15s76NOWspcWiG33Ko1esNx1LXVV0Z8mWHPsuUuEw
QV0FCdS/w4oiuoqmJ0bR4dHk44mlniTn2wOcJq1g6d1D62U+ISPkHhEl4g2uQC8+Kr+BVAoLOMZi
hnDv7fXpKHW+30JMKbh6Bep4ExSbIw5Q27mmCnEgtwOVPDWHBtmh4BL1pSmkY1MxWXqE64OMFxVp
r6LZvkdRsAR3+H75GhqyoG6beePQW+INWhPlQ13dv4Y4MtkWdb9lLmOTL4RHDwG3pV0+b/UzWkaD
VpQ5tnP+p7idNinGArsab5u/KM/2nZlycCjphtdsjMF/iOCzsPgRkBWl2dCHGinT9K8wOVQWTd+F
AiAHsabiINkHpVNro9eKuqKVgG5ZiFeU7iTubC+t6rr3sT6fppIJRKINMFkVRUSsYoCxkWcyeRfW
xEEvbBkUr2uFuf3npjbi8fqikC7BvU2MsKcPr6VD6RSFDFF1B7ShBB7WGPyh6yH9pdhkoe2NWlsc
xayYr6n0I+J5nNQiTh3fH2Ae6azRwdNeHXtwFeGZ41Z06x2N+gMd6C+MjYokf0thFivFud1nBNs/
DNU2w+1pBcJWb+3w0qyRa1a4ZPUhEtDfQ/P3nLBobWp+Dq+CpLP21Nik07d0CKEl5GpQyJ4tU0rA
0IGrBMZTVr+kpkDYhsDkGWerSbDpJUShLZ9niIbm8ty326FxNVP9cXHhdUwPMuElqZP3CWejfpMs
Z7PFy/6C7zRjvma6xYlC9ZurZBPAEoXjJVkQTYlK7H1gJ22h0wSNg7vQiaTtBYRgTUm8TI6+cBIx
sGHKartSSdTGFbdj0tULn2YQdusN9xLjI4ZPLo00UdKQ4k1xs8yqSu1oWoQ/aP7EMMRFhsoZ71qC
RS5ltBEb55DG74e01/C2GTYHVozHG2gbIDRxSCkm0MSknVpwK5YH/3ktZa7Pt8zwtedXgdIEg2+x
oEhQU5Mtgf2VMFa/e7P2j4Oj/AGHx2+ckqApB5ObbUP4nna7sE5duknQazF9SpBRGeQ/LZr82mcH
fNnSI0EFRZQ2EN9/3xhBSMZ7uWmEZ+S/SptAeGpQeaKJCuhbFnaRJJmGJHR1p8bVm4nbGv8Pjhm8
mXCqsM0WKHli64tz3JFZ6bDYSmx2z3VLzPtirtH3Pjf1kJ//183XHbBa9qpCPjpaY3m9y2n3W1hP
S/tS/WqGUl5PqPjgz0AN6emmEfptX0kwI9JN2KJLvJBLOVTllmHzOf67TqCa6uORE/7fn3aPIUM6
hiUXcCxW1qTHokUzVYRAWyOcNzImuUCjpkOfJ9g84TgoXzXniVOK+5IBiVPNmEtFXePKzD9ZQAuh
9jyRj5CaTzujbD9cg3PKbKfOdFJvrWA/ry9Uvp+CDWEFRqeBij2Smy9TlzfGLkjLkki3DlAsNo+c
SNfIxoodeREIQJRVGEJGdUKfNtMh3ZafUMXpBgVidv4H6wh1586XQ2j28Vc1xz7zb61vRAgTOLUF
wDunZHC6xjuet9etrUoGY9RKHvgEYmOok6i2R8tDXb7gu5LAP+h348ga7dnjgYvqQPtc+hKV7U4d
QCl6HlwbdydLmgVlYxcNO3j8xJVTn+91PNLitA5EtCsBmlf8s0TMJhMOhVfl/qEQ2eT6SBq7n6Rj
ci543/ctiT+Pn0dELSxgybJ+rAA7U8gvfRU8d28I1I/N55gMzToinRC8Owa5EutC3CuvJ27rOHJ7
yYmvt8/ZKK85JB0t28D4Rigyhm7JhAeeWKDvNEzjtn/yuIyAUxjWbQqY+DOwI3WXFVUj19LNR/lW
vNFC+ho00pAX6Nrk/AL33TY3ANMGZT7dP/yMUJCDBm5KdyF9eu1gJXUpvMyLNq5t6CgMG1/BZhOP
/CxHJ79pItjhUXR0zzKum7uD53VHBZ/RperkH/gnGqBU3xhaxSCBIi+8bQST1ewXWbXDCtwBhbF3
Es1AO5pz2aBARba5QLttF6fA02CWsX82gbP/lX0kc04RXy1vD7xbLGHHYThJAJDJkj8QHnbkQCZt
lkO1FyRG//1XJCWr59siQ/lCrtjh268dgagGu3NEnM+S2/9kmFtOutN0sVaitgd1YSMrCqBX3sXH
1R4SHbwn5l/GOcAqwY06nBWkCpT9xpdDDH8TwgmWMF4MAXbA5mnS+sVRcFP5dqTTGTMHmYJWB83P
F+nTp3HZUrSAPC151wwrFOKNcySlQGNP7ZG7UU8FqwrubCcFdsRKqEXwljFFe9MSXHl4RNKoHj2c
lw7r9ykPB6266f9KrTC1bhmHqi+Iy6TjJASFLH3ApFGbkfPNcNOUB+BhuS9NnfiP8OcrE+3kbeg2
OxJZ0hHMNYjOJCNiSZnx1aAIn0hRLB6KSSNMBhlXhpDlDyyF03IF4VPXrY+MX/kLnO+7yrYGZGWG
S6Nx39uVuvLKrOQYkZk9RfUFFbIWRQJdxLiY69daCRAskT4dJkz2aiB49xEIdCjHdKdgbUorDEUr
cCbYZR4LDIKUZCTFLRFN+2EYmLOAXcxG+NZosLSYZ0pe7pM5SFjo0ztIegnOYr9cVIvZPC1Xr6dD
ZAZlcJtV2BZkDW7mtRnxgPWMhmRUJoh5Vvyotkxd8+u2YaQE+Rcszp4BRbjaVTwMOMRh+8nvMomC
KqazaGRKVuKYQbnk8fslWEhTlGiVu51sVL3SnKcL9CCOA68e66chMf55vKPkjCxkFzfC7xbZflG8
52USyifH+KVfBYTOu7rIj1YJZdYC6rKrEjTe2CaRVqP2Gik72jUvCUaDITlm1+spYfq95sGrV0JH
u732IET01mwgOZwMXShHQm2yxYpMSZxdPKqyOEXGi8JiAQBlhrJKhYdOO8dwqFGP1ZOYjwlIYNv/
WhaNsl9PaX9a/eJ44qb/RaZ4QPKzROhZ3zWjhqJGFjcx5keLWSBrK9ZXSNDiEhVDKE8z/r9oCDjJ
ls2R8rN2d/VvkhzuDLXy5Y6R9JX2GqNwe22tq/rHnCkSzksAfZXOiL5x/HfCQDiFpl/eO3s9483f
eGfrQgoK1z6VO1D0mATBdHDchFdiOz2bCEEqseD3uCFgSyY8siOA09+TlCHKXrdNJkTAH7iF5ihH
qKdfD9CcsOqf5it9i4B7To/+pECL3qSWaDXdAy65VmkF5GOm6aIPIwP9RdY6fWGzKQN3RgWG7z0t
FILLTxwsD3ZvHjEdHNaM5ASoraaaoC4ZIso99RK6WjPsCmwJjG7uVinTTuyW0ibRITTY+aWP9Fj5
2SSzU3lZ+aOO+tHD+10Aa84xjDpKT302258dIYokBiGa6h/4QyeBZ2EXS6ZKA6NmQgJiVPf3goiT
betSQseMN/HGvZL0Jh54HmU4DrVg7RqFZyEobIHXBpaX2qs46DPFtoZ9hn2s18Ro42GczRU3Tb4B
hSI98YyHaDUdxOok6OB7cqHIoR/hi1TRFuxgOmLe52yW79DjwyOivt3YK1pYT4Si5cYTjivNx8Hv
rVt2dipCBT4JjolF2qQqB58f8d/9ACK7fonNHgoOO3SlEbK9lTUw7dcn3j11LOZnkAIoAY4Efxnw
idCx2tOgVn527wUsGvtw6XAJ2Rza5dsa6sJ99LPu4EPftknMGI5MdU2FdThnSpFoZiwxXkQVuGZQ
lnx4ulN8wt8A5GrZfS4hi60jHBA5ehpnPk2CYN20F/mmzrQKY32RGWmw5Gq5DmXsCT+GTHlmldsT
0xIyoLAYIvrkzslVKKVhwKkqBlO0wMmZ3nioze5c+fAFaQSU8zBBV5k6IKKx0bIY509Pcsy+1Tyh
1wa0ece/r4VuOtkqJlIySRdZ9rIZHL2L3zW2bO95+REB/042VWdzgUVXRfzDnTioDaebM2PB8WgY
lIccrI3m0NhYg1pFXZr8SPExUgXKkoosn/V0N7D5EbbiehSVhUkJIEqofHygPQhJmyljB1fxbbde
uoo51MZh0WlWr4ZwWFMCWZrb7bPd5Tp5/MF7nt4gx/ilMLK1ari2q20Plhv/YRtI0jQtwz99Qgxi
rk+1r2poxLSxwNBCbutmBNy8UGF3qcXR8MxFoLHx/ITenKrGizmkpHdxB2HtCIjGKZGfJU5d2EXN
uTzL3BJ7Oo2ubOb/9r4eHTR1J8RkGm3ftyMse0VF3kRPnNih8niqe7cnkVefX1rxcRbxYwmx78nJ
U//kOEYN7cLqtGUi3Wa7DdrdEKOECiActBqqIYLui/zK0zGFmtP7a1SrSNnowPUHsbBFbAemG+jx
WyAduy3dZYtBVgYafXX5q/O6LFRlk7FwQnFK9mcJ0IYsjeol9LnSCXH1ot4eX0e4Z3tZ3PN8fZrn
4/HDv8okya/hY/qKlCAv606UaokcEgEV7WGgRQ3AfxFAJb5L2QVbk3LUOT8ZLPc2u79g2lY5gGix
20YXFVfEnvnihtSIdNUpH2JjLL/ZtQynnaX+H9jxWmPX2eRW8Pa/JAmZ5jSCJWSLeiJTzjxzK1LL
eyX2hS3JZnpX95Mvnsf+6iA7NX/GirvAWGJo63yFM8XzQD+mDn8W+96sZeu7aO/gUyXNiAYFNFJO
Zg9c4V8co4lxJliSY4T2PTDYKDvDyBstyA3oYF+z9VkBIBwqwYjfVZzmajdLRViRiv7FIWTm8Ei8
+/QTNyq5K957Q0xQ3Pl7D4iBD/JI9S1WHM5VAc6Cp+PG1JTsd2AcOtmqDGuupEJLBZAztGbf4cr+
gxbm7xqRrY4CZQ+b5LzZMBifyfN+LdtybmVBw8qsGLoJhlKY+oHb/Q6w/GHhOTJBofba4qiP12o2
ciSirdbvv9d1E/qsBelZOFqbQfGZeeEVh0l19CWS/AHJrFrmXKDjhJ3JPPF2ohprnWbJl3r25Nwr
R6RmJUl2MLZA2+miuyk79GB3f2BW19krRA0W4n6Xgi5EhQeOQN/LlB/I+1u5wu56nBkqfTPq3SFa
47Lv4Ftsa6YLspAPG/bOAoSjEpo9ulNYdEIDIGGR2qa3yuT7cwuoKtG++kljbieVqbcHdk6u8oUU
+XmJgxiYmJuMRFl3TwymYAw/qTyU7+KUg7tMdVs0552GVy2MQnPZJg0yKQiTjTKgVB6/su2zpU3H
/1ORTDovC1B7mqaAGoK4APMRbtXg0yJPVWvwTFnx3d+VFCbb3dPCg6d1TfLs5aLsbIBVrUcMJUdt
l90kWAg5ld3w25kKpA0jgHE4e5tlYJGUJvBbOZJAB84+dqYwsg6ra3ehvev7SZtrMqG5/I+ImGEJ
+9x3+a2ZET3TYfcfTmLETHFQp4QhmwHX0yhlTHRA1RpGrEZF+UOHSuRVPuklIxqEyizWa3Ts7YYQ
97eSLZKGRaWB9OwAhkkxDAW5SsICpkBYT2jB/aq9Llwe0N9NRtMUlnR9uE/fhoA3Op3+iBxWOVcm
kSqSX0girG33hX/3J2vWxjB9ywKW5Juqtu+qLDjIZ1IAokBcw/htaE1q0i8duraLgnso/WjYXazo
bgSMQuTkm4tNRakPlxHc0J6Og4933+BuCLZ11teyKzmpzqdLuEDD0xHn/Lr4myz99g4WqVo5QvUm
92kwzZKLn6jX4vLAomL2PJc0bF0kqo4kKF2gjH0JtijLO0DHim+huUQTeVBAyxGLA7NqFgtEQo1T
RxK9sqTL3YOjUKbJDDCn3Q8xp0BRJB4td07879YWAfh9X/mEXL49d3zseFEPL6Wcz3A6Ng7bbkLW
ES7A6PWhGeJM1mhKjZfT4sHC/xfkxWiSt3C8ALeW8bD+gvNmA7RKgEeDGvbZE4YWqlVp5kpWfRJI
cCgDSHbHycGaS4rG3MxwrQG8FYH3ZQAqa1iEnh23epsJs4kRqMdz7wjfFW13wsNw0ntxbTePRmPz
4BriqWL1GUQGnKQci508S0WtJ6q+FxLrm5N6YF5X6RPxMeMoC9AXVu/RdZnpLP5XMhUc4K25pIPG
HG/go2eLXUiRaxKqk9Aiek3VctNZxMqqXrdLFpTlmFRuVXIKDrvsTdBKFCFlcRRuTzQEmPk+eRYs
ChPvv50N0Vjazj3z+QFe7a61FdmMcwpYubmHpLqT+0RhOycFl95OHUxbwcTG+TzDHnmsAdE5oV3O
RmXKNXENHlM2ccPoEaxHn+P7LsTgfcIEAQtiwegc/mGLhFYBxFxhErtywrD1KTySpDaxPk1DZdla
9RtDJFHlMdoFzhQGBtE6XyJo/LaelDbNl9jibQZXjeLimPuUnNBBnSaFps41o3xTxBvnN/RVvx5Z
7aZw1AM1rcuJVSnWEA9OSGfNb0f2sTj+EXcGkDrvRMqPsTFM74SSi0XsV1NblhdqTXXZ9rtuIhFS
NXgKnJv5FY+PkFE396jPMQqbt5q2/5rlggf7VdrFgX7dEfJBIUpazK3zBrtSIsZv1EZjiapr6Z6F
dGYBZ8ixj8HfKjCVoY+O/n7EdVoGjLB2n7Dn7urmD22HGGC/7F16dbb7VQ8+oUzyQpvEm6ZZIF3t
uaQf6qAzX5OXRZBZjHr1agFKE8qybjavTlKRBDrJojXE+NHgOvhZv7ygW4epEpJyLY8YEH1tl/fa
lJ4+x5/hUeaF39fggJh9ugjL3ptNP7fzJgi7iY7xyxLmLFaJBkt7YgWSfCkD5Df/AzUuBLxZzxFt
S7E2xXaZ5CO6A1NaNrjdr9MYnLT4W/ofSj9PBjh03+lsRqUeVgvdNvCQ06DLQ5PRuvWUan/6aBR8
ko5Ohu75vM5x9Fvc5DVxNxtULuf5MIbBHZX3gQJpIAX4n3wWExwUEF4EJ3rG8FoonIxjdSasL4dk
6YOVcmTsaZ3F/z3CSYpkcpNVHSSwdLNoMPFTLJeREUap9/aVZQ5gDJsuiaWC2XStXoxK22KZRC+r
CylXReBqiyLvgn3r6Z2898nfAixqNxEN0tifkLo8X6nkcFn0VckxNzfqs8e0N5ByI4fieatiwLX0
dmYHAyoNmwygBVkjUY+9Hvhkn8DUTVTjT7NAGE5+gUgSQIVWoUfJNt16U1yQzDZ18BhWasSoMEi+
o3gQomEsONw9AI9qXlYRvpQQAmqVmTrDfr56xo5WxB59FDri1awng0Dd0xZ+t8qo+SE9cEUw7xiQ
JcBc9WCWGe4mHdtepIvUxN26OJffkJ7X6KJcZ76YUwG0k612DonTCkgtTG9o9gcyHLNibP2t91TG
U12c2laEHeNvMWRnT5EU/mxlIDQyVTqotHzz0KZA2W8godRvU/hxjYggPX5bvMEzfi6nq0Febp9a
MD0qVWS2fbd1wybsiXGubAx1gZVn6g34Z99N4v0xVWMm/p0kLmkDL5Hn7W+vRBvsqzXGnq+cAqOT
k98w+0Vp/dWKsTJZ4oOfr56mSPSU/XC9RHeAQunhOByXiZrUQTS9XV7+mPz4lW1+UOgY+1nqiO6z
5N1L4NppPiG8XnTkGqsRGC8Km0E015R0ryoF3aRdFkif59A0wxomz6ZTZYHEMApTOMDBTCLTtdGd
ypqlrUD6IObpFoJ36h/vAjyWZICDViKfFbg2I8mcq9Mst2Ha8y4zSPofiaASWyopqS3lpF8lSPX9
r2bfbgbAxZ3KYT0HL3IAdeqDn8Q+JdNlUj+vVb4gtIMFJReni93GCTZX7QK9LuMohFK85nJ1OJ2v
tk1ZSVQApYJa/Ql8NSyglmQqhEc6OJl4DFcTDo/2YhQ0ooBSVdWkv5aGg6hBUUsAkOlPfDPhb7g0
bgf84KdBs3yRRlxFp3nt3DkcI3w/ar0S14FzV9eVJGm8f202M9/VhBGyaXfrFrrWh3rzmqd7+mgC
RIwwOMJLUl03EgbRzBmq4JsYiN5MomR/7cl+/jCcIYgMKsgSkwtnb1TzYOuYhwJo6VRON7kaohG9
t27RLjzVRW/S1PnqPAJSceAODz0rdwO45I8OWU7XSv8zbWGdwEwTotAk+cVFpmyRFPhFlXCgeISK
tQxV1VXQt4KzGUsm1nGv/FD288y/87Agi7LYh4dtBNyCc21ZsURIBTD+pmRxZYmUtLFu5/WY0MW+
4ErectwgIMV7l+QBFzkTz+MSAgojuukCAcle2b105pZJa9HxXb5sbKAOCh2SpoBuapHLj82/xkoR
8ktQ14We1V+AikdqNWfx9iw55YCwf4kCG/Q2yyDp+LK5Cu8HQuIUVJ7CMydd+1w9IH4HNTXYvbMe
nOb8XsJa2EwCT8ExabYq1PNOlY4oRrlntQ12UnoIOTRlQWnK6B17Jk934svSSDjCy5zzMYGKF7UL
XKP8duIkrB/onsVCLM7NQpOqVkVkhJ6xgOkztdrs7TqVTaNzOhOEvQnHjjgxVjlKYVE/bC5JP18y
CYePOrin1G8wtRrD5PnoRXhL9IvMORzsDtuZ1r05qWE40gVwczW0w8s3QzG3xFg1/arAHMNIOe0N
/gQuqXzXDMyaPyE02hRqod0Ml/8v7HLxDKhzX+34cVFWE/BZaNgBUGXQOf2tH1AFtkrQMexkryI1
Km8jYFXH0cLRteqERaSynnslV7hA4v2GYnpyXtQ0YWPPt/uLzuga47+Xn7y/XCW/4+BXAx1prBBo
3lEM9dkEwWnGvdxXySjOeo0gPptWAQpW1kT+b3CX42BnKwjJmqRACav0XueAxTI+TWYZX4PedfW7
CeSHP1RRk7+dae9qASJ5UPtu8e3el0PnqCL5JDGP+L99T7R0o7PAGWBQWuB8syGv1ygy0p5is7s9
F/DbUi8oufq5ZlFq55myH/D/ydOLho85L1YcZ5uovlxHDOzdrPSNhm0V5oplVDJ0IZ3o+b7YVD2P
mSpPt3FCavkkjVeOI2nGOh1wraG0x5V70iavJ6M6X29tSFQ2HuuYbRBBTdzREpdPTmShI8mdqjpb
nblKwmdXUPqGNRIiC4o555RInE5glILWyycyWiH+HwdS091bdPVki7lEcqEuK9sabJ8JNmZ1bGPk
GlxGSJHEh6UQn0UiNjC/7SQteo/Dddg62QHpzC57JPBBeIvJquN9XJ0njSe2Eij57dZvyCIA0xo8
Vd9LnF/d9PQeFG+Uwd5STswA+xTzjsUMkVNN7zepy0AQ9RgubY7ZSggH/X0mI2ygUuCNAHPTsPsQ
o3rZIrOjO7qmHxSS8CeQtd3NEm+jJgfRVuedKWIpqrKn4hteKh4YLtWNqyTpio8CjKXgh6062OsY
j48Z/JUMW8mstq7MW940Yqpl3boSREYVgzdo8LjvAAzseU90+Oerv9RZ2R0OfMSFPzw16XcUf6D7
jAJ2a0o5KMQ+kRlq25/dnS0DT8KP0JUKMbFplhjHuh4/cGManj17itpv00hZS3plSTNFwSI0HXM3
nshSEp67hmaiTLFaW18AndjxYZ/6K5/+YA25um40vUAIxp1BoawZ9VC8cjphEDabEzblaVXZheJr
9AHHFbuyirAdzXAxFgDpuC5bRvF1cBw58mENubzdE5Zg15IzmvDS7vQEzm44UIBnQuLJ2c1oPIDm
mwCHy3beOKMYehwCvitVosdgFt0nLf+WGLMICq2DO2XCLrBFarziVI6CXzX/1VeH35b5KGPNwwpz
DtSAMnjhYItDAa5OGokCVamH+wZx09We+Mb3gRtU4xg62mw6HO+wbJ2jisZd1vW0j4X+sCJjXwEw
ryz95CdnPqTLD9dg0Z8D0m0WVQNaQBqKWtG3LT++CVwYrAWv3IklYWp/YTriDgoYDy4LL/DcTzFU
tUAC4fKScXr7g5937A3+ilLdHuytChqgKkfxJYbDHUGgHuyikItswxM8FrOXEtXQHmyLSc37pFGm
z5rdqMVjFoJzJN7rxJuEPu4gOjzXT2eIciakPzgU2YMbum+PsBoMd2AIeJSgDi0yQS0zPMH5KuJI
3wniX0kAZzX9mrvRwxZ9b/XAQgOAUgimRpKoeEjuOgEaln8cY2RSvXGEQIrdSvA/oaRPqD/Xj2yC
UTQkY/UKAjkBVufTtEk+9KDlSBOCc3VRrosi55Okr0B5bEPWv067BgnNfCnsqacFw7VhfOWHrGFv
oqLruOoNGvuf4IxSqQpSY1qTlCYdHSoyPkwfFP5AYiWwM37CEZYTHcED33YZdNe1227TIuBMurGr
Co0jty927Hf9paHK9HeWwEp8jhGPICqhYSuW+AttW5OMeXJplpwSukooDUOxvQF+VAYROViqV8Yq
8VbBdvNGiU0pMyLHdprlT3NPRcHd6ix4WfCAGvlnFT77jhiU8v6F/VZ4HPjqQKePA4NaCMBmmrSy
z4B/TgZSWBw8d1sYd9HmO+IAXr3AwKUxMYCYv9qRSgPpcbrWhO30c7gRBXU1eqXDJja/eVmBeqn1
yJhK373PfrNGKZdxxzQbLnD6ak0sgEeotMIhEtCUjB8tE5/Vin8qeESLnkkFjHzm5WFcxwyaksrw
y6lHWJRjM9vsur08x32aCTs4ue6TcmpxGZV34okNODz44lEPl77DXXTsIXOrVaZJvXfUq2iBBow0
kOuXYRyJ2BFwnHEZGTGa1OBWRafMT18NFsn0w7RZ5YFKGNSg6JVBPpaHYfPYnFC0lF3uJxoQ3GFd
6PHWQmCAjbk22xTB7YBTTGq9vLSMvu47eJ5SBaTR8Oqec/0fAl+eQF8iUdU4nFKdYzU3OY9gr+vY
6SJHowdmP3mPrxGrAqc3bvplmzhDtPUPA9fxrvRWKj3vqvOucNqecKjRx25z0ydcSLKaXn7V5LTE
JraEeP21GVVjv3mAFnEWHUX5TmYCdXGzF1RnR1miLROyrxgFREmtDoYCy3oiQJli30ceaYK9rhBX
0PoLiFWUoxeRcg9SsfaS4ZUk19L4xk00ABGnd5cfIwVJo+8rinOnFdipJL1eSVnMcLiEJFMPRbBf
4szl7ZTrGhp3ueV65sKy6QrXdDlEkBpvq05CXkVlXRX36vsq+bAGO7tkndYOLPp/lgd62nEFPgUe
PNDnWbnonyLevBlSbQKnxbuuB8DpfqqsUd2wP4U9spE3tqiOG+K18gzIT2NuLe/Z157xo/nCcFIp
W9yNr8W0AthLi/azV7sDEq78p0RHZqX35tQZRcdi68AQD03r+Y3l8xnntpWaASp1KNe+MJzzOaMJ
17WZMj2uBqMe/7cf5LIVK8+KiuTTrLWZ+NJetUmr/ZcKBoEIIYaN/ysFbD0G9CqzJdL+7ZJPKvLR
qolbuZmA/KsnxYMethPVc4H/Fx7on1JFhG2dPQFSuJXX5iLoEte44b63LE4P7exgtTrEc5rauT/2
7W8ncaBjDV6UM/W3pG3elpQ4GztH1Y3Z3n1aGqvXtOTGrySaQfQIuHGmzwx93ATtbfSMLUdE+VZm
6Wj+h+zGuHWgirHp8C1OsHx6tXll0iongMW7VCYbqn1MNNlb9nWSZvU8BlcMwsJRCq5oLvK7BK+e
Ruc/h9eVvFyO9I712UVCXmeMbrYudcokClnQWjSmO/caOuaelyQlxMvR36bDBnnYQA0/hu6uRByF
lW3zEds7tRq9NO0OlRhNakWvHGEZhbwEpxRvBTpKzyCC/sNANGQtGWjoT7b4M24eMTLcivCmdoTn
UBAN6fofXEZJN2fvKaIQjp+WgJEHvHCdCIiqFMR3VcUTDmTZQFE9fCDyhXkCZLqFy+PROa6XaT/a
NOni8XBtGlCHJTacPe380yn2bsgRQJaOksZR61IxarFc0l5/1OAy1QyY31slhoI+T73sKCnGWqzK
35edGzqYSoh74sHVfq++Jyylg6sERVgS8j5dDIAixfLq7nN8S+9jsC90r2cw5q636XVWXUyk2orS
qmY0oxykqZO82tLv8nWwW+kzvLHKLED+v/TXtsm+vau/BUJhUUNTfXInpr4FfHrZ0s8Ay7fAsmac
X8ow0XZuIxPfA6R+wxfa8MmEtij1vX+XJe9GfObbf1ZECA+X9jUsSR09uUYW63zQierMUKBFgYEw
Venupe6DRUZpj8jLxiUPYajarHuB5F3rkC3BM3fy8Z0GyDzSV6I0tv3UAwS1m5oS5K7tFXjI0bP/
BFDhIp+revXviKLR+qB8NYMm+NR4o1vJz0nz4RvzHqDYEbhrzmTb3khKYshUiC/q8IAYJCY/FOQ7
nHk9HLgVALy4riN+tKCcMAmDZZEVOkb690EZz6ghcD8dvXR8wEGBj8ez2zeVPmA/BNJPAYwZF16m
5ByRPCLPWqm/3bmErG5kvAIBfxYA8XDFUuqJF1r5aRi/xfJds6MzuXHr1F/WRXwPYkRbUtSdeDKa
N0wLrtFMDoQj3cAZ+fLNO96sN5Pn8m5oZwVMRhDCsfT7jNgdd8Gr+g71QBT9WTIM3OBETD54WiBL
JFa7pPy57MbSKggSDybQzD+oAtXzas/nTALsgMWho9V34OyyVLTzRHfqhE654t3Tv+IxVH5Ns0jP
MsXc34/a6OQywEMSNuFvby1cJY/3qPXOZv1bpyNQJuCd/b8nyS1C6Q24aVun+DV2gxB0sjqgK00w
go3ZGHJbPLbDHi30DHW+LspBP1xSfSsQBJSikaGHxbm/IWgUF1Pje96R7y6M1FFO3wVA16P7Hc8D
eEKJgDyis0cQ0vqzVWaPzxOYD399ppYowjF0OHFR6gI2t4k8N1C7DnNN8mmaed53EXJgxZbhHIjK
A8GbSsmbpT+wZ5e4AbYNBnewFWOry3ajBdj93rFwt5pKSwQuDKYG9NT8O6w/jb58TQVYqXGXPZnA
pmqUdE3EZbzli/9mHcEP81eSkRxmdYE3rVI3hTBLxPdnzxjGH/sghSOR6UGdD0eIKDD1snBklJQD
iyF6sp92l07X8fM/GqIo42kJrqHWGhDcflHPpKmmg/uEISUbweOE/K3QlQLbrT72u1APsZrHUR3e
lAppMohziFneAKQYCX3Tu79GOAukSzLfz8lMtj65XF6IgnWc6Ag0MxiiL+NPSeo4ocXGDjo6NdTL
wWNMmkBg4V/X/DoNt+owoZYOjwBfIllBbYsZFN4NxCh3Gd4kDyK0Ol86MBRrtTyFyTbrhSPfDv/n
mK0XJ/flaN5bfeemA6vnFIhUIjFTzpK+0i6DhsbQwADyRaf3ru6y7GcnqkM/ezdm/aCRB7HQJDIb
nApTf112wI0U8eiiB3Uu/41zr/S/sXjkqPO66nGHDQD8dJttprv3CWDOgDLrezhN6l6MIXZrT+jK
p4g/xoc4hl/WptQrcxzVaX34gXaZsRN6jllFAflGSpNOs4dkQPWVARies83yHZx0FduMT9nN0rDo
JYfXNjK8jlAgtBw2qA6SxeCSq0FmVABfN6OSnKx6gjSmm0ZIDIhKzH0s3rdzT7Fq0/54btvFY23+
qpB4saeIU1LqWJx2UKMbELvvv4QYMAfuoSPZtvqMfzqGDjuS/O/NGdsfsX6BqZkVH6h1ZqUT8OFO
uhAihDgOOci1ePMYzTA5FjXUNL16jWnVjCAx4QmWdrFmh8yljc+Z4goqD4a8jvQU+sZ5pukVKS8q
E92AZavIuEDkCPXGzmiuuOPFxdXe0IQQF2Z+LevQpfyol4yEKfsQbBvoS9S9U1vd7sqHnykqSKpH
FZs8NEYPjbWNLO0Ie8IO4S0SUT9uhVcn2Av8Xn0zXRj4OXTdg5Ox/2pkIjd59o2YmUlVqF7Six6g
Kum5zCUltJV1o/8YE4EpqDOU1fhraSkGtKgVYNMsN7bNmJz8VOA1YbxOX1HJWNJ+fMB95EVN7pQC
ZRheLKB6qjcujebk/PAZX7YLZ/udy6jui47AWQqMLUfiRoFmxI0oK3MQof6aU0ScdEXq+9mOk6gi
Ozl0zM0vjXwert0bN2azlVjEO3lTAM/8zpgB2ZtA4cCpTuyaNPjWUAM4Xp+NBBzSxCzpb0FJmB+N
8MnFwUKN+kZdO/vk2T7/MJx6/syCzSPi14qUx4zJ2PMaPyif4e7Ms4pcBG7+ty4+u2wJs960Zi0u
ZOPWl5OcqdDQQ0hj2NdVKOHIAOcqfsUWGRZlbVTEkZNvtdXHhVGp10qvxsD+WBAYtwKLmb3rtGL6
Ggl1SkDp9kZfywgQXNJEXs9fmD9H3SQApbRxRvtu1T4UedJlhthhWAUaf2jbx855w6jR37aq3Lox
cdVdIZNJPiljDeJ2HKK25iwa5nroGTszYoD+2b2MjcqjJxYhRc+fiu2SYhWLX7WRi1ZY8+8havtK
25mprmA8sU3bRDGqyi2N4YxMxwELlxq5Tf7M2Z5u+oR36BYia+xJIEPnA0YqT7tKpE36DfO31bQp
O4JmPGIrR/891t4SW0/gE3Puk0Q7YJH94kD4sHzrujdZ3M8eluwN9Zflg0VsP/28Gynt9ijf4Hy3
Y+JWk1vlOk2u6PnrnOVi+tJTLp/qB7Bdx3GsZdLwrZRPuQ8yNo+MwSUvVVzblHsCVrqrdYo1ngk3
kTvccvgegRZQw7U+Rb18rGkIJHlPYzB9eB4o0SYAMxJiyHV9QNuGoGeGNe21jezhKb0PMcUQG2ZJ
WQGbklPZTZv6Ut50kmpMrAkpRaUzqGAdool6OMSuBysWPyoq40RSdx6jNs6aEyBuqV4GJNjWWZxj
aeitc/4ITKflmzAhgOywO8RK1WhHZikdOzGh4BFBvxWOkMXhTUvVYTT0QxtWbp3Kx64dN4ST7MgT
E690Z0RaEXxWb40LTsyN/UntxtovP6beuSfD0r9o8h1IeN8/Jai5bB6R43iY3Lj0CAGv4/IOqEbV
/YMyWCImslK8XF268SCdEPW5wI76JxKc+a32/b+IMMyUoCnGPvW454OlF70GHDlZE0uPPeJbXz3v
12SiHL7uKqtsweU+2fAL5iKA3y0Wxdgb9tNY2aylJ0BLuyV1YbOjTYYzLpDFnZQCfjBNk+3z3rmi
xGSUtDpvLkDq6e5r6gCc90N1/XEh3g3wD77+K6kLCyH2/iGmZQPUGuSPJWaW/YESWpNiA0bp1aUa
6sN1wTJao1g0HnoBtMuiC74yOnOegyjyihfyCKMpDMp3O8dL+5xpXWtabpY+/UkYb8MqyEQXwuad
XV45TSgP3N3CE5S2x3uCux+iEIgXMfZGV4mRHrW35B84/3oM7kWkyut+5eqIX2XX+NlR8Yv2/mpr
cUXLFVZ365EHhZpmKz5+V+V9Zf2zxyppFr+Jo6ffYzAzk3PW9is1gRaG/DofVz/3k2o1YqOiQ98a
R/Y3EZYRvy/zyt/Aa+pGlMJoBiw//MXn1vy7vKLMUOgC9aDZbI/ncVeV2JeZxFYwwvOuWXO7R0BZ
8Q2WDDZ+0l9D+Osu9kYz8iwB0iqpEZi59Pm0NFMYUKwXn7gWPZiEKXIKT26C8N7hRclET0cRMODa
J5C4LFInchdS0URaIvaAo3HMmj5k2lX6HKupLmg1IxWN3clVircDX06fy1HSTCkbXOUdhbyfrpM0
uHayxA+M8qGy+t9xksaxGSWklY52ztToODeGTaWREFbUGnyEnEjLKhrjYpeeMf0tmI8ChLFzcT0P
DOnUGxUzkNGfKQyI7RiZ1ojQLUTKVswYxqLcvBmyAjzWPHYDgaxcJk/jYJhl7Dt+Nc9Nmk4qqsLv
8cmfHMfkrlz51nv/CX54eKrA+p0lKAR2Y2ylWX/yxcv9ID0SYeFz8kEOSogAP56YI9otGOdvsA2O
RVsOAiI/aZtJN6OvrJzqZ5NJgDVU3bmMzPXuSJcszul1HYafevOvG2lisXF7RaUWGjGuGijbOi94
k9x/d/9x0Mh9Z/8jKTix789rOqpD5qXtCS1h457FaHMxaQdQaQINsZ5GqEQ1a/HyeWZ8Hm3cAkyk
CrfDX+pMHLOjaAfTLjbGygiKbc2ZJXJUOzllxeidMrfCM1Ml/soJ5OxWosQFgPCMfMUbE9wTtYzb
hXk2Nkvw6v7aQbkibZwLU82+smIhmXdgnK/o29fEIeY5mQr12AxuGhonhNxludGbzRolPYGuHj20
P6G8Yf/ApaQ2dMdFcRQ9AK2E10CqRLOq27DTZsl18jU8o21668EDlXOjCO3x+R74w8rqMdhw5sAc
JzJtND1BV9flemviwSJQM1ikMs92tc6boR8S9xUtq+NWe9jwsUf89Pt7Q7yOqR/jGUk3e0PUMs0W
rK4n2JpgI9QxGnMJ0O3a3qruf/STPeklGsLEm0T6WRbeVzeN+BZTy3Pik8vf2ozsPSgni3K6/LKF
47cI9mpSnwQRaArPGoptpScTqotVKmeZ2H6T1t537ZkkpFO6BYyJj9Rxczi5DyK8PeGn1rzPECL4
7iCGa1rTBu7TTjcW7xS4dfSKsRIKlrcIc6hGRJEjjyMxr/NqEOIWt2hDIZUcj3VmAmc1INv7fL+k
SRx8KSzcTRrHw5xa6SmaFkvO0Fzb4/XCYRm4+pGTWTmmg0E7vlabo6ds9KGlroSb/BnKGRNCZwt+
SNVlHQOp9HnXSdrvUMVsZX+BrSYeAYKUsTDtgr21UlPvdi4djiPV++uyNvh84toX2KEnv1wNQBj1
T9l/asHzDspeMHNTNopbcnIy84UYESLL6urR1E0rndUEeFwpCn7o6aMllVQaJknhoxUFksGDV10d
JlrPGtpWsXcYRgBLKJHSesgXNCzItLnGeZZaE+E9M46DpULbtNFXZrPw1U960u5z1SiG7rcEPqf7
yDjL00z0gtnqlw7/HHR3MUX6mwokioauBF9Ym8GsY0JHjWzL0A+Jd1F21wMWhujRiZZAqHMeLIbN
vzJmeezjOfrdVWqhKYDoniyzCEe1pQJRi0t7lwFJP4CGMI3r/bgq+dPb0OBhX7FSVOiA4Y2Ijww2
s9tN9E5w6cBN1wjWJWTPzC3lNO9VOwuYqR7uFS4SngmynfiT8PrIQgf/4eZh892rYbmjp3Z+zj/Z
DuXjbgtdgXaiDh2Qy7NrelkaPIX2er/NeV6FUaJEWRug9ZpW1twe50Ygu/4xwN1OXbHWleY/z3a2
K5zTScRKH4j/54dFRLIDhAL9+0262hcll49ZJp1RyR/NnVZqafnUAMl2BX1tjeDuYMa2+RHaD50L
afjHX1Zpb8X93C09vVQ15IYnecQ8EuvTFINffQhnJSNev0Df8QULK/J2HGIZ7rJay8BLMaXkVcaM
QWL+HfGIQSZfsGcJxwi6yRAdhEzE3A3v/IJu8KcV1CpJODnvvyVKIFch7jKbJZa/l51hifOHWvla
LzCLPrzMwQxzdPZtrrpXLhknfRNoz6FwXjH1SLCEJRlLCVlvt1yFwQf+Pm1mTWGPuUVH/KEHiPIT
MLgqp8VHIS7Tn/BgbMv5BJn7yCRdBj+boZi3x7fp63r4cJF2ubRnJdU+EXSg+xS1jJtySlWUawW3
2CqQ21wBlK6FGhUDABh0/OX1CDjOI1tHiMjPwaDxI00i8mSoiO3dEh/jFKIQBkO3Q3pnTZ1RKg9h
WeX0W3Bh0LmD7x6rnBED+GQEdcvGU87wSvcwrwUpPi2tWvH6ETajirKU/Kl2n3Jt/bRuYGZ2Z+l/
fBQcrF1PvNfKyJKP4LJmR9TlJ4xEhif5mCYHd1plM+KrpLNW06LPvoineNHBNPHP9AsYoCODZRYO
/sVLIES57wqzGsTHNukxQos5hiaHBQAGGOC6Wa+9oqrCPPmj3JxNSEP+TMs1ZH3SsJvI0pci3Yja
QTMIPKooXPX/yWC/MlR99VgCDi7wk9UsiPw5o3Qm6amZJnj9FMX/KUR3xOh5Ezd/sfJDNdhJl43Z
b0qtA5S1oi7ofybt1/sX9hLAvlqaGJZjl7iZNVon4yDUSyf6Y1XiMhLYgVj7c3syJz2BQXWv7QW/
K1UZ1HA1Y9rHpLHsaWXaGp/z68uVIfkmv3kVKDMeD7leqv09iZHVgkQSZzZRsv880KRfwDNzuBbH
wC9HiEYLxVEN60XbCdPo+VHyxiWTw9faYQSW1wE5+eE9VHqrsLSUuDRIAkD5kLMN1MH/wAwn2gYi
BFEXhbSNUHq2QSqG4J1lr1feDehkXPOrJYmShzoxNMP0Z20yFdP84PdazDJ6S8U0qQ9UEfI4WKGi
15y+KUt3wNU8NhcICyTko0h4uaO9wHV5E4lbaHiLdVfSwX4Y3jMxMwM++2FAqo9bjh9mTH9komM3
ArV5I/C9mmtctxPNWMF31rI/NDAlgTp7o+Hve1pa0s7Cjvg09fV2kPX1kpVbs+dlpaEmG/E5rCnh
/L4dlXjDoR2xt+xVxFJbVPlB7Gst/4LuaiXwNKC5Z+CSVz93jvNdSuLyWeK3IE38KhuhG83xBpPr
suFAu78uuO7djw/baqZsf5TNOjrhEcyNQYF6etNSaqPVVQ3XyQbkZy9Rw6wDbTRogdrd0fSv8CSZ
BdN1KD3JbuPUCldcMcoAwRDPhz4jTyWDw5/JxBsJLJmR/jZDkWQLhniLhwxB8IKPQ+lpSNlnPOTG
BFbO/nlb6w+GzskHZP9JL3PMoAU3lfVYhV22kWVDoFOjW2pDLBRM9o+gmHWvYzf9U/NT/OPjiX/Y
hTSTDc0uC8Cswsl7szJP3Qrl7Zimtx0P7WCK+I73VBLZSOyN18Qp1ulbqiOvyNZXpJQbsdvhB9si
ovQ73ue6H3RUlY3W0xTGsxMcvdk3WgxJ3Bg7iLJ9fD2ix64BEerKSoScn3howc0WTlol15oV8iBN
ziBET6RBvG7oPGgS5lbMyrCtx5pxSjcdzVM0hZxIPAFRyUU9+yyqJ87V5OLXuIk7+CdbqDN+BRSm
EF30WgJ7r52SFPNyJSRjJrhchGOJq2VDsSmWADAK/gLl5wksylcAZoPhqv9JkGVJ1xz2tkyGHUae
E+2Hw62sygWkU5yx45vQIdcx9rGiO5kdOjcqYxzFOKYozqHXO8Zuh2lPEipNbw1csI2QBNbsIinb
2udrz+M2+WGK+PFH8LZy5nSyFf0dQlJS6FKZunW4SQAErb8YY2XBAL/RhMw+CT2q3aeo3EVj/ntG
nosJhA47r9GRRl14eBMPLlcCtjI+0TLt/mJfvUL13a0Icdcs7E+zWSy6ZnNX6s2AnJi+OfzzU/mL
IJLixvYHrUQakurC3G1gSN7JEs4OV950I7w6f5148ZyC96O4jxaT0In6lnhFZxv3SXzm9Bx3GMz8
FBT71sO+NXa1JfAnGs/dAqcmKXi5xcy93S15HhUmdQUm/HacQg3xTgRYNMhrL52+/HQspHsN61sQ
mJt+DUzmGDquq65LIRlXHBBPyWdk2izsIkhg+ZOofiZsrbqdsLUixgQDZqCciAGXp7YHkHNDIY8z
3Hsu7K64LUNeqHEQEOcQLeFT7k9aiqXcorHbYgjKSgIsTjq01+x1I5CDwL8mAOo/1r782paruItO
SrnSiU4w8BEXKDtCUUiCE7gajUMnC7Vgx3QbYyGOBsjUEk4zuGVZcxl914e3pfjUbbS1NkUcGexL
tNm+0fCl5YExRLAKS9Tse8E4uAJzrWeNa9U4AVcUAoKHRtqLeAFev4cbukrYoafFBZHQ+xvYsyh1
wR34BTF2s/0utC7cryzRfGvP7zPieRyN4h2CIYVCEHET+RKC6k+atDqBY2ni+RfmiyEMAMvDgNP7
eMomkzZvQqtcTAyKh8jtBqgFZIViMHvgkJ20E6wZFcEzj47dbcEyo1EfS1TqJdqVS0Xd9aYo3H//
hxOEy5qnmOFsj24otxlSX06YgN3dgml7ddLRsPs4AoW1JZ9Bs0Y4lk9h135xVN4B7t5I9zTDGEzZ
Eywk5Bv31SDywnGxrH37dEIFmIPxJHq5LIr147NA+LkNePCmN13ldQuSJLcysAyBcrK1cBrXY5DP
rIoTTGEvyZoJSoY+TMY49m1/vvPNSX7MIN8jo/4lzPAP/J29japW1Kg4wlrmPwHIle67cNgxuwtY
Za3OWKvFOa5sxvFQ8TDnPdISy1gflm+r9L2Aab+8nrkgap77g8+c/+8EtfJsvbepodXDJfN0BHlX
w/O+U4DyR9DOfZ90GsZDqbPPvLYUjRMTxMjapWg9zr7EQELeyHFnU3h+IB2mms02MBy+H5U8paHO
3bjup8vSkNMtnchpqIwMa0xqF+uUCcYsei6zbCRUJMYGT7ED54Cct9fb2qGwHYhxKCj9HxARrPjW
ZuUibRgdYskxYyi4V+cKDO5gR3SqXbjqhQ574eZ9DV9dRnJM3GGz52pfwXtYNjRHhu2lq95MPMvI
CHwEp9oLnEfiB2oDsSPWit6q2CjFC5CDTo+mhUKkUmDwcF/+dT7bCy2Mbd7j7vkzCHUcfHskn17T
PMy1Wy03IyexSSGMfn1aDFZihW3mxZojhz9BwmgaRGvPiUFEH91wjEzLgPg3vUvo2eOELGdYLPTM
HlmLzVkd8+EWaqP9ptYxZgOZlm0IPrcFzrYkzNIfg2cUwehJjukxUt92qIoXKjJvEls3vjYZqbMJ
NICEozh+iRB67fe4AkT0uko3I7cZbDWncJzms6m5J3eDxiYGSLUoJDI272IV95J1k1cuTNLrfy6Y
TwGO6fQ8uYjnzlE/7566cnNNrs1TbKZcMlxo/4/+XaaZeMUZdZHSAmFPrC2EO9NcXNwQgPU1wWCx
+aDmu0Kt4KSc+W8WVkqwO/Mf5+TqArn2EwpOz1XctwxcXxxOdYRh4tBLtqhivCjNq4MLQTf15Wzu
gdbmikrvD13GeCzPR2GFHM4hZOhutuejxfUTAUH9yY93sp6Y+vI5uvZn0vsUx0N9ODpqGXpHvEKM
JB7c2w4Mxw+PRjo6/H9COfOUxFBDiKw/FsU14GidE39aIwedZuWfl7c/PWusHDKMMMj+6kpaUCCG
ICGIG+Fjl+RDH4CtTf0Hcj9GwlDOhQDmg29mLVPC71V65NM02lyd9iUvOLt+k91XIj2y78brvATe
H/TmNgU3d7iELJXlofG0PZbf6eRbs7jULDwT0AF+30utetSumeXJ78tBdFXCm728f4OLeg8pGOLV
VkcOUTtEsrQEuJcyt4fM8Z0uul0YVrQyo6zFhlLaEZK9IEzUQgqBQe/Y+FLyrs2EZU2nDG9k5fKj
66RRFj83HhjAwOfzoyKZSnt7pMy2VA76L44uAhYt/kABT//mnn3mQPUBXovn6DsCtaN/EfSwKLwl
LSMQbQrCJNvZPK/aeRJH4Qlq6L5sGgiIgnrCs4NdwIB7wVGgw4XRV0aK7ibqiKLD2mcYq2DFWzuo
wvTzXOx1aHZ8hUFOQSfVUA2tfdufYwNgZNs2vu7AGxn5xZU7WQWu2+T/KQBSwnXvOdxvcaoH0NR/
ZWwMjVThYNbci2V1sCxbDeXXCFBDo1f0jyUD35YdXUE6YKxOdADntmAzJ1TZa5pvnrrRMtsTqG1W
IX8Ov1bZHFwJw402h9IVCB/iFT+va7MGpdT9fmXMZhMVx/thiaMNp7qEJtwWq9XY0r+EHzaOAHCg
eAwxaI7YRI1qv01LOqfgKJf2R2nYu/is1da5U1Vbr6vbEkZ0JK+QHcJtUzaK7gvT3xrIWwICc/RT
ZWleICz2E8K7FjrC0651qFKTxFYIWLkWUFOmDWZfFQWAHQzOXQFQXRXhhYQy83VQD6G0IDH2OVHr
8TeKVFSQEq9hFsAw3mVyg4rriMd5izMFpvC810sD1GkkiNMMWymKOJZPuUt5qFZJA0bAI3lyK3Su
qZod/CegCOEf8zeFcPrMFWYUBzBnpXpF0bWbMDiPnZbZ4KrdWTpme8qcobQd44s6IApCUXlXLzKa
Fxk8QARGE4n6TLHvUx+fKoLnAd9J0W0pwOpOk+YT/qsNcsNoYRIJ3TS7oJkci8fpV48sm0p50K1K
R22ZN4N1d7hTVF28dSoLU2mjNbBPRjengtEMT2/Cd8nrIBOYAvf7FmsdiDRly+i3t+WJJRQPaM0i
OXlenhsYxW5BZsVrEWEuK3WYEqabbz3XJ00m6KDIaCFcAX47mBa0tkQt8R0v0jTHLKo8mAXBGIgU
ghZ+4kKD86iB9b5dzEV1T6RRgLaonuwmmkbdeqcpQtyHBnMrV4az8yqq1FBBSgV1yk2N/gbpPNWp
s90kmdwVUAmnpmbhjXazfgxz4OMuKh2er1+z3oHB1XNewSjemS2kdnJalDlL0+N3YYu0FyrB12TZ
AFIJafDroaVKUNNU1Z6Seg7x3MQIXc5/Q0X6Lk5Ly0kpVE7c+XvQSBGviDOmKOiYBGL+EqfH8GSc
FO7PdqvBpOJpSNrxSFV8H2vRbPqTJx0iPzPL+HzFeDr5tlJM0PN+2q8K+DKFa9/ebIdmYv126HA2
eo5Ly8U9Q8ie2hmzoNpCJqCGylKu+phjjvh+wwJ2gIhtuzP5yonYOc/nP/yEmHNLasN5I2OEMdcL
tlKwp1OxnWhUnI6FBk29tKe/2lFl65fZHnKi7YOCqbai9NGC/Y5gNNIPX1HPRXU/1G/jJPBvUcwy
X78NQS0HvOqXL+JfEEA6/d+9sVOEQETabUneWudjuQbqbaLo4cO6/hG2qJWgCpZGCl1RXEUdn1GF
lCOrohg9SPiRt9DnUQc3QhKtTbyDypV/4EofbzFFzC5aCLMd7hwpuWKg4/xS0JB087vVdJqokvRx
mHowT8mavfntA56JP4LMjxXLSOPiuOtvHJ4I0Sig+WYyA/nyKtdjW59zkXRa3nSuNXluD6gUDZky
94bC9aeida2J8e7UQ+vR1JZM2vcp+PUIsmHfu0YvWJBbUKWqPEJVNxaoZ9wT12rMFOcx+0r2Ceh8
qe/V0V9zB+z57u17+CSfUM1aiaDII70M1W7q7Yp4Vb0Ma3IUoQJ+kh//KeMtZoT7h4/B9tvg2xjw
iNOGB2mFE8l8LzhNrPKIxfShTLmYPdHk92AfQfQnslOXl0xVRBqfFpLjZZi9rk/1dQQtdANLDep1
otHqiIdQHFp+u7JGkqzduMw9rE8BP3qVZnRMX6NfLVE8hLt0Tvg+6uS7EfuLxdUSNp7PVfrpnCLV
xtZ/y2L6maFjYM44LT4hxfhRCHidzHFW16tEYTPV08udYiq3pinVPSXDIOz7Hj0cHoMyaa2Z6k+m
i0yRsFuPCJ9CPMwcfB7bMV9jQ+Gjfm8OSlE0OEGHnp+KhtJD2+siApv+GVbWVEkZQAWc/m2ncPr3
o+9aI05C0v87hvNNz9HNYeb6N3SaM2S0AhHTtCqTUF81bxm/mvxCbI5xYgQrS9BTdVNcx/HmOL4f
oj9Rovro2G4NULkmn9i/Z8tZVcYumDQGK7LjLEB2aJB4I3SYtscK4QPgvL5pbCiEWO8bUKG+I/6A
cEv+CbMmunhNbY9+UpLfJlfsjwi0lF1Zhf7203rD4tBR/xbjUWbgPStxvNiR3qg3IN1ZaGlGTJ5N
sPxMuHviulylOGlkNpyJxS3nNCi7rYbxAqFN5Dse59ZZD4041jr74rUT32mhdePtlB9GJnD2B9YR
2U1n3yF+av0E7oj2ne4Vk945YjSknk9JHOZjcdy1QNs0grXZN8G6UdJ1RS1Pm7DPYCDrqYy2vgFz
biZotOarpffdUDddy2dGn8k03/bIJ+WxDqDiSoQqQO0LR5IOJD9PrYY+6/Pw1E2kCFrdl232juA6
BGKG+71TB5g6q55z9th+A5gPheMUcr2G9e044ScXa27L0NVG+loQrtm6B+H+09C7yJeyaqi5vDCu
O0lPc3/YOTr91HkTsM+k375mkVDpyoSkKjIxtKxYN60MTw7Go+66587jAq71KLhMGTIBepjZdMcR
ir9AM7r5nre5DkFw+J09ihJbzb+rsELZCehQ7o8CardaRwu8OihMLRkZOLXRc75lMYmcfHUpZlNC
Yi/ZRlFr7vnE9zBDCPeMRliYC1pBnVA9ag3EykpcAVtNaT5VvSvDv1qnX0gF6LhUaZCKVfd73vhg
WzO3mBa77gZ1GdzqaMzGimX/J1g30+x5KISaHZVuu1UqaTRDRwWiYnsX+WrlSrbYXqO7hbSQ30fA
D2T1VPr+JM9oA6UHUMzTZMAvxUM3qZp5NjGbY0U3tBydKWauBROgbag3OHG2RGyqVoy/evFFDPUX
SYcwZnbZLR23ffVSJfmivW9cQLpvsLbcatRe9OA6GVTy7E2gpQytf+QMsk2XyzM2m1iIuFuO7zoG
PsMp+T8sYdoPEA3izb4wtWbkMno53ziWqllrgl+0VVafW161ZdXpP70vlLqYwfZkNwZneHf7uhwM
xO3uM9C+IEE+bZVbfc7CDwmdCSWda+fYXcFo6MWulLOh2UT4WJHfssFi0qwPDg8iH+TU7Y9F2O4D
fVT/GQ6rC7rvlsZJ/PEGOYPzW4fkrPubimKTOAArYijPULy58pMi9Mxut3fxUnwBLaFsosQ38M4e
9s/K3meiYBeQMSkkjiHfZE66h5k8u1tieyJ+/r66vFl6aH/e9dKwz2YouGU1OaxqaZx9HECk+vZm
hRvnbOrmYPQyrA7yL6Byi8O1w1GMWMSOtw2C8dl4mCY/jxYkYVjmAB04O5EiWj9RsBjIHiukD9D3
Sq1h4v1UPj6VdU9V2OGsa8zxBjXquSFEIc9QHooYQj2rgKz+HGSD2pcxxVar1S5aNlU2LFStoNFa
721Ka+abjv7hsILQ5ENUTvLVUBbm8BIJUA7YHxkYrte6813iSPxtgqSmtisHxQOTi3Op3oAnuy4T
fhfv2RWtzMBRjuVm8RRGEZlrkfG+rIMILk8oXVMtgfHVISwEweEufKs+oO6H+QivjU7SJnHEByzR
xpQE5D6CvPJ5rEIUiTZ8XJ2S41oO71D3UFl8XS5iVmOURQTWbYa9IqMeD/oB+PT7kr80spd1pz0l
jobZ0ZESkYN+7ZuRuNh28O2J4g6s2zQU+YmCIsSDXHHNbFezOfejS4zaPGGquVjmYjqURBsNxUWk
XCqvPyTrOGIduVdafbnlxDrq7toIMkMktqoJAn2PraForJZis2iNzYej/lgQJWQYPttC/OPSFki2
hOj0GavERpNjk3+nAqaaW1YjJxhjykNGkeZELNdnb29iaB1yQxf3dvrr+z9+2Vn+5pbsr/Gih7aC
i4D5ZesHFO8iRYSv+8wVAYA95X+Jzww1po5qkHYk8/EyO7rBgbMMBIVNifGJQkqcKNWlVd5R22rw
EU0RviWNdEDR7LjvXwF3YlTneZokoov8GjRDXVsRcr8XJohvv97lyhcY5ZLyTjt09fmm4fjU1l/R
mtAubvxyMthosPXGHq4J7IDXrl0u8s+KbV+4wcJ7WCd/s+W7hnCWjNBEZz9sfPWtkylY4BP8g1tb
6RwqnsWVyE10Ysl1OFhAma4bfZoCLvuvzBQY72Xdzetz3am2KuD5yUNCf0Ga8P6QhTlGPxRgzWXQ
wmB1Qks4+fjIgLlVxTDF36tqmtFQY3bx9HvwDb+e5Q1/VnFR8TbIdzBrV7pUDvxmDfamZt037mpy
FEVBtBfDlcs5jOJpKSD00lLN7WzQw4Hp0GNlqpQKS8UXhAftCq+klb8aQYOUtdDdQmqtxcbh7Tur
CinrGN4FJXPYUmKEqzwiGNFEzJmxjuDJx2Y/R41cYPLyvXytXLNfljIwAuDguTrEU74xn+N7Apbh
DMOHXN7eXa5XGeUdmf36ZXavdSUMaat62wm8AH2xU8rJiA0q0xP7PU+NG25jTY+9o2NreDSuXpyT
fyXCdfxyI4HVZDrckxW00n3M6vjDz1wXrTNp8SO4XpNo1KRdWxuvdCZwBsp5znySdOldb1LVB0KG
iGb9hmlo8kW+AvQmP5Rr3w54GplaKN6yhdE1AD+N2SIHOxjlhZZrHM5YWLBx/vrWfvH8tqPBFjWG
Gulwu8ktgTv9ziZZrKcFiSryclGUNZThTrmgMggLZKc3vbe4OHvlC1W5skb1x9/6VnhT+gCuFWhR
CCqkDQYXqKAjtX5P0oPaav7w5jCgwkUJ+NyoO2N9Bml1rD1A8Y5KGujnIjvem+wOD7oN5aCsVwiS
U6f3lBBsKpBFG+F5ZeRStXzGrvS+QS+xMx90KeOfLGs9Xf1FpnmDHZAHzbi2Q6tF5P3TM7PNAzHr
Lt7gxbDBpfciw14C6k18ZEcM6R6Mun4w5xAQnN2uVpEpeIvdQ50N/PakvkOA4XD36medtJ9saUa8
uSAbBr4VLfbM9TOyHK+UexUMcqcDFrJB4sKDkJfbRnA84gx3bkZOM5TKif/5HhlmHoREMnW2wtHH
o4Xn97WNnMp8/8Jpmp6jHtM2bbct+SaEkVxHBF+M/YsEkYYht0HPscLeBZxFh/XgXTL8eao8IYqy
15YKzRIylR7bNwnUGG2K37mQi+GN0GveTiIwEF7pn0AJyKuTT/jPbgXjU0/wHajFc6mCck6/zw85
pi/RanHtYBxlg/97WRMBiTvpxYz9mRn9Cl3QHGsEWNUOqr9yESzJN8qja6ix6JaXe6GSA21fti/K
Q1BPxeXhIs5Eg8Tc+5hpvU76VHXjSnNHEqZiWGbc7aupLQHUkNgt2Rll5TsPNKgLx6jGgIC1RksS
YHMPD+aQ2TNKODDYbGUJRELWbd8Civ8mUJAYyrrJMQoEQVdr1r7zY+681KPZs9izxPncbMMBYwUW
j24Dl53vpFnysNAFbawgmz8Uz3FZXeuyczauU5zYNYoEsEDwCsEjA9JTcWJyHcE3ijGT7R9A00W8
l79c6ENcfaHyPRQ+l7AAUo2VPyNWWkT1Tk2ckCapBHtVWz6VQiWbavsHg11mNpQ5+BDb6+hLxqEy
5fVhrOV6e4WqtUeL/EDKmpl6Vk22rKCGgbkoQSWNiSf6Q9uOa4OXRuxXcVDu94yaHdCIKkGydEcD
coYcVCTs5Grdk4xL/S/4v3rub+Q7TKTIg11R9MkADRNydOxDQFkQ5RbF/c+FVX0CqNEEEkgkpyLn
HhRf+joJ85AkZycZ3ineiVwVtccA5r8eyyPE4xDbyvmNCbKrZVkh9t2cSWNIjz/0/rUjrr207U+Z
T1TSTP5THzDuQhosfKlCB6fjHbmM8qnExTmdju96+syx0Uhv0xwrpOTAaDw0N1LnF2zQV3UmUwDf
lZkSA8sDbxyVxwfPm3ob8zRD1vgpQDw1VTipjkWP57eQPi169e3G92npj7eLITIJVUXB2ZLvaH/u
1QLl/YT7zkQFyMSPNw+wf9QPFFTKPQnpVe8GGnmA+ZpuMq7xZ8jILLoawZhnXtRUDV2ZMKFxNHkp
8vty01j2mYEP41BJVVZkO3TZNyw7L8UqC32HqvHvbS8sZhSsKQe3XM0/nDsyc6PPuY1+BNBfpng7
rYxrbf3yips11k+D2OVt4lmAUiojzXhxnKkKoN4e82kd+Whr5fgbHbWoDj4fZ2m/sQ+ohkSGgOUL
Ypc6VM2EU/rgIgP+vecoFY47z9IyNN9mNahGUgVZf9G8uayRj8JxZU+6+xygGJVI+EePC+Vn73wa
30f7kW5FRF3ncMH178by1GCOEfp3odFkz299glmqcYk3xQS11kHu09vF6fYGMK+uWiF0mqOS40jj
6CTMlHl1r2yTz4eqmpOnhf37+Z9pwGu50Kn7eKkXN1dCO9fx75KqQXs5HEC4vDEkRnOptwoW5K5d
Vcs2JdpbETq0Mg4wF0zBdZkTkFRXuyQ1YGuvo0D2lsMZ8B2yKSjeTq1SCofJPdFLWiQUuhBKwYvP
BiXgltF5sCyeNQwUwAQJTdXXt4hJ4FyEC4+7CDPOC5ylRWjOxoYYbJI/BdaVHdFj/+8CsFwZuNrb
ENtcpldNVUNAkC9VqLbhQNqL/5Bj4/bAmLRbSw1yxeMEwLSyieHwLvrXxMcancagj7ycrXvL3qPJ
GJoHL9GO0WrJi45Jr+SztYEHuzvXSHhjw1IB4jHTs3grBTYwbyW7z+jy+vFYixLqX398gzucZ8Rm
sRdLljaXWpgxVf9QriBiV0VMJ/vNQrhTvza2oKpIZMfTfAnCinEKpb3GRpjFqa7ReiSUouSWx+8t
ztvCZrumOZT17QHMNavKCRrpEf6K3+fF6AVDhwPVhr6+K8q9D+8S0VA7mRng4AXIb15XIwKS6w83
AGSLnPZCxBpl52+2xcgUlidEoifIIaqTbvWqRRhaT3v71ZXlhrkczBKSEYFRJUytd43gxPauaBrT
GjPvT3CgfOktiwRLRR4a2uN0jSd7+Cjm4GsU+aDFQ6Pd3q8d6rCbN6brlPHx2t0B6c3Wf4iRY2pi
Yu1SVH0KvonA0XeW+D9hFIiQJC/gizNpBSTDJdOc+kTTjZTGwTKSQT4ndIxc3ZnOYbICrOwa4k0h
17bNjo2rumBxkUuSCN0p03a76EC6BxujyTaEQyDH5ww7x0Auc3AZ98t5mF6Es/WVaAf7T5vsVRP/
Ye3BNDzHwxXFWF5hHGy7F2hGAY/TQ49O84Uy1Prz8hUSB8dPtB0G0/s9A6n2en7ardSoVfnyMCdj
WunZrFztxmgnq2qv5wFieZm0b9h4lup6xjyzpEb0YdHdPKqA0Uqkw6ACKMFTJaa47CXy4zr4ZO4Y
w3eZV+gpTsD4KJ/0z7mk0/z9dZYY+Hodb2m6bVxxgrYpUIAbhIg/IrucvFiL6Glfll/yKO3VpFsk
Q57vv/rcvm+S7pATgUU17LpSrWdDhhqXw2iFTvC3WVo4rWWAeLNkFSpuzL64Yq+1dt/Agddmyeei
zciNfb2EVul7IYfrZC78nOTkMbcHL6AkKmPIsk9NRyFViBdu/Ji3u1UIjv29hd/26Qjudewotx8S
92RuwH/Fieud1+TLLFFHPwrHp8aWqVHRN7N9uAG5CiDylrAKCkac/5ZKSVXcaGaHIpKnKHHP1Au6
/8iQhDqgmcegi3UGLeSYzDL7zf7iuMXeEaR3PdjxWa93+VFcQ46mnf5+9w/zY16+i5d1FT3wPthC
BsboUq/HYk43NMozAiKA44M/fY64uRzILblhKWK/AdcifZe65oGM4LVnKRzeCSRJoKFSoYvNEg9b
1KidPM0RQIzNeNP7MS599uT0XDEPVs68hohrDVFttXVV45TdBLnhQAQLaFGPhqEHggu5HUjSt5gx
fTXC6ZtkggzDejLJ4zoKBFNSMR0ooDGkUFuaMmzhMVsORcqVuYtDT9/SuvSdxOiUis7uGJZ/550i
zVwODMM0bR07kkeEbZQLy6sa1BM6nu2KMOvM6NrTRLWGLm7GyTleXCjX11eI45gwwURkiWFKy94t
OuHKJjwe/pDRrvqF9vWZRBvRPmQ2dD86jgDhs5YbGHIPdXq+zUCc3iYKSi2Bea5QjiZkIzy0QXo5
tP6JEXajR/TIxmwlmmBFEvHv1cGQEhvsn1Y8aRJKmy5SRke/6SY3g1al2LS+bX9/I0wCVpBdLIqO
MbKlx5ndRaL4w2KKqFMDmmNxLz4O5lbkLEFePnGna7PFmIcWuXn4v4CFQ2PxKHuwPYb+nA/eyKBD
esMK3JM1sxJXQhH1gLDLuJBmqxmVrr12p+bqV5FOKnY2wWxULPIVGXi7tc4ytMn1a57mlisKEggO
gndgERpEy22o1JKKdsyO4kbv1Tt80g0FUPDtWZ3TAWwQqvyxcOAZdOJMbrvWBVykkU1zfU8lNVW0
iWylGUI34RwWzKE9Bdc7PUeHoEcnL+uzPNpsh+OKHBQNRXR7mKvdWxffDv9UxRethYa5yC8reHTR
hI2+EH7vqZDzf2qgTBaQVkl4VfKxrdRzMNNkwU8nZdENvUBVB4rgbXgw4+wZ6FSMrovalkuhHMGJ
QnmtFYEs4XXiHPex5OIMOc+LcyyLy0apCs5zN1/DNJoKEQCc59k17/kg2p9EScZBL7miSayC9RX5
C4FBiK/hl673deyuqvHfD5VQ0X29LAW7J37Ww2VD7NeTTnfEGjzEbX0zs4VUOp+FPn8rvcoyx5FY
3jSZiugSGdYJBnz8RTjXWjUpq5JqSjn8KkriKG7zmuA2ifNAFLrzyicSd1T5uoGfA4SmooWjNl+m
8fFEGDHLh1CrCcXEIATQmTERSqfsImu60juko+3N2+mAOfGix9brjaMXD8OI9IBFRsAFAdAZ84WG
d3CMPme7wblw9Hq3po2kEhrg2BMZC/WZYzW5LtSKhXApk2kE+4QN2OXsXCGXqI3WfzWcEPBbQ3b/
mrD0anxaQfFmh8tAgq+n2X4Zu3zTXRVqf1lmK1w3JExyhdYhdK/HaULvprgilLEyDmb0h0wawBWl
sHo9xQNjjZIDkl1eElos0tjGCpXBcAliFlo3wdQw3w3Uai/I5RRtCuyyUjHwz2Kvj+7Sg+nFypNj
z60P1bVEbeZuJubQpkJIYsfGWzjSo7gg6+d51MdO2hnp3+Jhzr1EmOmMA9VJhRT7u1RKgiS8/Bj4
wra2g8WiRoZhy0RBO7ome3GDyipoh6N5LD4SymoJgWfkmN9/h1g7KJpoBHeoYvdiXOk+8KDeXzb/
9MYCqKmyl9QRiqnEThrRWSPVaa7g/09PEcz7zaE1DGxReD7emMefY4ZZ3TlmISbDJYMWK0m+IQuS
5T0H+kEEWqjTeukX59nH0w8sv88zJKM2DzK2F3L0Xx2dX6T4okDKuRuhdrqCAg9F/cT/6ziBrKtQ
QpK0PN/CWe644XE3r3uuay03yLwyVj4z2JY1y4XHzzghf541P1j9NuM1dpZQnP7QvarXgr9COiad
8M6sIn09eb8qOTK3J2MCu6WK6uME+7Kwe2Dso3srX4jtbfSmIDNXpGtMsoMkvfIhErYLQR5HNJnh
2q5m5vQlAsZ1Y5vL29RUZzV4ZOVnYjISWI+6hLIt0Kg9dZzOJRkgJ4mbi3L64GKfD2i9M+AsXutP
ik3WAIeb+ABtG3+S9cQ1OXauZzaaNJ0OY71jXGmgkyYHhThblM1Nqd/HR40tAKGd0OII2Y0ohe9O
hxhI6lC7MLqKhL3/dAvNrWCPo0PolvMHiZ9Ck936lKPvL8cO5N3XlEA6bcZsm9cOUjbiybtfyth8
O6qpv4QfjBfW09bCEwG7ECczn9nZtV5a9roVfz/yc+8EzFityqWniroaczDFuRjL3gEJ696GJNQM
5PgZF+IFoGpFPTbyPETL3m4b5Yq7poO9aEIklzsZDDX+FzUs9bCOln5tk/PfyDamMG1icSRMOBoB
lyhH/98Vx9aH5IzYznijVW/Unwehhr1Ex9Gs6XWQISNY13q2C7DQuAT/bNj5TvorMG2BWMMjDEck
Ugl/B/TDNU3gcgWTCQL0bNhTg3raaav9LuiNC0KqoBXhmhB4oY2lGTJemjCi2IIVcqu6u/ylIuFC
LZoe6Lkhx5MHXqBc30oqROk9ZDzUBkHa8NicaN3O1usi7aG47ffEgduIqYzdnwsXNXJlW83q6QnE
cDx2LZFy8mILYY1h+Lg8QCtrpTkZjHtkrjTQSpaDUnWzqxReUfNPy8rWZjlRl3aHo4NKUCZ1pKsI
6ztMHRvKmK1qG7j0y9yD+voqKkK0cJ2X19JpMdASpjrUGm7jdyOw8uZ72o/arfichjmjRLVXyw1t
79BxaH8B2kL7HBC6h2FgI6o726L5hx5JLD2VoA==
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
wOPAGX/3n6PtrF5KQ4vyv+Sx8F5mt0HMeVpUOSWWGnR5Ny8gHhwozJ5vwUrijfui6wYzBlxAuaeK
EZv7rBgW4PfnBGRYlBHgfyjYxc4MgRLqwxyv6tkL0AbTRHnriGu/b5AYoO5BZhgS+HvrIxFlGQmN
hpqBy4cB0afpXNHqRLRAk8y2jwo3fgBPZbBSDfzp1lk8BjAWta2JoEICMu+RqYUBAoj0bP+NwC/A
5jv2tbt55gaM1Of+hRsVFEtgG/9hNlq7VQGb663wWMZaN+PtRkM+P/jcz6gggH7PYJXNfVtezHWO
yFguA3fvY1ol81HQLVIAinbPwtLdmDd/xXVX4A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 7040)
or0Yu5F765iW1LZ6fhpmystIu/5zk8qR2bUn5UrnIcf6nlgfBwCLPHhVWINDsHB7+7nDDF/2graT
5N02XVAGZMUxrwDUy5hjbJs274+kRwNDfY4ZfcMmT4/9mgZX9i0XOwQ7cESaHgMCD0EzRDAnhBpM
M0s/Yf55tUZvCGTBn6SvxRFW08eVKLzNocAursY7QxkbMqjAx7V3hRoqe+3laZqWXBo1cEdrcYbi
N2eKIR+9CvQ8JOQObzDNSf9ae0Yr+LPsFKu2P6gLp/ikCmkyGyaC3eRwLTZQ1+rM8sFNaZ326/Re
e9ACkaHx5Te2w5OzIE7twPnAIzBW9yQ4WEmHm5lE6IwsY+/D2VQJVG0rCkW7cm5jzlyHPSOifKng
oTO3QhLZ6LWE9sRkSymMhFONk5QEOC0Xgjw/G8X9Sv44WzmB/Rse0FwvLigDNuIf+E+Tbn32IpQS
eaoo4cl58S1YdZOKXrgQiMZDDNrcBAZv22AE0t1yfnSukM09ns0WvFDoPriTEguae0MCdg0Ro8c2
3O/ANyhPcBVVdDJ49Iev0gvkeUskQa+mZLZife1Wrk559sw8TCpihFKl8VSDDrlVH+0yIAW9H67C
0gqBGXUd844RYce16DzZhTYkzRXOEms1rIF/VF8odIfFahQgdb5I5rLDBBf8sn7L1VcmUiMN2q/6
QvDzzQt5jiTSwIZHioOquj0PaL7xzwar1Ui5K+/mswyTZQd/g3BMg56VN+ZPsDN+GQr3VWo63iwX
19eJXpzpAAeDEu8K1jn4toYdMq/ODLSyL1j7l0M08s9L534j2aXmOH4I6lPlaLRg40nGlnifvgWR
8hoNiXSY9dvuv8hobyoytrrJZ+2ESYtUFXgh6pmNIz2kAEbWe6YdgM9Wmn9BZDxAN4sPhMOz5XNC
8fXWSwt86VBDMTJn3hNJ05e63yNwI2JCwquTIr/TiUbhr+/FqG0eoZsxBXvZavv+A2lN3wdEmBl4
7oNBn7fEjFdBkDa4pcWrewW7ZouS/gnkT/KUa1pvTOM1RDkzPiGk7prdKOnxxzwWbxNrSrqTNLmO
mSJmA4koc6/eJz614m+RPNj0ibw/dkcljaEmdc7Uby27rAlR7TqSsHNVSkbsKStRaxC20boEZVl5
Unt6rLD51nkGr0kdypAO2AkGB5jzNg3EMfU/6UVAyPM3HljL+e5i3X6O7cDb2damU1YFYGaKyyJV
DeLJYzO2ywZPp4j8RYYfAMp7XNoZfHcT7ZHrmdjK7FuU/MYZGn+R79P9ZsS9R+qGgYRQQb95UdDx
ChNrbhvCiGrJf4Xy77ZBfkiGs6NM0thsXdz1gDJ/4Ptt/9Wjl4WYZBhSn0LXg3wU7l08Y6+vtJbh
o1Y28nuPU6CKzBuNl2tUNG2M+PhLJknsLmk2TlVY5Y2/+aF4nJud3VkpgxXDqaDDqwid21ZpIfK2
Qra6ZXXNv+/+SpIbRst7DhUzfz8WUerQL3j3tGzaWhPV+nIwHDdEDc8chQVLOzd1RwhUes7a6zVw
ezh+nCepJV+hmz9K1jBK9s39px8p9Z5EY+m2sfJbDYQcDSQB+Ds4qeEVsP/DPrhw6LL1Te+2TVUH
ACs9sUUldjSxOwVYFzn1xypoYH+uv8TQ/ZDdvPOihmHU2GpYJ+ErXapAPnXbBJeikbBjrl+i4szp
UFbm62nMF9lo2cVIK99tXNVIr1HYqKw8nGvKRSbvS5gjELmbZU+U09BMm7sb4qdyEyJ9oqpPKsZn
0V5q/urpUdERfwKls4Iihqd2jI6feF2YP6expyhp2kdm+IoVUr2WoeSTCauLGvt5cW8uRdnfauw1
gJjrhpxnEm2JHQN4WSAFgLIZO/c1Jna6PIx6GfX00l3OPEHGwb6y2QmhG6fhP38luwKzimn2wPdu
7UNBwAx2c35K+W3/OyL+Kx86C2BGO237uYOexdkI6/eTV9XJRp+3I/RXD7RmbPkAnrDK3tThVNv5
SL1+2gVrUrq+osds72XQFgGddHYqxGR6sWmDRKv9GfgF+fwDE4htqGDPnYdhJUWyCetwLYuBCqCs
ywrBsFKHYktr5hl4gUwdG8l+acl2m10PCjWAyIBTIXQPbgSJ0e7ZGN027nH6TQz5LJkgu7dJpPrO
tOK79BPEv8idSqngsscjRocL+wiKM0uFap/hQ36A+YJkdxA2Y12pOwbEJeG8JPD5U2LC3jeyS9Gc
5RKoAD9u5Biu+GFqnY11az6zS0zUTJQlDbn0eoQmESvCmnqOcajifVAxIovCAJhXvEe0ehOipagB
mBZdHDVPm+xxoAS2VcuuULT3qKTFj/1d6XIJDWtsDfJE8KEFQid6vcAiiHwGIZd5vgZPJbWEJ5O5
OP+ihlg+k67GSfBMN9NQhcLR8vKKFnp4fWwvcPvuf1eyccXzZWGqhSgdJ0Vqjp19v/6RrMzrQ3IT
+htnW5BXMamxVmvPufp1bf7jF2B2VSNJEQEvtyGZ5N1mxycXioOR/ze/6ahlPzi24WG1Jq0O1fZ5
MzJYJyrhK7BP39jNs1x2Rt4s7ocuXpxtpAMOsIP69gKPIravbWuriq4XPVXaxjc6ZgCAksIZj3XJ
TkMz6leQGpvo8Rh8zdN7+t+bUJzGf30Bt3vEAtlFQKS6ya/tJu4sA2yN6jzVjadEMZVE2aPm5nsp
QqhYL8WWJcwSbfY5Ykl4xP2jY9KG4mjBw8fhz8PTdUEu6lL7NBkGmemJ30WJp9L6cKVF7JvvAka4
wbDpE2jRSInSYPGS88uF81QPtIdv1ZYp0NrApNglGz43lj16ELiN8mrElKFEkkd+H59R2sRN90ve
Gn5xI2ecG9sIAcpSRlGs4VaE9op9URLMZfgW30ZGtNeQyjOnZq3wUf1ntlxWf69as+gjbJlnk2a2
GD2fmDPqN3kBjZ8CfIiGU2XPkQZlnOISSgK/2Z61WVXhyz6lQ9K9nO8JT+HRJ7rlQcXbC7zkjX3T
ItKWJ5PTszSzXLF7v8qvFmXeym65U1b8W8maRhyxAWYwZRYfpo42+A5Jfx1vIFmcz0noiwNT/1A1
+SMueItXhE6GEsaCfF14pY65tMdFHt2GZ4L/wUo8ZYpyrLejk/M4cETOqqtsQ7JFvc2ezoZaTpqn
svkrv/qSI8vE02vnlYHyc2umxEG308/ZXOiLd2SC3azWDTil3kzRvhK6h2hpuWHTOkCc+gJv6oSS
gBIWSN3KjuhjVldvwBxWKeAlWS1puiFFZvsxtYZyTFhVQmaFhK8JCQdTP+Hz+ActwmE5bCBgnvRN
v+yov9j6/jZV6PjLfDukssnArNzy2TzNFXH8CKDLd1YuIZJHFfwgmz6AmEQPpRrnNMqL5HybnLVS
MdId+eVhXGZHJ9cXFB+zylKyEikFn2mZbQrIP/Q2pqA2ECgO4sI81HRHun5tcaAA7qAaQDs5YUDA
/pEUPHR81BF6XmKVmgc9ETl/wQ6nFsGvluEy8ITNR2kaPi8VHF43hC78wQiPuynXLto0wsQqrFuh
GThQYyZohiEovM9NXnBTPQf0xUuas1t9JIjufqLmikJtwdItQ3EtuyDGqwKFz8ja2H9OSmInWrgd
5PsoNj4Fm9rl/KZ1gvqZU+PUVSNZLpeIXa+0GLysHgZnZXNytl8D+gRfdjJfaFtvE4hvGBt1bo+9
8MmbcfqYtkH8JRqzd3Kv6zGNUXQTdxI5YvU62CsNM9fw53vk+LVM33FBitvL5e0nPPsUW+DgeywI
+cGAMhOcD8kIzxejKnfNOh4syC2viQKdAx9Z47l17lyN41J8DfLyEGFsvLFWvwlvs7+1Repa0JZ5
ip6ckz5iIqiAQLAHhrow4oT6By6hVwtR2UCuAX2iWUpxU3Dnx43Ni+s/4KsDYH8nqjd7FlGWEHgO
5QdDm2TeOENe/wd+T/PF5NW+fq7HArYxQfo5mdonzuvvst70TWEQ9avGwpKzU7dkg0UZcUhjjBO7
dF+TshwoU90z1GK/nkudxBh048qRJOHM39oM2dDQAIKxPEdLgpL/OpB1SzlmwIQCaqwS4ouuAJOt
k74a3J6fRfbSVwFbuNkuScllN4+rcrPMUK+kLMfBpHaV7BjqJFz1uOkJz16223232Bwv/4qe2ynz
blIodJonNWL7deLXNGNPaSOtTzLMctfs/pn5BzoClERnSLNqhNON+xwSg10JbQWZ0Bdedp5vMKkL
Gd4L0hdAfNzCw1ylDpuxwokpXDttVTBf+y+npVEWLj70FBs7gCFyeAZD0CMJ09a5vkUChtoKPy59
Tc+LRlGIxrsPZSAF0ia7XwahFlMLNGzRd5aXcImjAo8UR2WjBa+WJvfpmRBzFfADWECOxYywfFfr
hzdh80TmGH+lwfvWWUZVEvMZEf8+6nG7MuXcsaRfaE0wJxBxbr3vLb+CFUcyAAGWvpb6ica+ga7d
VgWT8+zbw3UOHlSxwwN6uuLXkyc6mm1K2x3MskRrMcu8iQoJFWtw/PB2tUn2/WLoYMtChG8z085t
y2oYWAEqIdIIReo/5y95SJUKhxVzjSCtlKdjq3PFhePsLZsGG9xd0httIiBVm2HB4AzBjJJ32FaK
vvDmdPxPzSsbgN+Eaauj0V9a55aKPi53IiqhOEtWHRcJ2n1J1X7GucvXHRZBwiiUT9cvSeDeReBa
FJr+yuGsy5nfTaz9zyuBlZePjB83sCg6UA3pm10/o09Kz+cPN8nvQhnLXmIsZpbVGthYUJbUxAzH
gtjuQIm3bJC+sMgPg4VICzNOfMfng1QGsuLY14D8Yu3s28F36a+hA+rWT85pE5S7hLeDgdFsYqzx
9xN4da0a8azh7JZdc34n8wglOxStNvfh5Q1CdhVFh3rdfD2Nlg4IpAGZXdK/7x0wJNRo+ilNaar6
AnXW+NB5zvbauVywf0opouT5LSo34be7sk8QT4OLEXkVbBbYIyGGr7YSm9s8NUITBxAKiXu7YVTm
MzZaDEb+9dbJetPEjgGCJ3+bthaG+5I9/jxfPHOc2Oi/eTIYCDTZ4+RGntcwz5tHCF/upno5eqij
nx9BrcieCpg2Y9ZRawAAygU8foYvbBCmO+vuQfVyBLYkGDW4LaiLweROVAVd5/lNHxHxveVmUFqZ
iynqgC/tCD+6gtM6M4b+uv7SoaX5xDvk3bUKUFc3Y8UroqWpdGv8ZeWY6OXUhovA0LkXCWW75Pg0
Fu1XJMQKR5EZ6R+dYTo5WncUvVnimwblEqzXkThaD3MzrRPXg+O7Wasjxdhk0N8iZjQQiDA6r7bY
0ah2fKa3CuQ8u9VycaJuzqUW0n6GnXoXxLyekyP7iQebUBo6lWmqSVZ+Q6tUfnTrqcwYj/CzblJw
nkSrAfhK9KkfrgGs8crTZEzEd6uR7kHeReaNLFYbAi+UZ5k4eJCNzVgMo16GVQb6ozBhuaEF57Y4
dOgArFYPCRB+S7GMrYamJ4dOX4grqDsyQmc0a31CadH71Qme3IsexhKWibAbQbc7JytOm2jQoyjm
egNQ+u0Yh/5LI9On2xlTUBmpv0yuS5pJRKgkj79IoCqrdCLce2zReL6VmZ/pkr7eDoAMaJd/O9kw
xGKVko4YTQ/eLezds5MD6edBoOcisz0k7vD7t+IeN+MFlMPHOlkGJaQRqeL/zypwm3mYJfln7U3p
0B7UmzMFRlprIiOePlcZbYnj72BMJlARV9dXbQpV1TzpWwBV7FJIyLcd+FXttec2TZYRIYJTJcQt
+laJCUX8ft7BuAp7pI7tVFpdzIao3yskQWToVPlrnimPfZnJA33D8PJMd91gECbE6mUeJbLh9+1G
n7aijKtqPoZICqS5bP6PeiAM4VxjpocUyOHC4OPYr332LiLDSgURrOZ/UIftQ6RCz98TAjuHmNH6
wy/6c2cbqXrcS+iU07vn8wn14iMolEbKmmdVEDiDkOS+M4FDzh+AG6ia8cTkcLK4zl+ukR95k/2L
xIHMob61gJDT49ETgKB6uV1Q5tJqe4YGnGCZB1jXuARbIfB+NdqJr0MKkY68V8mcSGWoAfDmQyf9
IrNEYqyQN8aocHLBXCVyhI9iyvgEqeul7ctxtDLCPwRz5+KCEN8ReIg6+AzOvJN0LvGYZfJnF6mf
uVL22+cMCyxRI0WQq6pFYTX7zY9EWtx5pvIZLmQcXa8dseSGcqPttQv2LHrG6lz9NoCJ7zZprJLY
UR3yf5jC6o0OzRlfMNREGE7jxN7kCXe8OYFsGmv5SIXwiA5QrtNxdawURk5ewpyRNDPQdgyPNgEN
XI0SU5BQtSv9OnIW7F967cjxgpuezfUwaCGQ2zRpg9xmgkGXVcqkTELLW8ra/uZh+2hCHAkMRuEH
T6SXeAYYDUSDbFTRxdb6GEUD95rWV7iTWXX0q/9//tgMvK8HAeIZmPB0QO+sFAzwdn2yvYheuuB7
Xmi7STTCloLKLIecJOW3Bzlf4Qts+qKv6zEbo4EN8U3oXVRJ9Ydqi3Y4aSJO29CnuiiU8B4a0gud
oc1kAdgP+ZnCuA42sie7Gl20mDbAd/PJzqa67Nn2YEgE6VQ/QzaXaWVFntzqxJZGLxNpemuRmEQl
5SpuCeRgVvrSSUHMbRzmarghUSDSzGAlWtDezkZZGr2dk2KbXOWKzoiLTZ8Qw2DgIl5Emsiy+ZMW
F9puqcE25tzKMZmJRMQbsz4OyaawBzA7CemnSvfVyuavEWWslbq+hJRLtYoZ0/6O0j4ImEvI+w0P
WDK+A2JcjJWrdT8J5y5r2+BovPXjOhn4AITUbTvH1KLYiXzhzM4KJ6196NII7womVGB6ME6LYsJS
nzi6NwvAA6Ewk2nobnKZ8hM4j+gNk5WHOG+09z2I+AR5GWLOmZNtnLe4xx7CaXB0n7eNmgFfwnL4
xp2rPy8imqurOJHUt9gnBQj+bO6sHildXj3Hbnd82itVt2V4FdRFXwspxZhnEq9FN2nATDUis6u6
/FQJ+6cped+Ca/6W4YoE98iXTv06SZkHH0T3ki26kRQOTEoxuyR3caGV/+vd5maQaf2FlnPq6RMc
KbqD3Hdu0EQegPXdQMXvCS1zvFm5zHgbv6TrOOpsGOKLD+ovN/FV8rAU3WW/rHstmGJCnQbN8UFU
TBpNQ5fjBsUGswb5No5lAUAV6z7+ljFtWc/f70i/1QNjUd/DXY3TBtaAKAE94wmwVDsO0V4Li7On
9RWeHd6KLNOk4cBPVnn6ABccXAb/f5A6IWauEdiuhPd1MOAAXGQbjRf7JtlrIhBSGUufqk46ZXWm
yf6G7tpdUL5PnDgpBm1X0Eea1QRlxi/30GgL9SRg2bPwwz83qFlsBTlroV9g2AHxOfKk7TIqicXR
n4EsdvTvGET8qeUwrs7Kxly5bOacDqUGDneUwO86YM4o8SDRiu4nY937ZnEh/DudhYnwljP40ft+
eoSbuCiiLORv6JPga+bMaToNz6TX6nkq4BuxFKQv6RQdhjBwVohECj2whvOlL0kJywXH0JXQs21T
GNhRfU8sVn3AeTuKVG68F1Zcf6chtdqMiHb+cNvxSCQkoiaPhVoB3Oog2F2s6Wls2doRG699IsoQ
YlO4DH7EAcr8/9kW5xSKnPN9kem8z8524TJx2VYRtTKlQijTv2UG317c3cRAG75O+NO4zzC31Lgn
0YvHWY393XwVCa6jp9iwDnNbbio+RkKbxuKcZjEQj4+W8UJCYeAztLbxbRWKkAp+qhHLnrx8P0lG
uSsqzU8B7wH7fuDm1bbJ9XSyY7syOr1c9EKQ3SvwuiMVOxdYJ2MYE7H4c7nSTmF495ijCFLHAOpq
kcBLfVsJ2KmkGZ5jPF/yAOWtco3KAeDjxjQq99EQjjr4x2BvlEjxxWbaj6jgs+ZIb8W9ioK5YPRt
f/5If1WE1CE9C5Ok7bedSsfbcvxZAkefJkXGHoUvuPkbpE5i9RNX8Ws5F6T/plxAjtc4FzFJD8HW
AkHDEuU8l0+rxg4PPEmDhUoPpZTofQq7H17Xe0BRGeObPnp0UJhxrqBMYK5bNzxB4i2qN3jBT3le
pK4FLRwfq9B1Fiyocd5OEjP1asWobjMDBa+YqYWXcxuw+48aL9z6DoTL+lzA4LSg7ayKcbcE/UzJ
P3AhiYfiK8op5icgZVPUmb2AgRdL7kwLkwh3HfSirtn6QcKE7eWMpu71lv3CpPut8wQCrQOsHoPV
vO/ay86NtrbthQ+Az1bVqq1yW59awtEg9HFX8DvqXLfbGzpE0pkRHSrUzOezddX/nU7Lb7f5W0Iq
yowUUU0U6G5+IvuQRwi1cLTiYHCWB7pk3BCxRsJnjgKt2ppVsIYBugiauxmre8wnBwaYY+ybSUpM
gM8vhglH9z6i8KRUF+nHNykfE5VgSSwn1OxB9nAcDemfue5xqjGTgnQEiNZ4CBSOoFbE9sACTtkX
DU1yIzqIXGq6457ckkzLBVdSi4uLss2Yu/KLA3D0PW+hN25osBrDWuFAXjBX1jZxXY2wijydUyNu
woJ+91PX1/cASUPotcNAgfNxHOOWvebYFEa7yS9t+ZeOK8la7Ube3SA9c2nQS98oaNOKwpafWR0m
1cEdYulQJC2ESMqa2lAP1TLJDchgzFw1hVc8Jj2bSKUmKOU8h81MxaHgcscRebCmr7i3SIA8WtZD
cXoWa6OBKrkXBdLxdujvNNONQ3dn0VcpVe0vC9xhCT5o9SPU12DfC3rczDh0bSAYh6ILy1RWr3yr
x8Cm3mEdh6pi8tvxMmsyR4FSjAlwRf04wA/aEaCnup0XYXAKmA+z9Ao6rA9dOuImZfTW50xr300Y
ZLygYlxWRZKrV+1ILNCMoJGGnvnNC+J9Y8AuZlLX4tIuoTdfJswy/pGmqHeOA90UH5YTrCfLtkCv
fg4tM/7s8ii6LKBuzVZMPOplA9r/x2l9+BJE4jxF1WSpeNltWl5aFoqE73HM8TjPAOd0byRrAJJk
Xlt+YuFFYU63JWjBQBO6vQre80VAXohdLryJoKmx3iJKCxiFsGkFVcJsxqNXe0pugYdWKAQ8NAFk
CllPL7Ul9/fr5E9biahxADAxl5CoMJipLPi5G7bsRuG3Njc++oW1gcsc2UqEdKMXSxb/3QQStKvL
zYOSGvqeuQZcXL9j/CZssgB1wxNpJm0hy0XwnxihGnn8sN/ijWwhs2muyvmT5iJebVEvqSBzRimI
GaBHV2uaVzAJLoBN9otmDORgVlvvDtL8OSkrCddMANyLI+OA9IVbnqsgm6r2g+OLn34wqQvRZ/KP
SqvBJqU0NOxOjuA6p/39DQkMA1CnjynDrj2r0TcvNvzMbmm5iIPcBdyj5aQ42OKi8RWIDCVlPAyk
OiFQ+7vMA5hM5KSca4QCceJaL2xt0TpZLylJvXKxyzbStnKaBr+JzlbVVIW5NXsyGWiGCMWzmS9H
gGHWmU3piUjyVu4tfe3bH5phZV/PnHWUVmhrKRQ=
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
zFOMR4ErT3GxQu16/UyHW5WUaMNQw13zKu/74115k2dLV2MnU6scTudVqWcPUtCirN38Yo3qEeIM
MzPb49c2YrfYIrp2RGjTo2O5tkSbbklrM/pvHco/9MG5GhoJJHUduiLzKmKgkHdbl+Cwtvj4gUKC
cTAE6vlN7J2Khy6gvWfnLz04TR/Ws1ldeQDBWEh1m2VDCLl+mOgQDA1u5gxImCy5QVrEFycfHhRy
i9jOaLWCMaifENQqkoI3Kb1JyUQFEC81qOwJ+NKrKkupj7NAnOUIvqQXxuE6Z1yOpmHYFlncQK+y
cIkd0jp2rcFf4mNuf8OcLNa5gyWb2uFBZ8sVaQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 10784)
QRQetL/xvU0ePlYWHBpPuz8aKAI/1xJdbhB4XKs6iWMwhceDuYlbQDW3xIrZGl6XC1s5R9lLr8M8
XEi8OtKXueHHxWDMgP/59DfwAPMcEvM7/ox5BrGrt0ZyiD/OFoqVx0vHcJ/AxICIO3G+SahpTmNk
WCDB9Nf/oFF+hOo12lYc1ViUv6Tcq6fcQSAxkd2lY0WXp8tRG3I43a75YL4hyJ3sF31D7mF0Sk6p
OVMvd2KFvQ0nX6VXw5NteTVvT34bTl19Bax6WrhuVMjthfCF4TW9rQnzWKM8qnlzXz20s59raedS
cRzAYz49mup7ONcelUUE3Z0p012sJ5sDOST5ZtOgQJZBA7qFRiSft8i2M391gueTdazI9nt9ZtDT
aVvDf8NWg17dibsHOGTFNBnoJZd6BHW08b7IegMVbuwMILkX3PmE7pTltVsVe4Ov+z07hRd0Pfz2
h5cFQBdxqTuuQtZwMtm8v/eVOJz0bx7cAPxHFCw0dQB/LSEDJ8gsgF5473T/C9ThmK6VIhgpV92K
nT/Xj0q3cWhBZDjPZXph4zCNrNDraCNPCLxGlV/9U0iEaNZjHNMD8jDO7vVFzX6+HDj7twlCmqtD
wzuMu1KMCi6yEgGUsjuLVdwzaQzMM8n1V07sdVbzKq+/fk5q79El1++XZ67HdW0BgH2Vg2skDbwY
s/jLXfgXadxbJ8beZn9phX3v9Rjix4h7TyUDtXtc7cEctd5bqZ9/68UrIxbn78dJCrj8+A3ogST7
fMG8f2cSBSRmpu3XTXmAUb5mxrh1DlMUO5aCt6mEdWhqxR143AgmgTU0eLO9niGKQzA84svx1OiS
PRY+r1+2w5+YX/lvs3AaYuFYuM8mYKV+3amm44SkvYqpbw+lwzr26BUJrai8Nry4aocyQpJgO4Uv
W1xvykt2nJ/opXxtah8vszGXseVZTw42vok2QvK9VljZpnpDxGOVILfBHU7dE00fxGzs5si+h3+Z
EF7hMoZxw4lJm6LcSbbRb3jC+MxwffQ1Tzsb5J2tljSyfVWXVfK/yn34TVg5jk8ZhRG2ooQTejHo
IlknvcTMEfTUDXjlno32ulv/M8VaY9OPZlZ6e22mmbN9Uejp3uF7XY/2qFZJYKeAQRNVCDk35Ct2
CXkDs88Qs7NGhvNiEEsPPgTGN+6U/6e88OXAHTPY2DPmieOEw8Gc21HLdrsH5SnoAM2f8695S06J
QylyW8ZsryMlIrr+ewgldKILLTJptBPilT6gJ054vwIsdVJdwqgVj0EPiiXLQ7YvmFdp65Oh7Wy9
AE2Tp97oMO99duCJ8EIRQFa0Lus1MRkhVZzT8eYR2RjEDieBg2neDbfs1b/FbUrwlfmdK2Q0S64+
QoMKZOmaWXXEBF34+/qUSq97QAB5N+/tNFkv0s+CNHyrKEDyFRWCndvFD1UnSoVKArPTC6RNyfsQ
+AHkKsSqXxlvWKZIH7RNOcrELHgtzYto3DmhDZQ2/9Lp3suZ79Ynw4jLBrt7rSCk/FLvJxyKveMi
Z7epeyftfiaqIvYZQe3ZvqSpUcN0G1NSFRbQguopWVoCfWgbkBVEvgEeBcjeBMQ9TgzTzHJ72aRM
Sr8C9/Kfp0z7zLppYd4w19JBNILdIhOaQbXwfKzamXK9rbmMZ8VBwYC+Fst4lNWgt5J+kNhZxxNZ
kC3qxUzeLwziNUVky/hjDt1eQ9BwSaWwLlKJAfsvM6OjSt2w11bLk4WYilXoUtwufr3xf+t0V8fs
+mpIG1qoZhV22QlZ32IQ5Hk7i6RyZe2Mf/Y9ERbShNv6HvTGCtS1l7h3uedmQTNpThWFN1TJ+GnX
uuhxCVdCNI16d0lgZzhHr2Cw3io2AigoF16WVI6aP+5NZyl5LTsIlp5C/zBWkcmjdexq3S0Txg8k
JUWC6xYWF85ck9kdAf8sOxeBV93ne2KbShHxWm7KsYCs+8caLpdjZwI5IXwZehDpIkuEbXJzxHMQ
GLAmlEJ72ouBYKVkM5hbXgxx8IPl2bHnbFrDZdiHZ6Cdnd8ZayCW8TtAHRHYENOeoOIEtjEkOuA9
5tJCxluFqnZgNFi+ZBqC8dxsXQgqSYH26g45FlyZJE8Tk80Lt7NTuulYZbaisgE7h5lAA40ywBXq
zvjXSkFhdimHRgTD9RFktUmycpT2k2VYcbkaIhT69XxUJNtQ20mRvDegPXcjmQODKGnLj6Ypr9zd
L8EzMrBd4yPxeIMHC1WUt9FIVHloyGH/hEDxaxuOa7wgx8arQT2z4u1X4xvap2fhBEKgGBUQsbt5
UOBvkhouJtQjqWoiA8McMNgJfOYF1g/3ysJ5vrp/SE+g1Dpxc5cAfILuIktsl2tefaMCPQI8bMoT
fMYWJ7b+spApA/Y8OEaYrfVJd5JVcvr/RL3HsKpcziT1i7jpiLs+QK9FPexE6rrOUFXCI15rnJHg
OGpA1EnvomPLvmb7vipj8AsQwDz6a5bt2v1snJ9SyFq7Z5+IYgSTZrXj5HLJdD/PeGmEU/5O1zyz
1zrQiIiAa2OWDDLI3lk/eetKeE2mQbQBgdeNhWTE5ScjRhoSml+33nTFpw2C72M66wAxrYOLFOpE
KIExAJxHtbwbQHY9BhXc3a9YvNNnZv16RGgi8dVVC3wXSuUfuA6y0sIKkeRL4DsLezl6pF1hrBIm
hfKb7UeZOsSMYpY/iccXbtrVOEa25pvyZQFIUkB4JVYcMGkwp3RAMjnZh7K0iqkuDxJwdadWtayr
Hg9nzZCKDRoG8dRoE4ngZacV7y4upXlqEdC87wqdixbiACDmDGiHY1z70iU+V2FeHq6Gzv5HU1i5
Rsz3W5MXeZDLTCd0PoeBx2pxjVwOUttL3IiDAjmFHMdFOwJBxjteOsaH8ya5lrtvwc7gg72aGuAY
pGwOA2vYT/c4D4vmkrej1e5v4Bp0/0JzCSNeMcmyAR1LO/3y+7TKZbetdMfWnpbT48klBgtZwp6j
7RbOAPixT/NqSA/L7M/g3dsldVRg+U6PrwPeJ527sb/Xi1W3BnI17eXiWLTto9w5jKyr64SO12PQ
pN16cviis5kD4WeQcJuU7ND0CH8/++tkFehzz5CYFoAvDsXJo8EloeYYziWaY5Fx1eZJM+isVmts
4ZMaPVkcd4bRWKZdH9ZGmbc9gu3VYEXD3OzfEVwx+2tqQbcAsAEPl3rTbq/+s8QVOdsBDunX3B79
1YXrDnUWfDGqEPB1AYq1NiKfpaS0XLoHyqVjFJ/QCXYw9m3smpCAcUNmhLQs/r8yRT6kzjWxrT4l
HNYh/dar9xAfc871FuksHDZmHLLT2XnD7/iUBYYNUUoU0GR9yw6SeStW6gborsMi4CYdjxsMIgq4
9eec8AUrCU9gWw0kKKkkmjg5628HJrqqGwSgdnzu1tFPFFlm/jLbr6esZD8VjvNDFPYOVbeidrUk
V/b/WBKIwAL9rE1+N0FdWxy6F5jHckkj3+ZHUH7zoCVFrcaBAhIE2Qw+dwN2jO0EwfnAFqokn4pi
Etl9HKfya4fskjsAhrKnkMUN9DTKm1dv5d+3BpEXCbuzvFMEYFQ0rousDEhu+OP1RgydfsNs1mIJ
qtjgbHiB5ujBfMxJx+lb/y8APzpnyeSc+GfOyxfSt/mkTl7R7RSPWtNlWik0Ouk7WzwTotIkB5RJ
HAZHbASV4TutRFMRDF+PrDlrSKILoP8bfK/ItLVNEzsR0nUG+Qn5qKfJrELvPAggVGCmMXzHjS2y
4fwpXvn92NgYB5bVjJHI4ZKBnifjl5pqPd978M2Divl+lnPJ/p8XD7qZildbmeCQv2qTla0bQCE7
QtbpSoIGZSIovPgTLUMTIxh6rD0ZrsHxZn/Zw2fYSJknpJF4aOk2BrHy1UG4XWAp4D/s2mM/HF6K
RooQWUa6ZApYwSyfAkbg/Pn3eqpuhdYGtigoET/CXIdgKlZCSidGF5a1oWbXUkfkDRJK4AgMHJHp
B6IgaY/cx3vK4n4WTkqoa5UmtT99B8RQAV+15yDq+SHZ/9tfihwZ0ehJ6KnR1KSopSVP3DGPJ5Tr
XgZLyIb9ni1ym30weBdqwEeu0X8MgUP2iswxvnWVDvIa7gjCKlMEIEarlGsuXhvs9fHkczIuEMgm
rq9nrtSFG1KUnkJuiLA6Wi2zjIyaDi3jWdGOrQD4wZVvKeOt5zb7elAEvFk2b8W/lOr83mYNQTyp
OSZ3CTrX16+7lg9UUATItncSaaJoUSsvd13+4wD/MWAFf4S5MOLd2ddLxgoIpjmklg7R/TjEOjoa
4p+3Jza1kBGJVypU9DHMxdkyfD+f+2qmjkpGg1ELiXhtWewL4Ckl2+HQx1iu8UtBCBlnu2xzxZHl
IBGweO9dhz8EAtScA6V3JfV03jAiRDVDsn1NhrF84DFztJwSxJRjGFFp5a1BRqZp5/xRFdXeiIKR
szihh9Kv4BvkW4eFNB0TIgpLAnKziepUVnyO/gd956yNvzLVCyUFlpSeUrcyNkZeXziDkOpl1UdZ
qXXR6GDwgujhfbq7Cx5cuh3kDdwTr5uk1a4unjbaBiR2upkVYcTUu/dTaivtS7l2Du6IQfPu6mKV
QueMgpQUFGpc6LZd9GLfq/DFK97r59GSIyLbjo4H9Gu+kZSW+62PbsDF5IINGuCp0Im4L0yVL50O
ztfspqoNZk6buib2rHT/35022RTC/OI0g1zFKdfxsrrxF+zoT0RCzhHmOOwoAAgiEbGfgrCM15lD
6cwOT7YvKKlYeaEkhX8pp1V8W4cqzEzHnoPrfU6Qc6KIoq8Q+fGz6gcW7eURBbjmnjHae6ZxkIao
n6LVwu9k+zYzSMUohJhECHW/tMpfDQni8SmVin3wucrFpdvHaf1IUZves4qq5uaL/ou+exXPBqmq
2QWS7OeKd8Do9wrpnnFb6t0ykK1L23GzRYv/Jfq30oncuKmTLccdZr1Dr/s+qjU3kbSaUBaMIPfZ
ySzlrMhmeR8bF99R52J77jiczVMxxBoWfh1iliYdMdKWjXPEaI7DbzT4fDBliOOytAEH2uR0S9ze
bwHl0HC4Y0OQEN0LFd9IbLmCIpsYLFCf8GuupDYuMAQsWO+EWm3K7xzwhMzrr6IISBPPGKZ6mk0l
xDKz7/9UYNsTUKBpzQfPSEO15FtWPA3i2vLRYqrqx3ffQAplqF0PvyrXE1lB2shYof5fREp9anvh
FuD9vYAIA8blGZ5Z97kOTi4x9SVuED180yY6iqmz7kXKCSSIwNoMYVE1wkYUkIe03ik8pXdPVY0G
wrHuceGMtMaKIjmc1jOKNu+L7f6jkXcn9z2Til6ND7+CIJF2eKBAYUlE4mp3KZlfMOzcZNNtq9wf
PH7alDluGjtEpjkMgPRjLXiu5odwBt+yNwlTUlQZH+k/XIzcN0Bl5yhMhOLXTio8ErKiS5CO00Fw
fTESXBIkG649buWIv+X4gcjBhbQ5ewzvcH5kdZBos7Lls0etd1ruBHimrZw/GTpIY2oWOHZO+pCi
uV2Twnx2IcVm8H2lylG2LJN6eCr8+vvXZhKLZwEZKl1GQa371zJI2mHAYuT+CatH2BypVlC32Yo/
mtuxC7ouJPxiYWQc64Cx6woYCbHzVVPEfUJsvWau7wZL5Oycx6fO7pZ4SiLSnRGTyojlOaEXCYBl
18TxVKZ0dByGRMSmtgbk7hOP1yNmI/veuonXUj9tayinmPmwdhNnyWWZ2MCnOeepgGhVtKrrSf1j
SQDv/d/6zyLo0ieMu0x4RWCI82r4HINUyevFUqtdGQr9oQ73HAphErv6e6X6SrThC/cxg5dhMOpe
K9mNEEAvRmuHjTHHEIXHw/K4CkzzeLGGjkhRr0S2fqh1J7RsC5vudPeKdJEUAvJqwdMZp+tvKAHx
IHTqxbljkWigK5IHOOF6dwcjj4xEEM0xbiqex6o8iOx63X8rBIWtjXjpZAbkmaESwLw464qA+eRu
G93eWwuCVjVhlrjBpxUGKJx/PbWn0wTUj98AbVRwON6RzMlwa5Cv0owCp+r461kXw2/ciAFTpsVW
zbbc2l3DaoE+J8p0zkJwdwj5YAk91uXCLZ9Zgj3Zj7ITd142Opm6U60Jzpf4ARH+s7xqR/zZi/Yy
5agLirs0BXAuWFrSh/GaPgamZFI3hNzKs/9p1saUeBQmf2afxJXoLq0AayWykyJGwaU7PSaQobIH
LYxKfDW5+mbE+RmYxKGHsiPQ5N0gIhPFaikAHwIRUPcIL3oHN/xHkYwU+1gBWNX5658pMs5Wh+BI
Qpa7ct/3Fyt18S1SlYuY3/KE0nHUVNupFTNOhyfucRiEpOpPW0JqPWcyxuPMLfMPXF4LgshFolaH
i5DAM3cmKcbcsbB0PFFcSZdyWF2KLTjhLpFLWgbK48yhuJlE1ZOpHlN4JxCdVI32WaGPUzRVgeXV
RVlyHckLxvCPMBz14g4BQ3rD7SaGAsYue40uAsUKO02rfA2o0y8jb2Xv2Y3iBaSqjA9/OvbsW8PY
I1QcOlCCbOB/B9FU7txaFT252KTsJSBc2rgQgR2oVxtCQEsFMzSxck9Mf5G6wH/0X9/eZrc1TZyM
m2Y6K7I2gNuBIbzHN3lC6EKB45gYF7gvmkDrNknnDVnTlG4M7MYMt67H+WPetK7ae+lHS+WlsCOo
tbxZwFtFoLY3yy9zXGccY4oYPthQdgv+vVWLetwg8xuc8RIRI+K0yGFxFxON4BZ7QLFt+GOe2Sqr
BI32TYuZKzOmWpQXdgzTbmnqlHpBzGLj7sj2/aH7Xs65eZggc36GuzF3V8xTwdq28oBaKjMHTJjk
oUVP7tTCCYgT46ie1dfaeiQPnHuQ8Ctrjgbl4enfxDUObMdyxR+dPWDlTKM3ENHBt+FvpKLH1yPg
FFTXlC4Hwna5J7l5469+yCUeXK+tzqmTWa8DezG34Fu8hkrs9wk1hxGNS3ph4E3Vcgp3XZ6lJkHC
14Q2UvALOcS7OE7loGjxNNn5MXhD7Hx5U/7au993wzMVfqs7kylMD2WDVY7Y1VeFam7cib8HPMmx
AS5pK2guKeNvOgPiatRY+an5vm3+PspeJGoUecGy/fmfQmivNCmVAAutUHAa7liVfTaPn7kwexoF
Yr1dxEd6omHVAAbAY+eM/8z//+gJm6T2SxovL/mM6wJ5ueECHDNfLvqUkKDHi9DB8/7SKV2Z9w0r
2A5a3kfGLW+t1jAPqN1/tvvD+CuGxnJ2myqaUAdhiaduvGDHgVuSQIITewXs2j9yI+eHnvlZVpJK
jvXoQqkj/Pkg4ATRIl8VpGxVHb1PiGoIYMIKpWZGOuxVrXfj0MxZpm8zsVRtu4XVCYDXDGarBzCT
O+ZJP0hPbYgGaHcFOqi1u2PL+4DHX/oJ0UWd3tojO2AsWErdQ/HM9gsJbHLfcrSZ4vsleKeOQ/GY
3jR4QCPimZfzKit7PLQ+TzXmy8yhvCvy9RoZUk0AKrQZMEPTuZSqne6NSi3LbfJyf3N/oK9K9H1z
C4o/KUku9YOjE/hYxFgB699b8pR8eW8edxvzTXlVT6+jZ3SS0KNpnAHIYX7x/NncoiWf1OSotiqP
pd6f96kq3OpMD/KvexqWqxvA/tyC3eCk5u04NwfWTK7UqpWxRSVizkHw1Z9FguqS2lCUil2i33fW
dlDSi8dsNVeeXn1yb3JSZ/+pyrzmw2ZgrDP+2I8g6rX6rWmXlAOpFw/u2lqhfzY0gDp4ENkMFOm2
IR1lABSSXgpnPLVKhca5jaC1NiOGpNlBXtzDO/qsSGMoFb54y7gjZVrn1/W68JbgRfADyC6H+0bF
MkOKQgn73UXa5LSvGLO5UiRSi3n/3u5QIceVOybhE8co1uszfcZ5RkIFVXeAh0qilXSx4JPTrsSg
oOqZ9+E4xTUmCfybBweP4v+NikRFf+iafu9EpQ2tI0CklfyiOGcGckcvcFnq82ofAKi0J4bA5zdu
Re5ZoU6FEhDPSZPUY0tVa8tzNg5qUDu4PvgAYzHaHzcCsoHea/L+woU6bvdxM9cDtO2qCmh/5ZpI
wk6xvTShLSkPBxYVdulYADaZLSt4Z8c0dHLLl1L5B8SfEXHKRGsobL7pHz5aD/qn63P+YJCoCVh6
J/7Y1faw5gbs231rEmex5YeA6lrLgzsuJ8gCglmsfiU6bEaY8Z2mKYVReuBuNskNWa2sYi2Py4by
qaR33I+8aAh4ATtFVtHnfE3JNPkuW6PzvcKKS7RJUnKyKQzKlcmyv+6dmgllOWXQ/u4GAbFswmIi
Ku3I15Ffj6x3ZtOqeU6R0Ogqbz1K2UyHL3Wu1iZtNt2csiun1+jHA8Jd0R5AdZxazNXWToLno4+r
L9w98P7Rw5l1jWjHdvOfIk2NJlFkTLiwdgjnxqsv32OxfoIozfJx5KWHaWuLVUjlRGWQWARfD4Ut
pp56QR5lKvedynV2U6yl8vxyjpJ7mGuE+eU5BdaIORy36Dss9s+b1sZG4o06DvH9zYkX3/WATqaq
XV5ITqxPdUJ/rntbMRONBJwLGYBek6RJ7RlDsjRuMZ0c8YK0IsiLOqqzJvdotEX1FdkUdbGsesLi
LpqcfBlIOZEo2my/sxryb/S5hOVXDXHc93rxa7FnrWV/b4koB0e5f9JO6U9dLfYY1UZ9zzqvoFtQ
cJ0Lhf+eV/wk5JX9KQB23EABJ8RuEVCzY6o6HBITs3PkM20FPzFe1yXTNdYzU1LT8Gm7/Q/UmtLJ
P+cxv1i452HnVT0p7CWdSpgL96s9yY9/IrZkhke6cMO/WsA9z1xYHw6fhZrfjvo6EnqxOm7R2Nld
thWiMY9lIIOjpCMwzk8kOiqryDyKqEm+nc/hBdUrk8AbE/Q8NYskirFU9k2rqeXK6bGA8WjkmjCN
kEDPamGtbWYusAEwKRV8nYk6B8Ge6TtwpRGQlykMnMDhhBOXeqxfT0xPqSP+pPbGHZGz5UgiQpe5
A/u8ME6pUZ7fDBCq5Q6hmKPoQoMMwcjZxNh0O4+D40cxcXDG1eWZk0t4S68krr3sxvV/JYGPVp0M
9u/g84+AJYAMkAP5xPl5wtE3AcyiY/vLUkK4BrldAc8Wrs6pIlNVmsn4V2MG7CDxNxRzymP/hjWS
wDsktaxMTn7WnjonpLdPlnEJkikw4/L7cvqFEs2GOxfafv2h5phqE05LxNlJgzm4GpGqZT1axk+q
U0zl8iyNUaRRmbaLvMYZIXfRHZPr0dClkjoUHcPlmfhQSHtZ2Wcru7YQpr3qD8d+MI/FFVNDGacN
T17p0PpA2BIcDjyXkvlXePt01/Sws7b4QHNxKBj3m2EwGN7zWiAiURY7s334qwjpIu1vhHZ12GLa
ECdS51zfEPImgkfR+F+x767UV+7IQ3YGO7rjBRFyzo2aDTvty6q6930PYl39iRpnS/+wLFhJL40f
QDH/xEYsnLcSAkRpvlCYmDhU4SY65n6H4vmuzHuAjEOxUzTR6+NpSUxsvnL4390PJXN2jFEgB+Kk
mLvsddS/G6XekXj7gYGiHCKQ9fePRYVcIaDRWD4CviH2jxp4Kfsv+ZUTPCCMpN0UDFXCjUwuk1Oa
pZo/walc2Mhtb7R3plUe0XJwUwxXaW5IT4bYoPOutsfODE5av1NkdxuWbJh/jq233Prq53rIReGH
b9rmHx97GiGWrHQlfoJ2spXgXZccLkML5cJ/6JhBiO0ZDx4/7PwpgqZ0U4thBf675zsw+XBvOY9U
wpgQuct3SfMYvKJWWceOW/ZCEzarn3nX30VlT/v0zddKsu+SBdgJuLmcdu34Ciw0Egc7gDyqF0pM
3x8+T4fRYaco99GRLr17TbbZSddpJy3Og0AmlsACydgF1bfZZQYQRPB3mfQwglA6MTTfq3H/GJHd
6eR6/ZMHZgXE3glqRsA4jfnOCZQnS1QtbT0CTIxCFAlxHOiVSJRE/DwjPaoFbAFxncMb459EAk0J
7ofr5EV5w3KtlDkvoKFZhrqbjDwWGxwhFmwyFHqRFEJkObPiDF2iNHOrj8K7705FTPl0izt47XIF
o3RecrtOM9FMe1BbejIEYJRO1iAoOs/bCihFzIEG5OknvfTUYUywE/LMuJZyNcSlbDyMKKFYpnsq
15Fbjosffg5xXKK1WGpWjJMMlAtNDnh4E2M5uwNdW8r5xlbtunJ4MVsxY6s9njWvxNz7mkh/waFR
CKcHyK8hOtoesrd1onulqldtM2AYC9zliAKuXXv02HJqjG0vX9Doj9ffzuMbFHcGeVZi934JKG4y
XaXmX4WQkUdAK0yJe0zm7johmCoNadmW/bCSDquXLEB6HSiUEI5b0ctzeDz8C9/G1GrjHkis6abL
QTcwBpQdbuTgGJZkPi3krHnS8rUAg4nglCNNDXQUX3+F79PVlbwygH/uJeEw6rxYQP/6gomqtcVf
pPvwAOhLQI3gxz0DiZg3qkYQcwvAF45qWTiXaRtZFvsQvBPqwQibeqHJ99AvtQHNHZthAKHEuXHA
dg8eon5J7+8MDrr+gjbDxk5UwTUPIMp07oIqsH7xddWWqIg0XAEq2HrwUL1OImhdjJBCYyDTK8Pv
qcr2nEcRO1clnOVG1/yfLFDU94k7qq+wT4tIbhOKE+DuuxXgfjM+0oAvn0YrS+tKUv3bdeZIeEHc
ySQpXZ9SrqkngxBLl0W+MerXux0h5RYuFSeL3NZRjrXOSZFjAwQwMerG2xEZGqCdpQ0fc9s5cI1T
3SdlRBDqIHxqML/2DaO9ghXIh9qdk+xqIp6qjurKu2h76zOEAd524MnTpU7dlrWgy637060BZt5E
OwKJuvJ9Y4NyzLAmGqmIwJ+xZ6AFgeq/n6fteuewrtjh2Qu9QmrWZXi88XkQu8xWikLXamaW5iXW
DQ56LuRenEKRiZ0HBVSlPO3MpSfc1UE1aD17V9jk+Slh2AViUhPtxGSLpRmWpuPjeVjk+kR7HlYl
adid+ewuqnQUC/22gtRSOEVnz6AHU0EHWogOGugBOQN0Oz88TivopCc0XRfsLG0Ea3tY1HZc/evt
O3CLOn6+1o2PWvrLM7K84/6A90v7FsSrk01vOWM0MNeE7pDnTh5tfHsj0NA0ggeMmR5QPld/aZfS
AlZQtHkewJua7fEhWlJbt2pu/vQHP3UNW5cBV9bWPomS9qon5GuN0pc2nc2pSdL9/RiFTvCPoyZZ
Ucld8soj0iLU0l8FYCEslNsOFUzj64ZNgDXOBHo0ia4n4eVtxfLtMhyQDjG/9umt2N9jhI2PVoVd
VmZUXCM+U4XLRV3ubi7bBTKTjGDtPSN9gChG6ksu4/XBYbxZRd8esMSwbCO9OTG29bA0XbTqAykJ
wCEIQKQTPWlnhlYNIj5KdkMr8UuQDlQF8krhu0tvtrCKaUE6ZxhPkCJ/Q37gN6Fpdi5Ly6bR7fSL
Q8BtZc1QDABlRz8A0zU8YOCzRrGdJITdGaKL5EwMYBD4CB1wfxIsg9Lu6dX8XAKH7fnUoGI9oxtv
+VQK6T+nZMy7umObh9hIufTEdGuVZTIpdNWCDep5vHcyBcdxvQuCwTMTLObqc23aDt8LM1rl69d/
t6Ti1ITpJ5wdet29pOcaEaEd170hnBhG3/q/QfF6hbgaFtcXX4N9UlUIEafyLeu027oP4iAhw9vt
B6SjD8Eop5KWziPhE07LtZlhWdcDvIrjCpFaCxke2mDD/F5KRTma1A4ZeSJZQGVTlAiDrb2WmC+6
CJSOS6EfSC4vZszylf277kuzDjBE7useMEBlLx67EXPRFSTtqXVD98g2CxKFJx3GfeIKUS/cpgam
QgK3BVzmiyp/RU69/ek9TDLmJGb7GU7BK2ZUh7WQwDvbSTfH1giBSkzk0solqWe5FU2MCQBbENJW
geeGyEJxkR7goeY+04pgWitiKfooh4AjNQ+QaKAo/h9qI9RdXCWZKQML57v9nDo7YngRxie9TyfG
O8V3sD+k6xP/x3VzYK0xeWvyexEcTTxtbVX+I+iVkmVYGwUoZSKb8YBakQN6eYf5Wg+SJdI73hSN
rk1FhVOidxQd8YOQ+BzW4KeyHGTJUWcq/TCmipBopX0vZwcG6jbmmULxlr8MQSf8phDX39evB1jZ
CcizzTOojtrYD2kck7xACxNENKfQiD14sDvnfmNapxQclAT+S30rspcez8Dr0nenbIOFc6HLAR48
Z81snQ3kBMSmzFifbQikggU02h6QQ9wucIyFeZaQGI+zuGTi6MYrqw6tRsa6i2xncy3Zmgb21jMu
C/oCXyq5O+HeCY4HoB9BseRyhmpnqHWe5AmqKaw+YCPygJqga4QJsUnvNV0Zui0A96MFLwT5c8tw
zW8GlxXGaQY5V+/ZHSAHtM+LyUUL1sNknYXSpbDMx36c9RXW1KEM2SU3a3fO6itVZttoKA0joWQY
rCpRNKFmlEs9BErL9BxTvk4UwPViNxjpXdrBaYbpjvSt/aXj7v3vFMnw7IWKp+toosEP51rtUXAB
uwoskkp1nax7qvDifY6IdgEpt24YJnZTow+5MWFPPKpXvz+3B6vrCLZnKTbuCzuRm9SrFyhb3dH4
5CP/Kc7xORdoEO45RFeYndVLZLJm8Eqeh5TQ7t1w9fut6wiDm89nlEqJYx5uwjq5Zv8BjQE7wN0L
67l8XvzYqOr9gfllWqzmyuibBQHpYRNccfAYtifvbOE4sE0lTvX0MIE8zMvLuwzARGadkVqF85ux
6j7m8qaTCPlvXTPaOYED5IjaOZRMwSedDZOq+1ilTe0c41jXkueLpEvaDfrYKT14vparwJjuJ+mW
Z8rj8syk0zSbiRC+Cg+EnlZr8a4pn7tU8QAjzl4MkLlQYkOAwxQM1P095OI+chb0hlGKiJ2Wu6E1
xK6YhRSNeqFESu0oilgH+xq1ZXrLQqxSZcc46FAjK+5ONBeHXc4tQixFFUfuwPYrCNp393jYrNDU
Q/gXNWdKHJFYpzXbrMdMvPDL3tFassi49INxc9dh/bZ8kWucATVz/UF2t3eEqgBUpjvpoVbcf535
p0FY7Wm2dE9jGTOmm89Wfqtt/O+z7ADxcgIy4D452YD+vm+2VpAwCDSGbD/KmY9PU2Qx8toFW0YU
xWDP8a1Qn79thEJ4YAsAW4dLbsAzLb7p7BzQaszpUm5RUn6H8sl0DGI+QbzoOfvbHwXHWNoQRXms
6y6oqE9NATFJ4QaI39aVKEdXm0zZIbrDoq/UUojOdysSKWWz6FTPIhVeXfZHYwZWuJ1jwfc6YLKr
BNMgWirlQ4mnZs6DY26ehuAtWOLDj9I9XQ2m51EQxhNStS74v1Tlpgp/tQVj1L0AjLDKBwegmWMi
AdTFCl4z4SsQu72z/O6HUCkKojgp9eHmWvFzYDCTyG5uA4MrqJ1jmpMVFkiWs2WFW1au/WJmuHYw
RT66Kv7IKdn5eTXHOsXTDshVi9tLXJtzi5qeOGgv1YTFkRI51y0mYbcVGwefRrxA/6SCO0DotPU+
GhHlEH3Ubd9PcrNRio+QK/j6nTsDBC4zL/f7+ZCUrV3jJmvWsnDMYjwg9wRUiDCd/SYmKtSd3w4d
T6ghkuz8Y12em4ihA4OfiWBoB82Mihiuzk1uTZHYqeYN9yMSP/m3G9qyuS9D95BXM3X4ZfPCEUHn
oRbPj33l6FiF6FQzgan/fyDxPqqCgJjih8V1tgbcdVub6rBMiw+C9f4r71ZRZIKakaX4bWEsP+AJ
JV3etUbSLSHGWAdrvYZU98lsyxTKSGi04UXARYVAa1vUGlnieSEGPU/f+Tg7MZDBbTeVg/sf/Q0a
KwmRilrFL7UCW6IqcNcXiYzXIqIZJpA2n81xoVlCjcdKC8/N9wepIfu0kKXYx5wC26A8o/45G/qY
HJrJwaNZzimQ5G57uiVKkVOLZoNJDpBzr+D//jf1p0GwPzoBRNST1e1sWLaFeWmgUIbpmFx3BylF
2n4O4CNIq8hWz3ft4vapj5wkzljjmhyrcb4PiiiYY52qNb3wWm/Scje+Pyc8Qx0Wz4O8FR2x7u0h
fxKUVQOyAYiedUYgsGu6HvnSBknx37285qVIkX7T5b6fP1x32INFrnkvtgNbb6YIOKlRBlUkfNw4
8IY45z4TWWjqx9wyuf42XfPjiwywr0hKEXYM4A57RNGQz4SGNMlibqC5VIgFbJBQvmZ3S5UHy/O6
sN3/J7hQnwqsP4q5gdqbykfcgfFzY7ZzZfIW0e4CuGU8l5rKzHuQhr8sdDPXJrxEi9MfzTWdf9uo
uOYYVKSHUkt05furijFooHtGnYJDRk5C9iLMHPH6Tc+36SjOAiVneaoG5qt8CJUNjtbk1m8p/v5l
bXD54waT321xjW44DZtn3RtG0P8YRKN2sB38P/hEFIt05Xw5PJrbP2V/wm/wckdkNwyxo2GJfzR1
p6cxAZM3UWKLTY/IFA0zMAQ4LnW7/cMWLG0ZO419bV/sdq26ttQVmDAJobVZ8FPrbOUmhEKXmqXp
AHIMyjn1xAYfZUw=
`pragma protect end_protected

��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���X��f;��on�# ���5"0 �T�PL7T�0����Ǿ*�Յ�'x���!�����*��w���0`>���M�I��M���M�At�YY?��w�/��
��D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��Ěכ_�fK[��Q�AU[�MQ���;�g0t��=#b�ػ���p"��oД�̈��P���2/��$5�%[�.4����%��Ղ��$���*F�F�\�A�"FЉ05�!��1���[0TdP�U+֡R�y�*{w��SjG��^#�t��?͈ ���~e�\	�4��}��.����x�;�&� J|/���M�f�,3��}�Д�ZmR�,�Y�Cޚr����z�/�Z�Ѹ���������\�%�sz�HI �2��M�'WƉ_�0�b�{�̃�?� �Ms3�(�\��]qS(�c�`�1		e����m,)�!�:Vӂ��t�Ǟ�mY�'0V�xs��D��u:���~��5Z#�0SX�=@/^o@�w	����OA��ͩ��]���S���\��Sp�I�NB�+=��ܛ�;�@�$�d�7�]��Ҥ�"��sێ��FZ��s�?�|Jb�)��Ȥ�u!7�t]�T��6�G�Л�� �a�~��`����=�N�~���tПI1�̐!N�Li�}��;U1�>LS6!�5'^��}����
g�p�D%�0[��H�X�,��e����94� ��s0��w)\JU�/�QG6��F�y'ol;��O������_��&�%L��Z�#>q׏u� �!!���}�ʽ����җ��e�����"�ă+j�+6e�ĉ���76�A�!���=�9o�_v�����*�{|6�Jr��(�|��f'���Wp�R�����&%>���?i�
辻��\���q"�a��E��d��
���8 *�ϖb9��H]��H�W��|}J�yK��R4M1�g�����	<�yؑ�W�P�)O��[k�	>Fm"��x���k����������q�@��'�� ��J�����|�{* t٥���\;�uUI�!�@_x ;�<&>x$�8z1���Kr�W�t(�de����F;]K���2�NF�} u���^���bȾӍ�q=��� ��R?n2M��<��Kk+��ٜ������qy�5N^��?�զ�w�(��&�B�����.��+(�f�W;�qNU����<�nq]�<;�|*j�Sቯ Bt�Ї�Op
ŴpH�r�mU�[Ϣv��#�5�x?�_i�~�$ѭ5�H���e7����q�8X
�  ��#c��Q�����=�I�)X6��|l����G�vB��UJ���)��9��U�_K[adJ�))�i$��7�w^Ay��+"[ӫ[a�1�|oS��.��,m��u��8�.�k�UC���6g��{9�n�F��b(�uO�����rTVZ��Ԁ6d��&��,��p6eێm�W�g�����H}{�eL��I�}M�:� ā�x�I�86M2dNA�����ϝ/ɤ��h;,�'�
{E:d�(W�nЀ�)�՛6�5��Sb_}Q!r�i�n�U{��vNU���8w/���B��PYߗe��|J�)�<���"}��@J���x�!��P���[3U��|�#X�d,
�9V�d���#�~}E�hq�gɔ*+�.���M�hX/���l�V����Γ`I�|Lbw/���'[I��\95�UX�DZU��*��Dh�䆷�'�N�\U�u�OI%B{\��rlvƶ�J��t��T�J�����LT'�o� �P�+�IQwY�k2b�S���9���&\�@/5�A�r�Ǹҏ�$��J{�WmNm�C�S�b����*����Adf��sOS62�VT7$D5���I�m*�V�qZ?̃ZD ���HƢҭ��ު���59E^�Ⱦ�F�.�9�\�TP���;Wj3�Hɏ�䕬i�i��x�o�4�|b�`tpIGn�Ƽn�]L�/�,�ȴ�#Bo��ζ�_�*~ +C��/��g�����qܢ���0��x� /���z�f�I��>4����j7���c��~�Q�*^�����g\`=~w+*��Q�ζBD����|ԍ�^7�v��v��x\dm\�x�D�p=7�����B��%S9��H��nbb���XP1��*�4p�����z�<��q�
d�y�H5����z�Tq߂Ƥ�Os��+p
Ml���a�n����SO���	IN�80H׿��ڪ��^=6> ^�����Z�*�����0�⩓z8����������p�����`�h�;Z��t��ꨚe�he�*�D��ى�=x!�{�/�q6�Yc��u�/��$�%�6䑥��KfthX��G��py��w;����¹x������1��P�Q�;	�q�������|�>Tk�q)J��� ��+�F@5��U�wuj�q�rg:CZ[�K�����P�y�U�N'��X*���J���:>^U؛��цF�y�\j�H:�Dp�*T����
�R��}~�X�"��,]Ǿ��G1�r�ѩ�
���F�h���:��߷��ԩប�ԇ|��C�^�C~��ШE�G��۰����ZT�ٳ.��$�C�U,�gQ����n��O�: ��uHQ5m�u��L�m��D���ޑ�T P���1����.FG渀x.�[�2���L|o�]���^uC��	��8}�YY�ԑ!�μ����#��Ќr�����,��p�m��K�^ۤP#�x�^i�tPq"U�EYEA����A!�Aٌ����>���S:�ȜB����c���H��m��e��y[�HQ�ws���lC|&}�3���Ru�2620�b%N8� Z�s�E�G�����hM/N�/dHbH3��U�`r�G�>�����y����u��P7�)��
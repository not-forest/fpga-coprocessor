��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���X��f;��on�# ���5"0 �T�PL7T�0����Ǿ*�Յ�'x���!�����*��w���0`>���M�I��M���M�At�YY?��w�/��
��D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����P�^�Mqap)%t�?�&�Z�K�*���~O��in�ÇZ2���RG����R����k:�H����`�E�m��C�H��Ё�]]ѱO�UFH�Ꚑ�L
��"�0dF	�b5 �A��Q��+�	-�eD�4W!o�� �@G:�� ����Ͽ���˱z9-�n#��V�G~i�u^�L�������;�q�A�~��4�X�-�]Yl?/�Pa�����4ǱT|���G4'O;&�;�o�u���i~t��n���4-BǇ�aM�ݍa�ڗ_�bF�5�����
�s�c�<���w����\�_UN�΀'�D���+�qS�e-����@�\�By@÷�:K���F��W��MV�p'^���w}�#��
�VﱫIT����tL'c�>�F���b`(6$T�j�{���x>!���4f�R�;�'~>P�V���^�-x�v�:F�4�>I���Qn�0-68�jfb,:$�9>�X�y��?��vLr}p$?�Vw Q`h1���M;�qD� 8���L�-���1�#���Г#���J���G��Ș���H�������I7EY'��'ϝ1�UREcB鲱��|"8<T#���-dݣ%�*� �y����\��|�;��郫#������rC����n�D�x0#�z�wO�������F��{����u�$I8�m��y8�A�s���D�aehq�fۨ`.�
���zL|��˪o�I(��n�ZF�0��1����<Qdk����/�n^�������u�ڎ��$�=�[�[���F ��������zw KO8�>���X����$��]�JȀ�(Dm�{�̞1�ĩ���9��Is�;�)���D�˒%p�8�@5����,3$Hء��uEw5Es,O���s<�})�-��Y)9EW@��g����=���K<�)�k}A
�����r�1�c}�;M� Y��:�x!~��X.q�A⿓���R|�(o��bS�N�����$�6�-��D�J^KC��Q��A/�%��B�c��b�ϟ��Z���"z>B����wl���\>r�����Z8r�\��*��5���q%�'"쯽Kxid@�|`�\�5�&'�R�ѝ�1
�����-dLz�K�Мl&d���V6����X�sH�XO�nH�Ⱥ��r��g�2	�L��Icu���9�ލnv�N\�6]�w�+"c2���h�8F��Gƿ�]wR<\��_tnOI.�מ��|��s��4)p����������v-t�.�4N!�-��eZ�(�1��yv�~�㑹��Rݖ¤�1�@9��׸{A�b03LO�?c��\ ����]��ɶ��|2:�"~rE>!����<zoW��ؙ���G�]��}&�į\|����Z���K_U�_f׾�LȠ��
�"����p
�y���~=���?�P�V��i����è���sĝ֦9h`4yoJ�\T��*1k���)gW����3 XJb!�bC��j�����;L�SD[d��7�6���#�a�qMp���75�aȷ,]G�^��Yq��Y҆'�g�E�I���/���L����/��}� ���K��b}�b����؋�j���[8v���IX\������U�Y�7�#��+K-�tT.E�w휃�ɲ�~ARS٠?͉�T����b�y�XS�/? C�	�W���Z�5������!�g�K.h�&�.� ���n{�K������/
�//��w��?���jr��`m+�o�e6�ش�K�E���0��ˀl�}
����O�`Z�o2R�_�s�2�6�t�2�ퟮ�$xԳ�+�{Wr�L`L���u7�nr���J͑�H�UT��Ogے�¨�|.ekT��ޞ�^b�.�<'�������/�5W�!�u�4�9�\U��Ma>��đ�j��%%Z��Q�L[��f����֑@I3S���t�<.�/�`��
}�{�:��-uP��T.{�F�p�	W=8��Z�x�9����\�C�WI+�����|�\ɥ��^�i��%�Q�A0�2�)����}oa3`1o�(߄;^���=�g��99����	?&�w�[r?�'w9��@���(��J;�3�M��+W����w��7g��X�%��úh�1�P����jOt{q����M�Qavd�����zq�19DN�J�t ���L3^�o�L
s��V�Z�ƛ�6e�Xț5z;���P����/�U�v�w��A���|�պ����u�D�`�zp�����i� M�!j	{�����G�O9����0�OEI����1��}��DÐ��-�f)�:i<?h�T�n.�{� "gSԾ��C���@1����8��5f�����X{�z�bb�H&�	Ƿ�cM Ԋ%;����u:������fg���N������3�����f���Gt�E�i�csf�rnkP�y���T';���,����D+�.����B�;�FoxO�F=�s�X�`z�l,��iRѳ�G��"����C)�q���K>u�V�]29{�?E��8Hؤ�Q��O�>��}�!�ky�^~��.%E�ZAb$���\�Zp��"%̖C�{9{ *��*���S<�h��=����+n�N�Q��M4��-7�Huc�&��*0y��vؿ��W���o���w���l��� x�Y��6�@�ª��Ҽ\�#rsX;�:I�Bcx��S-L���8ؿ���78!�݅���#�7�ѹ<]�(��UI�Ǎ��<b���]VXt���,7l�^}���������y����u�ɹ��$S�dR��X�H�fz;L(3����f���$��\�9���;Y�v���J	6ƍ@p�|�)/+삤'��OV���z�i�Sq�\k�pѓ;&:KL#H/�rƷ�����ƛq��n}9U�s��7�MDD�.�}�+�r�$2˒1bSډ�_�WVd#�_����[uy}�pE�d�as�w�\�c����nx�=5mfڄ�p}Bq���s�����'/��)qdJ���d�*������5
^�`K/b��iRU�R��>��5�uiu���z����O����Ŗ���UM�Ȥ��'�g����"�R�K��>Tw�vr�w�Ϭ��Uo�0_�_$ʑ����]Ɇ)'���~�Կ�����KP.��?实0�$��_��b��9���W������!C��=K\���%�U��ZjHSo�D��/Ro�{�=��8|9��z��j��G������=���a�� ��l	U��-J��ԏ��$����A�f��~��=4��3��۬��I2~�Re�<�`a��p��~R�?�3i���#��ͱ���_t�>��㏜��N�E��G�
�A �݋	�u�Q��A�K�U�L^�-5�ʾ �������V���fƬHoO�l診/��>K��soq�6�
X�L<�R?��-y�����>��h�Ч aWK���P�R1�_@��p�U26<ր64 �}�[�hp҂_Qw��k�&G��s�����$~��+��C�9<(�����B8�^�n�63��P��_����'��%\�$$�2&�}��� �R�G3��R0��|�(7�BBE1�=n�'��+��u  �p��x3;H��H��E��A�/�N��l>,U�g��0��Z ɼ.���j�#"����Z�=�ɶX�)q��z#�Զ��1Y4��ko���	cOe�h^(�42͉��<�]]���*?�(�oL�ͽL�����K�x\��O�~�k_,
h��sW�S���Y��4[���C��$���  oT�1b���Yd������~�	~�����h�=�Т����2B������!����Rt:�SrI�P��S�i׹6j�&B��$�ʐ�>7�?mћ��(O�-|df�<*�;�-�Ex��'0��餃�Qɀ���c���:���G���ks���N���A��X%.�����u�5�p>���`x��O���cŸ�X��\�	�
fA�Z��׃\D��0~C�b	��n�
����Q����0>ى�81
�(���pg�}�K_�eуZ�WA&WW�fG@K~G$ʂq�۳�. ��:bʅ��X(�|��BE�}�<�E��������Nc�J�_�]�����}pNb�[�|PF*Wa['˷�ԩ��EVR �ٚlZ��ik�E���ڀ&ݧ3��xaҲ��K�v���MIu���e��4��)��Lڧxl��A2�V��P?����%]�&��ߕ�#�؈o+d�6�^E��i�*�Nӛ_�����TsL;��.�"i ��L��o�;�m�6/A����Q �i/[��P�=��i������t�	� ���� hk���s��Y��9��lW������MS�I�ɢ�+k70V^��Y�T�-3��?���9�N�o"N�	Í���LEڜ�	d��}JL��&5k�e]�.��j�б�z����o"\M�-�X�:�i��L�����w��LJ^��A=E��E<ԓ�E_�p�J-�t@ϙ�|���	(����IXy�m���c�8x�Bs\�y�J���v��!�f/Rh�;E�������>�$�D�[�����Ůe������?eH�e�'6p��0��˔���ee�B�1��[@s�T|�(L@q,4+���CN�;���(K�SJ˩;�ע͓��3G�(y�Ѣ�H,�ٿ	.ޕ�ip����l�,��Bs�m�h.z�{|y:�����e�Cr$F�R�f>�F�r�Ɇr�b���.��<����ծ�_��N#3����K��P}�����/�*����RȪ6v�^O�R3o��v�TH?���{n8ނ���4�g)D��EX�r?��r��C�����z6N�����S��������N��O��P���ؕ��u���"��:�\���oz�͞ ىt[x�jD�C��T����@��S巫�-�
W�����̦����֑W1.Uob�.���P:�6ƛ�>1h��︫GS����.�W$����Ԑ�Ⱥ	]�p�-õmB��=���1\�g��lR���(�����D��ȳ.ԋ��R��B��vm���bS�1H�u.��|ڧ-�TS�w�HD9Ǽ(�#�k��8�R�Obfd���"���%0dG|Y�f�����7)<���E�"���!?���A��´�����tD��	�l�ӓ����y��ZYM�]~Ezb�� GМ�b�1��X}�h���i�&)%��cv���C��%��4bu�\��W<W���t�>[�X)�����9������o��R��Pn��
1�cE�{n]�8��H���d:�T:'E[�(��Hbx��V�9:�
�95��#��aRǑb����`���W������Ҕ��؁"~�dkӸPa���>����:ϟzD��Uȓ	H��h*��,�>s�'����	B��,�����'�tta�K���!��Cf"_V�G�q�yh%�@�r`쮘��M9��h�r�i ���_�~�)H}z��˒��ƒ��f-���h'�I�t��*[u,��e��*���@�u3������w;������7�
d�,yq��!��e�+�+ӑ��,�~�jQ6EI�?��c���5�k�n���UC�����ں�wv�&;����{ i����駹��x���;��I\�翕v?�4Q��t\�b���Ԑ)�L�c��J�O�0�q�kV�Ho��/�a�Y��,��d;�vd���x滋�7�k�.t���,?Q*�u�hk��N=I��4��S��X�(s?�R��g	�x��G����"��#{1���MST��#�y�n�E����v@�����.�ܗ����[#-c�&}�TEA
�L`AePI�Zv��>�4z�����ģ���m�1�Rߥx�/);���[u�f�R�&���������0��|�\���L��,�I��:�<&�?G�/���c��7�Cm�u�������x���)�,oyV�Y��
�e8!��k��F�0�������_9{}#t��&h�f*�IЈ�i�FkT_V��;�iT���!� y�	V��O7���ur���n2Rg��*�Z�W
�?Zg}麑u)���)- �Ҽw����:R��i��j�I�kȸ[}�Xs�ռo��g�Th��IlO�15J0^��>�A��{\`�7P���WWD�~t���!�������a./����(�,i�DD)"=�*����8�D��%��D^��i�P%�~T����Wd?|�ٸxy"��y�5Jy����PYv�����|N�v�
6�k������u2�cݎ��@��ntD<ND�&Zf������c�]�Z�~3L�`���䟁*=�d�E��Cg�[I[jp�$v4S��F�!����|X���Q����}��k���CwZ	m��v���{���#����J����U�Q	kWmN�_K�D�8���� �*V�yQ���*=�'7��dқĽ�L����K]:` ������{�5|��qM���p�K��
8�I��x���M������0����(a&n_�f��0=���m��F'Ah����K@�Ӎ�)N9���� �͙��Xs���0�S��l��B�c}�������|n���K�θT��]�Do�DhD[�?�Vj���F�{�F��vx�[�qZ�&<S4X�Q��,,;8P����C��*���@6��䌘�տ.E�O��Q��͊F�Nd$�U��72��e��;F^�p��X��b�>	����S��z�ê}&�(�x���4Y]I"j����b9/��ҹv"���#��h9fCVs�r_�(��<�qL�_>�s�1�ސ*�6I��w�Y*|�mL.�����!GO�a�A��-~n����g�/V��/]F��������a�̔�7w)Y�lIX"`�X�� w��;d�j������C������Uy7��&Q��ݗ�`k�5uk���χ��Z�Ȓ�<��G0�\�$%�y�A�e���Ɓl��2|��lNدXVpƯl�qr�
�P��HPԲ�Hޣ�+y(�S�rw35ڤX�>�"��#��{�Yp�X��ӧ�K����3���{m��>�`-�?t�Y@�鶞"��,� ��E�x�}G�z����r⢘��J�ţ��$]d�D�K!i��XԽ��E�����1yH���� }ҞK�y����5�d:Ǿ���zt���ލ�"@3X���8h��o���x�W�F&�L�tc���1tJ�����<^l��oT�C����X��<ޘN6, k~�|�7���|-ou=>��wy&Čy�n��w^��囟���FB���p�:��"��v[��>#(�+F�)�� J�Ŷfm��hOYz���v����tψ2���Rp� ���#)��K��[G��h���\P�nJ�VgB|u��᧘G4ƴW�D������U$Y^� �pk���H�V�_�����*ǧ�~�Mw�&���ՋB>VY^�$��_�������W�
-c�!�<�ԋ?�|Bw:������~��<R{=j>'��6�f)�j�r]�.�e��g����[��=�e�[��߂��o�����|�����H9����gDt�����qc�لBDD�=�#�����;��t��`e��z�U������S!��A�8�ZEZ�@H�l�ui}p3�&�J���@�	Y���Y#W���*_0^8��ft�1#F��䘛cl�XI��_�@R��No��qw��w�('�J��2�K�m��,ڶ�f
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
miX9/A8o/YnS8SvMGQjLFAE5Kyp9MTD/TsOI+v0rOcjiRE4ELWW/zm6e3LNMhRBc
A7M/B04d3mLygLZJ37UjtClaB23Hdk0585BhxKpn4lL9ZP5rpDatZUQIKVTZQ4wc
U0PgkqZuemaOHxFIxNSScc3RQoEWVZGG1zKVG9W9p90=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31392)
Y3RzPICLjHysaZACSHLdbJg+9nDx7RtpLm9Km71xVm5LWIHkqFxNcT+9S018hT0D
Yg09kBJgf7993YLa/bcYDqQwmtlTrctAzUZ1QwUDR/d5hgjDVE8My1ngJDkkQkII
c8hQmdP2qZpncRbmLoc3PvtkfhZDxhR43iSeZOu9MBaSmSYZb3ivmUW7bq+0k5dF
L1HMTc57Px2TbaLfmfgwr1AqhJwIMoB54cma3ktk4Tsehc3zIkdsJas2ujb6bBpa
rnxxnW8GrDFux7md6GpEkh4kaPJxl2haL3PnBm/lmTYRR0d5K8bQWLvg4ReH0p9l
xpyFi6f4TjvFb+Cx0rs47ZYo2dqMVi0xtU8idy7il8h2FQteOLSW0rftXQDoJbJt
r4/7FBw0Dh9ffpCbdiF2CXVvmIz/x5gzBk0kvfoPPjv1u2yc8KHbJi4sLFJoSP6k
4lLA3P8PfuL8Nk1RUbXqeZzijJqSoCm0cTV/buJYisZ5utxjFtlLhfe2JY6izcng
80ozzwEmdWFVOlq9g/xSqq1glmlb4xklux9TvtCh5vElCVcIBjV/fXUrguo8Z0pg
uNXOQw3HGeds+ng6vD8xJq27dts1zE7lFBCy28E1jN07vBYQI6Zt790TlxAEGKFJ
ZWperpmy7D9+o/ogEkwt0/JWWwnT3cE+xa64EcguikVXuOPW/8g9cRVnHUxi0dy8
AlXA/w0yO1+occCYE0tpTcLmFBugt+Jae78a6onVdpv/VW9elczwlHbJoblBnRcZ
5vVHEVTayYVr+QMQMPVouNa5A20HhaYMJeiUaTKSQAeKviyQ6xkuKE7ZOj9l4AGy
UW8nXwaPQjNDmIOJvFtEznz/dcXuytnqIog5LQlpBLcd69Zthz0PGM5ND03Z70rl
5IUe6mi681GaWDL6FTo1k9c3ImXin/rLWqUdfg2FUlZs6yI9Gz1xPb42/xPDxvaU
DflyqiKRlFcDr0FunkT4XphpEeUaQP4EA/UQYYxoER7+yGKsAhC5OlJuwQRgrTTM
JW/JrUYj0DdBr0xIjIgrStSY1BQbz4GCvYoZ/sSJxTsQ796Pd05e1jV1wjnCLrbO
D/IvB1E9ZiV8kn8XYDzk5bHIrMBfYm1AXGVTZveS+3DSoz1Zoxr0qqp5h7NTbu5M
/ATV2Pkyj0f6ufuQmtfatcRL2HVj/v3AyT522m8NvYcPSEsqiyLog6L37B1V4tWG
SZBEOf/ICowGKjB4/rn3c+XHPP6jHjpKeR66RiIHzL4P24zCRXM4WiwgZDJ0ee7V
xvfjeqYzzs9hKurPh6Ep6QINdGdkXUXLw+ZZ0c8di4btrs4MVP49G2mlxmSwVs8G
WEkyqGq8XlLtOOXMoLZzDBl4qngJWtTAiXwy96iYAZIX28uzOD5SFc9/pVFyPDE3
5Jkn40YFnYQItflgFjcceP2UG/cEeUc/8eIhlGOOBw4RYQmgYwK8OzUOsfj1vSV1
/fMCiWMrDVT+Dg48oqbB9IUkkVhGtcQD7HLzN20KkPw9HIyOeykKA0mm8jG1Cp2g
6tGXYZ2wnfNF/obABCB3tpe2PvJvpHGIATajK7OFvD6ZIEZpN7TGfvdoB05pFwkf
7z6hYGjhwqcZ1TL8MOZTkilIgGiHdue7dHbg//Ue5AnkiRblyAqcuZlPSssrJYFn
cVbyXO06zCp2zghGwQK/vseS/tCEuspxhKi+rPq0W2JHLliIwTQFSCrCXyeoAr08
KWFK818fc7rrcnnGT/vk7FCC53jv6tIcMjVgKe13eWc6tTj95Hkc4zoHEsPA/95U
dh/e+9N0lTQ0H+8sFGW60luMlcAgpwM6qfmuThdwZ3Teeuz2DLQPicA4HeDqvHZ3
sl2QoLM1A6aq3XcNV7lusug1tU9fYfZUN5aiBL+vXo90W3zuIgoV3JAhZZdapkor
YHZVKXWFZC+y+EKSJevED7Wa41M2vH63bHsqLzm2gicKMUO2gcKihRKXlLwE99yO
EQ7RZ/J+Dwmvwbioy6Kjb+PyXhLruDzbNjl0T+bqcS53R1KtJ7SIfPnpRw+ye7FE
ok07qK00JXx/CE2FNBnvEJxhtpC+W2h5HqlsNRfFJW0aj7kLVLflp5sP1jJmzrys
ZpP21zPwGkB/8qbzPCCl8nMBLlveAYI4RD6t+5qX2FYvd3WSlkBp15Dpr96SLUmA
GAAC1COKC4n7gs5QfQ18+VHBfiVQgY20lxmXAVE7R5VmpO8bJXpJVLfcvYsorEDi
MTyfSZuUCVHR9Uc6a1s4a60O/dNmuo68yZFEMlYNpcoc7cq2sc60EEJcKVyp8fxc
tme3Lw7TIw9xukVmuf1ioD9lwcyeFn9dggkrabmV50NdvsrD0/tKdYKLbWDS6vAy
fers3mNrbcWnMHzsBjYPPcZNBf4CrxwYVUhfrLfkcr7h6Ww+36XxuIWUqdI5Pqma
c5YkdaMfxel9hTRNeGkLjH1eVAgKDDIOkmjV5Hnl2YV2o4iQhD+dze6CUI/9aeEL
CchSb2FKxYOXcTOc1f/3u7umjtDIVRNTUNEmV3xelwWS4UVgDPCoE7serhRAE6l8
haBUwHlcN5hZtFWiEo6hQHk3xazBPGVntSrYQi4RFN7O5NpOXqTqjxkMuWka8+pr
JcQLYGHUWc9Vo+APzIattoW8gylPwPTbz4pQKp4KXiWWRBcjcoNlkoUEYPA1nXmV
WnwD64bEXFGcQDT0nR3s/r2e9Bw1TAZmGuM1T9hbJsrh0msqYNs1qvlsDpNBNXZ3
VBHtDKgItzpeN4ZQClg/XAM0CuO4CjgQhcZLDfagylMzNes30kiRSYJAryBzv0cF
YQj2vpUyKjFRRrUZEduzEXGtEfCuDa0AT4NKcGfSAf+yeVq1sXA/isBhH1YaeM62
M7omNHY0x+aa6gTet0SZyhYGyKvmbJtuOPnHN8YVFK/etOFPlTSptE5d5mhJJRP0
uCRvBK6o3xGw3ruO1dD52Bz7gfQdMzURnpXYoZGvcQxBTIFGbfNA3O3zHRhbQa9F
nT08zY9u/1jTv5wcsKvp/ByKAii+pb37xu329yiAWAKF7lcsfS1XMREKc3yjvU9n
kfRjs5KZJ28moPdIaMk6DWJ0EEkeyfpzU8KFrYeC8o+tNREqfXpTsqfFoguV/EHt
N9JZv+KoNi7DOLrIrt3MqT2zYMBZ1FgTIpKgg9PRqjMHYXhX9qCpP5jbPyHiiM3E
XZlJ/dzVtdjOKLGvUEQVt2QE8Ipx+d3gBoKvywKm3Gy75SgLU23nQSS1U2D6cm2h
OfR5Yu/0r+d/O/q+YRmwnjbhSKdqP6sUH3rHRHLy/p73pjr0puDOF6NN8UFrmbI2
BX9Al0UMm9SqqbZFnFp7l8jeO4JH6Rv0L4da0j4HiIq5P5uN0a4G9/a4NPvkH0iV
r7aMIW4O3mB5ZrH7mYzi2Ta+lvnClN53q6Qts14WzrxMmmVrKe4ebPpBHyH930Bc
CwqkhZTOrUDBpvEWLN0tvwo7k9q7pf3sXgl/XWDFHR1lJqu0PLmyNBuElKT3yw1k
813hubXNRH7FPZ0sRU78LIZ+/eSWxXNgZBzaqdOHP+bPlfWhIM/qgQYoABaJMcNg
AQLminnAu4K0ymNesAbuw5pHuW1Qu5spxQLINt8Jp/gTBAcJj70NAhIqf3vYiy7D
5hQOyLG4Umt106cKghJTgR/zXm0Sym2q5CBhJJNXjI8fKTvhfxeit0lEGLN6snEM
9Pg+OxQh0BMLeZEmPut89bfwGPl1hajzzjsSZSBaUYuWSsGyp9tfIIjqVzwh7shI
Mk82fHgAMDXp3IifgIU2vycQaugk6v6cGF2JXOwAMDugKN97Lnq7A2iuucAXiB3E
E2DmswveNQlBlL6H893/d1f3Lgy2y3mNbwcEdEpr7e3vygkBYSV9rrC2KIXAmoxQ
3r7u2/fL5MkGEN1WUZWhoqXlAm5bSXIgTgb2arJ9FmKU3HyT9lrHC5maZJKd9Wdr
ezHAC0yXbgQpu9OUboollCyDYIi/uW5ys6xPfpgw/xt3e65BiEFbOmww4t/GoUBG
zk9zRkjwsI51esOchfYKJmNc/TqVmNwWVWMm3E/8GkUdVFuQ7TMG9bYy6Co7Md/O
MUp0Lg1nC3e/lnfmomVksaZggbuyEutloLhOlVbsbh0eeOuPH3kwiMtCiWsdSAhz
deMiHloOPD2PSjSjJc5lab+R4v6ygNGbERDNStAFlCh356/56614ADxxGlFp64wL
S9nhB37x1MjK/IyxDLAonGzedLxAN7F4kavpcGZdAcXTAcUmdYljQmql61t3Fi3I
+7tiJHl7lFi0kDwRVvq/ka4psapKbnQVXv6YwoIExYh+5Ov6CeCGMR2OrAeWBTTM
H76UqVm3TJI6A29cki3CXEKk8gefAHA923e+0emoQLyJaL+4oCHIO0Uw5hQoU2si
5MjgqNEOfrlpQgHzgsMKNrdAKyMYzcjy8omR/Wxc6LdED/ZIMxnpWhYs+Wr52abG
tYQZFlXyOnT+eRSdo4yu/vxPMWGdrzwDJhYVT/knkmT7j1PRW3QXtBrlFEg/1I+7
vpo0OC3Xb5HptKLLedDdel0/4sd5YKMsboLXU6GG77DX1DQ/9irltFoeXdCD7zIN
G4OBLCUvGyS2v4p4T6VyVKJ5maRWSCWZRAbsVoK/MA3uyc6w/AhZgF+6L2/t0LjW
VDPShP71HrGcoBfXObEnMQs43QE1ohl5cKOYs7FOFxsSbxjrGAElYPPaBnUxlw3z
NJF2M61ytlrkIncBFCyBjRTiJyydIBsSk5taA6bKEoYZwLr8GmaDX8Z4H3V28sRt
3pFdXBNGXT4Jr5/EPFE8F8Z6CHRAaQUllntCp9a+aP71Qqa2eWW9gbsW16Z5gg81
+koCoSV3AufS+WvhwlM3khMRbcXW7ieh9caKoPQ49yNNxm+dLv/bir8xB5zGAqQd
EkYLTYC69xKNIl/7Ptsd1vBu811LNal4prH9JrgiHHcStC/NsaPsxS3KhuAX+sD1
j5x4dpJBBTDtDsRN0m/glQLTNr6DyyERbQTYi+BPFWF5y6KUk+qSCrphqDnJIb47
GT6Pqluumcdq3eIK0TGJrRM78VII2rDFtakFsaWYEyK0Xu+8+Rt9H+f+10CLnTom
OQmjRtiNBkKZ5EVr0kQOI8BJ2zo8yBdZF8bxkr1hyPHuJAruj2RNcZPR6SwY5kYx
pEo4IuCpvmhKsymQaNaAcC3n7n2BA5wIxkTDuf2mzM+I6mSBdDdSHcPSCZNGtHFd
d/5oDf2uL0H0M/rMHx3mdhCpFPZ6M0DeNZQCe93iDJEWPotlIx9iivQHLW1MQh6R
bnd/K5AlmE45F+4y0gAzlNab1jTptaP/QKrkJc1NeFK4ZezuS2EFgtY6Vzfj+rhk
IhUmjKgNqxM984eDuek2bqTmKXLWcJomS0QTjWOTt0cPNhXc4mJRpYg1qbRww2i7
QUr4mDenttRE09/Zp3AZ3bSRkPhN3j9MvUTpCjeCQlx9nAxGPffen41vPLLvsdhr
8PCpLkwH/HYTRLXqr5Y9qT4G6iPG2847RQm5FEkk/Q2m8sBe2zLpUgvW/0VpBYI6
KErjb4nI7H+97DVt2WAqZHhWcf8AR5SxBpqSacncXQDZFnJqzIvrpKB5bg/2oy4s
5OetxTHIMdXPTp4IF9ZijEgnfqnfNVsRiU7ynq0EkFhIZezGJabj0VIQayhW/fLW
ULYiaMlUJVrTZAn9+vC/qwj+ArNa3iRKJTfJju+g8IdlE0Aig4AaF2yB5yCJuWV7
IgVFhwNNUcZwwK+acQdUelxVx836HJxeQzAnANZrHqwJPpOIUS9w2npTLx0n3NsX
m+Nk7TdjJxfnN9P137PdXTeXHVBuLa8LsfdAcUUSB/4G9zLdDvb7nlfV/LLxeXhm
lNuH0ANu9Ud1nHuGdZ0qHF0q1My5Ece6R+/7hAe9xgxKL5xlH8JHA+HD/ekIt8s2
lazZe0xyrtcACEe9hxt/QIpZhiuowGaNhb5YIUqZGyZXG8ZGxSuM6OryERLzg/y3
fTG3XOIBoy2qr0AWyu5IG/g3wxqBtYTFUxw9eAi8lWmclESk9EiPVOx9ibXykZ2J
guPdBoFPFEe54NOBynwBPv8Fn4rJVjVr+y/VWFjzN2rN55p42OC+YIYOCJGL3BvU
t33naBxG7snkpbSaI2e1n02zI6CMfj9/oDhiHPToPi0Yw8y5Yfx2MECIqT9iUq3O
GdyBRApNLfaRvFlimcEpT7H/5A9zLn/CQiiOxxxW577F1a937Jh2mzg2JdxHWbNf
V3GVJ4a8XGXaad5iK8rMsYFQk65SvfoaDH+JfEudUPC3TOnYLBSYN+amrd/OI+Yc
R0lpgaxMYomIprwHo3CS40FTBPxQOdSi5wAOH83Oi+foTRuhdBp6KQpvBQc6OsID
If+74cLYfmn6IRlBI780WNfJXNUNeOc8TEkjwuChl34+EV2xgyUaW/dmGYgspH7C
qpHOiuEaUnQ7FyL7+qBNDuuSMJH4fZoRIB8j6fN/h3sbuLFLdi9xJeXKW869/4Su
3k0HmUpKkOObiVjMd4iDW+n8q7BWDf6aj06Z+yuJoxpQFxeQIM0vYCNGRA4qokvZ
8sp+cSb5XDqrlTciS43fL50yr9odAMh9tR0So30nkHWumv8R07xVVt5N2OZa9VbV
2uv36tRYBVJiTPHN6mRnewZZ0sD3f/y1tSPM9GVDsCXILrIJpxAvQVjMHFbX2/nj
/tOAi5lOmDXAHuxuRp2dj55UoDd1BPHgDo3fhGL9WpphphxtGqKPu+wmQWxmtkZn
98uThuLz7kVt9I8Qd8HF3F9FqpN4V43pUoT08ft8RNoP+9G1InCto1BnsxAWo0qn
n7Tjv5CRmNdelG36iEdUljxP5RC93SRxvPRJkaeK4COkOtcHRS55ukuR2NR4f0K9
yAjVNo8GjRAi92WwqAVE/rU5lhvJjvApKjO6WNlnFiMWeYdhuJUSi26RFQPgQXR5
IV2eQQ+so1Zx2UpuiXZhaZb8GGo4EZ72P/yGzMSYPnnMy339HaLZR+SlxNTzLXSo
n47W5ntf+gGrRX+Vus0jCKvJuABuT6hmRVOXTHW/nQOM8R5YMzLnO1eCH7jqYeVo
AzXCZG3r30PMYuhHqfKWfutbJ0iITS1oaV8aX6OQUJVeJm10y0VZ6Xl/LxAWm3s1
dUMi88J9eoF3lIlDESkMiikSXUi1eNJaO0uGOT9PNZfozdTy7DD9G2ihFlWrnCAC
Zl2k6ta6YbNGL0XeoC2fvvGrypMhqgMz9TQXvttr3baEGd6w7/sSOjolfhu2YKAp
ftJPvLBXBQJVVRQd3SIrxMmBpKWhwWmeuZzq1gxFRDWqKamTPN4X+GzfA5INl2Nf
K+iYknVmChgPvWvdCGHEJerrNQoJ/w8Ijz4NiOxP7Tlw4FISyhv/W7/zzjQlwhIM
gAD2lGoGUFJLkhCGRfD9vAWJqSOhRsJBhqWGytG1mzeFIX9bIPHj5nvfGUfe/J4i
0nTlb203zmvzKS94gM1jOkkogt+7KXYvT0mj3xYhgO+ENkRUPQbTXkskKp1Hm50D
SI2AZ+Rg3l4MLuNp2HBRxVpvINLkI6w17OFrlh78whsBuAivAJOEja9ZFDpidfbd
KsLa1dolRVALs+vr1NDpt8gJ0ZevfX5MiRVkxwfVewxBUSaueQ8ARzECbGQTQFFO
Hl9y+DAthFABxsF5VQH7fx5xaJ714aHTg3IstekuPugVyNIDNDHJULD8CXOVxdE5
fueYrNydymgSg8CM++tOpCLzzrXZX7ezoYk4HkNY5OEWHzrpY9H0/JRwEpkZRL/p
+KG2aLZmjqJsUOPDBzFDw8jj1LWNuLtl5Ct30P5v+YdxHFRDUjq1IWmkLF1pOW/Y
xrc8aRfDXci8ASN/EU1TU0T5UxjKWCpOHZHwDMazSoiuWDRbxuB4E59lB1287ygN
sSXmbfMBDoaHlciHUVaCv/lkwJDgZhiWRqAezax0FNStoH5BA7gFKDB4bawnxSzC
hgy9FQMYhi+fFAbGhXuFpUEVTq2VfgFiS3df8b9S8FZWFkwL/jAWXl9NCtrXKEQn
gKHRwKFzXYFwmcw6/npXtcvm3oTbKY8cFs8s8b/VugX8UE6HNBzVGCOZRKZDRg7g
pYNdQLeEE/LTMi+rNTEHQ8sRhCXaK3/VjL3/8C36HNg6CW7m/7ft59IXKO0y+ST7
ujrV0vDfesE3krhRsrX/RFKZJipon8wCZKg9WjwAVYQ/KwI83O9b7EGCUyz/UqiM
SLFKMxeTEoHXXEhtUaCTv4CX5JZPN9ZkNtaGkDHRBUOyLgx3SxUFajL5hix1fB/B
HpLbmftd+gmMlbTnuZQ/4mAfVU0dzo6LASQVEpHE7x1i7KRNhgZ5JZrKcJmObsag
bLdPWqVed/ysfp40hzmXIgHtddua95FoaokBIxhm51EJtajP1PkNC3ckHtZg8sK1
mFuUHRn+ec9hGOR7vZuramiPDorOKUH5OuBl9Ef8C19SEfHZmG36rIQzeiOjWek3
x4qcQ6twvxOLw2sgKTEZvPb6kREZsUvHM/xNoGlYtenZ0ZZO/eWeWRW/msR0fUAr
SOPR+jAt5qrgQEtxgJbNOypZlfS9fsQlD0MS76m545Uh62fWibDKi0K462+T8qVL
m5nZF8yVy16CxtlR/ZP+Ihp7eBXkRBrS2rlFXFPS/+aqqtFF4P8ZRHevDYwk7AqW
6/Xls744/ULWXfvwawsH5pXArs4i+VO8xo8be7UCeKkY69uCkMF+eMxBjoyzyNgl
nOttyLVqSqL2b82cwXDTkmPfM+9qdH+UYaGOQ5ZcO1CVc8/pgxGvsvBZJw9N+wYi
1ZOfE3eLbUx9Lp39vEH2hRkdqEJlOsc2XRdNcrKdJjluaIgtMXzCj13wYO8CzMw2
DY7FGt9iOKcty5z3CZBiQBpSIJlto9WMRdy4KMX6Be4zCCd5jdhxtLl6gFWy5glg
JZhW0cZL24yj4e6i0J7eyi/mS/2S1cb1ssWkfMA6NNAFzfhpEOADtKZf9wBiorn+
zLKfZ1pqlighRb00cG3Y4UsIAqKq0DgoZ7g4+idiGJmyuNhwUy8t30YE89zV/HM8
E76zq5NEvqC8GsamNj4bW1gFPZ5uRg5UVzqG1mXDCzaWCnyy2v6ba5sGXaXlAGTx
GbLPqApm1h+nFlBIPbBBAlHlVuFbVajZxXhgOj0mU9rbf8TAnh+O5L22gAZA8e4X
ziBv7uGv5zBNOXl4hrv2TjPj/yBAlf0GE6a91j3/PD2NueRxecKIXblhpEI+kzu4
27O7t2PWHWuEQHKmhx8GiX/3ewvZo70bE9Oz57TA0AdYUzrX4lhroQIxVJ/5trD3
Hs4f5gn5fsF2iOzymufXDtZQ+5C7aLOEKW2TwUf6swuYv7elZEVaOihydNUKP5HW
X5xE4Z5onMTh/KJ+v+0orb5YKH2v3tS4CsScHn/Pm/AvTZFTA8a5Nl+4v+Wzpf3C
nF9wgi0f2C0hVjVgfBloUH30AFpvbpRyp+xRV43oN1cQexVpPrHVqafeRl93ksLA
igPR5npY4MJTuHapGhojWjUsV2mbTtG4yIPX45pDpI+OFTH1kxbTlVpr/XSoT4GK
OohMW46e/YOXfJs8YDAXCXyVMNhnPR7GBWeV9FKzWgRMSNPZ6C3ScFHPIhnBbanx
IyLFK4Dzr79jSTsbDsalc026S5lmi/3Biw9bXDnuthKSOzvy9O/XbPRldivEP94U
PL/i6hDcKRL1c0b3hqE8fjWNhF1hFh7VoCmB4vooWr495VEDPBfatFOwO/ixjiW/
HoD5wgRaSoLtzpSI5Jy82sY9ZiXGm6gHJkyEF73k1QFsZijke70AMKbqPA6YfHoq
+J0DbbLNzCQkU/q6Lzl6c/bUnf4FSJaYK5SOB4sHuFFesU+kq2uGYci3UCzz0EYZ
tLIPQRqXL44Om7di+1qnV5dtyTdPMw7q+lJ4UTHjUmNlNCTu9LyYCeKXAgYnMr0y
BwqKSLXnx7uh0p9K+nyEoLOYYGL/zhPoXD6Yw+wnJt6uGi7Ctooxvtn6uSXVT4qu
HC9rM9X1KQZuxfUZvxPoFmGjRp8H/dvGcfnrvo9ECBQeLRN5rdy5boe4hl811GON
lyMxucpcsaYdZSYfmAnFOCw3ohzxgQXXrTZfiG9zKz6WEuBaWjrn1hT457aWzWOx
zPA5t246Xr6eoqE/Ldlmm8XabI1GM65dl7Rx22upQzT55/J16l5unxh9NKleW/yJ
oHF8VFwRgtzpoKhHgk7uOvq59aezGFB6dgZZvY+8Pj7z8wMSurVhXnNx3/WRoroQ
8J1LBO+T4JbV5J3AlAQWLzYOp/dYWZVZqe9gO98sRyfV+qW1+/24jA1ga6xnqn6K
OfiVW5fuwPELFelRqFE96jEtcyjb/yfDci3AtcjF4z/ml2qQwaXdRXUY0rxmT3RF
H48BT3S3JxuIawDxE7pXmcFCrZnlV2pYT1RVLXrneV1flAJnWj4imrAbzM0ZW3gd
luaEQobQji6xuzNh3psvbX9JcPmJeAZhPe/ZsTxk4m7V4EBQtj+WlbkgZ9TocFqP
fG4/YJQdT9lCkaAhOjgMx2t7mlnetOhUSYTpvpVQvkTLdrILnn2Y2+J1qicTFvdg
HDV15xajp2WOkNpOBa1UYxMjCNdI6HV7ef1PYIJR+auwqjvj1iWanr+CvP8+nAoe
xVYbFzX/gPYNlSpiyWeEJK4uq/JYFqiaKl2XzFe8Qgm5RaE323Q+RXRMKDvJjQXY
Qd4nzYWXWkRx6l7w6RPWuI7DngBQkGxdu5gKRKfBnllW/IrpZdZOOeN/5kuSTucY
VNsuJS37XgXNRhN+Elz8h2RAQifzjZXp1OA0+63RNiFmTq1xj44TGAQ6kgUpXwXI
9RDUzc6nKqwAkIfm+QkGQt6GKVgTOZkReD8n+9vDc8sjmcZxdhia58zwIhuei219
YaEASkI7hGTFEP+O+KSCE6/x8xbWxd3WEVGpFqzCt3noMlCkXf3xaMKHVZZf8OOn
Ud7lt4iSwQzzHNLxLOnKWT2DYbpSwAht+wE8LCRzE/Kw06OWvdWSK8LQEDWayGyi
31ZkED0ugVniPfu6eHbbdI+Sll410a0mzlnqSkrVQt7MT3Ugb8m9ZGIR1jB2XZwZ
xDSglCSSbL5zt1Lpd54RUsMqOZtdE/2GrQtxhFsYCCVXTCM687PRKdjB+Vn5kZjS
uo6pXSQHiH4LfliuYnwi2C9i7/eEawVtX8xuGc8Qtt2HY8yuH6lRM/Mauk1exZCE
PYE6ROPVUrxovGfdmhQqLqvpgZ9okTeSaT5BjyrYP22Tu4VqRybIOaDXvXsHbWqV
wWHzGY2rRWMwZgKCwaT5i6EB45TSwo1Ve1KoN3wmSIdb6kWsa7oQY1riEa4UTRDB
V0JFZ0j7KXFX4mhNhuBAIKmbW0854EXAI9xUAP9byBHARQyFijvkAMu1V3kgGdFW
toukNTUuiXi5l4BMgVjK+DLVtHB6Z7RAYVYDCkgGGH7Mi8PHj6Zpy7u8/oSlAYgT
yzplp9JRHPvgrPr4JVCz5vmNQabOqY+rjfF7Glg/S1TINwfEmUGV1AcFrN4TiL/J
/F0I+8quLC1uX8QWKxBaSliVskypAgoU9yM36ku5oQCeXCSu6egxW1BY4xtVOjt7
TF/ynjLQbbmTCiS/gKT7XylSHaUM/JBNF4vBxPxl1/6+r1xc/mstzqVnfB25WVlS
3vwZELtG0kTDrYGphVXDokXrTqG/3lMW6Q466ITP3jbkBGeM0e7JBwzGWj+UIqDk
X96sk/M/15EilZeGB3xne+NZwHhwEycw/8dWiDFXVFXvNnB0SuY1RsLL1xXdUXr4
Vnb4if95talY5/ngaCpVaqieoQcTUKzya6yZNcIQkVGS958HuRDgrFMmMxeEQ/Cl
cuZOGfwEjpQQ/0dmki4LweTV3o77FP8enqY6g0SNpe51AZVxzM9Rvn2aK+6INhnu
hCGlldw+Y4Sc3tgt3WXKTi6eVzPHbKBtiabsfFlwsQPTRHwxzq63ed/nIICbeu9U
+41qKEh15PL4iHQVuwTG5HrMnojeO7oeBZHh3OE+JWF7DnPr95CQUWbvVCWj27AG
ghyrhU/gLIEZwMd+IlEgfUQMuWUYkpmd/ZmJgEyNTj6FR7WLvcrVOqdAEk05r1Yr
oiSNXXIlENf2g1SZLZindQyH9s1bXZD7Q2TF11iZFPXJk2pkaAHTAG1RQfYxQunf
bisrNrFma4jrMsOhbNqlXvLN1G7ZTOghNlWr0JFtgho4ZijBCg2ahr05bm/R4+mO
FHLZqTVaJwdUl60TJQqbw+0QsWVbLIFheauK6LokREyUvsaNPabskUqyJ9BqmhoI
2FzWRim9T9YgEeNrHqAahwOSTI1I109xvQhZ5Paegu/1gx1UXQCaedGlyMV0RmnB
SirZnTK7eiqpTLzVqGfZJ4cUnfDq5tmKdqSuJljHyDqNxAUjOVWJABC8qB6gFwC/
2cVPO+LRiGPtPTb4Pmh5JS094T/hK6SFUpKyGLaIOkwJUpncFtoTJ6PQYzZ08ouz
huINzWC7xS6QG7kaj1KFWeilLw8cnI4pYFCdisH43sUsvv3gUvjuJybu5/HtRVVv
YTc9UQueW3Qqz82F0LUjwz0a20/qyvA9vtizLMPna8/8pbPK/WiW1JaH7zaS/7A3
8XcQLRFGc5jxc5HBKMma923722Vf3vEiSrbXM1ZJclFVvAk/XIPsCJEPQ92o+wIJ
3SXl37dz0srRVbzhI4kvMT+fAW/r/noleMhlLajCKINWHZXY40Q/Rv9kViGrI3e8
G1O/hxT2m8wSiBUOwxU0zqniZSdhlwBtb/KNL4GuOzMfdd1DpOtZU8cZOSnuK6Bj
0vzID5JgCgPCjyM9mfybkTsfX0UK3NERxkIGd4nS3WO/X4rv/+83ySfOuDymkHKw
RxQPfC/HxOBQNfvAqeySfozyhA7E3sx3/JF2xIPXeoy4QkuYgEEVyrSWdvjMjdug
5Fmf9vk8iah588O2evWsqJPUVTOR57QyBcyfUezFw2x0Hj2+At55a13RA3XAN+a2
rMu936ppgPvvTsqiId+mWJ24dbGqgmW0QbOmERQoA96MhDJklwtiOA3Ivc8xTes7
+oKY+nZLngo1oWVhdPbGmaKPY/pce0gl5u4GDEapSUFj8erHl/wNsn3vxd4wppUW
5QScJY30g+lycBWXhoWherZCaS+RQ3egEPkmVuec/ecs6c1c8iVa9b8jPtOSuylo
WK1DkWdZuHAenD/V7NC0XZy2OqA1hD7SULa+cy50yTIUyzHtZ9TFgTgBxdg0fiTl
UwwjoFqvH8Py+7ZiBbhiPKHQfnJW/LgjTn+TdljNHn8i4Ue8a54TljXQmSdqIkgD
1LaOBhvUcG8sNETQbNc2p6JyZWSrt3yvB1gjb++mzN8V4XTAet7qfKnAdxOm0EDt
kxQvoQRQKwPEbc60R5iYgs6gKEHFY80blv3ln4xV3Z9wT7pnjHsXqzORsjXIRc/f
sCZ9BcuLLjsNU4p+z1saFyWiTI6b1yBJTgDo38NwdyX6MBMYnqeGnHjCstfgTyQF
Y3xiMbctjqHZ/3oI6hFVsmbRUm+pa8oK+6IHtXFp+7EKixZ1kW2dMCZGlvfggY0v
5UnRVbGpRG2mcbXhKI9ThDFE1J+wzroL2DJTwZaeM1clMdXe+EGTHnFf6DuXJKxa
ECYZouMh4foIRwxLH5387HsK8y5LkFQjFpCd4sENn0qz7cEGUiVjmiibQIyCqZvB
iZHPAKhKKYMm5HfdmJuCNpQ/fFIoc6kuMKDkaua/4N83d6uugRy9N4JqyNsNLi4D
gGV0KWYbkqxteobOJ5mJC7TbbIuB2NqRsCM95It+h/zU0rrzMHCS/rA7BBOkLV4y
lxOiNy9P/RdhVPPKdYbXDi462hWwl1q5w7kRYvsCF2SzzHJRNwEFE8/YPAIZxcWH
w3ACuH+Gm8WhRzwdl2CLoKSeBVk8hinueXHcGBl+RRR1vR+avxl2j3OzCWyuqo15
1uGkppjAliYiAiADtjOF079QSZjf063I7aRnXjjFAiesCwm6XIQt6wV6KibVsIVS
NzitmJKdRBvgIvArh+ApRLjd9oHIxFfdOOP6hW56OhC4dtjevLmAUUruRUaKZsFi
VogPjyowu6oThmcs2ib16ogAD67akuB2Q9J6J7nyJEZQQkHPvVq67RWtJpk2EV1P
zEc6G9Un6w5esCBuMRbWrpR5jGlAykPv7lhsiybcd87IbR1yEv3W7g5zP8Qj78Lz
CDF1NqsT7SUk72Sewex/dp9eDashdY73ZVuRVPzZ+D02YaAtUTCgIo7eM/za13nY
1ywfNn4E/OqOCYs8uKVl8lJFwWIlGmFn+4Lslay0JCzCAIYSdYqSDASvPxQlznoL
AM6F9OROHZo6X3EeFK5R4yV/iRVjgokV3/mt9Mx8o4d4I+YwQiIykYoxKIwbcQLo
EhFFqEABQ9n3IOFoks4tPAQaLwJcfGS4EEz0305m/3KVIw92/YdgWaHJK+SnBl1y
xS2XFAltTQ/kCehWfayHQ/IsnLeaQ6tdMawfHJe9qEy9peDwB6ISrgryBDqqE3YP
y6rXVYRCq8ngPjSyvKkXdoHxQAqDtUwgm8zd8BoESIHJ2TWIqo217yzYwLLmr1aU
/tFaq9NdI4PwV/KRZOly8rL8aBWp0/ZgLnOLzCcDxQNmFggRyQlGcjUO7CUi4vB5
FXKejOIqUkK3JvI9mM6/eVWX0/jy7f+99y7adGSujRsiy7NlTBeIoBqjeIphlEHY
McjgUlQTKYZf7ALtxxjyeJt8hZioilupRtsfOUDYX7U2q964P/mPX0OUPRlh5UNY
RpioIDI22vUK4tEjtPVeWhabFGfo/CxRfwyj6j2tQlf9Cdta7d0+vbGae6hWl6RS
qeJGeivM9gKy/TVjonZkiaafW6j9fSk7QTaNd1328SiQ8Rqn3xTGJ+3F5O1R5PfU
VbwVw3vxR//mCyUIc5I6psrzqvEVzgQnt+yRvOURZ9L4Caaa35ryA8bJSD2oikEY
7a8XqyZAqPhEI2lvwfOZSgkJM6muCDPcZHEZhwE72CSvgc2Sh4Ura1Ne8Xauf7+a
t9hFf62g85oEI/UlVt5wrCc0wXApBXWvaWBYVTd+Lxi9+VHNNiN0xQJFkvIrR1n6
vR3ATrsAbeF3UHuEfFZ20uB8rYBMoGb4ondiGgSvWSmHzeAYXuQ1X9F9vXt1pLrZ
tzukSZu7aFEqoFcbPLqit4Lx9pYUSLe3KNjrU1Rca77UOmb1cP2icc32a7PUNmFV
Io3t00/Z6IVPFsC/BZ/FCbqGxw69WoyuVAkzYl38gDpFdtd4+oLv7t7Qd3I80jrY
dd/VdZfu72IU3t0jdSrNP2zE5zZLdTK6TlIxIwYJuyEJquC+fOu6KApnwHKYXRoD
EB7LMbiVkcKSH5KzUGPZwfNii8vpZ7pO/d50zMsJT2WPKiT5uvJsggPNHT3hUb9y
v2zLyPlQkftOqAjdHSf+NTrS0v9H9YdfaZf2rmF17qdyn/wTBTFFyPrFqeE15Uq0
RmYQ/hmmtCSMmKkvAo/IaboroemsQ3KsEZGAPRSI1Q1uje3ZTKuZpF6fEdGPgiEB
FpjNg9Po6iHnr1mxcXkMFsScxu7pAP95gjyg3XTTsrt+LVWJvpZwMhZ+UNXhS2V5
+rnV7PTHpDoC2SXUEFcpLiLsgb5ESdkQeoI2+ZNMtD6p9bjIoxZ/AIoJHHRdYYTI
haMm4kvwqDYuR6BxDaKEk0j6TV+WPCEP4wwCbgSYJJKueXvOXwEnldJsgw94EXr7
scc+kK1nUX6HcgVr3zYeh7cxEf7qaoJBpTgmUMSKdq7vZXiZGPeYckwNSd53+1Ho
OBMiyVcZl0u8gvWT1f67wIcJw6CiAeGEJsiwC45bU97mGLlAuPp5Us2LZVcYIG3g
dJJs1B8cMlKeMqf5dE/AyazttQnnJ9+9SgWBRH/w+1jg6Qg06bXXTdk4YVicid3w
i8lQl2NpXkLlM9gjU6k8HqbG7E0Dw/t4i+Z2XYyEIUUXXqoNYAFdO3cp+UlLF7IF
tXo5h9vn4Q+VYLJbgYtEX/mIeMO+pWF0559ug/ayuyU/UuRKPDb/QLrxo9Jn7wZ8
/hNlN0BzfyZ9n4UmKNFfBd8eIVN05sHabS2zuz3eScuCdpnuRYbzAR3FmUaA8NY+
5FhwKMmkRvVPlvqtTPcCBwQQmE7/DI+Wfa8A5jiZYnEuGm1xj8NNTeFbTcQno2A9
1sV6veNivIbgU57jd0x2ugmJSmnB/hxb+VgBGDFchhj+T6WwSIE3iTYirC84dJCq
yEh60bD5ok8is8QL6QCCuTTaYamVYTVFjKt8MdbfTaFq+dmsOa27RCqiH/KZwYih
ftkgU9YqNPBM0YwPj8ba8gRIhChwqcDB4TpDstvpvHyQiyKgTlDAHq111La24cWx
5DDz7KekGS83+74f5b4GpWWNDtIN1hC149rHXr/iZ4cBVaquL16rxJv6cIp07bvU
zNKW5ZigEcNVgme1Wlth8cKv7GtDrHwU7z9DVizIs8+1piu5GzpNntKB7Xe35iSC
IW3b00TOf/ZMxhCJOFnrrzIc9HHW8BEH4SsvLnWK35zl2bKsI0bh2y0M/TWVNrT/
fMnooq99mrZeu8OpIEhW0R4dRFMN4v9eifXbN36pTnn1LIhqM16ihgny/oEs/CJH
5x1cBOIEeBiaoqJiOt6BxCWQNuADGj7JVICoRZIrL+E832oIKp5Dtw1iDWOgS8l6
zi6fKLN+Yf45Ixq56dQ7Sh2ps394ulbW+5zKuDqRVIFMZ+og/Yc2+QC4OdcQArNy
9cjVKc3gfGMSZKDyumCICx/nlTIrnr7ORVGjoM5JVbbVOGj/4UojP/ZAXdriNSj4
RI97Kma1GVXLrI0pOhJKPQWMCzuaks2hzeCyQorUrX6U+8djxUR4rWeh91fXHwyq
fzyCCr7oJve0wOU+UbQo+nxuGTJGYRagZhI2IKU23xoDgt7ABPuGkMiMT3YyR00m
mht0OGYQNYyzhA6RdbhXxFmnBET2UUM0E3W9/K4NSbmgYN2abl870xPsEcxQgffm
Q8P7VjPtmr0qw/wtyMBrEqjaeupLAED5mtrnsDj3GqPG9WlEYkleRPaPKUDRNgQE
N4F7k5XndYHs9nVSiNh0K4jEwQgHfmJslVuBajR7cxPz1mJ03oCJADtqxKur9mBb
EurI7Vkh3RnfTJ2JcxdqY97PXpjhk8miArkEySRA0bPafqJNvyq4GaZvBm4yUE2b
8ZvTzyc/RPDZONXVPVd0/xGtKWrInT5rHEKuwkFdAkT1Jip0PpuhANp2Ih22aZjU
Hrwn8wciczuCBswAWSv44f/KRGY7VAo+eq2xhEN88iWmjLFyeCCgvQ3Li4D3GjDA
tpVMCS+Xcy7JR0krW6FLc2X8/1Dzm3aSLjiHFNPIn2ViptIo2LssY3+6iULCh1H1
nYIpMOjX9AkPEzEiA6EFx9iM4Di8mgV9F2CiMd6TvkMajm9lc1ZDIghWEY/w62AT
2qVYU6DKmlKoNlkyuGwqF54YIcRIlzM2z0vOjQPqxq/dFb/VvaJVSz49TJwZyIw7
5ZbSG0Z5ASWsWsySIghpvl0NEXiR/glDg5ApaOIGS/YrO2q7qpHY9E60MaLSObOw
AJDA69x6GzkfgbCH1TCdDRTFTbAg5r55Yv6/86oLcAMWlatcXdcoB576vGobs1jw
zS2iAQQt/nVL/4CIm1d4Cp/YpES3yD3ql2X0cKZsOeyHBKV5DYGbfpWMLx9TpIxf
Ln6ISkMQz03CTvnvnxHf+GSb8oalynkj42jwgI6owm3FziKm2cAkoxYH0PVuf4SR
PR41WQYsGr1UG/gm9ntrE8kDzS7bDi2nKLz0SDiHxwZ5ndTnHAwqGDI5S8oJW6kj
MMq+1zTdMoylfYe/LI2KXxGha0FLdc/ot5WR6QFEK2ZMAPYb7m7CSjeT69vQDM3k
I5iy9hC6rWyZf8poN0DoDEswVKjAXk70049KdVyyGa6uDgoLOW8jot51RAw8sHkf
MjFHFx34vmUqEuWtFhUGjbAKxtLZiW95oEuoYb7ZkN8/mtFgc8vVeVofGpL3eUi6
mk4lKnc70D4lA8NbtXul+dRgfg894mApGoMznoahO5Bc47an3SbvbW7Gl0TToEoP
L23mPCb6yBtt1iaa7jVTHbfm0AN2T6yBiyF3Wcxbn0zg4Yt+rPgNcSCzcwXticFL
MhuWBAFohYW93FdeaZSUONv4asASe6fNPYZSL8Ik0MDipcN0RP40gV352GinaBSM
tJ18nZRRDeZaWs0vn0RYeKhx1a6pZ9D6O0BIywnB+hE+Pq5B82mCTTCOKt8WmLLI
nB0ULOsByqW+Pj4+cGwpIX0+wCfL3zHbQEHaJONj3IeqxegP/BecnL2IStyl0iqI
NrRQXsq8BfAyFiO5u7iljkr+hy1VFPq0AJ7SalOlmQdlvH2dQTHRJic3Meht31YP
C9U6zZvrg0SYmCmDw88uwvUOnWMEqSR7fzzrLmSCX+UQn/ppmfjvI4zutqNuFC5X
a04ziIfEaCofgD/uQ/jb2THRoA+3yBBnivLzyf+uI9eNyvMn6WZt5zIYwgsDlqbG
W3BxqFRFlALLPy1Ryc6fCbvy06OmFTtkgnR9Zs5XbXtpnCNZMDZd6jjQgaOY0xxM
eBtP//GzZwzQ8+oyvfzDNKjS14nD5zhNBTLcp46BxLyndvAB9+2rFDugrFJh+sz7
YFDVRHfkkTzoN2bBGQ1UnbWZUKrlwaqfTfkwq72MonsJMj7oOT3UN5OSftugWZB0
zeuCHvHzJRlmOjEfVqGynHvOQQ2fX+tOMYZUZ9XakT9IOtqKTchCuAZqCvC1OytR
eGP9PkWZ09yiR2h0fOcML3vNO7jr9ey5wPfxEk2ps1ALYle5xSrto/T8xwrv/cRR
uFzq1TDGMu68HGORVFbCIwfg3i018SEtcQkujiMGVRxVSOlG899KxyIZm3qiH/o7
K+/6qoET7CSlL1XZq7QZCvKH7lDRQpSNlHDPe0LAXJKP+aPokrftKjnIcFAd7+e4
Qcu364QnDVuiniWqDkIL7fUBRrXgiXpcY/LsTA4IM3xQBpHIGW8jAJXrRZhG+SLy
M/lEnORul9zC3tmsCiUGSEgY4ZA/mmmX2QycHJV6FvpueUnfdEhpjkf1euVdwKk+
+XyPzXmswkl448sV1aKRKkkJkAUHRRMBasZSTF4T1iM/rbtWw1G9lE7Q2jpyKTVR
9dv5U6iS7O0DPV6zZleul3fA1skX08IRTUNxXMtAhTJC3fofbFfq5TB+IzY9vUVh
ip+vyk6fgEE/fQrWjaJdzg4C92396CgxgqXXoVmDUtMQEZMO6O9fKxY/GjgbQhjf
C7V/MQfvPWJ82RYsY9IxxIkxa2j10Z8xZ9Hvl5u+wnrxSFj7HBI+8L5q7Q6oqaaZ
hbnqr2LJ2tHZHsFyV+O1YtNQqtI35Cxi0X96cPLNn+jF8V1J2Pb+NnnQEKxMVSkt
5ECXWj0icd8xCVCDVxto38qyyTFaiX03mQn6dPKibSoLZuE7H5Lf5FpG4l5T2Kuw
Wp46CVqgzsEMyyyVw7zJieSykCwM/zKk+VGdg/VGqd5zcG+Hii/6WTu2UfKWDDT4
/noCurrSupH4qaTglzsaVh+73caIbksSAQl3+qM7loI3jOgKcnNaTWXEeY/OYifA
xzVZn+GHU+kSvECWkWTPKgXWTPOi6DoPfS1GdW+8OPoOhBqUREhJy/Xu5gI6ORMW
61bQQkkRhFwdI/ixOlWWIxtnRwKykLItAbYQ0Y1e33orHbBW9rRgp+d7xxVcFa5G
g8Fbn9zYE20CyyUxhpNpUimoXohTlwX7XLZDAUctz9gCy9ClmBVJFXe0UmTO+CV2
LrOYAGqY2KXGvx22QpjYHN/PD9xNiE2H/bNzEbQ/l1u9Z4/dehv4RiIvJ19s4yrS
4wvq3ez3hers87dcr3lOWofMz4d4GXpmUJnNAuDF1x0vWUSVPQFRacT6/F9jEs9r
pP269TbtKVsLbQ2lJUnKezfXfstt/QWwcoG+waCimzwPLA4q0EYIHiWcYkXPXkuQ
iPzFvTrdE0/k4IirwdYVsN/UXL0KH8LiwaESnNxPG+AAyu0itFJxtRC5/Jb6JeCw
b5WLncmLQlkxY2yEO2oHfhMXteVwv02Y1OGl8F26ekQOJX7MN2vCeZTggTSp+bDB
DpoPR5Y+rfaEug4B3l2D7VgWPETAhWJ9qrqiSDpSGZUUEajBrr0c3Ckojirp6ipf
DrIbBP43vqaciw+xVoZJAC7I0CZP1oGvVJtpbjvd1NznkpKhc5nVb0hUAmqvos5R
FGGmRnjGQQWZJzexG2aBHRX2iImUvSDeQnXHyCeF8Wc+NkD+CdPw+cbwS7NT0gZ8
uOSF3QM5lNHi5QtK2d0wIUP4t8Pf4LYIch90a5iFTnhqiIay0zgg2mgkQ2TDWOBz
VzoDvPB6MWA6uWd5n2xKLVe9aZSK7tMChNKuwN5UL7Fmc5blrXDLEFoIhuzhvYrk
FyK1BPeAksIMNcwe1A/ncJcBWdaeWQS5hyKh/o+jzdC+YlK9eEdcOLRPzBTbJLEn
IE5y3yQTvHPqA+tZ6A8xZa5315/3F4cfRZ5K8Gyc+ZJZy2QNZDVsmSSCIXq6ZOeh
E7xRQVVYWJRWLQVi4HyjxE8yFuArNrYUa2aiWLErmAWc8OEh/LMyKlDzWi2CYpE9
foytm4zsWd3AzOd+mDrkeSE3UtrHR99PUAaJhlMmAxS7ADTk5pafFkPLVj62epnd
SJik4ongLHrWUXa8CcJqnp41ibyhrcfKgN2DBwnuNDDA/rtLwT4VHFhw64TO6ERd
AEE8Zgiw6DcUSRfZ1gveL4xaZhdCqHZKfbvjR6N/ppPIzo1dg/WYVJ6eoI++LjL9
3+Ng/r2VMHltfsFVVuNZAnqsQiBrcBZmsJnKO5Xaol2qeyrodnL2pPSn74f3Rk30
d15kaayqzQBMYSN2VKFXGcwNYS2PG07F0WJQmjzdORnqB7yo3s1jf9Tj2lkyC79D
YaMCHjZktUcSfJfgKNdl+CCCMVFafIz+hGUnWeRAeopdE+R5ize3CqHm3GRMAqsA
AwpKcQ/INcVNc4ijFznpLulSOlg9katpyGK/yx7b+e8cynNrETCzjny0jO3TQKAs
UD7MEgVrL0rcC7MkvmXSh6B+CmvCoT4CXhsM+cFwCxkYIUGSAL6WQ9PWrf656Qak
t4//Ei0YOhqcs3vLznqEhUmKZ5S0iXl2mYzZcRMW/Oxpc2JUlU+Gv+anTCP0bMPP
ocvKqMwGmNeOrgg81qTszar0gu1J2NCvvKYRs0+0VL79n4n9IsMIrh8+Fq8fOgFQ
Sthy036s0QN+KY/e2INRbq9UzPVqDxRSQlDN1JxnYUPY2nq7K3jQkc1LKB5mLELP
+Puc45WJMyO6opDgIzDyaVApLJtev2cg0/ELhElqHym2KEHLjmN9CiGi5DOgUD/o
e5PXJ5xdm9nN3ZI374kqSjsUpsH9gtD+iHx4YWZjevZD5NynfarTFBV7EaOh/9jF
hHpwcxu+4t++yJxkoVN3tKKBLd8terlQOP+qfzETeZ7x6ANiJmFw3G3YKxqDGPSx
rC/pHrgXafpJ4DlBh70dZlhhDxSu7R7OB8X8NuTJyKH3GeDkvxa/6XiQ4gipgU1/
RRCm6mSukbMhVlpvupniVW69X7xxMUWWflkSuUNE74gfVQendYfw2mXpcdfQOW6w
5rwr880c0W/+WLRQA1FO1p0utmI6SmROm4GSB6FM6R7zBFFAIdfkoxWqYXj/Fgtd
FOI0vV4d7Ug78vVBxu8B0VPndKh/wIdcz90LTsmxy6yOVriEhXuEhJv+GoQieRsR
PNafdP0slie92RTv1PGX9TlvZclIl6U7bnYtCs77SLRuNlOMN2Ptl89PJRVOu2Ea
nMlQaqGyfBOUkPgJsNmbMoVaolhc39wDNsy7vDi4EE0K43xXYduP5/xSf+utEt3d
UMIn3gEy/tu5zSJtt8unjlqr1kdqxRBIvPDIwTnW94P/nfjJE+cBRqEvks8E0lPR
57Est1CQ95wDX5TbW0DXhyOj50P56WBiNHn38X4/m5xHorE6wQiyRiJLCJQ+zjyx
cMQMxJZvamRj44mMfJjJH2inYO6stWhc/pH2RRjzvyrfj5rAPwmMP9acs2Izjk7C
BUebh3ruK7v9Ocv7siQMy0dCRQs9zkidA2z0RK2++KFBjyp8c7WioV/tEwFPR1bs
Ubb2ohffIMekRsn7y0D0pnSOD+lVDy3gal6e3LvjeVTX0fOGkxSeV4vT4gi36n5d
HHqfN38OCSUgUSW9ab7DX9q1OgsqTPo3Gk3zkrSPSnwWn468zmXP3vC6TsHy+v/1
nLfKh/kCEjRTCtTkaYtyJ4/Iej1mIaSqdFo4SZgwZGA2vtL78GX4xM+dJvYf2Rrt
YGmnTRC+VkH6XGIgdm6R0KHS4TcUTPpl2+XPl9dswDEEhfYTXtoH4ItGHsspIDH7
F6o7LSp7/K2rQ8JEOc4sEvf2Yt061AbXLnHOnHj7gLrKcvD/11eXq5a8Az6AcKBz
4b8GczgoCGrJHyIvMPRH/X6kjFEJk/iNfRrNY28//dloGV2MSEP3WRyD116G+zSw
qvzmkBU+oNjFfDUP61c68z2yTgNUQc5RwYkjOP1+b05tzA1mUD9o/VG/7KDjJBZN
XbXxnrsPU0yYlq3v4UHd78pJbl8G4nwu4s/42rhHoX/oK0nlNiVf2DbizBsWVCe8
Z2qzAIMgKQP3kn4p3QCQVo4eKaWZPD7+1Rnpi17PXWm+sAtXhHpyHq1doTHJV4C9
88Xz7QUvUkPEOFg37zK752Ff7kBXNh35mvZY3w9skWXiRPMGrYBhZf11vmAYRJPF
KgKoIgnNcJYqj0CJhgghvhMy34MDrRnJjIJPOyb5/RizBAzSareOnOi+fU25E3qu
KNu7NrXbBTrGXPIqORGUBj1mLhSk5AfzPI1F2UpJP/yQCEHI7ySca30VSAUbcSgJ
CFH4GAa5A3ftj/0jaxZuo288LyN2r5xdRW/RqAsoblq2gPLxLgZYB393AFQvsGwd
xn6eKclCFO3d9i1/jHLMDvFOCMhxLS8X/6hD3PPbcy1aG8+pkChwy4Aj9vu5nkFT
vxgGqVUWTTpN3TdiSdOP1k+8kxCWFcOjMMErYCbbGU2CDW7O+gA0TbcXsoV+yDUf
gAEdnaU/re6RPAHkFdOYI+EsayGpREZv2eGI7xsZ5Pb2WDiBI1jrpcrt8qVymGSa
+AES8bo0HAfIK1ngZA8Qo+vAvkQ49XhiVnNZhcAMMQPXcyQaMPk5DkzgHbpgdQKR
Y+HsOoXzLtXmVG+TDVK6+/HeNGCmVDka2W91BgK2xDZi1xaz8hqVAfE2VhGQw/3W
sd0mL1vfnXCyAHr1X5dQar5NisjfT8OWo2P9YO4mWavzMkGYZyph7o4YFiVr/ZuW
PUW7vUmMC/wRVdPl4DC0newsDv4uudolTE42yQOhATbUI4OSrk8LzUTDfmCLLI1Q
ynUvwtkfvzpE99+rNrYcT8mPz2R7oaBbCruAaCSM4waq6a/NEPRBiz8E6SlIjLSY
sP5HXxfo+uZBZYgqTZwSv4kM4wnIqvcKEB2oEhaGb3VozIPFQsu7rjHPcsSzsZfd
5BPQ8Md8whiCKVIGG8VOCT8DNM88VhsGy5Zr4Gsc/iXqU1+cozRFvrH42w43wCCp
pHxh/M40CV4EfRSua+BZh0BvNB4gYr16ItXwocNy1TulkJp7CXX5YQbTbL3gJmNx
HOyMuAhX28BJfoQFlB4r9LJ7rmVn9CJjBqZERJmSoVjeSRF/Y0Z8PAY0QnQ+zHR0
q4xAWs75lCJl5qoiF36xRfDS0hmdVXGFXJr59EJq+pKUNb/ck1HUoQCq2DpPbiTa
baoM0iSIgkhUfx/HYhjt5UcoKuZy4vEaM3wpEQDekirHFSu4yECiertLu+bssEGM
D327qDHuW4zjk2azcEaEiQTVNYyTVLOvCLzL7pvl9WyIGZ7F3lAGDa8oN/AcTuuE
fVwJ1ztZpXGHXnk+yoVjhYKen879zSSMNLaY+++vrdvNBk+ikC4yU/o5OVTSYMvP
sd59x6ZIWqoOgwn3+gzgXkleFQ6CHw/apeVOl1ZfTuyxSM69HcfqDr2VHghtkiSK
H7VnmcLB82Pey175LbAZO1Y0X/tu0lWjporndLWFSdJTJcN8nDIudn2h2xdMkqTm
+Gfx1dmx7a4XR62bamEifX00Syfdp1wlz1EK01Qi08J+cTrE3auKFFURyMFjTy3X
b8XUihNT/jEMW1uI/m6knCkAL9ftSlX1gpYyrH6GK/fPx/yxCTBZCAz2AVssy/8k
b0rJvaYC8/yar+e8LB4t7Im/GBh6UH8XJGqBbSKNebzxaruet+p5hy8OUmDx5aan
GTnFtZEZsbqnb7I/QHI/mv/9nR0VpcQJM7VMBorDDpdDBIT21mC37w7KLJLevljk
vTlA1HEJYed5715sBneMmx4fRXrRaAoFqR2a6nE5b/owoPXkak73QG7OURBONRrw
TOB1/j0+vaptLHmcKFRY8LPDLofIK7nGlhiO/djv4cVnvKTJpO6Fr/Ild1d8f7aq
qefzkX5cEiFIKE4P6ayTxl7ufhQKUlUGxC3CUD/KuUzkCmsHO6Qccg3UauuneZCQ
ei+pjsMcHYGHfGvxzVhIrX7OzwbJ3A4lLqUgGgFQtadBcqzPE2qJsT5+eQSuQemy
ZTBQ3X/69ZZ/IjoUh4cMWDZp9LvaiXojKjrg3DsqyAHf81dzHweyjU1zKQxg3uO8
3ZtrRmo0RWRtiqnb3fxjDNrs72m8E1eOi2g9lZ59Z5ixoUu9vVndm7OZkuaCLBM8
LqcOp5g40F88gyoBoMey/aAANhpkydV4cA6yTANvFa+iDU0XTUAV/AIYpMDv/1Jo
rp5VP3y5SJdNOeBVp4ZCnh+Ip4bQdlco7g6voONAYYuzbaVD+vF+DtXLcmXgpmE9
MpbryHu9gUWjm/sbKPLsAqbrWH4AWnemJZqX53ryu3Fx6Nkd2qlg5qHV3jLKfT6X
WLPmlmA4bnsJ+IBHbKaT44spGmxWZMahFwr7TI7T6imGdzUqf6/o6M/ej+a4OkYM
QilJZBXd4GM3GgiIq01FWlHVQYTcaPHU5NRQAOgBAd86SqMGkQgPHJGJNgn444NU
9MpXUcpXjc+m5d/woFaeUiLFnAbUOG2Ul8AoDxyDzYQQP18FH6+uVTDFXn9DH2pU
2e6v5k1ekvD0Gol58OOTbFcknvm2rqxdO5nR9OV+KIDrFwdkKRBxtuOeb5xkC9AQ
vD+Yc/dmXggA8IAD212S6GCjf4rWS9s3Lle5yFG3rYNN2HYD/aIhaBc02z65KoVc
fgAf2n7TZGxCqyRAb1OPjjmkh8/IMnzcmVeFaboJTmgiFqAO3VkJe9mjnIEDm5Kg
SYDER0Hx9FIwC8xD43wNeJzolWt2+vwBf+WdcekLshZ4o8ObNVYXuk6dsCNRjPL6
KkSmXwHvo7N2bf4/9yVUPhOR6H8hul7Iakcx6AF6sQJBl1dgzmG8LOe3AYci3e5A
OBh1n01Ng+uTkaf1mL5LcL7Nssx59ca0+RkoB2Ln08I2V9JYPoGXK/RWxkRmTZGT
Ms/S1O0c+ePpZ+jQfnD2SqDROsonw5ropteoXUc6IEU3IzWmlFjAM355qNsgB0m5
ja1lgJcEcOYhkKeFJ1qWxDvalMVyzH75mb25/l/Cj6T69vYlzYN3x5rn0WxkPZhb
Vn8Xr9u1w0JAJ/XSW64X51cbmk++SfFBd3Hilti4+p/gyRrkvRH1g9FnwKBq/C9+
VIEbEokDiLyRiqL7liZlDyrjY3/JC9uaTdg8CP9WzunWjPltkkZQ8LxKj0juUje2
WIMeEFC8CnpMtWZloue0IwbcCAUVCb/Ks9tPUcPhCCQGkb1wftn8QA30FEvD9fOb
TOKp2E3j0s33S/tWFjGSoHop83+Ju75fyssiNdGY93hytXA5nntC6/tHNwTSiILe
0c3SSJLhwttCSrDn2rMXU471cUuL8h6VYdVMB61p0r/kGr8t+14z+/pMdrdkssMQ
BVB5QZNtVrR+7/H9m0rBrFBAk1qL6kQYUKSKT1Pglgsvq4wS3wqPhl9N9DJr7AEV
kVMFZuXi+mAq3+J3/8fX/CAESAKlLenoOf01eellCUbP1PWzRWFzNQ471eCJmRbO
ZBUErdMzGNxFovNZRc9L6tYGP85Pm9w6n0siMIBvyuINAyAaQpzznrPro9/1djcF
qEaTWuEGWmaRpvWa9W9v9smrl61U2ezWJ+Of/0BVHWpWwwUwtQrKFYpXXZRrg3Pl
skbj1L42lRdvNfINHtF2JEpwpO9hAWCxx2octq2177KbqrrinRpJ8Z/VqnZG1V3q
a1fSO7qyI1e65/Gdk5vIkVhoCSX2IrAEEPoc5bJ/gLSNzSBwrnKuRgZCsRmity9b
Z7O71fWOjiq6NGUrKfguCC0jslk+NR9CP3Zym3F+rJhas278f/HdDLOFqCgtxnj2
82WEdOVtgWOCYQfuFPjcC+rlmRVAvcLRao/DDn9IiAkIDZ2x7xeLnZjB4VzKZ1IA
Pzg9BlhPDsfsf7Ktqa8iyov6stgtUvkBslgknVeGxt6v7XXAU1ddRTrdvY3tyF80
/PsJPKYKwwZZaaI/sB8XRfcsC2YCFP7a5l1zr1D/4cj0ndDjidmoImIf+/T+gGLp
HradZu0QC0e6gWqDI2ySeg3BLx2hJ+Rfh+IqeJZjbM6NDQoPTmbRTvSudXvvDuCG
Mcg67X9NpWRI/EzzVRxr9mJUYqoSeHbn10bswUKi86qo15OdtECiygPk9uc0tFWR
FNQXwMVP3zLxEfrOGmOyLsCdxL7Eht1bCgwW9yJ0TVnACAEAKVgxDP12j1AcroyS
RotzpjuXHcjDXXc17DzFL/aEJZfF1ED8B8gMSSKmTnWomfVrqa2rkM9V0vvYRyXM
6k9kzhvCKx2NTubi+NPikvOCkwglCqH4Yc6LaH3kb9jwjZfbNo6lMsjw0wd7PyqS
DzWEtwbyuZBaZyuZw4Q4+LlFGKnh/3VIgdhlcHKKaf/inuDDTmQArhikwBPTsAZI
gkGGgI+dn5lqgiUUMpI/TG8xDd0gHFCRDnZddbkZaUJGVfvc8RBRUz5kcS7XdqNA
yOyJ+VzOFuM+vZuDKpMEITP2vNdLGwpjuumnXX3eliNpzZSGksVdgyEi3J6TvWJZ
PHufXm2vqe7TyhOCHF0tyFGLdJCzrh75uW6P/tet/KLgSjq/GiSlqvVbLfvqN7DW
pcRKPKWSJV9SnklAC++lIwmST6c0enKfBzfZukryXAZGJhhkbxLLmnHcf5WN8Yvo
iUiWWMzCofIUxDVNAwa5RL5I5DCiCCTF25A+BG9fypWl4XT5enlSH6zrke8rjL7e
EO4O7gQ/K1hpnVZ+iIMJ4m99T/qumC4LpPHZiJgNEHrdvGOlG6H60pRxFY3JSqyr
yja8S6hD6/xj21Ik6cq8IV4Z7/JzrGOQM3+G9BXNJH0X9olrixI3GSEMnqne5G7s
WlqXwXa8vwXzFb8Odk6CxOwYOCvUIVyzRuvAID3gOHQiGT1XnBMKcKaNNFe1I6hV
ZHhiFUkdVW7tnXPKsOxf/SlDdJyYN7POymzD+h2Oe6QGUR52yuv2fS5yqTTy3LTX
5V3gIAbSPxbddS71nbQlxt1TYSwgWKhlCKelhXepwnc9GdWgp4hUz43/suVzGsyC
6WIqSZi2vtYB7ArTt/EvaYN7KnW5j4ydMrPE5NqOZMIW+PnRZZDZtETgUgs3Zg51
VRtUzVvf7MqvTeez+GLy7LVi1tISfOckWKa2u8TEIpJpbIoT7t1eW56pyzxKabeS
xXPYERby66SkGK9zJ0rE7HkwK2dd1Cjq3owxXFsCGP8HvUWy2UFTdRuGVDoy4Q+F
3vZm4i6RWhJikxb2Vaba5EyW09pIlcWZHpUoTv/RQU3RriYeOKHeXbtrKUAEXgsj
NTLTGWZs356/qnaZw2/24HTFKsWpCrEJuaVRgl+KtEw4/o+rOTDw6z5xjIA2uSAZ
ArkBpONhidBrsciJA9KBsL++KybOJPHFTQef2c8/dZqFis09RKU7KrqEhtindalq
c7pxgTwORK4ADmSTgFVseupqvxvWGzNdW9UqCgQQdshW3CDkzzo6b2/1TIKdJKcN
zcA5C2OkM8ttZ4SkAtp1Er9gkYGuj8jcLEWVwehaJTis+Of8wEoEjbpsRgEzmozR
rEoelejdAwDcxfUwb4n8WsBrKDF8srdcCKQGJVjVbi30k4qkgPuYTc2CwTu4S6SP
ACfh6N3nWrpwYb6HJpsgiW/EcsDH3VY1U+flhd2QZrWmoGxeoN1G1b+qlu6hDW5W
p4xXi957rDYBEY2/K0YguqVssnVPqPa9Rl1gGPwjjfi6JUmvnZ5ktU8qln0R2qzs
nF3SFHE4r5R7ndfXV4TmlpdNiASLbVXbLOdKXqs56KPWh/E9yuGY2TA6FMNEavse
8pLi5bwmmJJLDL+kBi7aU3ErJzdcRB1ajKsvIBIgAya0vjzEUk8rVliFG4KMHq6e
ux8TdBrBowXUUi+6/+6RKTeb8W2pqhY1tna4unJAICTsd/CoiL7f1EGC/4BzwKvn
MJP6HtpHmr06gVnr4A/v5xfLgTIRUO8qw2sIlpgpg23u9tOXmvs8pNxvd2wO+wxd
foFSfypRzga9nVLux7cC7aAzjMu3pn63NNrnV4yK6/Rgh28IE4ZVw01wJXeGLWQq
VSuNLbuNdD+VnhG9q36he6wME+5xcQU7oT3atLZAY7qeXbHHz2nm0sIs9yfuq8ME
RxB96qfE1j/iIDSP1qPAiL3fBaUmCz/yWUhq3x0iXuL5bcUpA43RCko/iVAGj92R
vv3SVrog1/Ou25wTdRoDaqp+ZwIwUxQr7kEM7wQmI4DAoabSS+ybpmQNuy6WFpMq
8hLMFu02tDrNP/IhuzhY9NrhSskGNCIPf2EXpiYXmoa3zCZab977qfqB0rQKVUE/
0zntD86w9+RlEwodDBlNUZh1MGfIoR37V/gLqNsElKE3V2AyAd01MHUmLsET7pzB
GEGd+vfRTxc5d58qZZeZbuHrfRq+6AUf5pZU8birHX8WicLJzhXshsIXf2AGP+OB
v+sDbFW01uQpNe4B96MwumTOavcTL4UDX1qbRSIaP04f4e3LmnuJNAjYaqZJS1O2
Unl4tuChWZlbnaurHQKBHvwiCbk/FkVbTzmSF8HuVTn0YfrbmJbAfjtQYCuh5yWp
tJQ9P5Zw9io4eoxmAB+nCF0qj/FRoAHwokYMJuTd/XPZyBYXjKlm79/GBB6/RN4i
TX2QO+UegvtvdicfY0jRt3vpvOnHX0GCkMS0sNUmqK58qajZg1wT0tEq/yqxiVP+
XMsBFzBxsI5HcoS7Tx3iVXsZ9SsGSUHEQk8cUWW/6wHv2Vq7gmULWJRoRve54Man
rWNZJqFkXPDFuunqAKgHXxXaheQzonNxO5iEwAMctSLTphdpPma+5NYtaZiTsVW4
eXfPMhYhUK10IIzqOWal8cUS2NS7ReQt38YuZggDS7YjQdTQhR1LS4yWEj8RxEV6
dwLdYucgGtbx54pCIc7GB8ASItuKcEWNvi5sJgScCr6Cw7ONjbt1dfLgDLwjPyE9
R/BBAerggxRRrYR5CB0EQLOk5Dl+OmuT/tX7DAfRV0gDhcOB2EFuW+KbmRRukKdz
Q5LrP7fzV0/WVbY91SHww8uixKZRlT3znDkUV4ZbOi+B3RRqctYWGuv7+qIjmxq1
SaYTwFDE9+0Y2K9HVIIaFJNk9sdnbASApgMPOyBCWQhdUkx9Dy3DPklwi/lLcaqL
ZhDrL6Wdr1ttpN1t1EL6Z6gr+z678d9zZn27b1/m6B68GZIbyAN7AzUd+3iye0Gg
I9Yjort6cUefVe+Iie5GLoUOwoUKD4M2I3mbM8sDzHdzN9+CSe4rVxeaz5SPg5i5
CNdStdVMuBoSxjAiRFIxLrOwN2Z+PkysB1SXyfdjLzdvivkLCGU/S1R5/7+K11x2
dHLr1OJUoS4zNi7wz1Q5tMMB5naznmYraXfsOnIDQ4YinapjkoIe7jy9gYZrKb/2
vecTZl4axPoYOIycQUkFUyZ3DSTxSqd456iZ9x3iZ40KIkjm1zSYCn0iVMi1J85e
/L26bzKVvN3ISSH7bih+5LNIwRZ6c/U8SUGHQVyu8B3JoTub0iZ3ieD7ZV+SPGV1
7yZjwo2EAxlsBwZzbnqlQbbLcHgZ7C/OjgZWS7qgpYSNu/zFXqb3BfvVuNY+KacU
rHkh2k9CkWmRQ9Yp1baSDycqcOP2O3bHaNsBTM8zOq9/C3VGC+ahuf17D+ePLbVb
OZVOzFetjIWYXFC96gMZlMlQW3Nggjq9B2+oXYbIlU1ewF69Gzcg7BqY05IkuhJc
yWutzDZfwu9LyKuecZzpjarfexy/1i68vFm1QzummFjZ1zqvnlgQIuEJKUObeHIU
D+q7JeB1OFUhP0WH/9OKMw2nWYqW9jwPuqKjNIPMnSnNUC2q/oJc0tY41Z3fn3Tx
/xhQ8JBcRT8OxOiKC+g9sD0Fn4yyXCEmOcMpji6Z+XH1SVZF2YeoeAAITxHUkjKf
7TsmHhxtZbsSsooWVtbo3Cv7FS4r28E2c+g2MRYivDqqz3cCd0pc+Oeg5x5BOMw0
gLtH9cDCjnix4NeFbcQrn1ULi7WSVEL26SkSkz/ZhLIrNam6yJx3W1iqxBmGHydA
QVu1fp2Zp4t1bWz8dfEeZabPVjQO+sbPy4x/wCEcUr7gLkBquRXFX7dYKLiCNotG
tXAiIQlbSLKurWXho5yholGj+JxKUjrOHd7tO2IIh/YQFyGbSa4l2nC5/tT/HgQ6
l8+eVS9IdT1ANv2KYzPIne8NU5EQLyXB/xODb3t11z612G+p/tgpxdpwLOsEiVeb
MWsDkvcCjXfbLK339R99na2ithNG3z9R0KyF95Jn2+tKdUdqUPNYZYIBWCJs15dQ
gpIN3RiDB1yCQHLAGZlwmifOSPGtXB63fklQ6FyNT0IDJwyBVkC1ER4mNu0gCKYz
Q/aSS5TeMgBbddQaHIajOUb/YlfNyqDsUFBRF+tqsEGhYR3cuboqW+Fk0wuzhi98
JKOppd8Z392mcyOhgRsoeuzqkI3gr0yt1+DWXlsGBoLukZM9zBNutfUWZygKxtOF
QSJ5he3ew05BQCaPRCUm93WTGHNQ7sm85FVKmZizUHuvhLiduSancUd4SJG3zKYC
gI/LazBP6WRiDuv4Ycv9dD3hqGgHSVGClkIDDLOsqIL4okihJ/ilOzKOEziuIb56
p5Caxg+9/WyJVBt3NKNBHeVuZ/l0htJSuSkfOKtFXtNzpXyk9/nEnAbIaUbU3pmr
cZf9uQAs63UaOozASNskBev9hr9CYyLbWHsAcmqWvdZMvKcmGDRChAWLfUrnsEtD
H+dJxld/KmUZfxXxStCJ+8oxHRe02uHmB5uH7Mvh9W0XEWNzqUhy+JeRPx7zR0R5
Zd9tredQVUhKMejgB3LmmUhWo0Xx8jS1Z8u7EwTsWVMQaMSssVBgGgrXYoK0Trg6
U7WbWDF1GLBWrLkUxaXpiiweXSVyVurjYXfCvbgVqwVgnZMsgjABSaixTt+R1C5F
6EsTR8pCcqRdAPyqzdBJFJtiIIxIylI5BwW/IHvzWw4Y6JHR5J33MvKDnXMyM5wS
mLMYhM13werV9nuPpQRe4PY5rID+XjmxkgVAjaUtAbKAbOFIWDHdGmIvnli0E3IF
QyLaljeRM29EELur4hMQtFPwB83UY4qITiV/00S2/7RtcN4cMDnc+LZohvGCBBuO
UI5S8vDMoQ0gj7bJRjqcwbVpc9dK23pt67fx6hIfjrLDT8viNZxqOKXj9IgFWtEH
n94oOqbOcS3fupCBbU/lTd86FX35WzqKL+DZ8m+OGjRGF1yWiXX4Xy1IyodJszIH
Kt8wAoUTLkoTjwyg4rp1vOGMk8T6hAlFnP1oVMvIP6iMf7aGEGb6yt6UjdR9Hl4n
50nywCmGqnyiqkKqs1tc5hzznUXXgNf+SbdOrTEA52kOqMRw6m9cHHr1Sq4OSTAp
e29Pz4v+rSalAimwskyNOLFewHOaaq0J6/Yrqc5mdAJ1bCB/m9SuX/fF4AvGO8L/
QsOIClhdaR06ubsacaJ9pMp7Lsjee5mK+7jubZM1FjByzwbuEe2L+yd2rsylWgUw
oTc3uylZFQi30vFEs8UevetQbyovb1aMDO9/XE+jNGk2HfIar5I9o6IpAybH4yjA
e3R8fRhNrrAq/OzAN0WCthWFaHm6UfXTsyGYjXGz9vH6UDVZ7pMWJVc2EEn4rnwk
/JXSCz9qvKvRQ/bCDq3rTK+GdLPCRWjDrfXCF/U9FSRi+rISuHFfZSxJpf1fvles
76MaGNRk4dd/QXk/QfTo1iQFChps/C/omUXkCMGup5c/TMvWE5vzwudAntBbzCP6
oiv9mbndkT5ak9nKZhK7nW5mIpJzEfl9hoPL7sUBYdmLAgmSN4QrERPJSc/RnKgE
eU/zuiu9BktgOaEMvPSJ0oNMosg6ZROqqH56THrJYAXJ04kO5rBmlYEB2O18vfOk
whEH4NBXAv4xsUfXetTezCmTCLK7tQtpq84rl0AG3Yo6atwv5NcNNWsoijSaVp7s
W1QnjYygfjpw96oASjFV8juJIrN1LtVl8m+gtb42M16MeKVp64b8yDSSlZKHWdwl
+owebMk9GsQLltw5LigZtn+OBQAXn/X5MQpyY0Eq4F2mbnhFLC8f9sIObsnX5w+U
5OQYs/W3iy67I8ZmPsJDAITZ8sIFy83gwDsPETy0utCGWdnGZSfwxPYzoqpeb5Us
Qr5mxql8qA32i7alvAbjwG8KYP37VUAiZpW51/n99QIMLO6/e2E2zw7t7m5tkin+
NfUJUWN2uotKEBCZcBp9k3WMVI68H1iI+oIPo6k1B79A6oOggzZpdTGv7dIXXdVE
lnpQOQEVr0MCxy7KPk1tthJq8maZM5nq1vUSfVSb2MNAsAjgfz3blfUBHWnNSP7o
XQXBtnN/QOYIdl1kN4vkmFMBDkkZVGDlwWMRXsXB6FF/OQylIqmS6mCz7ulmVfc3
WrqsHRTgjaKpklslOAgkBfyqII587BDBLSkRpAHBJ9DGJDs6dNZmalFN9pL3ckCY
m1aVWS/wtu3qW5DslDjgF9aS9/4djKpOXCr9pOTE3SGTrR8Wn8GcHA5HWKgQjxrj
h2fOA1UAplYW9ii3HJ9oiJZOLwvXVrfgppQmwiARjCcPwvzVEDwHh25AVyZKYcql
dUkpnouPmSV/eLckMg7YhpkeErSYKdu2SNvP/V9Z+msX+K9NB109Sh2lEyLGMqhO
80VKY9+bu2+98mb65t1VhBlU7HLd628nBLxVpv+ADWMWvrLcDaiIQth9Z6g41JV0
DlaMTbx6o7smp4AncE6Ws6SH0qzloWAjMyqpHO/Ywq6TREJu51+YzaE2zrnFu+0d
Qg4Zb7X1qodbvZHHPcQMivgPxDZaC6zsAuPAemTHP5+oq1N4FC5RTG17KJ/30Lek
qt8G6uPksEvWAvYZ0vJ3H8vjxtM/HGZIRSe5AYaI8lod7Mymp6AzLwNJ3+D2ulWv
bDDRPWlVase458P4HfMyXmfBZHLGt/ce3zfnrL31+QIKSVz21rKx9FxHhv0ghL1n
+5kKRv9kRG+iHP2Cv/VAGtORwEOCXB7kQl5t5yas0lpbaf1vdWj/WcGkzVyRF28r
qOeKqDDSUHnabvQGkBw5Kldes86iaol4So8zS7Xse1KJbvBV+xqtptF/1V+6eNIk
ZsiphB8AvA5kDLgkXQilQ5cBNZgp8XfPH7QSZMf647jOILCVLksI7UGAHB9r9Zds
Mk669bJ6o4MNwkgnziYxO6dbpwoZ2vGGbYIP7e4aQKV9BNPn/gXvNeVjysSROcUt
wVfIAmpxF+jM5HahW99B77DWIfzttqUUWoddemwVbJNYTbszJH88jU6+jwLQtR6T
v3FGl44eiASTUZV36xAfJmi2Uqkzy5x/s1pNoEIDETFBHC0PwNEkmbZB/olWJ7Zz
PYwxp+fk0MKrKQCcJ6u3syyDsYm4wzyBLAprWJT8cmLu/cHrHkHlUzG685chmK60
Tg2kGEAmclEPwbrRbF4EsgM3351bI2pytTFq2dfnKXK2YvbkNu2C7uRf846GjpUZ
J0fQbs+pKpWHDwKLPLyL5Lbfsj/FSMODaYk+kRv0ODNV+HzuWjPo3frwg44A1ASf
/y4DXiZ1DvhUABNAx6jG9uU2b9HiZqlZOvFRcIEvk1klrahpBPOQAUI5QBXROhlv
rWvvQRPtzCAeTGRrikza50/x750YjWn47k1J7Xs43z0JWu6Dt24dR6Ue0zHw5kTe
u/jRGjScL5d3a3iv1di16m7HVwCYSC7OryY6j8Omrx0eItQOu52AUHNy1OBCjQCh
LAHyHwbzjSf8xFXAuw7D9YmV6q0hGbSAGbhcOUNqbRq1l8+ngIViYP9yolsLBtcr
i9gF8OxTiR+2rjjC3MQRxWCBe3YdI/ik+ufgtuzIxn3A3pfBxhX2H4TmAhYfPxeW
g1eC18gSfWDO1s4fX8AaREi5mLoGlFS+ePUUAgK7ZW5kbxuscsy2YZZXXozUlA0T
pFle2eAzMoV6cUjZWpu4myZdkzlrAePRizcmmWlE5o13W3tEp2dC238bVzBgnoBT
JppJoOcvGoXiWp8Lt2N6eoQCUE/13Gi19LurICDoOAB9y+SfwBxk42bcVqrOKmWZ
Y2ClJ6x+MPMIH7p/roGEA25SBQ7uNUFH7MTw6Vqdb0XdHBBdD4CjMOZ4e6uMyqZx
b4YmurzZlvWKPolWPyGRW5yMiQrxUVJ8nkA5Mq87O85I57YLpNe6cVKXfdRLECmC
S0Unh0mk3HdjSch0JnqePAjIZhiyyw9Sdkihzb4XAG3jLZTcV2VS2kNz4euwR7Sp
t78VivqnjXYAfG+O2kocLqQiAZtG+n854duDA86gow7OUD0OQwCJ01AONyU4l8b5
7kZ0OAtODCNm7Xlv8ZwsUmqclO/PsqSzziI1+SrCJnsX36YZCMzDd19ksGIFSPrk
5i+jv+/lWMbPWOCTxf1MmoGAn0Hy70LbvPQdBpIhx64bw86u7koORZ5+8ZiQCITu
CiA1kClLcj5tnPxAl131HWuxgjpQ679ypyLsdEW/dB+m2DIXBG68UbDQJVAQTc68
G25cL13GNo5zRX3ph5AHn9+ck9kYZNxk/jOsaB1LX7Pxss3UutNGK0IMc6BA63qd
3fQwjW2xB7NpkeNuW8U9ygGdb3CpIop7zFfrUjLTZX1WZLr0u6RihOrbL0bE3O4Z
+l36IirCh7bnfbVnoR2WZhObI5Is0v7d98kK39qQMgpKmNDYvb0b2icOLfy/JYjj
ze5g7qh3IyV7K1CrNruotlmsoC3GP+qHwQinJx4qsi88WoZszUWHq61sh4uHwLM/
2gYsV07JRXW8KUvIlHF7qeQPQ51E1mA+A2IlVvGRbTycwI0o6PxfEBZA8PNG6QH5
3zMcwFypNKxqb6/U8xMr6VRqOd0MNRDrJlVuNz7RbQgF/ff7hNRz7lWvJguIHfMG
JZpeVwEKMEsVXR4Rp9Y/gs29IILxck/BAKJHVNhBOKaFnlLwO9NpcqOc5cj0J9dY
/sITpkC7YK5vc5GWjMQ75K3PgaUbzQhZ9svqGBBVTWxAT/kEQ0fqdw+4z8tpBy5G
G0hKLWKxl5SVxuPMuW91QK/QEunK/4KPCCae9qdy3kzrkIYWfi0ar/voD99EMZyW
xmoqtt85XZmIqz1vJ8RtOopcmD0oJwQtWbjksrJFloBs2Kbol6tQpdVzHSMw89XT
ITO7+/xpWgarMnrPbUA50SK25L0qxQjhNu8p1mXY9/gwrf3AVDjUR11dede1VKl9
DUJbjLY3uglAQBr16kTR0HCKnwaTOkFr/3MwE3y9zJWw9cRREqussOAF7ukofPFG
d08lmY/uRsWJjqSL1F+TCRfPRcO028hC+V0mASAZ7+oL4Ecj7a0jNIuErpqDveNr
a7qLxmTFyO+lWH9EW3Hw3x3sI5Jjk47e49QJnZNfUAzkPKD78u7s7/yNJCqAlsGs
/ww1XttLCcSFDuAiCe+ei1zgWKmoRkTDab4QXFB2NmNjt3MkINoNa4uZiJXcyGl3
mnCdDtr7fZe1icndtRyc+TPtAXf+uonCyQQg8VbpVC9Cf7mvoPxKxE3muVZ05S1L
FNkD4pviHIEHcwo74EsiIPblKtI74jMkKxVy/BYeNQfTyqOe8H3OwZBDI8wiviYk
qpUjz+XEtmXkv+xIr6CN7xQwfxl/3j/5bMPZoywE6CmlMhCsNwSwPnkHZcb6WvbL
5QssjQTatqF/nhFILtp/lRxWc3ijp7TspY9FhLVrFCxghWMPYBE/VipMBSf8YTxx
AnIIXV+pbkaxeIZJMiKXui7Y/dQNOdz+LX1E3CsojzV3qFrtu6S1MA+Dbjv7d3TI
Ej8+wlUAkTogwi+2z68aCZhQCJwxLJNwXbrSPyzYfYap92TN9E0fcojx2Mbfk+0i
+Ld/J3Lv6F1Kp+OaTmGIo1+m36LhohUqiRdglyPK/1nm+9au+J6VOP2hTZDapRAc
rUSU+fJr6us+iVsyHgTDQOBNT8i0vypuK7wk/C1m/vxo4wBVZwLau0wpA2rJvnKb
gkfi+02LdEguesKMK7eke6to1FQkEqQmGr2bGqfT/YlEYzxCuwvzCpqALtPnXGMZ
Xsqn3HMk2lmtOxWhMgoeFlCpde38LJxMeENXqPyQVjPv3a4j7lNYpiXONH7VhpX0
ZT8nXlT6NST2j8jrMU7e2xCR4W+97p1GAuyo+/JDWdNrPg/xyoTQFmrxAzwb6tVh
SsmKMRKt2s+IMemnGJAgYWSRrUGWH7XSp0DxPCNC1UpljoLwKlDlSXq/UftvDoeX
51OvJtzhUAd3JEpPRdItShtqdObWqlHP5zm1tqHAVMxgUdR34zrxBgbWa4Q8uLjB
tmDMgzScrqRvbjYzuqzCaPEXLP1pqERp2mTntKNugupUR7UtoxB81zB05MTWjpuw
M4u17g+PuijPSD6vw2ik2Q5CKVARA1wrC2E6UI/4hIDpvVUlD3p9ZnqNzCbn4qXx
guOPam6uE1faIyG/mHYJPANaHRxVafPv0Ut5rsJQeNflzUt/89jnnJxUNd+9nPj/
r+gqh0ZEqrlM9V0sxL0QeN2E+SzDuKwuLUoAonvokO/w1wdYFb86uKp4ocWhYwrF
el7rcRDTgTfGfgxTFO9yYWYUKhpN3wW3DeWdlwlfcQfKw3aAGTA+IYniLJe8sc9h
w+gMHymu2eKzXYVX7ZSvG+E77s+ZCHqemBYfKFD6UKx8FHDJPxIi55pB8yaE307b
xLhS+KA9/t6YFVMqrEYqooHBHDZ49CIeZZxH/816lmbZ+dGxiv/Qkjifl3/c3gDR
vdtlFqRKgy7jgUFWNrUpZdhAm/cHLrXdbMorrdbYKupqQpIwWRSN29oWyfYx9ZdL
+EgW7SzBPBhBBmd0W0Duyg1Ot8QBFo0esqodcCCqeE7mTUxh791mIgN/DawuO9A2
NtrsxITeFN2bdaoUFuJF8NHTAUh1axDertJGRuTavNcidcf1bUmJdIIoPFxNnFxp
fqqAZVlk9BNelhLr4tI8fD0FizM1QkwJsikSp73Vo15Ro0Y5sjl7UPG8tp9i5S0P
BkrNwAnEQij1uYgJCpoNo2scWoo8LIWIoVEoKXI1/6gsDZ3nrf+SngaRz/RwjNlm
JoiKW8AZWmtQ2jpmyNqumpZZyzrbUMMhY1viLvZDLNll0yTzJ4ECiMOJYTGVcrwM
Wtq5SuZFAaMSzA08NNfGb/HPpHkC9Pou0tyAtLMQKM3NnX3jc4SlYnBdAX9JDxMS
CUBaVPo2/feZGcgNkMGE95BPFo0/i6dlMqoaO68aNCoGPcaOwzANe64MEwql6Djj
7uLlMWIGttVpWV3BNwia2qdOMRZZeB9zymss7xUeDJ3pssBrsxFuB1fR2d41OJ9z
/OzKIEDN1/tJIuz2GVMifs9L7/XLTBYt7jStjVqLxXddQTI7ZFBIn4iDfMCnVMUY
WH4QmcU8Kl1KSQRV14ASC2Rd+wNFJEfZGlg6zkcUzJH3v0b16NWewWz3sT/7A4xr
5eiVEhsiGFQmlmxAmnY+nTJToE3KS2WyT0fLqhepCyRO+zjeHwYiNxCQfpsWBbk4
FXRwuG0DLQmgXz1TFu8lUmmQb0veG60fTWTsTm2XE2u+bqtR3YlIIGReoFcO8/wz
GqCwGN/djtCsM/kNzbuDiDE6gcA5vod2qT/cQXpLBGa/LEbMgRHYCBPvaSlWWrpG
UuDb7xqO/e94Lse+D3X8K1hMWDg5RDYaQkFxiQY4BzbDpy+BLWw0ZKt3SCFF+ryk
nx2ssANmBjZPgH++TkYmvzunfnjWN66CV3ts3uR973V94Gyi7ObvNfiBLdzTzQ/l
9BSpivb/iw+P1BE/++LfLJpdW1ZADOGI9mnDEcsoaoL7XC/oSkcDn9hlgrAddeBl
jt7DVje9XqWyaXWg3cFkDYuLYaMjdXtyxtfo5hzhhSqbrBw7VPfKtjQAaNfHXQRC
2fKkJAwM+SUxt2yrYfbc95akNA5K3LhUWvDCBWD3jnYi2MwOnvpz6AJBf4Np2bSK
Sbc2NMfAGLX5nkSY73y/I3E2Hm4aCb2aBZRsf5vcg0u5zBrTWSlC6Ug6SSX9p+sG
6Tfa5LwBKaN+WrF8lkKH7PNSgOWRyozDBXMqT4oRAtgnXO7GrZVkOJBC2k+IDyOH
ao+wEPFKloKAC7KWWcfhky0zcclcBdhCv6jp15z8AV+X4PFtxb+gPzvsOm0bm/ZT
MLrMJYO/E914vjCTDhhJI1moG/6bvNmpR9Gmz8QTqAiWhf/tfmS15BsD0D6S+/Lz
O8pjrByOX+5NRYyBlfwG47nTNdOgh+elwjCpXA6ZghkTjS4S9+PF+Zr2UYg/5Sv3
H9y48XYCxz6zwvFNmoS1dqAJb2d/BkZ0XjwmgrdkBgBA2B0lzBP6pcWs40ky2tA1
Wgxmxud1B9YZOpmIi0ZuClEF3rLRdcB0Rl6Rey5IPeAVEuxo/pL0Swpps2XoeHv6
UImXEX2E8zeNNPCUxYls5nhB3xno9Ap1Daczcz4fY0fxJ/wFIodO1aJaLKR2U1rJ
U5CJFdt0O4g4yVu8kayrPNMRlGwCBzhfPGtcaosWW5nVK+1GpInprPaHFXI9ghfc
+gaq8WnAkQa4UPLvrYzymfAnY0df1af5KZ3zofVnSg4oswccg4j+5plI7454e1lR
6yXAdq4rb7FmdOANHw7tDz9GUepr/PNQvsU1GYTJ3LgJYfd4n0poijgJQS80nMpb
JEEP91jlysuDphEc7if+dWh4TUxbdmFVXhKeSHheZrSvW/HvK3XZmLkyX/3QbaSR
LrYu7pV050O5IFgRuVtN++ukH/H1Z4MMF/oO0hbbSXaI0V7efVEKaUwIYcp1XNRi
FPh6LbqDMsYFJwoa5VHRcaqbI+bhOeJbP5OJIBuGES75zD4CUk7N0YOx7ppR1dsH
9Ly9NyAnePbXGXKmhfL/1fGJQdSoTBrdNn52+nntVDIwydfnH6PmP+3YQ8LPHstc
VZFkYWlrrXsyXZU13ZGwMGYygq7RWodl75RDwGKiJ2Z5wK09Bl2eSLxkoWxl1Pw/
SPGxwTDsz30lyTDL0Ms9F1K4sMb0yu0qLRWFEHJvxLcr6ghKWjpUTBNoJL28SEsR
EK7dXpwX0h3GW37qNjzpOdXL5XHp7JRbQKIgyTMUaZl10TVZaIR5kFSzTIynBK4H
+YrQs6xp17Inwbi/qB3W23jDbpzT8KLD9g3tmMr/q2KNZ2pf4+Zs5Ugdk0MuuS44
pxEB2ZBxBCjvIc92yyYVT2ahDQQwwbaqO4GWuBPzYDhG2M6tspKbAx62q4e1jfhX
n37NRl8q3P78ajW2MI0bjr/ZH2QVpjxPrlq3VgiOiGsC6QKBbLUtyW+YoWLjDXCD
KVwqSV3k09O/O5JUo3b81wC1yqyKry5Daw7wNzUfv11LyfZM2SSLQHAHU9wBmOP/
59SpqtlhNO2QyRClMAXd7iwb3dtSLDlPaxVh1z+DTe3prtIWp8lM6BB4oPrlfvXq
3ZKHkczc7M+TcyOFXWewj2EUDYRMaMBFk2Pxj/b55y22DLL+dnIsEAEUBllMgv40
OhiBz/NlRWbaCSo/4YzIu/KKWRiGHYR9tZOc2PmQ7jvpFnncqvOv3ag5GNwxh9Wc
zdZsE0aQ5FvJ8sugBbpHW+AY4kbdguiA8iGhFA5yAQmCIAfwQHvdyGrVB0jjqX8h
YO+eZqg6htMHwnB1HMu1TdwruMiqiHUAj5Z9qtO0lkY2UoXXkpgik6yaf6MUDK7u
4PEd5mAv94AKDWutVCDe7JlPnYkR7LQMNkw5EKDOdnnUEWvjDvW71pWV0mvVaUt5
e8TLpFYe79Sre7ygSq+P9ntHhQ4QCk0Dgk6LzNP3FXt7obeUOLAOmE6sHbj7Vnm1
rMLXrRtCC0GG8TeFIMSCcVsnvNKeaKOfcl+Qr6z+yyW1WOMn5mNWqb6/LwPd5hgv
sOsB13etgrVCJ1Z7nv6Xm6yQRvvxZkI26z6UoAFJzCNeKLWWL/UI/AzQljnCtJ9/
84ootEQv7yQnOMSshLngB1U32Kh7MGuRmXeTZiyOi1+qIA4X1vAJlc/84DoKIwZe
UNsT0Chj6Rn0aJ7s04Fq108ZA63o9BexNyTrrkw0EPtGg8rWYQRJlyZjLKAJD6Js
zXRqsCnijGnbFPZqyMfKIjv+ZCIlyHscNlFU7/bhTImLAt8ghejMW+UnSvvRD3rU
B21H1s8JBhRMEVBFgelQ9Qg3CqqJxPDsfCpHCS9D/77aVFcaLd7tiIeO5gRxhHpv
sr7fOWteUPqqgVIXGkiCxR2yLFiIlHOOaxG4HE9YpOE/1fCIqT+UzOvIO3O8S9MR
pY6p7wWJOAaOvw9jJGcov2pwMhZotJtvDwfODSVtRpiG0eSWO4Wni4U047WlK8S1
ngdv0eIjH9bd0KpirJfBSS3LZmlR6yLEmnGwRQudxtcFavhoHSjpZ0bIqLMqm0Qz
kHhYGT3RhoJKJtFjYfjPrkezH+x+ieWI35mlPGKR3LrxwcBTR9tpVfqXjmhfpH2J
NMpRb/65ixqqHMcEacxuC17glmZiy8G7KilUO9eVpmqg4wYeTBenjYWXZU+xj337
nH+9Rc7daAAEomgftR4nVputsfM0qB0pHG7pPHie2c6eGDPzT49BedYxk6gvjHB3
48Wr+5kDrDLqkFZ/7jDIHz0JwnPXMgdmsY/fxmtKb3vn5nXyVH6hp0Q+j3IooP7T
0fC8YnFdhAtHtzBU9rMhjdMblHWp/A6keqOU75gMtNuknIlMVHf3iQl+Y/WIvChq
ptJP48DunvHGzRcD6cSiOGrqFPW/H4nF/JBt4qNbCPsu7uksgjYnGcQ8Y8lT70O5
eXTEXk+7zNNFR2YMrtq0yYXDjrg7BQzl0BlDXJCdfALfkF1II5JTtgckNXLh5dcl
l9ggrzMp95jeP50hsBXPZnl8IOKE4KQ4VAsSKkSh7Evj6sin1yOpoRv3ksU31TT6
0XxIHQhqWnJDMXsjZNtLm3uTfIyaiJu1SH4T9WxFSek671/vqQjFbTNIjvAJMy8V
Kykl2wgaOOEV1weV+OGESZ5R0UNjKjRw+CTXci1poCToNurfk8EMcM2/KaCRFUhh
3QVINso5oTK4GppP9a1T9jgWj1IvBxASLTNabxNBnYWttoS1HmCWwMe/JitXTXoJ
`pragma protect end_protected

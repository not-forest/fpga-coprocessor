`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
osqwYOUToZCTv5gYuPeHXxAB29paI0kkQiWNDMqlNcs2LvAUHHDzPtAQBb/dReFL
q1NWBYsGBFjsqc80L8xhpnzKZexhdeV/XOwFM6cavLCYFGuXUoMUmjNX6tUimJkj
BbuFnrncCqMqgc8566XLyecqc0vMrlh1UO+yBDUaLzw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5520)
2a68hY2wFYEU35xc04v0JcUC1j1dEuGXc+nBaaNhotOdSDHXECQFuCC3XJEskdsh
rXzBCowXfGZWDYCuic3e3OiyQGYlsxtZi9sHmHOpULGJaC0F1haM+p9kKlaiQhUo
xBfk7DCv/J/20sK1mJQ22d42JYKvsOc269q7Bu0htgTnMljj/Ovg65rqdKp7oJRe
kkddckHZqqV6UXzWuOi27gsUwgjrshHYj5vPAJ2KXewno4wk+ksNq+5klWXZAzfu
47JghO+SVXkjBTymaBF8fasiFZel82vs48srbzBprkXtwA76/UcPvleT4FzXYMCs
OssVpgfuEmRuRyt6CsCyl2FCQcjB1WZgBMh8ebxDICXD0/CobFxKIbYqwn43jS2j
iP9gaoHnVFQQmhFnPjRV/k0ebI/wvOv5ESni0wDBpAzImuDgBC+wwPl6Lly9T+4Z
2CbjJKvTBDRQRvo8ZMXM4vPniTC7JiGFeBNtRh8tlgUGMBrLMo/zapctQTdpdUP1
HYHU1JqpuIGd5lkzPVD/I9Oo3AnDLnbxwBHsi8lG9iixmST9pgBbwUhSOdEo3E+d
QFphnBfam+DtU4HCdha08agEKHxlRC/0DUmiIQ7xX8kFmUS/HR5CCysfoFt10Efy
7sHxEYvh5JfWaQ/+EgFIQOMRG3lYio/neLbEF8ASLNbJtAPPnXuLuL71uVo0xoz9
nnQEoSJ13y+UQh9ll25yhc9zGQQJSErN0H4P+A3UODxcx2wxuxoONyH5vux4mJ5K
w94eJu5PttE3yqzbdvHR9eCg1tgwqHSVR7Q/QvukFFm5V9Bq7aYVmPkylgMGlixv
swCSDcaHeEsrmrY2Q2eyed4MrQpecR8CgCvafdfqUw0FsMzMhSFwiAxl0gWDGiO1
GC6TEMj0i0XUfhRMhdOBnqOIraL6YtOp3ehGK8mk3uU/eO8+mb2NYeKjALb5Xcgg
T413ukQYhsY5kM5SzJuBDFWQHPrP5diqc/hp4NcWOesCPeyW/SNzAzTog7VuPP4l
uLquRtVv5AviVht3IhwbfT9XQajGoD86zv22lZPvSBXJBaBX6o4r79OH1YK9abCf
mvcyqna7MZtfOFaYqAsxfK27/cBdM/KmQYhoD3rJMk0uC5kw4L0nBt4Y90v0K0/1
q0lBEqNsy3GoqTXs8pXxz9QfgH6vBkIruRXMmuW0bTUD7HiU7eO7t7R1Lytjojpp
fTQE7iFSWZDNALG96hPTc+C5aplYlA0S4aF6A2PPkxYLjnG5dR59H0qbbXOiLQO/
C0rIZsGhJiZDZXnzPQfWSSHh8zSmGgP9K1dKNQeLCewsA9CD4hsbElzIfU26suVW
LpnKmv0auid29OjXV9BU9wqS+svi6tCcI865khZ5ve7VNJx30vLtqD5gxRYrxG8N
VmPUeXdQ5y0clkguX7d8zJdqeP9EMzh22X+LGhp8ivs1vlCdEVFnMZvUQV/oTAeH
L6HsxI62Q6uhK6vfscZo5cAjrxv+tnkxyiYsw5azHkE9HHfr0gd7DEJ/IWNIZ513
TTKUhR8uCX5hhlrlwFVvIXCPx8gBClQQ6QWM9+nH3OVlHiz4ism4Qe40ZU9AjXh4
5+h87eZIAgvgQjgFGxwaJFxAAN0gaYiy83PK1rofqpnO5AIAKckyuexr37eaVXma
0bcn55yXnKyt9bB5Rm1NIGS6YGK8YeGJdfGXiOOBsgA6W+XNLBf1lteOX7pLdmGX
NQR1FRySJ/wtVHSE2Vdql55qdLgKFJYZLG2dcXNNEHX6LQhqKPdvyVLb2cCJx1d8
7t41jL7chEXUymkCG8uIhUeiWCXspA5Mke1kFWzw29Z0wTgyxIQ2y1wVxpPT05fK
yUTVmVHlD2VQ4/JK6qQS8AtVqfmXGb7PrblS5N/1zBNFEm7/y6kr06mpDEyGGHtQ
mnCg/e/QUITL8heJ6HGruYe7yOn9Tc1Cc0hxl5o4XR07zaNBN9n5tEScE7vnfJN9
dWeFo+uOSfXr1APeWBWKaeBstKSGdapeC76Y7ALLObiH8B0TahgRdT/dgLik2BWN
TKDwWf8CvPdW+gDZLn9K2uczeLWs5unL/tcCZt3hZu43cFUPq02yaHEHiRFPGYj4
MBCBfbtTdzWgJA/Nlhm/BbwmWsqGTdQeuFj4eWm/3yQ0d8mZN/OCw98U0c1s+Vo1
m/rr4E7nd3E4bXbvtgL9sUwCG8C0WyxmiektDLZpB9S7h0iDy3PUkqpYgRMnXeNt
guQHzQzp46Jnt6ArMYm+9Z8Lr3YTalSUmkHccB+ZhtuBffQmLGxY0rd1oBalEvoq
0tmMVc2+0R90fdmBnIku02EyuxzkQxrYKiN1Y7Akvzb2hobsqq9W/iE2Lslrq6bM
2Xi1Ii37sqbDHQI9ogBJEOuC4AoItIeuOmeOmKDRrvOO23fmVSi4lz/52XZGy9ZS
2jgzBQ76ThtxROMmCwuzuPCltCq64UJZWAKyBH3bKzpdMHXLOpIf7fu99CEjBbri
9376RbtNH155lGWcAnhj/xlfpH86KAdjuVruoXc2qzoXPl6yJbMGOOtOWmVAxSqz
+G2uwi165WTpRLXX4mW+VFmM/Xb6GELv1YOKVjASSKtm3NJWtjFND/0YTjG5d9aD
dZJN3tuSbXjpLpUoT90xESB2jQEnM9CSC6dt6xoc4hT2bwZott/7aaNMEX4Sn6Zh
QHXQgWHTVw7v+ntS9d4D3GXfSeEOdAbp6aYlQ/iZOtS+rlRwtERv+tcKxD5IgyGs
0jIL5loA6qNliDBAI9QUXVSZvxXgLXeIYdrG9Xawwqf5KcW5BTh3nGb8P5G1GZ3k
4B692Ae3tfjaBJnMBSOjALfA7rmepuJpiwpuFT/pFdHk0DeTIyWmAGi9VOBGhAov
pnKEItPyrYRVmYmC8EHqhwGlTcEsHNdiHi9KpUjp3E9jc5yNGIgf5hSm89v+F/7q
1FbIu1uxkeh/D2lok1vlkj7J7plYnIMtvkrTI0Jm3EA/a9nX+1Aizog/5+XUsv6g
Jg5+lRy8MX2mNbmFb4oZM5ncbU0+BXsNMFmvWFYZ+l5ZlkGaAQA+vRfMNndC1kAq
tVrdkQSpUFHMf8ELcHaXNeW2Ef5+mAM0F38HkleTk5/H86iqTawcM5Gz+4S1Zwxs
J3o9O6FVd4hXOJk0Fw/S6PH8srjwmtbFAjtYqS8WFAyf7JAfT77dR6w3kkP0psNJ
azlWJgibuaogoPxPxI+YbSLyoyho2CR3JXo/uASpVMBbwJrNGAXZQwEicL4mFeHn
DeeJh8DpKiX83r//wR0BdZ74vInz+6MVo81gCLc4+ZgU++ir6ryLxaa0EB6o583F
g+tP8okbAFpo6DKc2TI+M+ahTMtOwsesbKbPceOV6GdzK1ZHSZOgwo5xbOEETbQi
Kw67Km1NZpNu2eNBYq8dkPj5ss1/3G40mPHzxh08WoollwsY5y9altmgLL67k67D
Pkj5e1ADck9pXMZdix2o5fWisVvrw2gKdelaqz4PshYjWnrYlHCTd1w+k9VXwySF
fBZsjyVb6v5z7+aiA5oT7UKB98Wq3qVOPUNWYxtJFXcVjI0IwskfoqPHIpR4RIv9
vNxVK6LPSl/KHzayynJn+njiEoRBlcbdEhVhXtxIb4XC89B94vFEqIz79WSLJ1Sy
tZJ4gBrFt6lsrnDzoVwcrHR3jSFiuOl/wr16fopDZcoUdIblfguzPhBEHQkh3Apx
rapGOeoS02qj5ZX8sIYL5dfDwRxdQp6uT3SIT1o3c4WqGFgvvzPA0dF6yc/18P1p
LpF/87iecaC6bttO/7xtOVcM4wG7FluFh5xOVJ22tqFyztG/rWF2Deomw97UMxgU
oYcQF6Pq3KvVRYOC4z8F63NqoPBfmm5GlaWHFrJbKNu+QarcJd0/NgEJCbxiWJUK
CfFl8aRdEySd+tpG6JDGlwsbhiW+IbmNDEDRQrmqgcCKJVmLwQucezDc4sGl7mvE
iAxP8wtCPACrao4iZe3oBG9Y+ICsfITKNeOqQPXqK914rQqW1Bz8QzD6g/GP1w3/
du3eCvo4a22prMzB2K5/6ZdkMQEK6tuZE+a2Jit25wtDASHAK/2fSzysLXKH6U/5
H3cbBAkSpULtoMuo6cE8UMEp3uSSXZdobSqyKGyI9iFGBbngfoDKGtP5d9vCHwgj
zGSrfVmvq8LtIpxToZQv3/MOxSUGzTBSmj0hKb8sdLGclFtqfCkBX+x4lUeQEuSZ
98r7+wMTX+HyXgXH3SJJxiWPPNtl4s75Tm9YR6A/sWseEK7me+sHefnLuCi+13gM
XlsJClm9sC/PyGENhg0Ek7NAND83kesqsSr14aSLKbIO9ENxnhpxfF7KRH9NZFPb
uOfaLm9sHNoTZsQIAodzYscnr/Xn5uHMCbR5wFnfStjaXDJ5qWcOPvAy2eWX2kSo
aTFAIqmb5SHzqPjqYaJ9AsVBGEaOzS9vHh0Y1JLqKu36Cq/e/fVXjtxZ6goSr+xN
rEkU6yT5lMxjv7oBcs7hCprMXowI4s0l+iEshgdtls42mNChepNQbKI5WDDqGgSZ
h+gzdzJxG7yyKlut7mtj2omR42cEeMILXxNoIE1fy/kH4og7mRdjWWrEHQ0RIfRP
wYWebpxghs638fUPNC/1QwRO5dYI4BvarRFcqxX0MnMlfRmgynh6Fc4/+bE6DrtP
b3LMCsto6p5t+bk9GaQo5lYKHyo+XoRfrxHo7Nc85FQW87qT7/A2781ayiNgxFK5
h6wKKNgJLIHKHmXX9ioc62+fN57UTD1glDa0tKm10OtGB93WjEz7QF2DyuPfZMPj
FcWRslxovfgodoCwtPrkKS9uNY4c5im4nvP/8697kUR9MNL6kKEhFQcbBYZrPEp+
2chfMVynH8Hc4so3HOhw3SzwajvTkLp3KGM6Mc3vNBGVdJ0MDpKN3L+4piLQ4DAN
NaI1bJCaVeExBvMTmMIIUgZHxF0vtWOzxpOOIvqdwTcYgeX+ry87sxAnYvvtSvln
9rzf/p+pwKCVODQkL2VNgR95xeA4f1PyZPIkKE0sLM4XSGj8kYp0C6807oGYcX87
g+C5VfTrV8IchFZw459BuFOhhxIlcVUxfgkbr9/Ld3ZFkHL0wKxxvBj4gEk+k8yn
lhP3g0jGMJy2L3n1wTyYD3VAXupWVG4dCf76ueMemQRGJTCfY8HS/JTjm4EsYqGN
V4UEdfqcxl8L/8TEUOzWQPoHTzHVCZQGrfwveG8NJP+0/JIm6H7JlHzZqQ5Yj2LD
DR3LZu6X/qo9+vFYdVWB79V8Ruy4kLTcafq64kzHEuR+8cuHbxXgOeWT+nz/GnPE
/6U2b4jJR94QadCaHV6HfhVGv+P7KdtdiZj6pLUbCUSSuSY0RafQVksJXrJH8UzR
8ljMfarN8qtJA53QuV2Lry3k5VCrurduIx4o1U9Cd0R/PEPRQxuka/9nr8odSVrA
uI0k4QGGtuelxrfRSwa/HDqRFTSvQ99AG8I2ObegT9vzlXXmkoqr9oQoUHlQ5/aw
2IK1siO2caOGO08S05m+VYPlrw8mFFNQS7PPtK0VybGd/bTmIJqZUYOXYdX0PTfv
AhpepsgNPa9Ct5ijU9Us2X8H/ZFYxdRVR4pOLhbi3mcM27RjjQvNpYUhFvLpBuEA
G/lJ/2Z4d+ujyCxaxib7pq817GBbvRhT6QgzNKhHrhptrBFhasUdQQC1gQwYzniY
3+QKt8lH8VU5bnAcExZxs6pID7+KJChm8bo2VqYQ1bEzdnfVXJgkLLjvuYxDbG98
CE07TPd8fdyRAHGIUgQ10Vs0tCGHkS2ncS4n0HlBgEELiMOf8nvXxYrkpBSMHvBB
1d6XYWxKijNkVAMo9viUECFe7QFBFUH2pFKR6VJOUBJchcCSAo6dHFRLpFtSi+N2
h1HDGnG+E54xulfynKSNVydx9kE97g6+FTDrk5mWipuE/vojkF0k7xPgfiPVIoHp
qdWdjxQo17WF5TZXqYcI3fakFbGBQfkvzfOLrxq5eymbPDDh9J95kJoivCHFgYkp
59C2b13jiOwdBzhhWxWTC2dphYjDV2Vq8B/LHhTSHK9h2CuS2ZfARTUomZ0wwKIi
RVqNnr8igIqMzFSwHAtDFTCRodilbdxoyKkagKtua8AWDa1xLW9MOTsRQc4tPwZL
l+5xSfNnWvIYj43sySbtQMOYKXtD/lY5zK8M87YO/P1+nM9pyBRrIXdYRnRULm+I
JJi7Rd+E8+kfaGk3fl4NO23FK69SGBN1UbT8mEO2CCs/0O2mCLDxVZkTt3Pv3Xaz
71r8SGHLn9H3F7hWJ3W79D8/CcBpr49C0fJDtlpniTzqrrQ4KhqeVeTtteO1W32L
rewRIBXi5baQhPjr2e88XNX8lcRwHosqAUlYUnbMabFY7UCXdza/KsJnlyjIOoZJ
Re4904ONnTohXYxu1ctAcVCnAnSDY1k4wKiJqLwzdBQjFhd4YiZOMSCKAmMoMpUZ
suh6kpAijyFgNR/1sMsqKaYq3ssXw+AkRND16Wf0fwekMzOEP+eDa0iYQcrlDu1q
P1FMQQqudsTwBypqfKGGRRsXhplwRaZQsOx7kT4MjhUxStgtwshWB3Gj2R6oxueZ
TK2nsGWFpAFqOj8FeK+bM1IZYSktu9Y+h2JhWgz8DSfi5kj494mOTJ1gDb7m2ALE
a68SeaVjKZGqaeI8wsVM+BbZfLGK4YNbapQEcyIBRK2r98Atmm5vIVwtrueqR6pv
24KyqdxnQD/vKGh3y3GBy+6JuYye/57bmiCKGoX6Brw24xugF5gLqITd2id25YW7
5iFMUIBpL+chJwHg87drBSiN/gs+ZtEcsr8LXD1qOF7UamALRAvzn2CNY/NZ7iy6
1SVFfeR19FAlARwLGjn54hyQluzp28arhK0kiPCOPotXrNSZY9d97PiXYxGqJ1iv
Lgl+HzXuaSS3CK6FO+FBjqWUVrMnd5WsupTcuAKPB4UJU6J8peLZ7IGCF1TL6bxQ
f0tz3L7cPwBCbEBWLkKXvtTgaVOzIKrKUDT9c79aWg2ZiI+IjXl2BNQipCCHiGMs
U4nJeAgv0HukQ/DLMh3Xhy6EdJQx61VnQAPmNLX2LJz2ahFzjweGsvWW8a2Ch+Jo
A+tLcVR6nsSodCA+6kvrsEQhOVrdcS/p/0q8NCm5TyrYZ/YAzBfLsPmTLEV+hZ+V
an7SJ3SU+khpjQgG8PLCcQ7z8oPb1MHwnm6aryWiqXv4XVKOJ5TO9OP0HjG1JIzi
015D9J4BXoZAanC7ZxugpSNf4GGxklA6GzJfJ3SByyCx8g43l2UX6gTUjHsHMiC7
tVXwCIdZgq4iHQK4qbLPEHWoMsAHqFNP9sTRlol1UNswmXDU9/BJAiP1EemfIcdE
`pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KhNwASf1oTKEF9V6MqKoi4OdBr5AQgeSZ6Fqk0mmEUtmFnv9t2b0C4BquZ+2Pl3n
35sg1wPivvD77fQziqzb+H9VeI2amiFYan2hs6IwYDJMNb8Xd2x5g94OFZtM91Jd
JKCKFLebFkroi4ZIZO6h/HCvKObBjX2V4ypGE0Zgjac=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6208)
ow4D9IHtWtTjm4+x+694pr6AJaqJ8camcGBDwwHJkaH8DNVEXWs7kWS0SlBhSRoO
rumgsprHtFwhuVFCIf5Qdl0d9A/YzFtr+mHIoLR+vKlva0ksjFzRvPJt/lBpoNuL
G2jhz4/wYq/LPYvW9jkirl4wbXhxEZJfIVGyRhX/4azGvylNr8O7mOlRo8tBfMuM
ZpyXAQ/yDbTGUuwIZMORoPJGtVYjdODkGDHyGZGgn631xnIH35joNR2bCFJ0cGvt
iTiN54IQQcvr4z9Vu9HkLK9tV5qTYPZTaLmzRrbUTAgRGxUreXCVZB3y45hLWCyi
awX31iHnUJvBG98HTeAjff/DH03WFK3Douv1XUNmsoHrnqhihkyVTcLK8qC9oyrB
bz0qJDCx0BUbg0PtgsXhaYMirmjopTkb0N8WxSQ8W2N3Y/456LHPVYWzmnxEFo3B
pNrXy7z2U0a4jyAytVbNZfMaESFPdg/e6oaCCnxftmkx130ywHpsNNSUV9RtpXQW
j4mq7bRJMYrqR7D6MBp2v2C2y0RjuGv2Jbo9+qMxlIHr56JEiOn09Hzjmz+Sls+S
zDCUBn9A2s0yi8fIzOPXc3te/JpgG6imhFp6UoImGuhr+0P5EnuGlTRxjJ+ymM2k
O4gWCVZJrEnwSEf3wOmSTO0nOx0Vg/lSe/VM80IGACBmhkMYv0UxcCS+TMDigOz7
K4h0xf3dg/fGds2zk19KZr9LKeixQBPAW6DOlwdBqxC7tMy2QrLLCe57CC9tGprS
9MooKqnDZ313UeJ9YUuN8p8o+hrP8q4aUkOtp5wvdJW/Fxhm8a2rDiZPy4aQz6Pw
8akzlKgDY4Uk30cMaDkOuZeeC77MoOi8hGOOpYRcBOvySDM+s41tODSjJC5Ke7wE
P8L3BpHQW98QxAt2NxfWmZuAG5aBX5HtFRARlpfZX+CLu7+nZcxQieLQZU/djr+L
4u2bJcSJ0Rq/5xiyo4kFH7K4ZfB+lxxHmHhlRGDLUuhi6UdzfQviNgcz0Sy0h/ka
wiGESeaQ+5CcIOybOZkOQ7F1zrRLKSOtcZ0UVjSdEnZ+LdbifECtsQ7HDrj77TsB
0Dl/znuRgicChR66zVVp+Sm2vEH268R2N48ffXJ7xtrU1cp2GRWeV/DA5iQPkIjM
k2PrhGCw3FIW+fGSYW48bm7OrsI7NXFH/aE2BoiyctdtWinWppewPrTk75zXQdO7
WN1VAaNz2It1hqfiSMwwDTg5BgfBGzB3crGD5awzRLhK0ne/JQqZ3NQC5jo3UL5h
+90nPStyFuOSj86G+n/mPwWJmW/RT2kYqRurGNuoKgWezHu1rjiQMjQI8gX56tFE
RdZZ+cnxmeosEBvqvqRJ3yNeOmKPFbwmk+z8bRFPXWpQ6qU631kt5JQ3Pu7Uw7wG
p+FQyCVckKYKUY4VMSbRO2ckfG2i//BNCNRKIeb6i3GhkvRsLR9cXHNGDSWdLBKC
kOEqLNo1PZ2qHDyC3awrvPDUzL5IzgjLgF6hTwYbXDXPqiaKCboIOd82NFMHtZi7
XNabLSb0uqyJC+XfhWZbvjP+5O6IQIjPEWwDMGQIMT3JfFeggTLKsrU4wWWHLPt5
X1w1A2HdwnY9yxR+Vkh1UJatetDHNM+DEJMDF6aDXxMDyHg3wS0BiQ5ruBIouXB0
7ArUCTURAyigsqawXlHJxnLhlPOD5qiDBNub/Pre1AN9D+g6lVhmvr9+IC7B/UPf
7h1PUr6/sfTDGvKpTZHp2NRg4JPY1a332Bxl/cwkc6qQy0pf3qbbBDYhSpbTYO8h
vL/Mg3bkjWrd08JOpODJp4SnapCPXbI4S5Zn7gX9OYUqRQdLqf4bhRZ5VqzxyCT7
cO7vsuhCoYBnWRoWngpjyBrNwz1H+M6vNgORuKl8m8NQ/EZ88B5SXVt+5sCO02Gj
rOpAjskHFePl48fWjY+eEr8fGKlvXEFKn/C0vKRQJfIHX8HxS921C80Gwb5OJpL+
zOiTsgYQjBh8GJzTnHt73tYJ2VhbfACll+Qxc40xY2kx0Ne+5BWS5bRkjK4w1r29
VZhlGTGMPCBGtFVKICmTmfaVRyNUOq9nEvHQ8OtqjuCKDFZzDlyHfDkzFGw77jCc
7AEatHN8b8rZKWpU+WN2UwWd9Uts8ZZaCLEs4f2pgK4vZPv1obbSNt32+1L59qAZ
WMr6Pz7K4dndcEOZYFMMjtCeYBfNrpBgwyZDLBkHCE8BmFo/Unha0lCvqVzY35SX
LJBJaFyOZbcpTMQZFVZnMU1yzbdnx34GmiEmBKTc6TK5Moqe9Unir13ikv0UYIKn
9OVqspOZvoykGnd1Tdf3UBn7eV8cqdBTsWmah51K+LwRTk+Y17Z4NfMxjf16Ht/d
Tj4G2bi8S+rxqEhHhse5ia5rxJps5TUfagM6CpwcqrMmueBZ8/UQU6rpyVez/U52
qh4MGcDw3CrzOjM5Ntalsa7PoEDjT26xtufjiNl1NZPnayyNq1v6ZIXmrW3a7rXu
TAEkbvAC79/0Rt30g5Zh9pnz80ByK9tac+NoAnK8s9RJYBEpccHghBgxujVjJnSU
hkMYRJmS8b0MVgu9MPnmDwXlZzFI6W99J5dBEVCuhe0kpG904lsFqurx7puVDOMr
kpMga5InUy56yexPS0dW0JnjBsuBs3CS8eyuuwYtg5KRt5z9yJ5yubhH5/52C29N
TD/486bR8EcBagNgkS+zEiEzTdVMeQtALsCE96l8CRfRYw5NgmEGI5qtopgCfOiO
5FV7AAcwswvAcmIKHnm1NI0aqZXiDYb7Spw5ISAeV4FdboeXxobhlyVhRyXhF0QT
j4GG6/cAQjBfPC/2Globsd0sY6rWyuMHcGic49LjSfg3ULWjtziuioO3YW0w1YDd
pOB69Mj1dPihMx+F2PYU+RiRxSOPUaD7oOAaNMSraIr+UvraKAE/PtpfrEp/0yhs
xacsRGllElVh5dMFzYODjmttqwn2l0v3LHhcC99KncXK1dBiGwoX0+xi2NXB1iGv
eiWXO3VC7V0YaYBXefBKBr7GNMCvB7pTBmuxm4hgIB3MHD+kiZiPF0BGhkYJbhDj
Y+gq1O3Ou3w1pDeK9KwIiq+J5vlWootgLNEcutDs9pSSh6l0unGneX8cnpBJrM7j
0kPqxX5eBpEJjtpK8n/j9OaaUZvNxyU1R7VXGy/yRwAZsOd2UpNh67QQR6u7Q97M
wfr+1/zYOT9I6foyqoX+KfJ5mtfhpvHl/SEAq7zz10LIgZXtqxv4WgkoWk7K/aqY
6pjs5/APsuYRJ5FUzjsV9KS4jXdOdDIGz731RxzScM1YDs/b67St6C6vM9mc5DeI
5PtZXCR8Pc/qjjo+uAj0j52ro71QImU6qDUb+zzfZdHwvftPygNYYZkF9o3QcPX+
ZwDGo3qdnfLR2vpg7ERuPhXptX46jU/rkNQstmWejXLG2oAKggGc4yDwa/B0AjFL
nV9u8u0GzlVJzK55d2+JE9QPoIOIJUqK2qUlbdYc5icb0z+NvJQ1fHN/Vpwg+kY9
H931EIIRh5QYiTkrpZxytrHz66g5Z5+MaDS5TJ5gqmWnuT46Oarr1dJIkQrQfiZH
uwgBIetpuIRkgEb0NovhXgZV4YKzmeNEG9jF2y1lrH4HndGmV7ehDYTLUNZ9IA7J
O52osN96MES6kQONnGDzY3FABw3552uOc2gJ/YgSGO4tAR2y69T42TrSPFzkaKC/
h+DejN3CfNQJ51lUzBCAZ6R6dd7w9JJIIsbQRQ++voj8NwIK9r9Vl80LbL/br34E
jtd1+0yUrMTsmZm203HlD4pTE/77EpIXvIHJsF/Ow6nal3mPhbckj0EiE3Fu1qMt
jA0BK4XS0iMZb8Lymozt6Umpbu7gFN85gk8SyoKzuHjyGK6QH/iX7YsSSO1e58Ed
Q7CDUizF6+mQBa7zANtM8jNC55Sb5EKiGEXGdh+AjUMP5dfkd3MY+UOKt1h6MGHs
OLRivKhrGnHAA6/RoHb9TDW9OZvprUAO4aD2W3ELZMSHyiKkeRxPFI1jusmbk/61
qDgLMbEeJ9WUTUnIy9AmgsKjgGW55Fn5G/WJWSy8a/9Wts7GWmTS533Np3zkdZ10
sUH4OpRZ6RI9owA8p5tlO779S1nKenhjjhjtFU9bNpGAY+qgqBGBpM/9dEo+PLuL
WHEMNaUtvR6ab4YGgPQSTTPfpw/bxHV3dC5XS0HaBGfpefZmYua8Nca2Tn9gEwO8
Hm2YKBlaSsvOP1vlU5FlYUVM97C14X9ex5SYfM+d/yVaTLAIXiylyY3YtQuLsQL0
69IkjKxIL0SufvvtXsFGdh45ndPflykFjbf8jP68UacS2tQDEAwmdCJR9msG3XIo
hrQKwUsrsGSWgRsMx3osnazNDz7rNAxiV88Id9QSIkFoFdm46hBUBDX7pUAJIkCr
/2AGOzSai//ygV3/3uXFoLC4M7SjQyZZXWxvURwcMnk/UnOw+baEX2Minp5QUauE
wJ05GV0muK05FsuXIrJ6Wn2MazN+fscS/U8TIxwVOaNpwDdZxbnCeOLGtyr8HOfc
I/hfNNUz8hCdi8sCK8T344BEm6yQHq/UELeNKrOAU3eiP7WcVCjWO34oi4IcBFIg
zOqoZtRaJ7gZu3d3IgPAR9fvaFYcx6og5Yip3iY7sq0FkqU8QYOc1GgBhT5W+Ykh
nBDvcaXWUg16Mi3OKGHBzgZLgPM5r4PRAHp13DzWIOA5fBqKNJDZrc/ckJuCHvsR
zGZQ/oXMS5jb63A4VUPl0H9b++1/aleNf4MBJY2weF55FAUtWpTgAuudlzmV47H2
w0QYrHTumH03O53qplKg+KhD7V0ldXnepb6HQZTHBdvymHTwkOiWoFaQTPW/62Za
t06d4/Z/l0vEY7d523Md8gh9J2BV4/idJMa/RhMPgUilEJteUK4X8HgxY/mJfmaO
cwlTJ69zKloj3423SQ8C6HUhuRsna7r11bC4DCyIImeGniOgHfrB1M6mVXand12a
BYQUyjuoldYbe/u33rVgVNv86jXLYfe7RRClgG0SvieoyGXI3hlkoTHAA5FsNQft
GMPvptTKnzxqNdSHt0d+LF0NZkR8RZbeWFesPdnJOiZny8j0sy7ZJ0hwkQJ8jKly
kweiCVt8ql1ln+xdQoDqV9nBMn6J0zJ/LInVJAayLEdQP6sfMl7+/woESyot+81O
wX51aq6RQTdVsbJgOlLEhZqLd+/POyuCK3T7W4Euv0jXrQPdgeEmB/RsrdpVOn09
LZaO78hqCcBb0rfGInfZG6Kb8BzLBy8hveRKeI3t4erwwkjT23iGoOcxB9jEqCf4
iqVw+4BYW8+KJ4IZspFupE3dQoPy9O7Q0BsnyyY4BR8st6njhMRsYKxNweAH8ffZ
PKKCO5d7l3/vEQpmUZvI4mhOB812HHm187WaFt0Ui5LooocK65HRQd8gmNJAIk+h
tD8xt8/7u8HbH/oTjJLcH/vBXPd0Zl0A24lmmPi2qvoIUEGVd3gRL3w9kznIhi4G
s9OwIHcpodI7M2F3qwErAlB30ZMG+8U/crvU/9d8/sKfIXwsx1QUCCogiHYS5DW0
lZN+S9qSHGmGJFaZA/6IJ80efoTRLp68jqapm/9wRMeBOiJ7VHAH98xW9mfNGErU
ElHFrYs7/Od+nRjdNwjzFoM9omQwxanoBicFis9DaYMCVGqrjQcQ0Yaf+cnUGyea
eOnSJL+UF4dpgGK/hVoBnFJJZRJEyJlb3mouP0Z8bfCkRNMEdxhWA43ihkFhiG61
NdUYpRu1VBjN2MKc0SifsfDn/I7KMFuas02oCblYbmG1v56csrA7Mo1gq4MeVS7g
lYnHQvfHCteHJQqxB3r7P7T0p8eMkyNtZpohUE/V//BMNBcPYSaToFea+HP9iSXm
h/8o7HgNrY6vuSn9/b6OwdxaSk//PUBtQ3l41LpKRj/ojzddfulgRKO7vQaUdtQ8
GH7uoGuILlEWpJ1tl1VkWE5KfDjaFZ0MrR0Jyb7zMRgwEUpYfNvSNbc3lVEfZAj0
M+PcApm1VD6W+0BpPS/W68/Xzs4ii/iRwWOlfYdDm3sPS7tGKcH8qt3l1HrAUXZE
ZvNZQzgmw8KKODk4D3JdxPbEJ1OQ8Bb7p1pgp3J2LMhGblNfhhp4snK/n9H0jKG0
n3qA9ILBBIXy49mFfZpNTBi6HgBvo73zd0mXjKpfkoeTm9oRulU0kw6aJrnRStbs
oM4BShT2YF4xbSEBpdyXos914wOetQmAsZTukVJ28puFKP43evv5C2rgPUa/M/IK
DyOlRxp4610U8fRG0z/q/4cfGHkk1gDSGX0vS6HM6KzZsmgoOaE+UL/RDzwBmuH0
Jho6zhmrqceXRB9nCTWzPmi0gTLFHiBMujK8M6c8/Eow2wM/wq+DPnM60xnqLweH
Olwbvu2R7X+zqXTSugbegBWHFqXhVmEDbH1qCUCvadRoKFa9S9me/BCzdxn01PTE
QOahbLypSxJwlM/LlKM00RlzsPWLsA+5jl9Ge/F3JJeOjULY8xj2XpVQcdSThcrZ
XoLXcApj4jBN+xh0miwfBUAehym/iD+545wcQ00r2t8mAxYBuVa9S1309D7wPjZV
Chk5mT7yZ6OlmoVX88hM8DZTQSQcwIdfOqGxOGcdE65+pfBeqt4PkVAVZNFXe8VB
stxoa8pjVBJMPKBTALzLsu6uMkXRjNNmQBDxqe4pX9Km7gVPqnI1MKu1H8Xly6/S
F5mp8tnn0ouyZ8N8Lt38YxXfGT3BOgIdBhxmH7ArQcoGFoBNuNJoQaseZfwR68RI
5m+oKXt0wuqvgw8iZHBH+4vFwBERDOrXj+yNY3MPNQBjJMBndFB/QRpmWAIg1VyL
pvo8/r+JyONoURdXWoS0Z+JZdlFox/jPaw0tKDwZ57kbFcZMHlGrF81jxx8Sne4m
yLI/L1O1jeo2EJWH652r3m3Cn9kLyJlQ2s4JySy3AwNsdojKtlAN+/GsgS5EjVOk
yJIGq+R/FCSFIhbmFgN2nL1UduY2dpGdo4pAwmPye+OQRer7dn/M3rhTaAED8M0V
sPitO7d9gaV421guSc7qjcOpKpoCqNB/ENYGrwn/+fVQFc2ieitv2TJtqoZxkkvb
VWZdwMG8WQqjOgiUkt3oeaaCqgR5t1vR/Khtf7DiaIOTaItV3PU94zrh1fP/t6e5
GDe2+ES7GQ1b5H3acQLbkenBMDL6tU36bmbKxpKrWuM7pAH3DLAkx7IvKMYyPPkk
HG9wzK155pVZDFdvUNHaENTmccpACzz2FIUyKBfsxmRkry1nV+KDb7WsnmCPV/VI
r7UkTbTdPW4PPX8n8WZ+jWdA2Spto12shzYxWdXP6ZRgmYlFO+ccp7FaxAAvl959
5ZJhzWjcaRwBoNJUf74iZSAE2pA7qYUBTbH0zpP8gZpYIOgSeYlefgIZLE+7jD65
27SSKFyFN8c+TrJPv58NMn1IZthnDRyNeQ/U65T7mruERIIAnUuEyB43pALybqAz
qNZamAirnDPA5xCtrPYr1ezQtp11YcDNocghko53C+/79YIz3T5u63/FKQrK7xuV
jpgBflUaiWdmDIxrdGaVi+h1FpvIxxywHD/YTKJ2Wo+7HMo5q0k+PKnLrV8LODpc
OJZuc06lo6VxTMBvSURY89stiIADFDJ9WeK8Oy5yO9cAccHj6H+aE6G5ZaxaOsgM
X+g4KOLLke13vLoJ0qsa9HEtTvb6pTadJO2y4VikfXyjfDf8N4MJNrTTF+5fnBSb
/oUBzzdDK7x2/cC+p19O76zWCF3E6Ac+o/AqTGK8eywxk+fybnGBz3c7eUtvOtVQ
WdOPGKYwBuIM5b8YhUpgR86JvTpnwzEmXyVWhbOyTe9ub2og3O7uG5W9tNatDI3a
NAVSIfR7NgyoNmj95vkq6Rnl1SS86j8MhH1KIg/1YOGBhQnaH/6JfAmDGvX1BCbY
6W2PzjdKWOINLpoUjJ7bJgdp5V5n3BE93mGwCiBr2jlFax/b6kQAUJPsNjmGNBhz
07ea/WI/br2RzgQ30moi5ZU/pqSN11aOixLxqGabq8jwTHV0k/iw2u9Tpl4ASZkU
J3XWhV9f3DILeT12A/wFGVLw/ZRpkaKZBcQlA72d6IZV2E6hJgoKA3uZv/IRkL7H
LXvlMdm9Vuub+jHkInHZqpTidP7OOKYtX+TamMBEI2FvxMK10gEcl8Cz8Ccpi+nu
xzI0OOlwW0KrY+24a+g89a3TGhkLqWiTMo0x+PYmr7TwtdhvIGAkle3Nyt36LTyb
s2W6LY/snzzzSWpwpft9wg==
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
naIcIXfWPDHyaq0eLGwlZnBNxk7UfGDol46IeaM1hrbuirgK5xeNwYLymZRUHcVBRiq8l0zlFOsm
njWvZ7F6bIe4oAJR7K+2TH6xpOC3qJEQnxkTcoGxBMsSkAs6iFFdDooFLmTRTqCZ90FW5OCnlL6w
QX36wcPJp8KHlEjEkyJUjbaunxTJ1H+/z352fxP/guBZEiZlRaZrcKhTsVxnYq+eNtqipgEskXFa
n6dJGxiT7SUZADx+Zn4FD4GEpoQdJS01o9/SKp3x3CdY5sWooig/b+WDDXr6tV6GBKjgB/Z9FEDA
a/71OZtY8qSgN1DO5YkPYvary9RwzODKBNQEmQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 4528)
e+wdvLHIGQNeIDo1pQYe2K6c36dA8wp/Kw5RJlMjcXxWAZpENn5yccg1Mm8kM1W8zZrrYk3z6yx5
gJLaKf5J+MVWhbKtGTKjCqgg2ExTgY9p+cHrN/Kod8VYUwEG1AcBA3RDMdxBLprFOuUXvsBepgX2
gxjJMMR/f6w6+Mayq4A7bU+tEonEqYHxDC6jcQqSJ48m3m7Q9eQLBna0sTzBkAxYOhXzlyfCBycc
DIQdXeOcCda7Iwq1b/tc0R9XyRAlVyNeiw1Q+KvYw5jQ+XfsLDywsxX7NTrRfmYTqzJXNQ/WT7xQ
nEZBnVu7DUTRZd8CBo3hGHdYbMwlE4USP4ia8cEaud7qzbrXInXN8nG495SXQwMzpbRQkIpL+hVg
38SwbrBaQVbsoKg+SB7hZIJeY/7Rlflvw0WR2mlXu764FGgSSc9k1/BuBsYA4oXTAqoSTE6EXexj
frm4rmQD4EGrVEWoSr8VnuDYeqrpxIfqRWq+UnRwmsCSDxzL3NLlSjvh775Y+0HzxiWgvC8729AG
+zAY08dxtLO4/hvx+VwSFSEcMrRBPAkokkcl9/nyPkkpXZ6DPFABEZnGBgYTIQ1O4/ylDufXdrfU
S72oARK4rYRH8Y4qEjKOVc1cdoW8ypoT+0U0LtclBTvbDubRSbSdUUc9FcXVwTNgCzYY9pm70DIG
QBu4egj/t4yQk86uB7o3HTnHALhMlNb6eYr6uYelorAFv1FZodp69VUYFTB9r5FCqXLvmVCkATwR
r8ad+fQzYAo2FW0FX6sxREP34DUUT3BI7PvcV3x9s8wvHAuPy8AKBv2mElQS5eIuEcEaR4wYsorx
KQjZVrsMABNPGROqkmto72ouystUjqmk1LFWLH+3EjlGJyxJgzjUH10GcBR4s89kJS9DgCEmhxGa
0QIQE82F8Tm/n/+cXG1bZW4r1XEz24Px8BJ0DMZn4GIaemfrTfsSr8rmP4eu+LQm4eUZtZ8uXwhv
FQECOdXSOnPuXo3T7SRUuR832ylJdVJqDilGrWMZyBh7k0xhl7pUVn036ICCFUloT8wADsrLT9TF
PABppZkGw7R2RiAowuJMbvDssEOhQ7Vos34Av1bMDZ/EIKAqTo7k3oz2ZQnyoz2naHJ+lZlLg6Up
1W7FUgIbaWMH8YP8EODUT2m9sRhiwjwiNGdkogFr7Xs9VVx4LbmxVWR9+ujFYAizWSD6llnMFQ8N
LkTaRihKTMR+5ZDnlC5D8LHvAHjXGKq4MY5dxV+fQlmvUjijblz0kd+LtbBOWDG4QITbOOB+lH3B
YR3+ecUze6oY1U35WwQckRY31S57Fb15F5suNLGdr6xi/H0+UdJLbQrwgUwMnbLXvPvu2TAZbIiH
2nsXXrsus+2rXABt5aMcysCjDV8oogaAKHj044wrTwYQkArmzgPv27xRVLgwp8FD6ga1eCZFuEL5
KrnwAR8TXWqfCTwFRtNwG3y4WOhY165CUO2jfl6YFdomg0Li2JkERKUUEN2BtNnjxqinvUk+fQ8J
LsWdCm5ZkVzRXvhnML3Dv0M5Nx8q4CNGeH5VQHZWyQRcuMLavPctrmWKb4ItqxJke7m2u7N+KOKh
O6h0onmFeqlz1wMhGuXb6B1cXaxL1nbd5fw0LJ7OAJSowmRrso65NnfB1x2Ly7E9CLaLnNAGkVI0
slMZur2t3C/rePsl/2Szxd+bPPbG07dgvZ3g22RCTU9GSvMgAcI0vIsTi5z3smq6VYe5vsjK+VSj
oHjpeSvKmUnQUoWRScUcIn4HSQoO7t5ZIdpSI9eJlUlozORWSsMQ+P1P3i5qGHjxBfwSUt/U6PuU
lZQU+c5gnahyeR7skvjeASPKnmrSNEy6zEIldSHB/IstP6zUFIV+kZYYO79xIRoDzyLNIUx+2y6v
hecH6RC2HxRmURqmUwBdlDqLfduUTFDDnjil2FYqLtGLu+hJeDx3HednfLacFDKDY5Ojd7o4dzQo
6K1yrGBaEUYjtaExqjyallYeMb+heC5M0h6MfziKyhHoyKWtVqjFmJ2C978t3Bp+q2Hdv5HnFQqx
EcWz3Dlz/5tCJY1fANZU/GxAxI31NRSPyHdwlRG3Lj7X72gdbyxsbrZ6XWXlTm5ztzPjgs2d/LkD
a5jqM5PRjpQC1Uz5kiblFds0L+ynLQsdyjL2kuq8OQWTbPz0J+s020rFGK4PC16YaGgaP9CS/Z5D
owLHUV7xUyLXa42fajxCo5KUtR78fyOgMQkpJpTNxIfzsx632j3s23N12jDptiewEe/I6FXWFIf6
9ftlGz7gzUrAQhem7RrdgWvpGYJnnzLFGyAgyxVLq2gIPXWyrStE/bU3OOJO2S+r03Va3lzTgjIG
+jlZWRYZhnA6Eq+42mlXQwH67R7yqrBvCbIAruiHhBUsp1W85gCJtIcLE5PUc5twDnTzr+1kKPOL
A6ZrG0/9Ol/qpwCX7stx99Gxy2onWD6ZVVWwbYRNZyEYZYcCmFI6iQmwRyD8umWqeGjFAjBoZEWA
DWIQW2Wl+q6V47IzNWZxN+Vyh4vpKAgLMvoz7e5WLBuRyl3MI8fJneRDt+xmACIBUMg7E3hhWmuY
twKQaEKWtS5pwkiVfoTi+xCpqHQfAj8TwS7QAat6k/LOIv4QPeGwZpGNvHI3nQ345Zn+lLdNXS2R
Srswh9q0WEqneI5Unpjozh37WOioLdzpP61p3H9ISxEbi4coDI7zUA+p2+7NyuVmdcDmNXORu15w
pi8EHKhuPf0JoxIMHzNb40CXykn1V4h0GPGNmYnsjpZPkCdCgHsRcwhVc/LL+QCJemOoo2wsLzgo
EzPTvdOG0rYuJdIwB73eh3BrMmztrz0nN8uXAuu4zz6MzYq8Fgp6QQ3gIA83aL5Hw47kYzeGIexK
Ktzx5IuVQkL+Rh65SmuX2BmL/k5L7GBxMtBQU7qUm05he1ebbLDHomWTgKCi6kPhdv7bKV68FD2m
+FTvRQhBxZvZpoMswquZ/xAxOKiYGO+DxjahKeJtlfbAvV+ZXJ90sPfo0KPQErHIjF29Z0POQ/Rx
LnIGFjQggATWEGFzbc4bNEWEDocBzdgUe9dsAek9da8Q+x1VQXNipYJx/FhsMtmVM8dlDxonLPPS
W0f7z2QZrKvAxqiG3kt9IqVZDfz+VYXWFOi24b9twucx3IfXEIX9Qo7NIsRRzRXE7zoeKKjqwbvw
UU2TZIQ1WOO18VPg//c+9BIR59hGSAoJfQXtOSr3wfGfO2EWrFRpMCdpMGj1URR/65zd5NDdBzHk
3uddmsfEoG4Tgc5DZhBcWgF/Gdv/w3YoiOn6Gvhppf4AxmZ4qTQFUBI4LrzRmtGu8RxJJeWUbI0D
lYUN7zRG7azsT+2X9kbnWcs4m5hACKnSu+73UAzODXA1UN4/8q7HzdRUGhRLpbqp5ZdHlscG3hbI
BmVQ9C+k3YropgJIonhVZ0uIWxIN5Z4r559HWBZ3F6RDZU62gq5bwabO9TlhHOLCtrz082JAi1iE
tYE6lCwzUM5/q2GmGu5ZdSIeKFnM0qAIPHeeuQK1R0azSI2PO78N+A/PFtjW5bjbTG/8kizlrO4n
6NhkNTk4JIQa0g3sP6Nl2ust9DreuhpVhPWc0Wb74kDmhwycs+2EJwP884IGjauC+AWvFyPGcvkI
z8uwWWL6I1qrmWzNkQXDPyQ2AG+yimJlzMBOVP4dSiNBG+gozut1QhvCHClXRrKtnSfzPkPKw5b7
mw5j0+LhG9AFfYijXyg8//mBqni2Kh8+r2I95H0vSuyB9guJhwd6adPIJYIllcCsYwSrbUiolVZL
+g9+NWEqSuLP9edgdrHRGeUU3Y7VLJSxX9DbSJ/LrOU52t3mKaSIjRWSW8+mkkF4Ne8skPX54xe4
CE23xCQijYlTe0B8fpSkO4OdOwZHmNRTzOTtQJAWWd4rF+L2lmIdlxEXgbrn2Nxd6k+7aTC+D8iB
XicBwrgrnZ7tOOSWhO9Oe86U3iySwnuJ6vjChmzWS9FBsBe4UBUEUxcFt0bOV1151bwmUlwXN3IS
W1popoifVCN3rU5MoNxtRR0fXD/mZqQqxeRB+UiGmhmBQf2dOrBF1dy+Rjp33W57mjOmclYOfszw
s34LWZeMK9zzmd1uvtJv1g6eNQGmZJ9kR6CgztdnnJ5UCd0CwUCRaEin64TMayUJQ4AwjcjTXSEQ
6D6plBvu4JlY/eAmBJVslqiOuzyUg2nR9ZZuocTdt73oTi/OBnOJseVDJ5sYefFPhUM7A0wFMUP7
RrnCoR4Hu3i3C17rAPYiyeXrIbC6YD0hT3+Bp3WmdconuKSob1Nq/s8wqjG/rIipusjXFHwaj8cF
BNNXGlpKFLRj2bITDwGx88aDZ9hQKni+KIA/9HGT7LxhQNLOzHAE8pYV58YI+AkrBvv0h/bPOtI9
LfQrU55LtHclgAC0/d4hjb7coEXWmcoUXRyMNm15qmj5T8UN74F9HvVnPXqBq51WbYI7zEt/kVmt
voJVSkUIFoTA16GiVzkarWfEwg2D6Dnaf8I5bcthf8oQoX6Or4gn1T4FidP9u646SYo2zrJua5A6
/tts61XcIhLLXss9fcAMKiYMZQqAPNJQnAlvuFcahbvccK5vlGMwlVBK2z9LXIE2xE8yDh1e78tb
+zNSbWbcA2xZCXgS1Te3UC58KbsLBvvJv7atEoFL20PLjLjXwfVnxX8yRCYZ4kfISKKNsOzc6qHm
g4a4rzGdOvV8DsBZtiYfqau8nmC3h7a2YodfPMBebZrjtG1ezdSNkWYE3uRzq+GHQ87h6iCcUY5d
tq3brGt/2o6522Fd5ig1ZmHiSwGFGa2Cu4PeN/9rdqJFWSWFZt4ulZmmE/gq67J74zr6qOQbtUTM
0U00gnv6RkSP/erSMUlFTQH9ATn9Q444+6FHhcw5Xw8LpV8utrqdLJBhoGqesRZiQR2xlO0KbAdT
bK7BYiFQE25/mAInkRSed4BEWOst/vZ8Dxdh4WmP3rgA3Y9VbGVl2yo877ZhuvNREyJTdnlAD8iT
A+0EeoKBo03gcXUpctkrrQ6eezFR01b0vXPKVNzqYdXZ8WjqxmtATZ202cByI142bVD52guSWdR5
2TPPN0DYn6x3VNIFoxX392TOlQxD8LoEmUteA6hDJUfInsP7G0QnX3HPXyTyyooC2rIqaBM3PaUy
PyTFl2rSLibYtehzgBGQApD0nC10BpnGbzbKbMn3CQinJcqe6/O3QiCdglHaRX9w1Knx6lon1MUE
W4GhaoSqMIgZcG97G8hCUhoH2oYA96f5tYUYOPL5Bf4sC4bRwUXjNNS+hnuxI/UJjzy6WDxrBN7n
rQ+gGyKHY33iv5wA+gfq0FnI+pDARigYxn3WJbrkY9U7WJDwObYxm4fju+MtIF/cSuSbtA/UgrbE
uMB2LJTzFXyd8l4/0eksAWsqgXccuylBHfur5QrWf8xc4duMXGkXXXCI4YIZ2ZfbWYoM4NdA3hR9
DQCI9Fp1ktMbKgs82SqEjPMdS6six7BfL6OFhguOyOwJBcrRDP13TBpEPcDn4LTWHeWaA2F4TlGT
Mer68QDjCatOUZx/mYuG+M4LcQBu0Q5Tmr9bwFXFL6GugUbUG3McvADYbvDtpPQR0U7EniIu2v9x
Sr+CUQBDEGJ/BZvbTHD5XWGrSMTRu7+BIzCFEduJjBcUTrckwu9LijA4KgT8FUs1QughGfg/ZOPo
DF6ScGxCgfZ2MzJREJuJ0bidwu6brZ37+v5oSbXeGNcb11aoHWCM97cpGtey3/BzCSuCxVsBttEz
HeXIJg1MZCAtz15XrULkf86pHw7awvsftiwt46zmOb24iOSImVYJEd1J44egjGq2JQnvOj9oa/MH
HCuctIR8F+Zg0jrf4FBV6pXL4B6l4bnCtxngE56bPJ4me0/WUnPXB3NCRBzFro2WnMFtIRoWb1VO
mOtdXWGZcFgC1mKWF50Zrn92omFNiTzrj7ZjXC1lOclS1177sx4HvRr4uxB43yS94NAoXbDU2eTj
mkFRXrVgpcMY7N4Aj9dKMqD0ypu9Rko6jg==
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
lxw9ol6x3JrAtILl0/Rz71Rb4g+CPjp6MjaJMbCHh34NcA0tdurWfsVzuhamoy6T
tyx6MEktr6KitzvruEmJhyJzsBz+WJ//7IZ4x4iB2r5qVB5b7SsnJCVb/big/tQu
2TUmWpP6WUouCnOXao28Gur6EWtBwCMhBsr91Tz57XpYcAn4LYD8FNN2ePkCBWwS
c24TcnUoxg85CgIxywprhUbPWis+Be8H6OT9GOh+YGq08XmFKa84IBvaYkpF8qun
Q3iASP6tk5pUNG4NajXu7lPb+lT7jtfGlyKRykO4lq0I93vQ15s7UDeGDsUxNcVz
TbIXU5y6T+p7VOb40lYD9A==
//pragma protect end_key_block
//pragma protect digest_block
1d6cIHCME0MAMGstIDPJt9y+gg4=
//pragma protect end_digest_block
//pragma protect data_block
3sBE1Ai7xWeBwtx2JBffLIqXfHEbqUimLnVahTX78sXp32i/m64alaY6ggbdOAMk
NGOF1rBp64kjP52KBzj32+4HxZ3B6f4iAEBzen3aUYAj0LzX/58xs1C26GJ23boI
+IgUpmq4ewIPW5qvigu3MHZyyhKJnkNX+l6hnTtbr7fhKw6d2vt36Ku6hZFnG/BY
W2gL+Eb7IXexMUPlNMjh8zMbVQLB2HYWqLk8cbLZNG4GtS8x503qoIJu+rQdxh3D
vibBaPLZcTWY2vNhy09h9VYRxvHF23m7zzYZ3SGy1WEwF80kJ70izIMCqCC7Yffn
Bp0ZxKx2nKIplVDHtlB0akTpPm+TBysbHByBzwyWehfF4KMVVs3hEtB5TYCnopnt
WXrIFreA3gP+oxtOriP0PlOdUqmUsocTosNqm3c8GckL/3BRHRD+wPsUuhFhlIus
LoWm2UbcdRLDJ6jgrRqhF6Ixn1JiYDC8manSyk/0/y3ihCK8wWHmg5TU44dKxWZn
JeNzJynr+YwpCU2jP+CLpnPl0i3sSYSoXysfUMq7AJxhhCWxKvOld5ybSIAclTxG
pINzGvub8vO+lcVefKxcChN6ookBuy22/M63wdbBAMgFA5OeaHCxlIiiphDGF9ey
EXL9AlVFpn5qHMgEDDPzIx14Meklk3ee4vJi8Nrm0phjPODsemrcB39RtJnVGitQ
jI1DzUcWm6ZMLe1h6YMxR+AvO/65ND5Uo7xN6RsksQ2olCdKPVK56cva7oW6jMiR
HLOi8K7J4IhYD/lh8BNJQM2wBtsea5KOTbZ5bHJtjF2Q34dhf5Ctuy6LCoHpwxtx
5K2sClxPjTjnHp1oSzybfWTco+1CIVYMKd7DkhBX1PxD1iGMZHi9Gz0k4W8ThJio
qIp2Mjg0nHSZWyOXK/U8MFntRFK5mEKbONoeWBt7uZ5+4pB+Qkllj09k44X0YOL5
a50jRzdRuwcfH3cL1pq5KN+dybLKZ+55nSc19+ZELq83PvvM3wK/dnTzGDfB/hpx
6ttBmiCaTRVaCmtTyOfktCIdUXSwf3cl7ctqSbikmdQtQuhLGqHvdwqK7ACdrvXv
9XW0oKULm9O+roEjmOZR9eFyzjuJGlIxOY6Nk7VKzCvGswpxJQ8p3+SCbJKrmABr
YvItoCmv9cXcDsnkdd8X2XWIm2NiOYZKXHwJQJjeVIZZcvHalIC1E4JYN3u4z6Ov
WGRYcX9JMUwhEQmOvVB1wrC2xHXRsBYA19FvtauPxAzsKa4ORLMcoNd9xCzbapR8
7cYX8LmGS1V5VkZ4YbyoFwuKLK8YKd7ycDA87JY7Ep3IzPpB4gt432crGKXlq/9o
ks7iZkcaKM+0Kj7g74b8Y3706PKXBgZibfFu4sVIVkEQ0jDlDUKm2f9dZEJKHH3T
VP2sIn2KqDSWDz2iaknAF40OnC4atPeyDCcZ5VEAs1UsbjSiYeEpUXXX3uRPomlq
4XWHYz6wx3cvbffCxMyxfxF34gzyDksA/nLLv4BtjYpb6Ceuyo3mtsGxh3486y+P
HOQGtTdu3f6XTXAUCHc1msmHdjbRCWwgRdIEYtTzOJhQcqg1BF/Wn2F7RxTg1c1c
Kwi32EDaqp8lgXHMjUj5vDLE/oAv0mTY/jwE8eIHEiUS9+KYvJe1ouJ5f8UB7pLJ
DZJ8WsYKo4OKFXtRj1NfW/E3AC7RCdK1eXdgHRzm9z2tn9HyuG3/NRqTuzjv8vdG
2P2pCP6aaxf8cQfHiATiEq9N2pYuo0Tm/SkRrmoxX/ZuljkNDW8Vv+DEYH1S7d65
As+8mY9dooMxCoO6f7vc3lcp5mMwGIoWJktH+z/hO9HYz5jtYP9zIG+AJ8bkUzio
NG3YGrl/J22bgmbP5K0z4rgHyPoFkcuK9ke1XSAPrheA1KI9WN6CXlEV6YuqQ1ti
9nL72qQKCtxxCv/nLAL2t+0gqdXAh7EgCQDoS2SUl0Kx8ZUZp8W9vV0bou3NalLx
MSSYJc1AWai+SbM2hKtW5NdLyg8lKGjoef+Y/LYetAWak9T8GiLSYr52Mv65MS2J
LMfWUc0D5Q2FwdvefDeVer0xFf9B9Rl9/08REdVWi1umu4AJOnIijuj4iPMckrhq
1eMKILFtcOsWJlv/jz57oPbULu7fcE1yrkwUYIpxlelxDWNuXBhbYm2Gyt7++YUI
K4msB+oIU188Kjl/d1e+qYc7FFtAduLxVcdQFlXvDFlEj9bnec27JZNliaS8T84s
pG9xBoUna8zf8c9cakQ9xNvsiWIdku2SVNhWsFR1VFx6PxLanP9SRQ3/12kxc5fH
GKmoC5qNb9Yfz0mpE5/0r9k9JgjxGMbar4rNswLLsVCHcBgaW3AV+Cx20crpgPDp
DjRrktZbshFnGHCbmpGIaZWHwxzv0PZTRP8/3uA9ukxwINdpql/GrJErC0UjEvFX
JsX9bkWFPnSDWRjFXO2rOQMde1ucVZZrGW7URKtBGzKxKO2fyXEB3/48/x2GyA/e
+yOI7V6RAbOh+RUYtaP97g09wr2kA4GwucQPFA+GxEjLg0vJbbDWb3ABV5oHsvHH
ZTMJXI/iHhLKqRTTRGcigWPcGVy4okmq1zf5arDTfdczAXDnMaboRGbIy+ASx5QZ
HHZaof/PDlsXEwUyWzBOkOvhOFx7UN8dAFxKWvpWzRVZJDqI3vNi1RHy8xQzN4ga
p5B7iHzuw8vLtpdrkQFHF2L9CktLTWb/cbSAeRGeoQJsdGUpvIJ9GaJANgcGJTr1
rErwJKdgjy6ZGJ3v21xLVVPUa5qW9rATZAo+JH6sd2mQHCx3mcbGbc7pENv7wPRD
xsslG3YQ27uMFd8rDgUlCY9i9WPnBkysmbCElXExO0ZU1nEGB6X+8NEWrEb7iuiW
3pVMZu3jqZNVDM/6ZgWBe2xt0rKW1ONxU5l41NZpFur/Gc+JdEZR4JJe6p5lx+2x
95uOUoc3jAx4K6BXZMri7augKA/8c4sHluV5QVaAtG7ag2lftfJf7X5iNi6QUL1B
yIny30jasxxZtSXtg3GPpKHvDkHxQvX+eoBpEiCy0nrUrWE5iwjRAUUWBKWbatkq
LFWlKxWbfuKKgpy4PSUFxD15ftu9m+bR478ogSLa1R/lDph2bJdfBGujV3imnzqD
S5rJCaTCOswkHBoJvFuv0eIEqp967tCtj8qABR6Dzmn2de+A6ZWq3lV8B/NZcrkr
MQOPvYvzfBCf93s2L/0KMp5/gdcDqtYmygQGehn78YiBftSQ5ldpWNYWTc1hiEZ9
i8BQEAAG0ApIrmcDxIuYfB0QSn/WMifVrbp8SFzDVO71qa53/s8XUmPnDfMlLFin
UsTjlG8QdsHJhg5LK9NTyQvf8bbGgDwf77BFlXImAL3g8vFAjO+0RszkqifrcVPq
DvM6GAjt4qEM1ZNbg/JAhSFUdvRa8+bbbPEA2UwNT3Zp12jW+fWKC4A3wLLen3Wl
4HK6fuX8DE+oZnVL/Ec9+3H2zqr44DayE99NW9L74335A/qRRaYsxrCl07RVy4W9
otVBL9vIWGH3ZD87+3ESS0WFFhX5U5kHZgtwS+ePJBXKXqZ33ddKw56fQmwOApLV
5LdCgYsoLMcm9lF7H38dzx/LwakeIOpBlfLBFfhE3u4E3UVVyK+8MkFBwGvIkfOt
stk7n6icnSLzl6k191wFkVQJ9/45hWKCBvDqAs/m7H+0jUAEEaJRm3sYDiEqHti3
O1oBzRGVVcMxj13Tcv9/X1e9ceogULIyyReVzcYNw+F3+NVjJKM/dwq9gfCtjBd3
TIJZGfltRXQM3T+E93R5a01t4G9IhzYmP13WedrXO1xZhX9yNtE1GrbTKlNokLP8
so7OCfgGRwgpu25wpbIvLBzcMHOKg6OHAm6XIbTUwMYLgXpmSJHY7CM51jqBJDd6
20cFzUiV3RuTm0E6DgfdKunOjn/jNJWRqoS4r4BepcL8DXrnttUL0E0YabTSUHvA
9oaVwxTorMAkPwieNecE70325dEu+NyONeml/S6hC0PS332Cp+cXFhaHouR4DJP2
tu0eC2oocP5/PWXFWzldslqsSEPVPHwRs0oM9qfWVE+uyKxUjfhT2samtjP56rFX
jIhhPUnVeo4GMBnN0GYFkjFlg/D+5qhWxDc9tfDV3R/+B+gQ/Iid1ibDkuKFSf74
jyZb6xC6Mm15W9RuVjq5wzawCaaHKxDBhd5FcAkv7hygslMqzb3aC6cbdAbdYJHr
5SS+lf55jcnBlp4T8IbN8TU6wruOalT+kFCEDNmjnxYbQjYfBEwQbsNZngL6LMNW
RaY33vXm3cme0c1h0z53V+8N5XI1Nj8w/bSNimyUFx4zLsxugkAkAdcHsBPmPoC+
MxMfJljiItSG4EStia9jDbJQrVYy+kyRuLPoWhSLDxUy8V8XG9e2mWhhbDo3Fjfh
CnljqxSUPp4nnM7lCN9ifX+Z9/U/e/wPdJ1Kso/P8tY91bfw67Wcr2cUt7TFXmpQ
0Rry8NWaPoRDHZKvHD4TV4UtGQMYKeDTVCCDEnD4MDRmp3OWWlI8147FSkL1fdbw
KKuG+XXtS8Vl+ZF3Ox64a+79DwNnefKpmrT1BMwy4HLoSJECNks4zWVwwzH1nXxu
RbJ6n+uG4jfNirJRhrSr7BSnqimrBKOYnccLH3JQk5voNcuCdQWwRpDCN5DoBkvZ
zwqwHEt2I0XN00BtIByDUH8AQqfHlzk2MQGSfX6eGnLILhlzpjWThs7GiDrebIbl
0j7n7z7EwzsThVZxgRukp0pRo+mJ/Fk2ebjXqJ0ZfYt5QjSdIsbnijXEq25vpo7v
t4l6GuBnKFV1DOCL0l1tu8FzEObOLp9l7zjQPziQCKloitXqMVWV+8YIijfueEDl
SPTh8W9yM2kpJbTMgT+w1fjB4EPdV40pUFnarhtRS4mBG+bGppbR85ZWkxL12nO5
aSAhL0mNqolA87G3kWpMj/l1Kbti1oU84YJCII46+I9gHV1i6IeIRYeGIYvaiCNl
EXpyAjlFqNF8i1qT75m2JCXO1laMJvGk2ubHl3I69bbW3OdWDspeSE3MyiyQwMH9
mhKgYn4mx8+5VbO/jonXMyfypQO65zS1Ll9dHz32LZ+4TUBbG0kHeY7qAsjg6x7l
YnR8Hb4go1EgJ/3HKL6nKVCvRDL/TrlV6qF/j6pTs5ZDPd2tbBbYlt1zO+zdcN9+
10HCWEMV3ZiwjCTGq+tGZ70JTdtJ7nMKM0NNpJlHgh+PkKF3uVGoKP9EcSCy/W0h
nhRVfQr6ge0GW/TkPmQBkLsgpa+1+kaTHOssqTVxaoO2HT4seTTj1vAKZM+4ynCx
yfxhwn7HXTDgGhzpNoZ6/lZC8+jxm97N70imLzki0fisml1skoLhIwyj+tEDN9AA
DQmVrgif0VOGVtxSNRUkFmI9zS3rGL8Tm7LkYrkUBf5ek/8gjYYm9FjQenGuErDR
sLl3T/W0nDZBcAOH3xgOeMVNjyFcn3vTpeiVWTA6K54P0FopQTjhehNBmJqPa0OA
hGysVrLmNehPts37+rkAy5pxFCFITGnVUHP6Ek/kvhrThQBpO4olNyXAWOHLVkbo
vWI3ySsVVbFhz38jnL+5OFKNmSTOb+OVqHmFaIrb3bpiyLY10HYoUiAi1FIV3VFB
3Yg0P2M4qjECbppopKL2UYZlyO9ohbTxZg8a8Fx7mZeEs9PI9uZFmpTKaDau0q7X
/x7ZuGgbd3m4F9AxVDhhAJWdG3FG5CRT55OKcD/cM7H/iP5WrZzrsz6uPnbeAUIS
+Fs8oEFIF4ZvpSq7Xlxb71z3HOKpTtWZ1rALm4tMSiUiewrBhY/lL1ru1DSjmuEL
6L3rwBwzySRDGIM7sHSn2rdnuN6TaJuW7s5tKFVXFCtMKHi2n3DwLtgyTKOLNtWT
1ITxLc7e8r1Vmqh3pko/oR4AZ3M2G2mxqljcdu1FXNTDvSwj/eQWZhk3wUuq5x8Q
fndRhdsa2N1it6ZYkmI5V1F5s0zWPBYOvObWh2gw7ci+f0dQAIbk6SAJpta8IhVO
XIG0/Y63o1waKf+BJ6QZyTobwExhZ9bnLUoNe21wNDg05hIfTJLjMyQ3RI+H6rK2
rFb4jzL+oXXzmq5KnCjl9aQhvqO25rX/LwO6KSLgQwZ2kh+tVbE1bS1oBho5++8t
oAZhb/Tgqimx3sznIU0VzC70NiD1Ts+CbETqoBPgkbK+az4yamHDkvAxjAQ4O5nL
QB6heADd/7n1hHbn1WNk8g/rOGZvdFr6V2L6w/XjESsZO4LOjq3JoZj19SOY0LYi
PIhanV/kiRp8V1mYo9S6x107lTIzpG5iy2WmSxE17D0CqxMsFz18nzXzg3qkHwcL
vFvIVzLMH/W5SQhbce8Lyo5giIpDia1Uo/gG0YixiFjIRJjxhSK/E5/sPGLoS1O/
PsQm03MYkibjUAu9hHco6S7MnhkZjbomc7LCIp+XffbN+3hadYHbnBu5x3Y/UvLI
s1crZYNz2k7JiBoRtrFlDDE/gEIc70ZZS0HqbnOqiKJFNGCItU7CJBxvusDugjYO
d6b3W7rU4pfTw9qiEdIfg1gPQvT7xngF/wwKTT13MrWYv8GlfaEAyO09ZAoYfC1r
zQpk3MO7UUeyu3x7w9o2JMYrLj71j+X3YQHCzHlc9gjIGFBgXSaU0jKP+2M6Z4MJ
G98F8b6ry4+c1CpDKcDnjLVIAmeCT9l9Wqp2sW29bq4EvKCsHXS2wh+z0rSav+3h
8QghsmmwTZtiM/PKydUg4+WXcaqIXnYF+txukzDJAHJaiG55kIEkX+vMeRDbq4Hb
pE4aVp8xPsT0CrpjoG14RUh9df7i7GqP2lO4gliNWH3Sj/Jx8gYdB9BMoAsmqAfU
ALmjiorpeIS2aqju+qtRWUT/Jcybc2s2mrH7yDnMjP2T3Z9UNdp91SZvl7mzdhiH
+BhUQaKQajpi8lf0iGLqoLPvPHfVWa+DClHXVu8YbKTPMVClATjI7hUGenvfiRs/
ATYp9e1e4TjfFgoEQRvglHjNWOuvMeM++BbFORMIQipyRwc5pKMFW3RMOCl8OCMS
vTi5sFBTFVxP/+LPzGEkFPS6gBf458L04UipyaDI6isCTbFTmdbVj//aDsYOHKgs
PL9laJJvTKq1HHQ0Jbc2k8QyCUnlo8J9SClwSMCrok0y+ioL3hMdblO2e8/FmnMl
TG78ZmxXMjtGUh2FmBwBl0jjgDF/pGIghxg4qXbjpYBzmFpM1N5HCmiloYclN+BC
PlCuUEd9IJz8LhliFvwRrJtUFlqpxIJXSBAbBHeIcTnnC4vPaGtJtMTPkmU8j66S
G+YuM3ILdjWoG+rYz+Um40aFRI0SdGzsRmQZVCps1NfMsYpEwZ3xwczuAwu9bIZz
QA924zm/Ty/jspvL9cmCoqAH8kBHaBU4NdIzNp0MvSM+2GWVEVxYz20+iAD+MX1G
Rfwvpol5fQ+h9Q0GP9U98aB1zqjQass7c67kAFMKLxSgysv+gJAuwGPUc5TCXcLx
yPkqvA2tY6GMo4pSapHDhQiZ7eM94wRV4/OvbqQifWB6z11lOZNQA+XFZSG+r+CK
baCDwt95hbSA019832ebJKqrdd7lUqgZ0bSX2v81lP+54YpwSVgU+DtB1Ry0yOVt
0yJIr2t1Wu6SOkccx6+AF/xGH8LIJr17vKmfmI1cPteBhgewQKh3BZxJHyvitISO
GhZMEL8b+9qoM+8k355kuMLCp/wr/GRVUDvULMJZAH8ABgVR8tuMrzWtX0IlvyeH
U0dqVV1rrktJ6nHGjQrQVSJXrttHI4DjhAbdzKiJPiDDJJjSpOvLP4DGQ1dpL0il
QNdaEJrosb3q5DU5nYYeO47tu4QJ35LN95rKB2PcP7iLpBSCbzzLr9P2Gpi2OXf1
HCTduHJ/Jb5OUEiAz9/InZQvDb/gUF+sqGAP9WwbfFIYfXLvBn1O6NEoz8lhcMu6
eHj6REYBwh31pYWOOroFD9CWjDHJtPoYNk+CJGiReFYs4FEeLqRdBJY2Lq4YYp9O
vqyGGoEGA414J8DtbxY6Q0C8RAj29QkWvnMsei/NhOsqJHAJzDlZZZZVQFEWdhqL
UZGImEvMOmSgJ/3N3dHR9seCPt20WyNOo5Sd0CL94MeSHzrNvDz1v6qOeTlZ4+/1
HiPxpAFSZq4sUuVTkErm1QNeaqSBO3ZDT2cZMHRnyJ/l/am/9F+le9nPCOH34/7M
5ot21JkLw5WoupHDRilTCQo68/2M0xOkZ1I3MYSvHz7/1rX0m3mGVvAOCCJ4zmqW
hS7g7tdRKTaYeYkQGI/dbcn2vgtU+7zYoBcgUnP2LigftNGB8Toczo+WfU25wrL2
Me/uo8o2Bu2UYWJqDb6l9ZX5T2duERC6dXU62P0Fch9X9OPSR7sU5wCyfywI32zj
OhKJFOkQFyQ8pFjedII19KSuxQoQMuCN3TGEveBoKOZUAbXuUkWmnmjPwR6kR5lV
KGCucWSfRwYzLmOOvrRnWXCl05zVdcRMpbvp5Chj3Oyy+M4EO8JQDcpA+cxQOIT8
JLYedNroUU7CQTAES+rz0WxY7K1JIAOlWdxBbXwis3pEaNBNy0wAhfRcU993z0NH
nC55xda1BGAq6mTLxrWLEJMoorZQ/8MpaOUp0jMY0Dt7Qb8TOa07/NrvwLdWkOBW
/eRGjFybnXKEs+uCSt1AbJ5/8eET17+N84uofxjPhVPVizFcEFwfT9h4R9R3xwhb
HkN7amM2AjykqG+MB7e2V6XRG4Z9Z21FxcYJTf+70sX2EDZn53Pql9yCiq6PkDb5
3Xu+Kq/cd+YpIwd2NcoVsPQdnK/yDfVrNDXcJ4omvXAq2n31C0FNMlxFmXz798hn
4BnxAUCZcS/9V2chAclQQNIkx3IDY6pe4hlosnLexClgIXdJbS9YL6luMe2O3AOr
u3cJknI/Na+SsrS80JgENjotI/eag7vAqgOTqOOfeJl4yu3PxxZQcoAuqp3VgsQ1
SijPrRvnZKr0S2vVVG7MmH+2UFTwqeLc8fFBv/MSbHdwMOxZeB1lDU35hk5I5uhL
T/l4FlprEHK1v+h35K9+u/Q1lSz2ft/af/yhNzTUnTU9VJPyExmIYtFVb4qzHUWT
/7UXqZxjoCmJXgWIfFV9uPKs0ImLXNq1u9tFs4dGvF57fMz0FOaWrnn1OfqjxE8g
DrpVm+p978fMX/rDMDiMnQL2yLIyVghJxu7UR0rF6iCgyBS4KLbX5Y3WigrPxEvM
1masMvwF7oSh74tBiIWIA3wv4W2H3Ip2LA+WN6KyABB0pbGmD6d9nKrFtpbAgAGF
ZDOqe3py9wT2Hm6CVbsPJRKRanLRr23XBDKPDqRHUi1KgldZICSCABOfnwJl4bZP
SPVP+XYQv4OyAnwmDb4YN8BfnYREao4uYjyECYVPHFNmWRpZxSjAkIjk+rtQ7uiT
e0KJr94454v6hQqDyNVqzXlXsWGGExhJpoXAxcdkM834zS3sKn7k7FKH4oIn6G9p
v3X3T7z8kFaA3VAkULC83N468O05HiCM/2NqH92TTaCeWFSnDSNed1ScBN2Yzpj6
Qz4GcuyqZPnq6FoF7vblJNlqGzi8YgD+tH7uHLtV4TRSOpq0XGkmyl67NyOFFosA
1/b4S7xqmKcHZw07AQsQzakThPzyQtKxN6z8JFbyQcWl8/6+V2bjipWeuYVhmNo8
xjzSxraaDKSJo/sYr74WkA6K/UfDwAOO7Da/MrCPgIxz9XAIhJ7nzMFnS6V63Vq2
Pffp+DXpVzF8eZrPyQdsO8cBqmsXyna53o3Yenejiz+wMdEj8t4K/ExK3ANwPhEo
YKFJY7ZUxsbOtI6X5waHw4q8p6sJ07Rm/eEVnWcjGdg8HtegDQfMQId6LwL4Tr9U
wasalmh52oZLyK9Q8NblTMnVl0ABi1y7J72LNyvHviFmu/fSFhS6vDTLPHzVz/UH
q+GXYgFS3smKvreUjHLuycbpHyaC4Yem5sFbkHFT5aY3sWePpKiNGIsTnQbfftev
U+EmMPpH/UEpywNBGQ8tYgXyzBFxpyIqxnI346rBmdSY0V0F1K3X6TD3z3a8R8bx
kJc6Jp6tkmtq1D7RJIUcOZtj6xi1ujlvqH03mkx1bc+ncYAZtYlihweVoAWAUXo8
fMyiNCMwn2cJ6Dk8fzgizs3FWFx3H6iqw8EDu5bNiXw6irTY4Db6Tv/JXwgiy0ed
PA4ohxZIjfs0Xha/Mqk8WPUMKQXafBAEMOyEQDbdy4QHM/y8EZLZ4R2iOe5+VvDu
EQc5/0BT6wYRZSmV3kRKoJcEfVPk5jRHvi0S96lNeJ8RAlFrkIDzJ/2+aeYvBADU
IkMN42xH24FuLn7en0Z8UZSAFzP1SVi/8CaclKd2XcSuxjAY/xPvMH6btyCZTHPu
AcH3unQgCPvsQC8+fVJszM/O01fNHgTuD308qsMaUk4/pXV9e2GqVKhwy5LFmE/f
60a3MpmgGk/XqwaYprCbYvQ5lMf3EdnS3V7osUrRuq+7LYlviQ+H94bBzYcjwkQd
WVGYNvFOD3dQ+SNXT8YQqLLTaeUNuPk+NlIhG4SgsvgDvnzPNbXKv1Eds/TFtWfd
W07kSNLZJfoM4vcwhY7Ite/Dj1wesCC04ngp33VWyK/G2Nxxwrz0os6OgZ+hsPZm
1f7lW1GcQ2I4z+5Eu3XMp0GUdQrJJ6u5BcZ1QRFc+q8/2wfw/TwSIAgLKs1m1qBy
/DzrBiHixXgqkU6benAh3zZ5vzv/QxoDsZ2MGTOwws2j8VIgfaYTDhtdMqwj0p8r
MrydYUtLTp76ulQ1RkknTiKi0Ka4ONuZuVmiiS2uPIXjc5YUIFtylx4ENYGk9/w7
ERTbSTTiVMA2hSQ6pSHZnGcf9Vxci73UfLu570kXtmZZzoEN+P/RxFHarWE7TcDy
Q9InzxGVKnl1RV7XzhUCPyffsjyxsx6yHTNTI0P2ig9n9LRv2W1vp4jhRm23TPXl
ksDLWjc0x3MQrcBM3uCckHst8xncWlhOb815oVl/fcTO+BpvMf/+THkCrIBOg5Ac
2daHOlYX34Iog5Sb6iBUOMi4fn+kaLKF17UeDaM/3G5Vd5qlLXvaNZNs99xRCFUj
qroZx/ixQuIMx3hC39XctmYReW6a7P87z1bFAH4VQTVnKSjnN2PK+/fJxN2w6NGe
nmSTsAaYeBGrNEYHsOdmMZKNNfbEjUg1JysJxmF0zPsxJsJkMZk3LOy8S9zerOAm
rut8/2V8tw/G8tkQ5m/OsTzih7BGsQmxRQBsnzIn5D4nRqO371vrYm6TWGtHHmIs
AD0sslvx5kHLdem8gt4Af6UdxMIIvK557Zi7KNhyVxS7qTXsK9CdHzm8JI8FuP7Q
t9ut+Uq55PLzcmOlQO6QhJW1Lw3noJrreCmV0gzsBO/a/Hix7HtNppnIUTYxZ/81
hxVKYeYqR6nEKYcIJzh8SlltVD7Byz22JWXp6ViCaZ9EKIm/ldcw5bfI5VE12P76
awO1vStbQpdAcz7blAZSAi+DOVrjw49tUu5T+ikQZrqH/4IKsyKkGmslJ9tI0Pe1
N8EJ1a0KANnVjnadFnxip533Xb0zWPSujG8DbXVOiCqzcXgw3xPQDmVn+Le9nN/Z
Mei4YkBGXNm483X9Oyyyd7rmbqdYMw6W7f+52TSaoVZCZobloiUJ+zvsJzsQyfOh
RFKJjW5gm3rJC6IsESfQDAHLgzNItcMD4jFjXCdMpa0Ry4JQmMVw8c2Nkcna/T6O
wAvNMvvaWt/gcIdvIsb5uQnxmNskj0Yjm6jmJ+V1TQ2DjmAaHnIOG9t0SnZPx/Ca
YqREafqmjMZmxvA7CJDHYSL2oRIxp++XnsHZvTfVlrxcxMAULjtqFdLMxz4K5b3q
pOUk7LK8xD2nFU36gBoLFjdglNTH3oIgT35TbEgFdCnCE8MqnKy2YryoHFc2BWFI
s31QD6krKwgcK18NSc/R8mPUTBjC4Ue9iXxtL34wSiE8hVo0VFSWEmv9vFz494ie
v2Xj8ZlcCmZ/lwipZ/tjsqhM3NsxJJqN0Wyof576gEs+IQvU3E+DN6+QppKCqPtr
O6FdAMmGalbrw3+MjQICb76qXcicbPUMGs6Jv7lZDywZoIANgCpEZ+4sdNbOZiwd
QRR5cQ7BbiGU89d4iPhPP62FKBACAohtgW9e0pQoC1U+bmZIqLG8juHwt0ovTs77
y6fBSgLhKBAFPeYaUE8MBzUvXgc6NkwaHp6jubZIsbhHLvA6qPg/Bi7/N1Vsei3C
d9YyGJHjjaG7A/nHB9tMym7uy73X2P2NPO+om7Sv0ZBvTa2o/9VJWIvax7zfDhSU
+t9RtIHdPjVGPNGtJd+dO5DkjlHG/wA/90yXuIRCvAO9IBe7suM00JNGyUO6Pviz
3IUvklbuh5KBzV4UWEYjJDY3PKxBBNxsl935IKhZPzFBt6abXfbBHg3I3WaP8XrS
b/vof+VrbNOvjbvkAm4h6IwbeKt3xmVmN63BidR9A9UAj48GS8Wwbx5EmW1DVxaA
PsKPXpJLAKckaVLxsejavsOnMV05k98Zm6qiFDRe3b24yXcWAqPHK/I540cJEtxW
VDNDyfjEZ9q/vX4098CAB4eDT2bUd4nFQXY8MqnmXhAq49Xc6ObBzoqdneq54VHU
JuixpRWYeOoDk8yTe1bzeEBRxLqKnt2F/KM5/VgNfu79ZyShY7JIDDFcZbQpe5Se
v7Ij+i8NL9j9l1LPC/zJHLF8AKOnif+uw0qXuHWJSJ0zKLl+DsB60V9Z3uCm/MwR
zUFj7DOYnhinx4JkjhXj5psWpPgJc7qBwEg7DK2njBu4ryr9LORNrW+1f0sXlRnk
AtWMnBsewfJUSUGdUMu74V4oOrSKS6QB9ymOJkEuiCrlLFza8nEGCAritKsXI/dn
ib0SYM6oMJgxgpeKZLYYxtGbuYFeZaWKF2l43vk62AS22OLJOklrQijJkN4zT1Gq
rplTVYZJZ8b6e1fLzr2T6l2HCDeVtD1SNzO6/OIEldsikcDTJ0BGsdkht+UTXuUw
pDiveBi4hnz6mz9nB306dlj5DrqMI3FwyKtQ7sUcq8ilHgG7HzR1+SO8uDh+tvRq
aY9vzlmSV9O8JP0jZK48rbc3hg6YdpS/vVTD1x3JIhlBd1XD7RUjtsbGvfnpW7wW
RnET0VR8tG9qvY49X25enDTaphN83XXPfQVXTp7NB1go0hYVgV30tUm7+8a0/8MO
br6tcqyTC140CaNtic3r7vdiyprypRecTPt10AoHXIwJBx/BjjulvJfuPVXGZrs8
ayNlM5mR0jJkqnkTGb6mUETVs8f3MSYmVyOpGQtfATsmWOCIQMUxI9FHP06Gmcdt
xyXzhob8sDUAG2+45gt5QLKPFvaoXQzyICSGypxG72p3p8NZcy1ON9/cOzoWciCT
TRW1tPESx9c3sWCefj1EwKP8S9YNyln7KtRy9cKHK3E3vza9g/Kw8qQqXX9i3kHy
JYh4xeBae/hkbGq9t17WtPuV5UQDAxSjuLjnfX+8pMQ+fdbWCkQlc4d6TSBIhSpm
D2MVE8pFNhNy/ugwdaGAoRY1XpoaSiHovrUChbOMkFu7qqX022nmgoJs96qSQkEJ
rtPmC3YgGAaQYOkN2ydyIJlFJA/PV0bKlMxB1DeD9o7BlJQrEiDyXw0Xqgqpby/W
yRBWERhczwgatVkXKjubF8zp22NQ5R2/immGsH6ukQOfkHmsgfetVeaiPFADO8XO
yLf+CnmlsfNgOjYOEOZhzlofUtPrCdk/XPV1vs+2Xgu3LunEg12EHty3xPv2n6VL
yzFVpDgysPfVomd7EhCO4EPTolDXJ5ilcbccdULdfQxxywtAJ5ExnJz7Jb/vDXvY
wT5SfLIZuW/D+PsN2YkOutlhG9AaHXkeyb/4liLNBTQHn8vRvoS+bVle/qoZNQD8
E7y7rNYPLV5JrD4MOeqmU/DDaWkRq/2LtFTATzm0HSPEc+xcqHm4BUHz6hZsffOA
xNZmCsq8qmxQ8IJC03WlxWVt6HDZTi6I/qSUnz9c1CJDgFFC5DkXM8begPurS2Wd
I5kXxjxEif9xCsAl+B6BBQ+6HKTPF0nT/2jaR8GO7cXUv8w7CPI1JGHVOgQRKOnl
xqBZvLvKnNsFN9/VV0qFjUCrzGNJdPDWXuNQrCLrakn+6tLzkYl/9mqitKjnhUK6
D5ekdaVo1fuWlmm9fG62iYjv4bL3sx5aEiE52Zk2uD9O+pysBuKIdNoeGt7JHPfO
CcQ5nakxyPmuLPenQMq3BvNlSm/PIqpzr+3EXixldlhZcMQ8qsE661x5Emn+0K30
UlwOvtqvNRia/GOWOr7Re74+XcEnmWECsRdeJJyhzO++L0tmSVH3i2uzaXXxy3Fs
+5OzlEOe9CbBSu6Mbd3NQC/bPJoZy4siSiaUH7ajgFQ4gvQ4Ko3ZcfiUfexfZZio
qZ7OHH/q5hjFjCIeezenqhn78UTnxsTYL+Eqsbyekh97h7VvF352NjndsXpzSfoi
08NQ8R4AslsDthPxSfZ0F7S5PyYX8Z1MO4CzH17Dvj4zkgUHzbBUl3DXpf38+BMg
XtQl4RZeqgeauaU4jlEksu49HzBdT6mB3y7moVC+WuR8kF9BQ5wShdrkNnggjF0y
6deq2Yis85bhkMBTCCC2LSvPSkqJCXDaRLYVzosV4COcmEJ3CX5vRomGBSX2y2RX
kzpL+xY2zxa7gnHCR6zKEhDdGRBNWvUR1qwXxYOJRww=
//pragma protect end_data_block
//pragma protect digest_block
EiJfEQzk5P5Hm8caf/P/H4WqUGE=
//pragma protect end_digest_block
//pragma protect end_protected

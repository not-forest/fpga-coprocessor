// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
d61vu0xWMqHij+fSwpNPEBhvK1mQ/2QwNX5Eu+bw8GJKYJFIVxvItRYLF5kTpHRf
NJHqdqHyNOP4Ww31S4kW8Iy3cD9XNziOEzvhFwXg5qntUBJ9JF6sxF1i8tJb7lZ3
EyS/iB3kRarb0BXFg20/12bw8nwgSHzLZ52lV6eTEw1Yk51jxbEW/Zb+BXN4exDp
BCoMOhbr+DcGF8Y1bea+E07IdsUqaMMkrkqgleZKlzkcE5UI3VOaqrkVOPcH7xwP
SHxkO2DEKtYyt0NBzzHBGLdwcueEg5q9iYS7FQvmIOksF6fczsc2BJE0R0/c4aaG
6SEDZFdt1BoKSIJS4LXQPQ==
//pragma protect end_key_block
//pragma protect digest_block
oPZ/hW94gLGgmi/CxTts8IAwl1s=
//pragma protect end_digest_block
//pragma protect data_block
P4WZ8EtM9K9jc3doh5DeTsOMNOV1dJKZ+okv+pScoW6NnH7CAefxbzUWsU+B9KnW
jccNkkLKIY1XlYSPyCbhRctzf4G6ZvXrm0IshrMGWm/Qo6dBCxZAecU1Smu1DjAG
BdnmdyNU8o4vg7hdQnPrvAozp6ipn3QrryL7mtvJSQ7TmouGHjGK3P90rg/AWr0j
4K/ZpwLF1QGJttyyZySJeLjj+h9V/kEe9pekckXDXnPm3O5rYGIglpRdCo7XggO3
vsBJUM9flKHvdZbht7oqEcQFjBMZNrGEDVcx4sIgshGA9kzxQBnu2D8LJoJq76d0
szn0ut7Zznnyft60uaSEu+oLCP8ASwOOl2XJOjONDaS7joSgKLGtP8leyKsTsaEr
XEh+DDzLcjC0hTqBAhWtS4HXnQHJ0pZxDkTV3wAIIyBaAPxHl5ZvLr0Lhwk1/EjC
PYYtp7QN9atfcXrw9otr88q6cheMecJNAk6AgE/GD+zW8f7kY+cQ6KPspnlflkxm
uo7+f4JtPlGsAjN6GjHiYnu18b2gq5IcIHVUOgIeJlkCnv4r8VpxtnlLx4ALs57t
HOUfLzMe0auS9gR7cQIFUZ1Z8ptIqFn0cDh+B1mUGIjJ0tmHfpl6jufyGFQiSgG0
oQfU/AUEQ1RtHBiNspyAn/pPKeLcJtSZ7NVLdjVNpryCPnV1bwp28StLHC9uIIIT
5gtTdvFcJqqNv7XXuJ/HdRe3rOyKOrgCNvxRd2iVTE46FH7hzNU7UfZkODxzrZ9/
we8265oDPOSDnru27cbfD74YntmsYCKNDLCTUA+zyrnboE7KEiOQEJxBw7mFAROC
M6DhctavJ29ADWPrrA7pyg3wQF84S/3plxsYdEU1gkJ7tP40RW99Fqz8cUUodEzB
Ol04oR5o4Xsf2XO46xwRz/7JLTRSihYFOUsdM5cBFB8PFCQv6r3lB6p8dEveYSDx
kArnNpvQblfVN9OHCMeyBRbH2w9CInvxxB7DRfX5MmgkUnyCeX6frJrDdzjJvYEo
QWYnIa+JwjjQa7wDox3VIBu63Rq7/ZEjrV9ZAhJ4EEpD8xTf/iX/ax9efOcPYtur
pKoPZVVHg/zk76fG6LXiJiwON0/+eXJix/e32PRGAIuZMyUbnOxMZnajHdLTXqIE
Kkq4RvM1BBjPZTTRAswmSlRJP3f0OWdFPDz0W7x+46PDYhjCXXMVKedN8cyEy+3G
o7bate6B7MgBkCYDFR6kS77HVl9QzSyd2/L/4EKYxC5E/azlNhZcHyPLzhQ9W/7A
mD0BP3Q43Ox39/C7mYDCb5U8dwsmSJWWJ6liBLjzck+5sZTp0SoSMh+RMybbv4ou
dEhI0En0/4a8GsOr1V6xKdlPd0D5eaDCxio53k5h4VH4D63AIJeZzkYCx6+O2Kvc
9tv9ivlS1nzoYrVPQ8BrC3K8Yv2ijmWYG4GECqpXZBUl2jmQ+RgPZZEBed8ocy1o
cvEwpwWrRyPuYpeo1sjxPBqwfnx0r2sqMqVSg1kfmN5o/pDOQRHLA32LKiFwBgs5
zRgOI8jRwEm5rdJG6gYSI4c1gwm91OTb/tyWyx7gUiCOwXnXtZYv+GMH64d8xhN/
69t69pt6oBcyAJfX5GmS7OBiRYJ57U916frZMXB0jIxOswzfGql44NIfm62yIZ4u
4rgJ11T+D2GEDrx4RivfEyFzKOkfvtMnmFUJhKNUghEf97NUjpyTsbBGNLxqWika
S4bvrCr1vlcvpo4mPPMMXAZJZYwjt5q1GLXC1gKffS/RbMBbX/CGBy8Qr4YbYSCK
iKluYqY325x/huk6hCApLP+hkS4OtK8r18atE+Yqw2pLoxivdOXkHtNfwHklIvua
I9U716cJoUrxHDAkE8Sj2JAcMiyxy+23XEqYrVwnhC1xI/eoG3AxcDVqYLgOA+5y
5UYI3qT9yiYzwjC5wpL6lMLj2f8nXJx60HdQmDvcghsIhcxwqgVd2UZ1KqDBJ6Q+
x4tOWVwb8BBREKgu0PssB1AAF8HRzy+ap5u0746k5AQSaZn6TozFSqesGfBUsvyv
wcoZLwlcrKVrFWn9n0w4804HP2VRB9xVtEC0yW2SVZzOidrZ9YbMJdmqF5CnGXJy
q5f+XYTRIMpQyBeMt5OhLJwHF3nK/BZfePejHcceHPt6xh0qINEKLAI7/vPATw6Q
dRrbQjIlQYtx0c86gxnUGMx2RRCM8jGB7IeaEpyvzuN9OGc6odNjOxgxFXAW2sXa
FHYKxBmboM7OFTyUQw/474d4r/VKYjMN5nhKZast7nNVBvCcucjJkngcDiei50ev
5rlQBpXvjkwEOha6ugrW+YpGcVDYDjkFV1FOS/L3wkollgBSvsqs1h3lsFxgBa4w
VXZphhQplTHAkP+Emj1aTmScvuXt6dJlujhGYwo7+nNW+kBACMB9bzUE/0Swi5DI
GOgpIF4e7Mw1/2IOhWqQKGpdu76oNjnj6c+T6xLTepJKph8XHNG3IQGv/Wu67FE8
zRLq9ucaH6TJT2VLU0mbtK4nyFfEEVfyPDU0vIB07eXTt4XP1TyVsK1ezK6cB3sG
g6cxc1FTmxWiWrbLrozxvYyJEm0wVrIPgptINdBwabvcHdnKOOd3jK6a8WMl0NFN
IgvikEH6xJJOxbNHdWKXuClHPjEnjbfXFumNVaxCIPTbQZUyLeZneYmB0jvSFRHP
MAUOsV+xGVmFrkviOFlt+OOGU6+l/XFRRA/Zc/5NjGRt2e+xKY1SyY/+GxDsowpj
NG7BTvZlLWbQzUMOdyKBUWZd42DdyT/uPwuICigyGTl49gzWC/7y7mh1iYmmB1TS
TJZ+pGPWSNMq04dsNSCLWMBt2YlVOwCMOHPQoZFLxBGP13mMU0aKXHxI/kLbBCwe
ORMExuBJpGpSRQ+Q4eqof3HKEHKMwNWiotArrgpnBVXiOmjuYAHqvxyMfG9zlNp8
3UdatUvXJ9NGu1wTicXVKRMZepHtw5mV3troWsBFrkLGTYrBGGOvvpH87dhE7H1x
DQZh7lTdKyOdA4FMU10jtE2lSOOLY9Zk5l9QQCKhhSDalRLsd0Ksa+UEtSRHv+xo
6GDSgu7kIfGMdxlLb/JSkvEdchbRW5HB7qB9E/NL/uWleA+a7CL591fl/wmzh7+R
Mww9C8Y4+z/58Z9NT5q2nQJ6Zyu2W7fuhbeYgB+NaVsiAdMTi1VBMot/P9PrJmn0
AAGz548TtbWBTTljapXtomsQgylgBXE2WxGFz86Keim7NALjjpOTNYsF3sMfsnOo
yQ/RD9UObGb+SGcBTKj0oMViff003rx46BLjB3lkDzhPHKt17tr01zeXYdy2DbQ4
TXRLKGGgwaY+/++lsWAqH9iCRRtmR3G1+2Dq42SOIClomP6vKzHim+8GvKEuWy4u
+1TAEFjU++XqXscryBSrVeXTcDqFMf5M7Od2nV7BH4aSSs3X/1NJ8TNtJy+/FVe9
b1Vu8KDInJwo4lTIT+XnDaWZqmpA6YJcP11YwtX0IHZUN35bOYws6AXMHIa4hqIT
b2YXY2sNs9V22qDOQFejskxFQY1IdKX2uiNHeE2ZKz6QS6T14NDmvUulO8h/3Cex
+IhjwTKOuhWCDVO2xMEHogoJg6ZCDFI7vnGy0wCRrqgRxIHTkk5s6hPvCf+jfpHk
ryOmUpvvUxO329cxY0b5d6Ewemx/FB3nfNJwqWUYvZJg7mjafAGuCbl6irBp0NXy
NO5sbIpHb8qwDDgziwYRRUXjtwdOPUymR4Xd/gm9GxXouRoIsDSca+LSSJhOBkcM
ke/mRG0EeQRr46wbnDaoT0dsC43pXT/45eRAlmYUZGr28T0jV8xtv37n+HwcctNv
Osq5Pzth1VkTouajhmxqQCBbpyeBeQ9Er9ZZg6ZLZTh8ag87gyM2f/+KjCEnbK72
dorADEObd0rQqSVWrJjC4+7g5b3yFbhZcKDx7PLX7k6ksiKFh8vdEM9yWfpajWC/
3kgLSX3KHBakhX8RdVyAPZ0dolUOC0g5Z2Z+bntqF25BBzQd12RjW34aS9P6MZyU
ZFKMYvOuBmHPkK70pmifaa1hgptbNeMXsnUDD850QmSfC3o/PbHl89mCLcTC06Sq
d7PXs4Gp8BNzGZrRNMMHmvIWbR52650uZk3OPMYLsKYb/tPRAcu3+wtUhJGShFWT
zRQ3PhoJUW9YiNqy9LFSedEPtV1bn+4VVyrtXnXA37+v9+JiqKu4gulAzlUpIpSt
7qzS3x0YFvI5Vn8dNTxGB2ZHhCwQkAYbX525NF5zllTQeRl5rizn8T8Wdifgdb+2
IT0rAsebu/Z0cb6B9UCNGQRds92WMTPj4e1VPkc3SQZk637VdmxuC2y5cyeATLiE
6YSG10OV2ybki3GdmJyCtOT+x5YdbgqNBMNRTuqojvgisB3QOn1Ve/kMXHSxf1Uc
OZDeLgO4S44DAR1I1eUWNtYV0bfLeguHVIq+p8CH4z8KkhPcpgePu+JmHMuyP1YJ
mnVg1qxQLakpPGb2n+00d8A+yoXSquREfgUN4pLRw8poURfumU8LCgw3G0t9qp8L
5vZCvs1zP/TrhnSquPbrhtOcfmB+8UT3lgZlYT6MJaRjZO2LgomwGYD6oYUccCep
WRAfEvQogGMxMKRzxU0hTec3U/nVru3bwe9yy1/ikJEadMidRcKUyFuOanaicSmp
9px/SiIcQPh/ObfUn/4DB+zx6LIkqhBTfYAaK7RJ71DxDrxijtQmLvwZchdv9plD
l7VwNHix9ZIsMbbohueECF47vUxrvfeNEMolH6S75ZZOJyHd+cbvmAocOd/CVPGD
g9fQFSdJzwpcsiH2QSS5oUKc/6KsbKA8xtD5IREyaNMBSzYGFpWajsh0iVugeUW3
Wkn6mYFc1sqBVq/UqQ34HayskS/SPpNExvd3wccZ23HBVJo88LXcT6XJO8tl7qyw
fme1vIOj256uEm3TTV4yHjPqFCFyvSK8x4RHBJtmc9/XuIaKzaTbATzo/jSaWYSk
YU37APCZDbInqda85EhpiKldMO7s96DEKjol4wvuDGCDI9uBICiG5pPYF/HCDFpU
I8Zypk3VZRI+C0i4j4EL3FuI82E/c/kSGBnDbms9CyKwdU1v8mkcQxMsqiZu3+Wh
fJ/Zn32f+xbtbDsEmBVfcaZWFhMs486ChQ0DhV4JXZykf3AgaA79jBlXd2ooTCtD
aQPjnFYqQWH3shooGN55ADmDHh+jgrH81BXYw1Sec5rnwZKZxHoRRF4ZXJRSIniR
FjL3cLzfI3e7Pe7322XJjUKn9RKJ4DypkvjIsDKGGLBlBwJnKL50SQdJYc8j8f9H
AVAgk+Di/6x3Nzi3mjFikfMBjr2mlXWnYmjwNT2TGzSmCCHb4YUGLb6A+fogXbr4
W1owL5QPwv2DqW/HryCxyCePQIQcY8rh2o8mt2fe1QrUx4fbfMtQ/n96v3Fti5+5
ZPJfIYMhzeNorTtj0ssm4kOquweoOOuiOL2V/rGUYF9d4uatWFpYHxY3J6iDb9qz
vB7z7SbTa+Jgkt6wmMfaHM9wG3KFF0xNoTpy83oU4Y+yyKpqGmekT+Im8tLIWy7f
G6I5U4xtx6uoh2HXxoEY1wH2U5ZmgT1uddnwTQF1rg1LD9pG6nDtiyo8REI7IllK
kt3JNifbfKmKIiShcaThUmljjp4Yq6FA9OreDUod4J4jrJkKrjZffq1fhFXrYeuV
MQMwBoj1xwaITfc9bSlg1lfLUVNEBAiLqXOkohH8tI3dntQtFyGOzIdlh0dN/6Xp
xG8epbO2bo4/NLN7a3dMwwnHlltHn1w8tvU/24eQbuCpx1wWwwHJgFPbicKKRT/a
ap3LJMOIDvznl3bdqj/KlFuGBqxtpz9nfvgr0o0C2GycMBnP/Cit2UXb56w9fmTe
c6QqtYT18TWHFP/Xp7mJkz6MXEabo75pRFEbKqMqOVcvw62kUSA7e4FgxPq6M/qd
dDQsirxICAPleazKmDQoAL/et9f43iyqM8OGW/2S92Fbh+iHiF0A7oI/A7y+q/je
zBUgnQiSYsMt1Mueowouj7dDPuNqZ+zz0jfvcJULEQQQ4w7oY7C9fsdr7lx0s8i1
8FhHL64oHzsJnzDz2vp0P097o/4w62+2T4Z/a8IJZoOXLoJezm4LTZU8fghmcDwE
ZUiG0Gt8tSIBhMXa65PRkm5dPtGQ7cy4phcmI6hfKsdnAgn3usdvz3/Xq9D60OpA
R9EmZ/O5xYIrDLFWqpfX60Kos/OqPjSMJOe7+c9gu+arMRkb7UmdO674K2YMIrmE
cuvyGxj4030fmkcKwDIJV6PUcXfQtYgnzvahjn+++KpVe9jkgHIYYqos6+w4VDxm
//pragma protect end_data_block
//pragma protect digest_block
2H08HoSIIv8T5RfUDb3PKMiAbBc=
//pragma protect end_digest_block
//pragma protect end_protected

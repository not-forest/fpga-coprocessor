`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Jkr+GrQOMMFWd2/4wDPrLSHNZvvapYJmeGJrho+Rz4EazzLBJdEiQhCZGG0PTZKQ
sz0t4G7SHaj19HfZAbXn/rISiXvhDb0hMVl3JC+7hHIlZWZHIuj/H1H9cGfsupY+
48VciN1ypS+30Bu8Ke2IsA4wPFWftwpqaJMvms93Y+g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8672)
mHQO1EkUeHVQNjI8u77iVQ48MSruYf1quKwHQOnjD1qz6O2NyQHi9I2kxBWWMo4P
zV1QnLvfBraHbaduN1jPRNZVWElcsIzXkNLgwj1QKFeTPhHNdDMktJeeF1M0qVw7
UmngVZdY/S0Afx0E1ViP/X2AYqtSkQ/pahlDugrXLXuXWls2HPhGtBXXKXVvKBuw
7ckGGGsnZq9JmnBxUdbwCt243qujwSswAXx/7YuaTYgenLiQ9dkeg7gsB8L3cuTO
oxCCMnkI/zVCEgR82APhGPQisCTSrLli3AP8FC5oxPaYd99EM1QLtC0UDIK6T24O
bHAtZ4aHk+ZcQdjvtkPH82A3XoU9Eq1CgASpfiQRHLabJEGfZyNFSrfs+47Z9rFF
YPAMgCuV2jjTbNyDMMAsvHqvdDPpB1kKYClTGfmUx9dXZ0duem6olfgON4uKlWdp
M/n7dUfsy+uyrC6Uf/gLaS1IsxDytbS8uXqDy6rF2O7/G4SYelKIpbNpok5eUdVf
i1+9ThgyBrMvVvoHrueylDtBFFYMcGngB66n2soRY2N9o41VSyvuyhTh9UmbGnwu
JfXgXktKD7c/GwwoYa4Ft3bEQr+HNp3EkUvfS4AvKoFuGir4FGhg9erA8FWkkPAR
8vCRLL3vt+C4gSgoDkh/UrgiAGN3n2IgrftqClrg71Td8nnK8CdCcNt6mc/9BG/Q
QZsK66FpB2x3MbSad4vbzIdMvUPT/N93CN+uC0ICh+sEgjp2mU/E1pKvCXWjmfxy
9zigqTqq+yuew3J+zhDJkUwqhYYzUML0ouhiMbJzFx9k6xbmEIOG3OdvnDO0HDGh
62wZyKG+7RyqhFUEsShdr8lXYSpU/UPg+oq8m58YkjMHme+gd2u60uSGlnqcBJGV
7LqVdM4PaUd0MMxAo0/EnFu+fSbh57evYNyjHnNpBdCzapuXyhW6t94n78nM37x0
C2Ij7uZ3PGSVqJS0NKWwNwQepmzk65l5hUGUeFIxKQM/iKQX6AkIkdHZ8rdEpwyc
+SXjIVYIirQQK7HN0PjrwrQSDu3gD4qmlAkjMzeHP0GCNqfVe6S0QkaJZBcFwZL+
XxkwTKQO9/+425ZTUF9lG4p5kTduo5scXn3OHnxi5QXisU7T1yuKiCf6RqhFvE2I
Zg1cP+DGF/wr5OQAvx0gao+ybkknGXoWXihDtwHqPac/GWtC21Y/XI1wKXbdH7oI
j8e19DGwKMuzX/EPM/HWpa+jS1+n5MGNeKRKpvZp2+SqbtY20ABRqD9QJuTcHSD9
9E90pu0/IzfiGferEpiDDKhmAimRHK7yrovaQoR0cdjdGr/us1IvIT7TcoUVoo5a
e9ZEVox7tlI+1BuYXB1okBrKM6A8OonVrIoqz2DykdKBSOPkV3WkofDR24et4eLc
NgG0xST0RsCBSABb+DtQReML45Ca01pBBvDe6i3NJ3Vu7/3C2JGjGmlMB5TJPeqY
uQRPdXUFomXr1qWP37K6v+bPFpV5T1NqSC749nCmO/KERLpDpEvG869RIe1BNv52
95VTt0Rz8xYVICIadE6YUEzHGSA5ZgtKXm5YO1Cxi5kOQIbgHGmwuQSqpVJiSb4v
78lVUhX8R91ZV7rEA+9l/xa/ZyGZs/tjyugj18M1iZoAeJTT3gLrHGXC6r7kX1lE
8gOK3cNx0ZIlMWzXqZcmJ1Kfc7xIUeYTIPopHsHCJzYAVA7LvRmvq1jWqLT4ElN7
AG26B0QyQ113LbfW2aRB4+uaTOD826bPVwl/FTktz0KaaxUrMhBHzUWC2AxnL2y3
rBu2p5eLrvV5SQ1AyEo5NEvWEo9Q/VYnpxeQazblPQzFrq1WUPgT3qb252SqoRR2
aja3dvE/jZiz8dgLw0DvF4TUFRXLrsbaswZXXkEfptP0th49pn8o3BTpU2SeoBNR
GDoSWSY7XXT8w/BPYYsfoG9K0LbMuKPo1GusO5PQZIxFdemoB4y7DycyJl/uk5PV
iUMlSBniulNxAIKsa5eS/ChoeVw+Zlc8Z/gN8wfKMqZsdHatL6+RUDeXzeOy/lvC
krq8TgtVMgg+wuCVU9+jxhZlGd1OygoGTylmRxgAoy8pgKdbt9psMlW/RYSqQsPa
UbfBU2Yhgtsew+BwLUH98v+l+QfUpAi2YbXPh3Fr6+qCQeUtcghaCYvpLOyIs9oW
AAKCHESXACIH12OW4JQFi2LC8uV4Qg3R70Fj6D7zEasxkiNIdt89Zdh0cL38JxSi
vfHKRyAR5veHGCU5wjK5oyj6kjjjiCoaU3G1L7iKui4y4Y0DcXLBtGpH92JjcxS6
VRSrGq9vKoODAuyhspHiPclXbWB1PmK7JfXVSN3XHV98ZEGycP2eAYpF4ZSia1Mf
l7qR1vWjQQ0JF0oNKvBQscAN4EXXIeF/rjIgd6u1WL6ls9Vfm/qb24RS2BtvDvjA
RKLZmlI20yMk96bOROGM1gcRJJxF3E5zabyWla+LX+0Ysd012Xw+mkESa2kQJ/xz
rUsBzyn/jNyZiO/2dt/fckdp1wfJM5ivxrfdTDhUz+LQpeJhM4MQNnFjA6SnuCYY
wCR4WtykVjS5+rokQ9ICcz9znwszhLuoqtkjegWDZnd2EJV6ojFVmnhhSdGeXeiN
fU3kmPdVge4oFEoQ9l56ekfg2Qt3CIre8PASMCW+Zch4kf9nqEdWcGA9nKER25BF
TjPZpa0NcFs1J02l5uwAzZWrz5YMjAw+qL7to72sVOVgbfV2dJakdzg0ddzJJaVQ
SQQAyy/eLboxWWxBUL9ysn4xL0egywwXMtD3RikDZYfT54Ea+OfopgFRjczTx7ra
nsgZz0uLRUk3UX+wuLdo4z4Yac7dALmZg6lb3H0cpWlJG4rKidDc5fC1/9ph9hu/
Az0qsGYeby7wHEQmelpGUA+MnzJdY3hVESjJjZOVsEbsyeOm/8pdGsv8YMFvYWut
0kTfFUymW0cGMMyvTkP65k7EdFuQRRVjXBRDsqOPUCZ9gNpx8BG+wiRznuBi53lq
XG9BdsDqb8Qx66eTxpcB6iMa6D9iI9cna9rfIlvDXlHvWB+MtcMVIyzim08H8rU2
k4puukn6vw6WTw9UmQGxNb4ZDMURF3y5rgqbLJGy4MAOUvxMJtsJ6SijP7pWqVmo
EZmc8suKZT7EnEN2T8eOFaA+MrC6Q5Rma94SdnNFvH2GBUG+tPo4mAJ+9tlpudcf
Fnk2Ovqzd+ObXscOuW80DeXAMxGNv6sL5BgE42Ult/EoImiuqR3IYUpycgwYTJMb
3fZmzlIzpjUj+G1m5fAvT4zTUMhy4Gz9/M4eq31ZxiV+OElZiVPHXEqEriUz+aaR
mQ1kLWjv3AdUH8N6slsj3/UmWkjkQTu+B6neFC6GtWdaileoRaWLnh3lqZ+gU2n9
JlXchtnPh+rvIvIGrtio1MoFnujklFAUpDmkqR1pb3769GCvhmvkMR5RYfeeTc0H
82fA97Vg+Tn9g5NlftvMq6cToQ+zO2/GfbOIHCo3xInXd0H2VzIkEKY0wFFkTI9L
dSEGJ8TXajKisx1SYEF1aHhXeizpD+xFYsKDKIDfQigmCma2Bjk58EJCRwHpBqZK
x4yLYqVBg8BnOH0y7ivePU+hY2vLfDRtAlCs+Epgxdbukkf14mG3WNVISaMeutgE
BwsxQxuXtP84hBRH+Grtmxf/vfTjP/O8Pb//Lepz9hJ2Y3QjPu4fwqLqFLYFMUBr
PqR+7cYYzY8TAaxegCyIV/w3n8iHkq7QTowTsJ2UFDw9JVO+prlIXZ3wiPrQHHfc
OmM+uLi8Na11L8WKBMuhzoFZIAyo/lwsd3OQJT8b9SCVvh7L54ONwynplCZ0Id0F
BkujUToPOU/clIhQmfkN6g2TK6JpltZ8jwO6225aLHdz2PD4I04laTZjNDxJmgap
RI7HiE2TY8Q9hZYw45CI9XY2kHrHEqHJ8ZR7s37g0NSzVHCKOj2PDvIzqS4sGkte
D1I3sWJTCdK+lKIvTgihcC27FLOR8EAaCHt3S6pxqsrJ2UEQuoBSHqjNVNYlkw+z
gC0twW2ZUf1mFaXaYAETzSnS8dszzv2/X+k5gmDOe129jW8dkZET/WAiSuODLLhA
Ibe59JvEdzNmdNrx/waljXlEyr+50ZtlDby7xaAiqx5BrJ9vrRQ6+QhTlqkqhd2v
iF588lMClE+hU2uRBiX0ci7RxPG/PvcrO7Pt4OrBY083E5SqAxL+FQrIsvxfEPvz
EuA/Z/9jwzO8DIJXPN7xTanx36WROmvrXlmNUUvwTWAocxuYGu0fqcSqCUzDiwGm
zBhbSazXflIOXeINumk1JLsyQfY7ZZZGscuoCBbNC3SoxKVpJ5uh5zAv1SikBqO0
BH25RglrhZXoA1JSyJh8zdhnTn7MjAKG2rC1b+rG1N7bCd/LW9lT6VWOb3Y9SKvz
C6i9j/CFNyr582mq+kLZDpyl3b1pnPEpHe8Z/kUiV6VUwL53YIUhp2xwaoaHKYPg
e+2CoBvtDzGdKPLSHGUWn/SsemZkzdZGyuxiEWy6T0eCjckMvGkc5ZEstgsMZTXq
1FEuBLNMQmnH8eF9MkQhG/JBg8gG0nR7ofpz8XdrCuCr9ZGFdmv5GCLUJ6FsFFYo
tFQBQ3Tzf2kbAaw2OfNuBEs9ZrqWvVwGzN6HpkWe9eh8xRjxAxdPp8lfmUil1/u8
SE5M/gRrRi2Js68fXSRw9nhh/3YJusAfEYdrbRmmM1AIXac1OS+UXl27h4t8GZp2
Co0gMjbOAZP164wmzbNZ7u+dqE4nmnZkhFle3o2pByqVmMWk6de8rLH1/job0/Qz
dP9vEIU5AERxO2iyPTSvrwAE4W1Xuu9VtavyMbe4SEXGPv7IuBQoaxRshOKvlAsT
tR2TSeGGkZ+1kye5XU5YXh9wzNdPqDDCZloSJnN0MQHBPIZ7FNpj817G+SxiamwL
J2676PZnTAIischGQBX6aO1DvZReazDZWJosbaHAybMZA6zZbpRw5MI5TFKV4foa
IMxmxRfEOLBYpTe1OKsvEAb2ArmQqH9hziynSt53O5zGB4uFPbYHtU7oPap1bal/
63Gh49kcjSgOGYTyym8MITOcgIUhnojDtDTHxpSI9wMIiyDokIL9kQ4zZ0l13EHf
5eyKKGuD68a6VRNh+SoB+6q3FHX796u9zZky1uGMlU5FVdfdnqjaQT1RxHMZlBHP
zxmPLQth9wa8ejAFHdC6QzqzKvwGYuvg6L/a2ipRoX7ej7vwXNEVBmPl2wYk2Ebg
KEFjsfOetCW79BUe6aMJkyqLzt1xknaH8qlrZvXm0QgH2AntJ3DgU7srrrS3ZH63
ygGOj0agKhOl5pKOR4sgX7RTzWV35WgeJfFkLQH/cDZQGzQOwuRegy/qboiR3Lcp
GyjylJX2XRDlaIM1gclgsEczZFwcHwM7qpquUduHMUdX5bwGyyT1/gczw7AavzqZ
lmQTWMHE7TRn4XdYG73XoM5lm0vtmtdkZbRwkPJVO8ip6eVEu9UQkM/oNMj+3FMP
tj+x9CGOCGJFIRNhjaUMxzn9a0wXAIdeZ9xnv1Zvk3YMpFdLWbOnadcTgOnwf19s
ivwXiBsZ3VaKV2/d7EgnHE91FVMMyuDJWVYLJPtEsbV4cm+gL4q6iMKyvPhh7p51
8d8BZS2JwcTwtcgce8jjGerBAjFmU5jHx1vWAHECCbdiqUbZa/glTsCymXMwBKiZ
DV9gD6RegM5c6zqSmnDPfONzpP00wAxoR5JVLrnhLIGY6hayi92WAtqgNyKxarGk
G5j6g8kdd9Hk+65JdzQ1UE4bw4Lk4oEVbyY0VofeRd1wkgqMyZIdzbeZfVwnqE7I
Is8WJJXJ/LSYwbhCpzUo0EuDgFRyOjt+VK/H43H9L6cK9kG7T26N206YhcqSu/5b
dHAaY99VA1uVh7ltZYRoaRCJfEnFNFDwV1aCSY6uqRQmz19Fphay9mnDZFXzxJuc
kFjXJ3B8geNjohbYVJK6KVGIKsfmkEofGGpcYzJKUBEH1He6om5ZdHu6jlKmJdqc
0z706zRzqaTUuRV4oIWZa84ejdSLupa9UUeDM9NNnb6qUl9yJ/rOgd6Chjme2jc1
+6S0t1KIvSyv8NHfVjQ1fQYz7j/QqwD9lLm/ckssTQu74L78BtqL8Y/b7jmzIP7I
2/vz7sl+IEN7W93zxEhasK+BnMexb/z/KagbcM1HT1TsSurqcFNCfv/Ey8DvpToP
DqjzM/yhcS5gzuOVrmFvY2xb766Fy/jbAO6edt8hE7eOPNsda+ExMYG8TD9FmzwK
Kr+DWlAiXbaVhzMm8Ob5LX2jDL7/sjm7DlWY04nhuKNMpCp1m0Zl9yqnU6qPPVuo
xLvke1aP/U6IYcd5HJdRMGaxcs2dtRT+7A9i08Z8mk/FbptWf5ZLIqTqtoptlOsD
kwnTNueOAQHE/lRYJix54lOqbGnJMq3wbZwci7RBp5kn4cZ+s4P0FWHUOsfHLoA6
lt1uPt2YF/hPloBw2glfy5o47OE5kfVIZ+VDry5YE99hALSo115TUOQ7gC6UyavM
tSewlPuODfr3da69a5XQynNx53rTB5dm0gB+zoYRayWww+NpQ6Umnb9G4OBJP+xf
bW9maYt/WiskrsxXr+vRj9i4TQHoTc/ahvDxMitfphqxgQSv/B9wMUdWXxQvuBMU
7OkpqRjjc5JoRym+7QZiXbZTdgwoRcaOdYxroS07Fc3xo8g7bNsptBNO874KwWiZ
B7MejZZmrz43aqaj2XOVBWKT0Ayb/RghUNyejwrnAnNcQEOS66IzZHMSmTRsoRRx
vnoOaNcb6K8b41D0WrWqOam0QbMwVpOZAvMGqWqKCpyPbtlS3ZuK+eC+aHtD7qIR
BbFEI8mVirwynp74YAB5+WNAoUe6xfsbt8gZ/im2TWdwCsMmRcBpWWhYkkkn4sV1
Rt+qiFaFc64z7KXdlFnGwbhoBqidb5+9fuY8xl/a6iUSFBT4s5eBT5bKYs27UMnW
Oz7sCsfqyEsDThj9pFq+779jLYahAh7c1YyHQbUkoVb0cb5BiPeR2Kx63nj4ZAY1
gt07iaZ9uXgPjKyFsfMutjbwO3PevbDZQR3WEXM7VhvyDCQ6gkDYQ5hlP3gFah/f
cUgeqiE4OsSlVyr1VpsQe7FuQ3vQL+w5uiWnhpTrQSgGu9rVqyinakZMNDjEWWMp
0wCfwWMgai/Gw91ZFRCIltPuNtFZt+AJJPjy09HqkUMDfTJf/3wuDkR8jirJt4wQ
OsOC93n3GiD1aBuxxvHL9WQz/MaBnb8okaz5BC1hJ65nXZ7+fC8/u8+oyPg/ulbH
zrctoMEMuw3Frnu1zQVjv2LL0KEIx0DvmY37Oru/XrpJxsRfH+X7p48n08LZrEmU
WL4oiDduM9b4hxEUc3EEDlc5Zj9+tcOck8ptTvkdoBR9cOgomkInpNkjAZTyZkAf
ez8x2SMk5a8VdhcCxG4rVYa3pUpfLAGN3Ko+trCY4Xeq1yA5j0ZBEV2jCWmxrGuc
mxt/MAx5ofqb7/fACkvM4D6e7ON535V5gxmLd/gt+6FB7DYR3tLbcaHxwxwV7KTj
NddgKjG/4CDFDiVmwXhpzJy75OhSadrqvOQ0sKiTdAzDAjDGUfLSJBlueOemSLVH
Wab+qdJm7D6RVTEo77/LrRbqQoFXqsFeCy6n7+HtuSaWXjmlO9Ym6b8yHK+xkOQ1
JUr6TWJBFZcU0GySK2L0SFMQUd8h2s6jTmerEejRUnSyVfwegsGksc1E7M0rZw7/
/V+lYzbBC4Jcf6j0Gcy0q/iFEX0/dZbdynmWI76ENQU1qpw5NQdeA9mXasp4pbYX
j+MtqvdwavtKuQIZ9Qh6M0uHS50JtlpE1JTsHYZndqgHkgvc4hDXcnmfIKEOsMTc
6NaTwBBU7KxrRBL9do80TbXkUZr0XXNwndrvsrpYCY60fy3jznThSp6ii2bUEKjA
Hk8axhhASocrwLQLR1cGFtGnPDo39rFwJkUTsIafJ8pFHqExXmovk1Dn+Ny8e5Yz
vR/4gkXaQ7FzwUTT0X68Fm8fer9jzrivDX90V/bGVbbe0uCBu1Ks3gqf7NNp0xjR
L5k/4bVfPo42GHoj79Ec38c0fvqogJh063lQs0Ddmq+EyTUZX0sS5PHnLt2CREQb
MmYpVn1572He4zIMAFwImkoxs95PO+kKbrtqwnUxnR6VXAOnvtxkOP/1oUu94dgm
mjEggHS4l+HE1lPJQZoEdJgqp0KbjINqIqHNiDzrigykV3zIfknt5t2CCvJse+SW
KxGlhkGe1P8f9vI/n5WgmVUSDt2+TwjtnGC8PvlEicHh26jgdRy+BMZ5DLQWl/Dh
IHX6TpF05JXLPGGZKZNkgKrqyyk2yxbIcXmZtPpI0KDFvZeDZq8QqQyNkvXWUSho
xjx5GddSFzDuwU56aJNRgpjkmlPkcpm0JAmQM15tLBdr94YjSXJYL/ehCgYpcylC
ds4jHKWix94YEmYb0YGTTV9zWLk5GhDUVEXqKN81N5xfnXkswizadJ3BO2P+EvT+
P/PEnRCoE4USCJQLjrigebU1ZJyTd1lxx1a61U/RjFPxooKK1O8ZGRk9V7jykoyk
UVKm4SKGvBzPtpt79xpQkjK+c/e3s5LwuwSPPtX3C5rgZzeUhFvYbxT5GN56+V/X
aVt+VR7tuzgpv2zNzXuBCOVgx4GzXfx0i3l4LHo6IPuq4uS8qxlU6OjiiNRZoZES
wSQr2wDADBBShBEupaXh4O70FOktbPyD2OVfxiTC2xCrv9duQB1sdhp3bU6GcKSa
Fa5ITH0mNXBpj8GHeOISiwP9PJbZT7U1urRVsiEU9SRdvt3P9ssR24iHVdF21OG7
hqdnCFMoPHsJQmESfNY/l/+xHWtPQv1pBPr9PuDcdn2UVChknYFVFLjDl4euqTji
Hu0ApB2lZVrlupIZ9+/a177PuiB89BZpXXode9wM5O3y/JN9LkqJL28GX6BMgNMS
kGPBIcODQzpdILvcvkt4CQZOwAIDT3QZDYCdNxjnLP2TJoeLNYhgrljoQUOMsHeo
0py+XDWv6AhahMU6crB9vxPCNIXs4b2ixN+SOU8aOvdkTJHxckCw6gdmpdUakidq
ASZdtAaUPxfts/MmT24RRDrpSFoLHaOEYgZD3VKVu6G5w3RLG/bKLIfFvA2yqHYG
/+7h1i7+/vaI3Y7694whW3ONNdNc+7J7FjoUC6Td1ffISscH3gyR5d15b4yi5mHm
lT8WGzXi9waar8xdhstV2volgZMHcFZ53A5BjkJcUzxe91aSXYBFIZsX59+tBOPu
QEefAYG4lHUUe5SuPQSG6WfcthmzWmKyPxZsLba41fBffhcmKZqi4xehfQOqdSuT
Gt7q1Y9V6zFBGl+DRZxogN09c626DUPgd8U/6hsXbDW803gg90WYB5SeV/6EIb9z
cef2Egvt4TH7LIxGdR83ysvgGSazEXjgYhxC93Noev4n9g0MSqZY1pOQduJ5G5fC
ej9VcKlR0cNitoybGGvX8L75HBL0J0DzZp3+pqfumYCV7I6B3PFoUYfICrqef+jt
IDKW7xm1Su+0rTv4PoaNaDrUigSquhjAMd5YtszBl+guzi0BBCtWJ8i1TOw49iww
tUQ+fVo2bZW7PxcUoxFCawIVaXaszYQvA0bh3K0TBmLYHLKMXHMLlmqGzgs1ZIzN
2pIkaO6k6LGsLWyyaGVLHoj3lniUiZ6woEPkU4kSd5gQNC0/bvJ6oRV8EaN6+F3w
xSy2GAePuX5wjtm0wWJF2NqUHM2YqyeGPgfNitT4Sj1lp6AUk2c4ncYLfNYPvoNz
L0kW6D8WI7Qb5CZTkaV0b4y2u5q1M7PjHtF4QTpYpV6JCuA7tQzgbLieiVulIbSR
KdiKlqjPvbM78k4v+IZ/Gcvvou337Jed8jwyoifvtp3HTWPvdd6dF9VT4UynEUba
WdAyBThv5dS30Ok3RewdXykbgcn6jFAgMmrs41IrWylNKKq7e28XEpU/U1wIqUmi
p8ApuGgZjG2Y3QAtAlGKIjeF34oItyH6khP43ExQCZpPDMcTPNQh6+WDTymgJklA
/K5X6JlqKx9bLJV5wFHQpx9Xai6I3vrjNTNGK8EnmDN14Eu8s2S3paQZpw68yHhl
l08hE+JxjUp51UbEcvNM3LLHmJ+MfrYEU+ty1RXW/nVlN0PjdN4ZW2204486GbIN
wrSzaXO4pay7BtfwxmIMGT27jGTQ0L305QEQwtsk99cTE8XPNSg1XYN2ZJ6d4EXY
p57vNMBATzvEGNTDopOZxoPkiCkkcUTWZAUaL/7jToTJ3DN5Ph80XpWr1VmATJix
/s265OdiNYnyi6D4mTtkvGvMyK3ZCb2fL1SpmwyhwvvyMEbZCXz6KIWA6O7gblKq
/FFLByT6WggbaKO+NngfVP76m70hDBmXsUV+W7IlgZtqbQGq4JdfGFhzNC4lHGTf
YRF0iZpRGi6efyY2Vy9YSTu/S3vv4smtFB2MyLuPb3LPGT5IjSyF+wQhTCOSDiKi
Xxj9P4orwNuQGoc+BcLrPHk1AgUN4v1+dva4alAp1UyoxsOusK2Nq/rkdBb4F3vZ
lciIJMIH21X/gmk0oGYO2sgXPuqLbZ/c/MnH+W4LyDCgvfdLLfIzKf9tYp8bNjRd
Dn/rSwFOAI24N4RDo9GCYTONH66gbLx8Zs6hKHCfLLF7YDtayEvvnvtaEgT5QYUh
/YW2MNH7PL0B4XxxTk+XLqTsSagnpPUJM2L3SsJMgKx+T/xYjx+Fis0CzTV1y2ly
C8Jy66tF/8vXaJP6K7J5SI8Ultwj/ETx8k+UxW3d48wxRkL9Y+CzdLkQComZuvC0
9McP/4E/MFPw6OGm4tcA9xklqsnGcDLfQPrfsvoTXURlVQf9bEPNhZsIMd3US86X
IlzjxzuC6zC69bCHMJSg6b0TE+cHOrAZi6J8mCp/ebRtnM2l31PMLwbz3sg1xrMx
wO6fB2N0DZimeDtJoKDqdf2GXOeM6vSUoUf5vBIsPiaDXymueiX+Rz0z00ZuO/o/
VhOc3BLX4Yqeg8k743LIz2UVCY1u+SrqvEwHOcH1whcIvf9+Z5/sSZ8yHNQ2mUYC
kWAiDfa2NS+GwhOpv+RMJIlk9JyIdGp3NahnuhhhIfSbFWWvG0BN0Ms30gvONrlH
9WwXqiE7AkmmQBTblj5IY2H+MGPcYH54MclXgCUg+Wm0TrmRsl6jApGMUFd0inMK
zsRTuBnQHH1ek2imGkFRGqj2W5HZoyLsRJOcsBQX2RjDZrbDJCMvoF21xRqrWsZX
Pp4v+wrUpxo6Mqs68RSiXiEq3C1/cnSPup1t1oDytXNgYneAIKxWFHJTJ0DRFCrT
Uonol6gDWL/UOOFUZnTVxZaUC93VW4dFkv6pQN0t4uwTmsdS0+9ycJeLfjF4EyJT
zQxW7zymEmILoD3aa4UImg3QpqqixdDik7WEL8ENIiR+JO2/xkx+urBrSlf5U5uu
cePVWbtDWXXLPddEvZ6uxfb/WytCSmW5z42JRfUYIMt/SK9KuXxyBByUFevnW3+X
f7Aekdmz47A6kskgjgB2n8LbOMzOlxzw9JPl0f6WALs=
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
o90oDl7zVM+M7iZcVt5EaeQsV0IWEI4N2QdM63dvwDzixxK7DL9eI7Lh0TQn38wz
15ttUqfLmqk2UuWkwp0kGdhfPHnLNwu0tJha+OWdW9q5wwN3+SyfHzdO6zs6+jkp
Q8jidfxXScjLWF7ZZjQ/yCtxxddc7+jBEx0ZvptXTpFt/QH3htUVprxN7ac94J7I
NJVSczag3n9Lei/JUp0uuVeNwIp/Hf6fk8AuwtfzW7aNbJbGIeLSB1Y+fEix3GT4
9dpDNP7UmyOWvu7yhKCWWUb0w+Xmf2sl4N1iwuselXauPFDUYY8z2KJrDdvznho2
WyMuCY5BW/+ZHb8vvKIeag==
//pragma protect end_key_block
//pragma protect digest_block
8p5rILoGPjrcpqQ+9E1XSER9sKI=
//pragma protect end_digest_block
//pragma protect data_block
+fsLCugdEEQfIJyfXalaSXIgabC7jLsxymvvdEoRony3Bq/cAOSrdiT2S54v/yIL
X3X0wdoklOxW7IcxXDjUxRYpP6FTZTLJT/vev3ZB33XqO8mQV/QppJI8TuGRoPkB
816azeOCX0uDRMppgYpmVxBMoxzVriY5pZ02E3U2fj0k/gvscSusERTqwNtYjs0B
MMiqvZcxqbnmpKHwtM/Q0W41GtHOfa96BeLy92qJlGWg0ZKAsysVcyWQMxU45HG8
9mHIj3GHIdFKqPlSAWMqK185bvoCsr2FE3ki6tNnVUvaLI6Yl0e4kx7KLvwmEXUr
e08csCn7z0lfwPRuGMLAgUnrbPG1nm652Q5cpyNRHq3lObIVd+L/3TryEcg3xaMW
zkgDF8pEf4R1psRoyJVSZDF7Tz0Upc0iJ38pCQuWGJ+jQgcmzp1Y1QV/2TJ4OX6w
8sbm6DEKw3Bg6QSDNPhg2IB48CWcwWltwC6IeY3D0o3N1nh/oCK225fI+Z2t0XHN
uYuefxiV94DvQJLJd+baaUjCnF7tiuJaX6QTWHzOkBN1lTvm+6AefV/Jez5R3b2A
8LbNVOEJ+lSvURitWXusDXkY+LReqYj1Krup99sxZYwiPY4tIomi9u5rQm7Wykmc
+AJ1Wa1ioUU+V9J3pQ18nsvfe7YGsRJrlPSjDpqp2J8hZRnw94Uu2ZwKBYNCMjE0
vF4YP9mv64Uve0TMCi2+Mtge7yVbgS2jvFJRyZ7KsyEsEBN3zfMBwKdUKLarIOhm
UE7HmUSTqI1ZfwvC+g4zkgqlKQzh4Nvqcxe29/kOM33K+cbTaelEQA4/uWfsoPor
GNNPvTg2lsKxFlmtgb5uzhjXe5ezjvXf1hvgtmmop+uqi0NgaJGQqK1Ga5llSXTm
/9sUMHQrb+kbgJqmsVXcuiI1Vt4xcMpBB1qTz52ggHvKt06f2hMpt8vnZrA6VvEs
HW2S/E/dZYdtmIE+Sj+XEms2qvK50I1O7znw3wwx79DPcSD8RH5yj7HkjedPRk9F
h5XuKmx+5srpqz7UQnPTodAX8nkEub0ZVTFe6QI9+2PVxQUW3GqUysvlZxcjY4xR
gNF0Ti///srmC9CzVzYxVD6QCGKg7yp9ovEIMttNrdKViSVsuDpxtItbpFLLGT49
Rphgkg+TDTlbHI1H+fbFRVRwUEfTomUnPOu0TowH0nor30RU4TeFqvSyKIic83xG
Khm2w6hrw4Hq3107EpQK7WxRn3dRKshoRe2xZiyUWzrpd1n5j/AzuN3FTtFnuiL9
ODPJQ354KaW5JsJxqcUkoK0wxvsv/kMMiOKdt2N0UhVWsWorqpN71IFO2nldkv9r
ZtgDGHsmM8GEhsgzTMy0ZfzqXWV6LthVHUP++PGj6HQN21ApadjL6fqmlUflbXW0
H7vGiugLxBXGH0+AlUcyloNf3PRIbjM/zpFojACEjADvvacgYXmEowjbvLDUShrE
gztdCQcLd4dCMO++rCrHUGeqaAVsTDs4jU6jtWb07NbTMyihhCcXlvXc91sTwZ+h
1IQ4O/MoR4RAmEzDjVcma5JbHCrTNRp3+uy/RGY5DwjEdXYyPZHZxNQfTLmD4IGd
kmKEeLxrVFeBfEaYqnFo23gBGiCYHrluVQYJfG9VxBtx92ghcEnhEhvYG53aeyqh
WRXqfbDjzjOezSxbZPZGo+MdCsQvqUd+kPIVWu6Rc3YhnVwqV2nnaMh133Qoyqf6
BAYm5oGXDN8k2OGFbzlzob5Qdn/a5kCBqqhZJ7F/fU+0Ai0rnC3uGG/A0aovbeIK
XhHXlzdeu27TyC7cmRNOiuGJ3yRf7PJccwbpG0ZDzQ3CIYccanzSYV318L/ntFl2
SA14MMniBqrCfSgzkAaPGVPMkJTEVEYyYOp1rd3cOHf+xxf9mJF1ZP9m6eDBHV1p
jesrYWD+8sIVLI3ppMfsgCPsiE+UIRGdwsmL4nzFb9r1pEUtfuccgE7f6NammOr+
fKxHLBRbh/Wh6oNc/xHWGJBI7qpUnEQc/Fm86hSWm14HCf5b6Q8HH5Vn+Jcd4fHE
e3p9HYMId9JPvK2eu2d4d91JT4de3cZni45hV4nEpv2s/j1fUluMsQr8GQwdlwrw
cdr+PUUqLCAGmC/ZOAi0e42ssr88vmM6oNXJ8SsddcK41V48WDgPwksj78KfrfEN
vUNtrgM/yQyzNwYxX+k7MUpNo4LcXZlqi4bSjX7/P+ztSKJPKDpy6zGAWgcNL3ML
jXjfbRw8BAcbCgbBDTa1R0oiwLZwHqhlWmHQBXPP69sz73ie2qCSB1mxNgZ+QcO5
O15gFwCunRHzF/qST9Xl0bMAZMC67rgqXdxQ+OIGaPF2fSOfXKvp/WjrQ+DeJiXW
oIe8xJiyadmfsSQsxtw05QP3RQQ+PB4Cyenbt5yshx8KY33TEALcmfmab03wcFM4
QZQU8o5jCwe5yjcPdPmVwAerKh27pliMF/OS0FAT9D2GM/8IUC8HqrUN2QQ+Fh58
mhcvkLIWBV4KpoHrZ/Ard+zmR/r+h1b439iYdi07I/6cZ3c07YN1BKs8QmwKeKxW
Ftt8valw9OmeM1DhTyos8aeyMu4Melcj/PhybkQmo+Es+ijgnjawx9kh+QQfu742
I9eJZ73uziiQc7CvU0qm+2CPJkipB51wLgIfaBUspDGy58FFDK6lhBcGWiBJKgsM
gHeFmi7KR8HZeaabP6sNVMYYKByuz3fOnndDvbVGborPT6zPhqZRFtsbpFPq2AVU
CW2q49dhi5Kij1arlh34rMfteb9qpU6mETkOqCnFajzt8n0KgyHlg6OVNkxCo80K
UXXMWLb9BiRMIIPV2ebtSIjUU4szp29MAk9Jsn95sU7/b/FvYHEDM6wiKaIEtJ6T
mpuwpKLDw7wfIKD5fpZYb80uj41iMD5fdUTPQ4pcIA+GRzhgVfwp4bUSOZIyLHTy
KEVDdwcD9R014xiVT8q4+r3/4LPkg3qAvALfXtln4Cm3hmUmPi+NmedjnYxTmB0z
P5c6iUBD4bD+AVVPmvCNlI5r1UPOgZ0HcROwuPVU33uKWzD7LzdEqba3NwYWhtoh
GQKOOoxG2PpErBYw89PloR+s0lJEOU3iP85EjdDXQSO1xpLpfJ64iivWDGt2h7ys
TzSO2Syu69zSRnJGEZq3ohOJreLTvoGKBkkN7h4dcGAQ+a9OFImJP2zSlGp3XgML
3ijNXUaIsdxiZAqsZWx1216B3by/WbI7GOuPvu1IdUEjmD5yBpuPdkGvnYHclG/L
4HohEwNZkAfEfVFrCY8sHC7vocyP2OgChSM25YPil/k6kOHqL9efMgay2XY3OKzF
OH8rETwq73K9DESGgKa8XcI8qvSijeCzSFh9d9TQYq+DmdJZrWqoU8nDs13Q5Aoa
1ScnQ+p54zBLpc80gR6CRprO6fULYaHa8vg4v1dhQlw1pRwYSBHwDfgGNWi09K/t
ZFVtOQ+o3d2bZpXd3EivvspNi927xVE82GaH2o9vXmsX6ZqkG0JWZ9ssACHEAPlv
Uesvz7QcaMPRqbRckkO+P8VjV1035OSKEx42ZLbAyH3JDZZl16vJnvOXrOPlpFym
aJL1nm6A39/NSYFdLGtqYFuF8duCG4TeneB0rSZ9Bx5VM0i6TKVmv3CYt9bDOSDH
whIy8u6NmKVOKo0qe1vOoWiWgF6C2dzCkhalmuoe8dPKfqFSUh89CnOEUV6RAXkK
JkvWkR8Qq7Z0Qz6SaBwA1ut2sp+lplHTcouke2daCxu1eX/cSpjv+ui3goWKvUxd
o3J+mmUHDZuCbiNtmZ0mlj3I397Oazv5NkKLLF1O1pVaAtn9t0aKs1Rf8KLBtosf
tUzLIMZrazRvRwOulGrwGIoeSgI05dqAVtwrPo9sOQ6OhPvTwwYlMRmNOrArVwdF
fpiN3E3gn6LSFL9IXv5pdfztsYQ/lbwH1J9svvQbTh5fFf/9Ffvi1vi7H8RKq2vn
S94fik4wlJpePceiwHmOIbbMZrstd3jIu1IiHVAHoCTuH9/bTZQl2BLw1Z4bLI0g
55s+AcHKuqylYpphKt5eN/VdAbduvb8ZMnqzaTAM3I6JDuvnBtQhPSnLk5lrlyk/
HOuvA3uk9oNxfwpCggKg6VhLeu2SN5RIgb3mVUCUd3H0kMNvlc/iZv3h2YSY0AzN
Rn+G+btftqaCbUGHTfnm7SHx8ANcFWWLOlpuPRaRgVYhXqAQwLU9WpSslZ1OGgtE
yKXQiP4YD2xsBBVwO1Zi9tADExc9iokx2nXdJrOM8AIapAlTBtCcCSkfOVOYkDyW
VJBfnWwl3UT9240zv7if0rYezPznIxV+4+U0akseivpfhm5/sLvV2ENHKUWTYBiZ
j1XYJn1//AnT/H4eF7of8I/cRl+578PHqeiBdqiw2bHVYumewp7vnsvXxSSIER1q
cYckiQtoeMbYKfQVxw0KJk6sKtuHJNxe1r622wu2CoQYHpadkm02TTg6g7qKzPRS
KPN43O7zbTtDjjbA1otp6bXZuvEHIyqopwUjoNRehqs3LIesfrrVMgJ8ghsQH6cz
pE6Qh05r9+kLgF5dEn6gzYaRnC/H8limR6Ihb++aMioGBm/Dj/7Z73QEPkqgFAQ8
vCp2PwwKji2NeB+UeLP7e2cT5YX+dMebfcAuVzyK3f3+nC/4O/oneY7+xHyCQf4T
okTxJE517cYqDKsfChNt8iTlhOqh/YKeuqI0avNUY6h9SmlGVwg0SSkVgQ7b1BkC
lyRT6y0KIn1QzdOS3s2s/1j6sWOgbPpbivIcQrIKzfo9iZ0DRGa+VD7ocjiVhtnT
DE4NjiPjn3INCzK5fBVsNfhqBUJ74m9whIFYeW4819Dl9w1hgS5PUnuiywQLaTaz
ISniy3liGYEFX1OqxO41IduhowIY5EI+1MhytAzUgtBIkGrUbNT8bPNqt5xqzwpF
MFSVuyPOOx0Lnf0AcxS7BRm5Ipsx7YnYEInXEXgqHdKh1nE+eXvBTLNDSUn73hfF
TD8G+ju7X+ZQzY5BLviE86uIFFg/NWD+ALmUWpbkdl85I9K7q+6FVx+HCFVcvLQD
3Y7zLt9gz1pgxPc/j0fZ6ZFWs2mJI9x2oIfyR71NvhTZCd1YrEi0A87TDRyXYkJT
uoPyIJCF4lk6MbXb1SK1P7e1OOYM6gzXxw+1C7jjRdKsbqxawz1EPoM0CX2bWg7W
pGCFXW246goEaGv/AkqcDflKYA4IpFlTK63SLgMMguKNwgNciEbj8ngA3em58rhq
R17yG0fqbrI0xXM1zU/8wlApoUodYj0HFjx808jvwSQU7UjE+jaJpBNlT2wadDlK
jY4Ul6vmFvXuXV+NQj0ag++pT/mBaXSwyeWMilKNXLh6D4dt0FZClD4xuGG6NTL/
4S2nO6mJI6MLGyDg3TSjyAt//mdB/I8eLa3sF5KZXA50I3exoByJE42/htdnCv12
CkXb68MEPZkjD5d4X3pJLK+YO7dr69vX/ETNmOhP/qtE+coV+c0h4rfUbxYl4Jd9
vzL2AC2js/d3jJlZD//u4A61Qs4x+Hhyi9Q0hE81wfFIDiKNWFw+BMMC1ayrtnsE
sJ0pDPsIB+o+2tOHujrKKLqHqbJH8q4Tekq7ZaTcC+E0AFGMID9zOPr9Mq/p3S84
hoBZDJfzhA//U2xDk908Fz9FhUbsC1Zmi+Q9ambwjojFLoSjSmTr/6QVoirKoax4
8dzx6HcodlJDjKCB6VW7ozdUIs9AbBp8drTiyqiaZsy61Lv1l6R2mwdVvfBtTWOB
sxuxRuvj8PUgo8cs39VZYDXYvE5dDwTW+NGNC9AixXQi84VIuSzUTPmp9UJUIOrY
pWAKA4YlFHe1cbw6INGIoootOUeNXwQVY3f6CRub53uHX46JV97FzgWp6WWPeU/c
MHfWLS6C386TQ0XNG5w1Pe3XPptSbyQ+UxX3/3HMim2yhiE8WVij9vWCW11E5ghA
WIBcdgaAa+xVoieXYignbhOyAYvtvcZYpnWskJSaJr/CADljniEFyGiyZmc6WEwP
vUfMl3fq8O96nG+Tx6NP6hUj1iM3kWWg79PTpcWSmh4WOfF7G0x4/06ZAZkCF/JD
xG9e2DSyQt3USJCAmdJgrmtG6EBYy9U1gQW0dMDFXQDXY2osDAMb09+sROD+tvTS
24r2O/OQnWQqeZPyXSavhGmycSP7NmPdTNWFTA8bhLrLQAdC1lw+bnnU6A3Shx7A
8+Tsr5nZW4nFBGXj72Is27zTw2zcWigMHEbANfc8SJ1CJHCKwQHsbcLJpOwh/yIH
Q4dV20UeMNZfPmSc9ET++1JErfnNNLrK4jHYHPyvWwRRYz4tvAOg4oMpJYlm0tVY
Or/mMUwLVZ6MTNx5IK3ysTCXzUbQH9XT83PfoGgopPHXbuTKp8qXNROlcMMq5mKb
0ME5xjtFrzEnlnp0NPVGGZoR+6bW89YeOTI5FGkhbCzGzjMe0a6NSrDZCd5Oc3d3
wwhjy5n+pMqOVYU1ORzB2dyfnCRT5sd3f8DlgD8FgtTDgeUNzYV6Agq6rWT34Emr
7g0uAtsEoo3dv4CmDLkXdlpm9cF3suNRCa6SvzbWgiticmiEjHgX2/TmNyk7GfTp
BhbB842TSFzh6Zm/Zrw1keEhuKgcUzhyzzmE6b6Dugy7Hq7IDTbzVPEbZTitg2/E
SqdRsVheqmhIrt2SYT844MpG0GduZwqz2368lHDd0J5OSQyu4FOmWQp0tyc/uvEh
5MZ7PUyRXM9fORgbYTk1upr4y3F8FcUQgoLSxbA8yNqlImArNtzeeJJdtKfQnAf1
8zwYJd90fyCQhKXYNk3XGR85WyYjZLZBB/FRJxMsEjBFNxQHQVykrVro1T78YpQZ
m1Ulwp2W3+UvkZ6e/D3hkvGdkMwvd0/jsINS28Nh66c3s+EHQHNiZs3TmieKfeX3
MFbmup4v9zyimCIpqoi+fDf0B0QfSLjkOSit7NG8wVTRlNcw+5FJv+Dqu3+akDmy
fwk0Ygtuzct90TKxA/b5ty1BLLWNJZMR3uku6J3f93L7g7X4BHz463EeUqKmAUhw
w2/zOSMygefC8LH8p24tAbVb4KhVsXLVYB5o8nWWAJXA+Fz75hrc9TWIdkD+SbvP
BfrNe80d8QMTzNsKqa/mOEMzsgAFjO6KdJkc3tRdFjZSDjCCSeQThZIKWzcqsIP5
qtz3X9wsryWKbMHuUJooGGoBeHDs5c7/l82T3lKe7i0Oq/eqU2153o28/xzRgqW3
YXkovqnLcGlpzIWeulKKNfwtt0W4nstqdwTOMHfosouhzICtpvlH0aaYQ66Fjy4/
mo+8kLkHvzBmTJqXqxVOdAjcrGMo0q07Z233Hutmw6i7ruvMo23xzdik193ZQ4BR
59rNS77Cv0XFihEk1zozlQZbaYdygL78lrI3Q03YaNTvN9GnmSoFen8/extzDc8O
UipejvvVlzqPpOVz35Y0rugwSN4dG45NAApHLe9PYGqY8Eoahmi69D8DroE/W/c9
c2mGi+xL00OodxKMe/jwqDGey3VztJeDo+s+ZEytISol6mTYDR6JcFCcpSzoWnv3
T4Sb8wwPSbk68IdAWYXp3/qWaYJeq3sx4cx1p4yoqyP1dwHr48YHRL3f8MygO69o
JD07RTuCa+PVzNxIKM1Dk7Qxx40RnjP8LhlixVQix1+CB8Lct8xXcQBSsGhnKS35
dtyIVXePSWwovs0mlXe9/of+vYsGNOhmAYHgtNNeJfdKLNC6irnmqhIX9pmTZndR
QhHxdgSUVc+HvzwQM9Yv6TFwIkJUtG83svf2Lm5As/t6nyPgSGYXNSM3DvoShjsE
uu/x+txPIU8S+hnsCDPaevWdTYlZ0R+zfb/2F9dwq6mvN67bBvtLiBDjNbGDMGsd
1fxVt1RV8AW7oxRE1qaKGCXb76Op4G0cPVIWxgpdgr9grPxtAvIl8tST/fL9DAId
7QmYKgBUHD0gyB1jyLIeCKbOYxh8WVmfVjRbgWfny9ThryWwOIiY32IJkwAlpCst
Zt4TYEX+GrFL/sASDr5nxs9U4FofSTe6X/k9FLn8nhIJqfhGj3Q3WH9X1QYUjw7F
sv1nnJrHsnuV2ItKSimkvoU9nq9pwX23VJIP+HlFUmCmOZyfjN9WE6uFTK097q6o
+e3GnE9uptTfU1IlH4oPNmIiADUEzOVaTz6/vxZDFobllWPaB4dLbkv7caLLf0Et
9yWK4qOCZyof6w9NQkNMivM7dm0LEzpDBUuvw9UyyVv3yCJwQ84tdn8XyFz7ZIB2
rf8qjuNDSTZcLf3eAroXqPQ0LABAMniU8+ZJhblrCRMlhxEoqKEWzDjdbpiA7Q7f
AUQBJhWsaQ5BHyTeK1r6oyGC3BBfLm1NoU5Q/5nJ/NkQm3Fu90VzZ+8X90ApW7kz
U/6w0UEBEHf8kGvgZ/3bhT7PMTQLwsE8ScQo5lhdy4x1UTmNUaAIf1h8+9PGNjye
2uCbMZ8QM8O+Li2YY1rwzA==
//pragma protect end_data_block
//pragma protect digest_block
be0rCc7XMLi5C3wTnCs7zQJj9Fw=
//pragma protect end_digest_block
//pragma protect end_protected

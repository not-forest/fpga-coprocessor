// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
w3xqazuQ1CjUrgxfjhHRVmq7fo7RCN8CqLXAgogJrDYw8pWDmL22AJghTJC0bjSq
j6B3cC+XQIW8ZN5JECKRo69ECL6e9DxoWYPu3Tkho1Q5m1sBNP2iYRDnoZm62vKM
7Vsk0OcXeXtQt5GowNpic+K9FRBLgZ/983x4HP3DSdw=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 31296 )
`pragma protect data_block
1PLuzGN9RpUN7fiNlqYL4AbdhkXaqThKedpzbnPWgqyaL7yhBz5oXYU9oEaKJD1W
JxPI3DQ4ncCpX6whKtVOEpCF0lTY3SY3v40w3ox0Jr7dKdOXpvMaJsr3EE455MSs
zDXvIktvVGNNnQBa3gQ4bdBSoIjXxkl602QSEnueLaUppKtREsexWKyXT0YwEhl9
YGvSQ9iGbIZ0g1B9ahJjGroIYxt2/orcVgt0PXn9vMgJQgOoq5REW/xECpw/I+eW
WC/LsblT9P4G/pcv/mi5I3ugsg55sUOVvJ/9Rfvrro7VeGsFsgGSDIu+GL8JAOy7
ID+FTcA8+Mgt5SSPuWE5dMJT4oeh0JBOa+iUIGJiJvBcbfyC1zkG9F3Z3j9Ar4/i
+XHbF32aVlysfwrIY/aXbJUCx21fHV0fucr6ZTydVMvE+LD7SUYgBV4kJAADnWC+
8aD2hhxm9+NJkz3jDfpHaq3bjA5cuzaYwPUf0i0KlV8ZQdrLJroLmt3Fqp/oaalM
gYwAhodmXFC+ZjQWK9sDZovU7/VaqL/TLUYhqBPP6bVGxHwaF3z/DtS8zP12e/Il
i3B7oIdHxusQPDLQ2QTT2t2FFzq/2SXprMNJMND1tbxK4k0X47CxqrFKiwVb+umI
ZxEsTeaJ1lDoNKlBmZ48aCvA8WgHoEXkJvQWNSN6sIG3fABKflfyEy8KxGT9Gt9m
6Ejs5HpL0eOLIPqlpFMxmm8GW30zyVkwohxpvdTb3ujqZpEOn+3TAQwoxbQ5LzNB
/6hNb8rM4N1GBnsnpzWvXMpaRUexCSx01WeTID1qLtATPcQIY91CsZ7y+W0kArpJ
psnxpDANuT5wWgx8Q1/XlhXMou8/clz1ocvMIsuG5Wr0L22LPI7Xh+1cse+WxNm0
BEqVG3R2kWWxkCaBFUQkyp1cwbrWWUx2zIJWgQlru4lLz4XDir0tlWAfZ34tKmZB
XIZnJEWMaSXnIrhO79VmcQy8vEmpeAf3cMBCqwKfNe/N13XJd++4Rvp4i7LgLWHn
1Tt/RX/EWi/BFeLrCw/6PdSfhWWiDngUIXsqgbM8Pw2f3/y5k3hsacKI013OF5+n
JAp8FyjMqxH2R0E0V4eecaUFDIPSwr0LzNULPyRLIq+smdheVCt5eKUn4hggLFgQ
DEqNsyaQFw6eKA+XYvqJmungeAwn6zYtLN544TKnvpv3TpoJPj3O+Qfdc2JDj0QJ
/BKNGhUEDECTpPuboELlK3zSJIdTIei3cLYzkmZPnfzH/H5kLU7Z8FvznXIkUGKn
MjJLwdkVRh+qRz6j+NWchf9dHHlU55m+pAcm05fKDwva6LpiaMYfpDvA6jS7jwho
C1MI1OzROfH1K66IK5mwFFhbdkAfXmHabXEjvIjcwdWvFW4LJGru1JGkG2UW4FmJ
ylVgy+EspJJKlHDMF3YAphzsEpwR4lS2N8Nf1qe/j1yHOcGuTbOwyCkuaSitrAXS
mAZkKSHnlmr/aWAegl5cVE4uWUF3uVbKoEOwf/i7JFn2x2civNptN7Cf3GHne7Wf
oRjI4hn1hJNreUi66qMGd96foypeZibVdmgLHnYOFAZROiOa0DnqNjHDNi8kxH+L
WaRqlUN95sMq9KhYg9n7t8HYcCqN5ADkqXZPkKpNVIhySbHwpN6AQrt7x/RYcrh7
/TXY0BNy+JnmZ8YBXwkjSB9YuZQ3pV4IBBEZURUca1YFNXcE36cCmUQ1Z5o4jJDv
0WTnTQbpis8AysiZCFvDhIUdYdNtTSSsVMVVvgytjMSdfZPJiyhO76GfdRYqQTw7
h0miEi3wQexKNghTU1nxLXBqxJD78S8PjDF387i2/M9KaHzEaCmtG35WxuVDCEVv
m+6ucp7WwR47HHvyjTNgMMkfBaJ0bjhI4UGWHdHpffrvcXU+hf4QFk1ZOCcCyA0H
AahRposEMVxdY3uLLiwrepKdyO6VnKhhC1cR4p0U49ckIw20w6xe5XIwwcgMUDvF
qemAinGVnHX7kmxhpZz3PksGgd4L+t1Mkh9zuf8M15O4q7sWv1acsCNleDWlmcDy
C2Q8IiSc7oYl6pSh6KrAyZO/1xBLr4YXkqaErF2QMSvJHBXFqsSwPqBXXlsehPN+
oIYic9XqNZPcxiqDej3/pUDB7nMYQc+KCzHWmnvLlyHRiBZqSfb46049BtOxt5ZQ
ANrjg372wBokvBAGznW8K4P0bbNbQzjh0bxgHQXt33YAqaHwqnTZqXZi/tgcT+7C
RfY+KQoaq2BF5KvkXCAxf4zcprFloXCzEOc1wKMIXDcJBqWTOzLS+S0HkKUjwjII
R/dfT8+T4dYqgxJVxqKkkA6kitWxfFN1M6dKp0o9yvMPt4VVV1BNsgNV0OrRVBQZ
3jIalvlv2r6AQKEhupuYiw5WkdGng0GYiLFzm/+S9G/2TAOHAKxW7kn1UVRYdRZD
IB/0t5iZpSMmtOg4qFJxPCRQt9Ybop0pv7U44ECtMifWGnHV5w0Lx6lwj4QMT3Vh
x/rWB1ImXnC3vJfT4Xp+CALtCkY8i0DISrQW2yazcOXRHN5eSDHFI6UfX51Q10I/
k7BN/6KYRdv9TAsYATQsNxCqvH2UPutkEY2RyxtPqexLsbCeH/z8TTXeF6Cck/MR
zpXXynMhS8fOc4GvpMG6c3lpxDjqJpJ8QLj32vq778CGRq/ulUEoGKgu9P7qWseC
EaPMbmrcik46+qR/MPl5/X+p6IceWvAR019MKIQYlAdVoBqHJMxzogfDI3h5S3O5
WyT7+bf+r7Yw++8tSD5INjgYoH3QpoxAcxYij+jWxyqZKuWyqE7btvuc0x0yrMHh
dI9ucaiUcnBWpXnG+f/ggL78ZV2A3WClYuyTRscrKFRHC4laZa3x0TQapY0HNNRd
m7vuZmvF3R8D7vMeKq25DBkoZvE6z1is4ISfStF05vtxWVfB4Eya5OxltkeaEzwX
8iYt9IVN3QUBmMaNXUX3isj7mLYttBqiCAdlh8o7stqzSaSd4uozJsaGfWg+gv4+
vPMlm/IMNicyhHpNCED9NDLM3JnnexKcM5EwKxcGfbx6P1Ig+tdVsT403/jRAS7E
xfboIMTlU6TY2r10rWqBYXzKxSyqGbq+y7biosP0OGdz62eezF0K0Bap0kwiFQMS
rpvhPlC3qCGmAbebjWCpqrNRdm75bqsBgnA5dT+yXQEaSbI0lItifEPQ2gbKpHMq
Qe6ylyoiGXtfxPX76ANJYdaiuUnYkwDgI5R8RWhhHWAsVc9IFOQQ7lSVGi1RzEL6
237JJ0Ru8cxRTOa9RJ1jLPIpywYtAKoUW+FalokcV8Pi6qpYcD6vM3prNJF5mfbH
LVgcxAXX5z/ZpN/wJo2z2OzzQI5iJu+AnkwmN1J6geN1Kn3hT6LSZApSCbeQXvzx
FJGH9G3ijTbrcY7hhvhX1n7hJK/2oqweg7OJ/viU22FB84wLLMqVBhqrJNsSCbPt
B7dt4kf92SLYjSrcI0v6yx/PtWUYl+xX16gpokLV7AwHZNK/bpHhOLWUOlmpTJ+I
7olJ0nKZ/urDoPZ8g+RG9X9+JvWaJfsqoQuKK2gQqDSvFv5hJ4a2vX/vtJVUmz/H
BVVNPP09Qx5D0Jgd3L7gn5cGBSaeXLAzsY8fYk9XBpDnx29tKYFrMgH4cxFb1qJE
gpo+wSJUdz23pDundkQnQygZdOHDPX0GMwaUAlPsMRnY8X0TISCaTEbPC3R1SzVx
V9oCB3n1SYIebqS9+vHspLQ8cuMQhMRTTGzqy/nfkiS7NWdasOUUndobP1mYt6Yq
xf1WOVNtgtphCklLV2Quqs7kNRde3BTQCBtjBD4uY0heyV3eDFI5qZaZQ8bqrKxs
gbY8RnKxN2dLJ72LjPAsEn5F8fAQEhPTcMNHQnNb4Y4hwY6rBL3gMltrl4Vy35+a
L5bVWEP79hdNKjirmdF0V3+D3kdU21oIvyTVnK3KrNtyAgVmVRJdHP0Zzofna2qm
9MLcQ0HRaPKm8KDD2qmFcLPRJ1P9Uc+dPWlPhb4bX+dXHcHalDVDGfd6gnCV/7PY
0Bdn56LtLRMkvZ5ox/eFxMYFhC/7H6e9joYKLhQSVNyXfF6qV3EQ/9i55ZITjsxB
7Ilor6fmWmYAxylnRnIw98vOh5wAajPv4n7CQMClcLJJewuNEb8stNpk2hV07wK2
3yLQQlZEPWfIWq6En6vEQ/WI2O4GslixcWxLRkL4L+LYIUAFCwNH30wfChQvdrhD
cdWkO3sXZ0BfoTs0OXEUPoGwC5c2PEXEdnQL81fMRRuQY9wR7gR/ID7nHGZc0VdU
u+OefCaepEK9n66EbBPNb4HkmC+39tSv7pRo+wxUy1iZQWaWDFj+Y6flf+p4zBBd
uwbmEeMW9kNvm+PA63v5UCVT91ji9j1ktHBIm5K1eBjfg3dresK9kws1OeZWnRo+
aHSsVARrY8v1+VunOBeBMMWs5tmQZJSkxxDvnUO9L8YGWVkc6sJUpLhsgikMY7bM
NsTmGcBazLjwig6qxfHBUvbjPzEJLcdTF8WTqhFI3Wh7uY+2ib1uDgwimFg6GZQP
PhIODi52YD1nIhdEasZBnpGdrs2L6G+YlUwZ5f/x7xmmUrr0uU7hgVO1nMTFRAYG
+IEQoyHHVy+Ox8AsWGaiQeLjCQxG3nWnYvmsQHtGJIkVY45rIWdESV+2Cpfiep4X
KMYUlUsxbfCN4vrfyI/G737+a4HpIaMQ6SMOiG9wBqCXK8Ph1cRwSG3fNIp+g9PH
lvAMXUUvJ9zfWW4uwANWY4a/M8yr2B4aYgrvpsVrq86OG/PG47fpKmYX1rhgGaWr
ClGL6Az0ojoMSFIAFAW2zXhwV9ElJp4FbTp0kK9LCMsHfGhYmKIvKIgJGhYnRhnD
l5NAMR4vDOsIxhUQdPaIcqamS+wAvg8rsoyHnLYfzxxKiWG6mzPwKQlK2OJ5RfNw
MbCTrKzZEDcCCRD/N0q/Gd335jiN35LohhEMfk1shmr6hS5RPCtKnvaNNIrw/NM1
HMAX1+ihdiM/e2nDUq2BKYF0HxFkzkj81W3XC0OIaGhnC0qZcvYqeUNCa+EdcM2/
wjjo3E6twwMS50N8GPFHnWILFrDYHvhk6Gs05Rg5vezJsG2fSO0Jsj63H8zyVTV1
VH7bzqJU9WbgirGMcaRn2/gOnTY6REu2Og6S2PcP6kH0mwUOZsR0A96YEtPVDV7S
CKNzmiCNIkTLzsPCtBTEeE8x8NZccsgfxcyxrUJB+xfTD7oGFbbBvDiBYYgi2Ou0
4n1CzTcUz14VZKHBhXFzp9oGZ0Oq4F7Q/oa2k0IW1pZR0d+tcQYor/NdfaPTS5KG
clOEKOqivvBYO6D9TQyelJBw0/Wx3DFa1Hdq96wj1TphjSq6W4Ft7Wme0qm4K99Y
7YGdLqBZ3f5rovMyIm6f5//3uRE9edT0I+i7/YEja669yh9LgqqDhyYNlRCs00hd
Uolj5v7KZVbxOzIyVOQd/yN+99PjFzaskFuunbwBJXlTWqC/XxzIpW18Yv781owi
4zdDDpmtMZjpvuJymFvlp6+/v1ZfRtYJ7fJ0dQfNl5hIwpQ7nQiebVJDBMH1xJco
km4Ck3RqmUWfVHD+RUoIu4EYj8uztVuxzDKHwOJtT1oH1ESQfHqbPnHVoFMW46LG
/WcJN5Z5idoiHWrBC1XgUCZm2N6n8t1C8zTQJlmujZU2mO/tMxI8aTDGpQK089p2
MxbF04WVzVC6elt++YQ4bwctWc+KuR9jpexC4uvEoiGYWpIIQ4XLwys+zZDvutOI
stTlNafJXkyZn45b5tgB4YstWu73eQHWsn4Hspe/YzYT393Z7NfUKvAwh12fB1+y
B4cuC7QUeC2uUqePzwm7IowZTXPZiMWvqrVsvDUZDgPhKvJCF996OxgBHjQzVhPU
MRYjvsngVanuLetFpDyds4UqTTIFHuhhp2dsV2tEW6ETxUMy6jlC3QCtwGzYUKZb
QR7SwM7Tu9BqTCdmAxb8pkewTO2ygZ0/VTxV1Zhh0F1CNyQQaaPcWJdM46TKwB1F
zbSl8L6LuOaLKBP/QRpsfGja5i99sd8UfCdR3Vd12DIEQphJuW00krCC1LK6Vitu
0jpvabwqKOf6nj6mZn5v5f2moXn4HrMID0IZYdnFh2N28hs1y3zziEJpRK9eiaAi
CTFe5TVjjbjbw/4Abyrjc9093Kh2zfEAPdvII4r/8Sl5eR5hnyrvpENmvVWot3N0
4P/2RhJl+bJVQTwKGsxdpYSMdGNuLcQ3uoCgb1gC1yiPvqiVwABdd2UThFBa3SJa
1ltGbaRPkoPOyB5pTJOTnrxhQ8m40o1s9MuulhXAHmY+6vs6ffxf2LBUhGighjDn
SK02V96S0HgZd2946hMg2lrzc2SOrfqZtADgRJWxuU4dWUDCKc9GYEclmaDCj8hL
ZRaWadUjwk0im2D+UlhJt8LBWb/EMtS9/rjbNuzyD8ZacdBKFytWJ/yOa8ebiV10
TfXedsEevnPHRAExdOxESG5LW6IvafmJXjio+gdlGzwPQAKp7A7wK5sZ5WF8/YC4
lEdoDAJZKtxZG/V1SuU9B1MQchl1jXir5PMCEVMcrnqs+tp4rppFbsmHO1lSgzsd
+Ni7V5uKWeOXwBgOPqbAjs+P7XXxYc9yLjBBVlTFBiCiAmIlyhmLIWAAazNbs7V7
fRyQwxnHWQobU2+ffSbLt6OieFmd1XEsQxMiDO3Xtzw8zW4gQMgNEAh2MbibHwYx
azUWcVNfG/5Ry8HqJKpM61wXVskvijwdgz2Ri/+R7RU/j7r7sSM2N3LQSGLtU1hj
IJz8boG3ac9APt2b4SJwbVn0uIBArMLghiix4IUBrDvWCykNQ/hnDUP5cV9hFSRN
TQig1ZKZRYFQOQ8mqrPs+zit76c46mq6uTzOiTKuZWhgohoOSZ34H9RHPQBhrSlz
nxTWFkzs8eH5gVbjHhlDoDxw2nJMiKyPPb737iaAxXRPgzrT4KE8CY+J59RbqKe8
3/yiqCOM7bs3PbaH3UAd0pj1O72JWIeHIGldJZKSqpUO6W8nIZMYyf1kEzYFKeaJ
3E3VXBN4573jA+U8Rgg8O3INgSTYDXqRKRVKLGC5QWXyuxcyWZYWWjAnlQ74PLru
9mMkfGNcFWw/9TxDIpW7Ka9eV0ceEQWDGQau3Vbx3ga7n8O4CjZPOqsRpopYlpkQ
x6A2OoZQYY3NJbtggYKzYwqMJ/C6o+aEBniH39O2s7k/zzTmw+c0BRC5qz5Dh4K/
nE3djMPvmJZE757tZPResb/njs0w5DZvTfuOH0G8WEzHbQicsNXwoOWcokajszej
7z2YfKVWgrtIONDkl/saSERDC1v9jCMD1DJ5U/Yulp1f/G10UsK1Yw8RLABo7MdF
iV5rajGkvitiqk10mvj9+mM5hYh0FQ2E2AUmpMS6d9vRn5m4e/O6rZqQoAKb8VFq
6Kg2r8kiBgNo5TDoHgFPy+45gksXetzScnMdUEorBWqic6TxJCz0w6lKSI79aw47
Kvb0Ebl6EvvorkXiRiEtYdSdx+hyejv4VTosbqrGFoIkC8nUtVW2YBQwebGUG6xe
5PkfViYMXl61lp8h6n4CD5rRSzC5T8DKUAxhtbR/punh7ua2h0YYqLLhZIYTbqA3
Njd9N3T4xGTsdHMriAxxyoqotD356Rn0V90hmmO3IRFbNYEJtDHsADTH/p6I1z8U
D8pEAc7RJreHbQ9YIq8KSdkrVnilC0r3j/MEWgneUfiYlzokjHx9DgwH2TbU36BM
OSUoZ8xLRcg8xwXvyHAVIO7LsRtRfQ6UHKwLnIhST/se8SjtOqKI2taXj6AQHz7J
YdfaBnqD1IoNuK6N4kxn8yv/J6QnmjxMvWsg4666g1afRaUwWrnhNm4EZtxEG+Fz
LFLHgKOSum2FRFZLT8UUZw7uFCHD6ijVcOBfq/K0i04v7I8OFSvXyKgoPXUk253l
kDvkcPDw2gjhq/Mrznp4tAULoTHt4jaEJYIbGuL5Oq9IeWKpBVh739J5WKxSZ8Li
60+WxgT4o14UblndI9LRQi8SG2H6i9n2YWkpj0LnnB6fGukhDnL80g6DI3TKTITZ
RJimOlp/IoZhLcyJI5b5SH779aXfOXtvrghNeTmJN0wpfRjQBkHgaSZbunjFUhJY
/jynM3wCebbqHvgyIK4RZODANSE8RMv6YLaSEkv1/2jWQNv8b7tw5tQpvhKLX5um
S37niuEHXXPqvyL+Q4vxqPgNo1a2YKs7jLKmJzIad5nUt4WEKS7POxmsCYnBJyLK
+gnfxFf89sMiFgXOYIwGtzfkPRwzARa2/NF9WQrEgsKo7GBZEu/9DvQ8oOb8PQ4f
r3wxhmX4YFaJpVP92jjiNay9NQWXSLdN3B4Chgpb23iriZ41S2f8RLljaW2f6IVA
JbQifDAWYZEnBMBOPctNWMeV7irM01a1CBEIBrV5SOZCyAHa3iTypsZ03ghXTVz5
5zgR2wLEs2BUIrQvuwaV//H89kKwN52xkXk8RliVccDhWpTgnyYp75PlJ/J6rKQo
jbuDO+e92QwOUALkcieSVSPtvH2J+5DjMNozZ0rSfbe0RpEX5d/9GU/q3mTLIcVk
MlOGqKTd5uITAUGvi2Ap2yB8WbIWhhQAFQ8KVz8bdslP6n7+QQujGPsnqznTmrHg
qjOB6p/3QIbfYUeYR4716sMON923cHxygKG9Ng/pMIpw82hf5aWmefPDKxnzwytj
6KFvFabUN78cZVqlM0wQQm5XWSzL1Xo29MnNgem4Pak0pkebrOab/lDCJ8juq2Le
k5zLMKQ28GRGb7EZkc1ilFCn3oo5aKefb6LA6iAAtLXmdZSElfaVf72PDH/n7gtG
i7QpYctLDyX7yNMU7z1H7T7T/L/Vx+K2oKGSuQqdfRX7ZJ+WLZsufdEjEydP1vh9
ukqZ0S46vcIvJzf4JtCdnuAqQIzENOyjhpZ0QD2+TmIiWY3VNuqNVj3Ke8wBNkeJ
EZTCfnmqYu5Ct3hSYXaYGG86jvd65HNRIQ8decooF+Aa2yx2L8slwR/Ib2+hPWta
3cf4fkwVezBTLBIkcrMiRBoFbzjqPYw8eK5NvT/TibW9fOUtMzxjKNUyxJPOtPDb
7PGIaiUgosgEEli32/5Rv8oQ8qaziu7vt8RocdJBhfOKsJiQDaIA58IzrAd/BhdT
/5ES0+ZH4FnWXR6kCsy8B6zOH8SxK+lbMe+RJx5L0yW9Eh5WkgzH08U03gRGdBr3
EJpevch+q+wdfsBuqqxouDHeYJWEd5vtnAQITqydhL66dA6LZ14HTKkTRUakHOKl
lU169l98b+Mvz48YdrGj89Hf2N1l6pWJhz5vr0N1HCAMGHdt7looCOCu6TRJDO6h
EPRCWk0ZVAkGzXv1H0+qSlZBQM9plUqTVN7/bO9JDgF36AUZpwsCeDVadKZQC3I2
1yKpl8m0mrD6RLvD4PjG4OfmnMrkGvqEBIN6I8ZZQOBtQ0Le+QkfPN8pVXCN6CpG
f/Cgjc3BML3JhYuqNbLuxq96rWi/CXePsLX8TGPgWZJnGKMpuTlfiOOlladCbqd0
gaaSM89gFgzblCLziCWXu0gxI3uS5Zz2w6suW8cOAFmj0qBb2pTOj8ZrfQ3IZoKN
ZW98za46CwMZFdcl1Nsap5+3Kq/Jt10iFT8MhoiNkNDFlLbtiwPk5/g5OxAV9z6k
otWcofPyhVeuidRYJumMf4j6tFooWqxMkSk40vidweAwn5Tapu8k6PSby0os7BBD
67dWDaTQxKgOXjicNHsJtjpKLv9RfWfMZrrKA/yAzWdlKn/1rXOwL7FQ8uZRRd5y
cPpIkqfRQaqh4wVTAw5zqYzH+9TNUsVU8BdTbDQtnDSXFOmJZgc/ynRhTdP3BpTM
iVs2G+SuLbi+FPmmP8hGcSc7J+XfJYzH1NRf1W6tKi4W6wbmZDpBIFF+2UqNJQQK
9uwQxgACPQOSYVtx0DpMkhZT4MWtdSUPj2nFYPatl8jGMOKx9mAIko7ldy/FVXd4
sCffLiUUFAJNhumc1dPKy2GVSvW81cLl7wBelW7xmM+Kr2BurTEqc8m0TOvWIbxS
IGoUNz3SRX087L0AMFUOjI3pMSbNRjEnCjYLPuMJJAfPXP61M92+HmYzIQcNsgvy
/PW6ncIGVJ8cVvNDMmBdWWGoQtnBJoiTQCTo1tU++kaGW/Uzf3MDONXVYfd3xYBa
HHrAsR+IPnABexUb94tWIpkNi2Yr04A09PcsCSELTGXZZZBiDthZrCkcy+R9rJ8o
8vLvCAMVciG0MZi2qUprYghMbjLMqE/UFJnrVOdcfXhu7YPLRCDz695vt1dJRcNh
Q1j9auRcKY1DX5Ii8wA5WWFAOnmltz9AsgjxWoO1t+Vuu5ZMuRAH/FmlFJ0vUg5f
wytz4rTz/8aYAmmKhXxNTYoRnuQe7lQHo98a+LDFQkV0AtKkGikHW2ApCmyA8Cov
WthR12rqYCTcd16ixadBW2JSUPPzjvBee/UJEAMGJ3QRcwI0IGJ5FIU/31J9jq5a
00MvWoyoOSNUFLyYTr7+MHLu7tSy9wZivs4ArEoh1P0PJTQntNPb+4JimCLMZ8AW
/22HOI8fc7fC4KyBG96F3rIk5VcMZ4F/oNPjTLeWk2l02vaa1KXdesoQ6EeoCyx9
mcefkbtIXS6dlWkZmQTZkdB7sSBbQ9PXAC/LyOkN1pBVJ7Tw/2H6mWaNN4HEttjd
oZH6+AlJWiwXruEHml5AFxeStW6r/B8A4HEcUEIVlum/WGDmdTu8qyJisBgoeOAb
gmwAc6MFwnBuBEzTfugFwSR1pbZkyTsTMj8yJcNjOQyJ4pVPldB0+Yzn7JcqFHhZ
poYkGIZ5BhL/Hpw8yfWUDsOxUkHkwowGBEwInv5+ls3RPUvPtxuXfyaDuXdlrfoC
rBFdZXQvQiIXOAjnnKMNpP3xZsYU88wWBCUVTaJ3jK7A67os2K0PYwQt7v7PIKMY
C7LqFQemrQJAZlJZTBnySg/vAIqJepyd4gzlVKXGFllYOli5qY6AyzpmE4L6jHMz
HtzhWs1QDnO2u22yk8z/ronaWip4Jw3yz/RpnIpKt5LQMK4MDdLwmOlc08xbC7xr
MtHHzWSaYcjhJXW4SafJ6XdG0d0ree13A3YnAUSKNLK29gswuxxM6AidG4Gm4qxF
ArT7S646QPGRMTVc7zprjzmTD2rRZuOs7qD5jbtO5PgLqYBk1W/UglDH8k6E2ku+
9RtQk09tV2ixxHw7XCyNcKooMmSpiDuJwnDdPwY4R9nrOECUArllVpGALN6bHxqH
bbK0E/XC+Fc5Y5ZRfEJZQyBquKFhkK/Qc53/UR6VGcIjGMxvxjtlJ/l18TJIRSL1
7wTVYsb95enGACe9OzAZedGsVrbQRMXCtKY7Vw1rOGfjRU8WO/bM9MIeguzIKogc
zuIjNQWzaGS2eOEj+Rfhpz1ZQcHV9kCyx8qBfebLxfw8c1RZ5cjVzGr3Jp5k//T4
F/sEuGnZORI/Lu7GJhxGnAGt+7eGsZQwVkYNATStQLk5mDUo8ek4TnTizd9ZtKSm
uPisnWG4uoo9mfZEmjzllWUaD9OhC2M3kMW7e+U05P7uDCPUF0Z8JP/259gHUIM7
gg7450Ff2UjXUAQQ2dJg5/4ZFF9zZAijByWCadHYRSgm6KnL9G11cD3W2RKpaUzV
9irta6c82WP5cf+Qe7Q/psMFtEDpyqSXKWmgSNW5Q48/uUoVbv3eQB80DB8WldCI
ZEZWGH/hishC/cq2fKTvENrBIUEmB7N494rVAGamUG4UAg607Wpkelv7aC6YEL7t
GwaBsp0I5c2v58GyPeEE5GUlc3od1zNA1FD4CjmXRT4Dlo1sY8ipjPtLDnY3nv5Y
IGNGWXsvnZFAvC39YotVJbmC3E0Qkd4xR4f04JFg101uB5xsDMhMlL4YA1nv5Mkc
3twffy1pxS1FLPWsUGf3qjIsy3ylB/8+gwb3tpuQG6qKo+5NGwufQ13twIu+8CFe
GYsPkLsQ30mnBrgqbG8INnqVbeIYqI54rYu7AjZyL9JTv706Y+YIzgfwGrnkgNsF
n70YhBbou1oJJ6l3Sa/CvFOkDVOkJ0tkDfwqPXm3U+BxIwN2Xza20lPIezSfZnqL
ZRCB4OuA232F2T4aJfSE2uI5FsW3FPt0pmoJrqdXLXeez0BqerwhoRRuXGQZ51nN
M0unwuLxgOSVpnA0pH0FgfBkPnO953/FwFSkpI6gJ4slAQ7A8ZItsVRcCpe9Wi8X
f4oB/khs4HNF/guyPLhMUpPzZ6WAuqzBwqBgKPbTCpccdn6brFD3Dq2iul+STKVC
sXtWqNKrXokUv/aFsTZTphmgprBTTDAzdDeoU8KbwN87jSGR8U5ziFWFHYB/lFZB
9IJ64AjktwEt916FyxXkG0UTB/VDt/Zxtk4dhSYbmdFTf42BLS5OzHUQ31/yp7oH
lWeci7GDC8pep6ToJFoeJ01k0fyzZ1yYRV2OxL5gQQ1DCExcNXOUoRnZ/mGLI9GJ
MadJEt44VTWkwcPaereSZmDQYymbd/uRLQnsh/ahY+zAA1kWiPr9Gg77SX91ApG3
JsGjmokUdvjhZu2/KIoA/pjOLdGE/XMaLXGERCgEFTGPQkzehvay+LgV8AlG4tzF
++PJ6Tm+5EJCiYzWZLsTPpDiwjEi0oqIb9YOggGXooqeX1VehnnnCUFohumAjTPA
4/QrycmdUiqOOVrBQmmn0EvYPvcbZry9hj9CSuMK48/SbVwSp4VLBGC+TlBOlpv3
Se+hT1W5zMeKmnD5/41Oe2JLSnCfgeSNnYyp3CkyJSixLXs1OOSQjzYyHAqmSqi3
AK806jSwb4G2RTROiixy9GrRWW6aw1bpnLQZoWiOs1DckaQ20G89Z2kHyCAmLyas
NYVKP8bWebvXPzWgODdjbuEHqTykqLJCsInrVmsQnVM4K6tWw30cZpHcMtsd+zBV
GXJcJM2IScXVUkAgN8H4DVSKwlAQa1NuLA7DejOUN4PGeEreGQYksQqtnrUkoeel
KUqxVxNRGQbQOK40LXgBdKEh/gwciq71QFVRlVauVwX84p7e/gdZhaqEks/YOaFG
eDT5njtH9005PAAwseZsz/BL1EiFpBDGF+vKj9mFRIa652srvC5cG1HQWeEBXdi2
W/3EzSWlEYILMrU8BD3W/spDNzZYbUAUPqyFYO/NADu83SRN28a6gHjWv4LX9r0y
zUWKy1eESuT7j3Qu0fLlhymORX7lpXLEjUqoZtpraMY+rI+g/GSqVYNyw/QlGZ1a
BvojsBEWBu08ktpCIxqKoEBxjwURXjOl/4WLHyk+opSeLMjnKfrvZi6UmwiX8t0J
n66D4kDrJA8588MnLQWE3miQ+1PKuTTVcE1iwXIKhEZzETkOSw1VgIPB3eDnrQbE
i+E0fdsWX0zNoRL4knI7i9kKU6CUVYterDXN4MubhNqifqaLE+zMlOoc5Rn6G6kt
sSyvIOS2V7mvAG+j8KxyfX9+a+8+tfD/QUcfShHpvVH0vUGnHF1sTh9dFTiVp8Bh
8eoeF3qjHGy/9/MThLiysv3WhisPGTAaBnT48eZ7RD70L14VMOM0D2VXwJhfKxGL
YLNguGK++/iinx79C3DkXWeryqBTZIBTC4r34SNRDUmkRgvE9sg8LnGZmaYrFhOI
neq7EhEq/zmZZwV7jFhEr+rDx9kMzZHznpxmLYbDEkL18c9hZkpeT6MWM5Dfv96C
gZ0o2RGIchItilao1fdF3qquF1WXb+Bvv4jaNLU/Y0Oxp8fb/43z2wXKHyrFFX5g
88Uy9sbD9NMEYysffZkgz6iq+Z4GjKn4WUWyxRsKcges6NQuNLTawbureHNo62SI
QSkxogIktKsM5F85AZ1dN47P7haBfqbUjeEKhSClMagLNfzXoJrrA3DFyxB+C0cQ
Xb28nrhfWShIXrVOh7WsHsXCYUH9wKREE+01IpwokqJc4EKXljy1OTB242rPgXI6
UBjaWDRDF4KMzf3OOZ906LS2murFWdZtEJqPtTaTPqX8jNTCGirODHgF1bShspZP
UkGl4hfXiuQHH7cUmrhBl/7PJTuM5cvJwPxVpE+XQi3qlJZh4uoznRODOsN0KIOJ
KclTKUrWL/0QISI3LhVthF1GiTu4v5QVtFA63E2nodb4gtJiASefKvQ6L1t08CgT
koDJUwt2A+mh6G7OORsOCmzQ1dI1cVoJ7/HNwcqCnBu+xM4d4Gg1+uFPk8gSU0Mm
X/Gv5m8wTZgYuQgcog/Y5XMZrL8Qlmq7bbVKoc9QQvrNv0lfmB4xxRSBP1V2p0eT
5GdeQU9X2Oxw/InDPhXtEZT6ireHXX29Zl2wCfWh/Fieqrhqe1Hp8MnywciB1/EE
eIAO6l4DVVqLjmLPLEFJE5c0nNLh0COl/QRe2v0yMtYrreWQNOUiaoL4iKUqo/GM
vTQ738awA/FTVqiKa99LFHzucs07g00uOijZ1RWVMODvbIwVAzHIz/oJasxJBWMk
uihwHPbnzdO6rdm0YZqfB7b7e2TW0IKmMvOW5sPgQonvprMXgm4bI0euBpu7vBft
SGznjDxQKXy2Q6E39L2e9YaudSJgc8T9YE8h28QJrN8oYZSVwuq+xBo9xfqjYc2m
iHpGR7uRMm0BVMYL1DtaNVxgznEj/+BCVjk78G+Rcqr0L28QePXUPuBUsYtUG37N
UQoI64WmtmrW1+78VpC1/yGdCDMb+AlvLoUU22Aym/necZQoHKIzCWOc7RI6AAGb
OfW92G9al0YUGqJYi36RVi+Z8MtfF21Z58irqxOEVnmvCiNT3f+7oj5gcJ+n08RL
I3LvPh+WZzx0fkelA97da+XFayLGD8ae9wR0z4OvYvhSvLGuSNkF8pJ3T1zcYY2a
JiTonAEaUAj+pgCIAb55/WNvMsnsst2kABYkC4iT+3hGjiOMeqj9gIbjStVRMaN0
yjPZ299tnbGIQkduq0ZVvz24KJfyQtqK5j7L812tuv/CyAu8QqPtNifdwGzElTrr
sCMvEs49sKSxcWH3/Qg3STWa2SsHipOF3cXvjmaaldrFGK5PPRXwGmN+nFGJLsOX
oWFClusZfVY8BzNdG7uWL8ay95k7bqQBIwOZKitppIUUo5Zo1rap4NtaRHAZMAR9
Xbdw27ROqXpwATWyOeq2LBnEWyKRKUQMsLfcMcrtXYeQEKPdKY/0V1v1RS5P0EsD
DootM1Pn9MD/mFTFeg3WvgiyQtq7BiGddCdSh3gdFV11EFJW/r7T/5Jj6T4wbuRR
oAfYVSkv5joDRqREACiqEHg7Zv2coSgzcoguWLxVwwUTFvlaUKS5PMeixrNpWDu2
UvE3uvI5uq7BIbK8oo8+eaLPMojMypSNKt0bQNz0LUcHAXfYikDxM8ago9L4ofZG
6WrW8e0blHaiZRbF8G5F1iZn15bzkA3WkOXAwmw11W+ZBW/U7RIOOFSNzy9oTMpZ
m7Uqjz7F07Jt3aPmAoosVcGIkVLxi5FF2ltnJ0J92y2k/zf7RsRGbKi+ANpXwj7Z
VlzrFxHlJ3hYbAJSvG3Lfbt526sp4gYTTdLVmXl/oZihN4X0h0dWpkPjHVVZ5Zpz
IS/DP49vw4oBKFy9aQjUrOeB4I3aV/T6cvSaJ2JckWT73Ie+Kk8z8canK1QRdB4g
EiyDl4viFUZHmT5OhgoUOJmvRpPYLeS/PVv6ZSKZ21RTmSnx4koW8LtUUbsdSkVo
TfVHxF75uV3DfyiiBYLEzc9GM0lj4jf3/HHQQQpe92+Fo+MxpZeJIZyAfJbPwqsX
aisMHs53BM6FTFCJ8bEPi0MVKBp1YBsfJmP8v0RSe2I1BrDLEo3WDTQqzsneDd9U
lSbH4GaXauJtnYf3G4rO/0Mgup8pOllys21pKTmBZbh9JrHhchrxALY538b3FaUO
n32JG7CzPnvBVjY7fnxgjF9Sb2RgvfzuRKNskgcxkUwY3qlYFZQUwVfvR/MjvbH/
VfgC+B/CA0sI6M8R2TY1h9GvmS+tgbxpYo3yIgTTLY4ebAQFNYvEGXq/MwW3l5y2
iUcvkSQVnPCR+F6+8m/00bTA+1GKnQaTacAfiyadOdOGj9saWAuAFm4IcvkS43Zt
p64xCIBrJWKb2s0BTuxA7I+V6oxqEte/qXFKViVwEOR2+3u9QIaTYj6j/lSNkrA/
pRR8RTCkffVaM0H08UzDDR3P1sGwk3cOE093u6mljFBFvl+TAPaSLLFhE3Yrg9L+
8Dkd4CYq/qNrouTaR8miCVu+k0GmhO9SV1zTfP4L7nLMX5RtzwjEIcc3WgR56H2k
AFIDF6OlJGLOlQdWiMzJq86r6fg/2x3hHXPBfKnupVvKcIZD1h+ptrTwTtlHAN9m
xzfJTN+fWf1dfyDm4JeeuQ5rh7ZnMULj/Fn+KYw8Q+Td3vzoZ0NNyO1kJc6kRIIN
MUwi1x/RZu0D8E+d57/oqg2nm8kg4PyrMhwT/trXYcnEhvuDwOFjQyWmmCrEvwEs
+tsxVgLs4ESqrGJq9kS466RStTbdx5/o45WGPmK29egI59VBEDDNWSBIyOyQQkqS
OjChn3YL3S5IjKiavozmgQdLYLKIkflHkZZSqWhiosspEJnm0eb7q5nUwXRFf8KP
5LErPKOS42bFF3k+haHCxdZf648GXfR09W6KskzZK8mYV3BrNQXUfFo9pGjDkMOY
7K/n/UE5WbeMtkHGE3hNLmFuDE6aES1DHSn8wIr5VjGIQKeJ9BobM4J/10SJdseg
9Hgub6eXEadWBJKzYq8OuXrHGCwhDaTeAxRdxmdWY1k8XD/+HsBJVbBBtVwApWhq
qpELSYMUEfaKdVKqnm/hCPxBDSk6oPAObYUBf4sizpZ3kdNctSkZIwfh4bJ8FNpj
yPALgILm2p9pG93x7iGwUJTMTz0txTKmSiFKxJps18zdfAqFW/Pk6Mu9rkJbHhTe
i8SGQNsJuiD60pk6Vve53pTLS3uDWsIPuO5HbGWXpZM8J+4DJUgEe599meTnVm/+
Xt3OlcKD2hF+IEL223KDMwlfktx/SQYxjB/8O+IZ888cZidjkw6W6zX4Mw4cpD3s
W7RLcEUQDn1OlbYTYcrhNC0TKLzJJsrkey0kD0wweTbNp4RYaluqshZH623heOvf
UsPp06JktHNmiBHKQateW55qsYImReUIucDCydvrbLDJAsi+AGbKmfV+JBAk2vzo
XtlHKYOI4NXbSl4g62gH4N9hUHLTO67QI28SBn/WrmtAPQi6GGwNQFcRnAvX6MX4
XjnYPbHEBnb0s4w68C++Qn5JTBGhPgBixdQfRbe5ZXIZiFY/wNVqLEpffGw0Vp3f
47JB8pyoq19jLoAEi/78kBZTdTILLQQtD0gFs4LnhVIQuRpLxO3+Lu33v0vgryie
EsHWVy6VL3b2YWeKWCxEUaY6TRBIGig+W44vpaaVX+Zy5c7mdrONZKg40j571aO0
Ap5Uc4IJY9lGAihwTpdyUdW+39iezMrRnrv3C0gyH2j/L5pcBSqNS60RTn1vjvTK
yrRD8KdgNjVJJl7Fw0/VSHl8zxH9dGhQkB3Gn4V0R6lmr94DOCkQ1o4nExod0mx/
8JTvRtCJ48jWIXGhoBXsMqpPGY1bX10GfwPniPFPq/5IaVSsRUG71rxHRz3vW/73
oUM4IaPgB3FS8w3GuV0tJNvKUds99R2vmylTBMUFBiRQyT/dkVzIpFySMb3ig1Ce
5gxXQPvHYEESozz9/zIMzKijZ4TymrJ/B/m8nBu2rCSV+rnYp4A1jw3h1K3wzLs8
A6tanR9GMxh1or2A74VoZfKbBVOAljBgGYoxMFsWwPEHayySZTmm4WaIvaYHCbQ5
cY6+iymtnLnAna5H8S+y8kIv6dpA9miOeqZrPKw9Jse6orCuVqMsXO4ucmVY3r2D
DTa0BRLYdESbQR/b9+s6tnsbOhrez1j5OU7HCxFyNlvhksDxY1eJcGi86ZtFUCVx
Nj0L+SeA6mDU1W8Q8zIdyIxhG8fV6JPPppdX8MlN4Y9E0qfGi9b9DanZ9/x9agkj
JDkWEuxcBfaAyRuK1UvXwpvWgGUw+8K1sTfRo8JjXLTjpag+tLSdOcnpPK3U/4v4
RXI3FuPSRsrV/cUl3Jhhrcbvd9Lz4nOHq7l10LbJrhFuUXOkn7b8QtQJYJbOGsqj
wEcHXaCKZP661twvQbIwl4m3k3+rioEgXjfsUWCjP08jLZsMLOK48nPYj6EzX63c
gi126rfwC2liDhXUuhFme9KkU/fNE3Ael7F/llqydO9Ce6LJkylOeRL9XDqbYnCr
1ZaJw/cwXh8ICE0cMui6BkPWc7VJGlVpyA3IUcGgBmfj+tysFvxf4PR4RxOJiR04
0Gwzzl4mJubHTcfJO/cdAW7dCKK41KSiwIhD21t1Te6cVHmeHuA5/lu8ZA98HICL
UtwUWMr8iIayuEd0HpJbGCxeC8p5OXb2sTja4f54FE6PkCDSXZ6UT3vaDU6CVHDZ
ky925RDSqTCLxmDKsuTJVI9kMUYOddfTbvhFHFDvaDBVniEYv/isHG0ISprfrv3w
/FW1Zou6x2efPfwrYUlAZou8pgryJi4DebhwGkyuD7FxtGT9SSw0cyKBbDtfc4D9
enqwrEJC6yfjKaaBJ+lblTUI28xZyeP4OrwNmEPldO0qqYXp0lF87mg9hjodg9JJ
/UQeOrp+FXGVGgzVdYCrkMboZaJOEo3c2R86ZvdiRqtWVGWNhR1oUxgdjJGB9Vk4
o8sxs0Mps6CQLo2j/5z1QWcQncEMYwUsNiwjTaMaLQVemazOdejQvMHhrjOCXUo2
KJeZOK9JOz02MY6lQcJB/t1HZZQAuFt75xWQvZFm5uYg5CcNtqvxLbsj91eMIgft
R6GYnU6fn25qAioz7M3xHhAwyfFz+vwfcfIAAGSG+4HIO4IG7MEBnqtDEE79cHPy
YfYHXFOLf2I7m9Kn8QwHsCcdNqJK5vfBZtNvMqkZ0ko8vLPl9HWDF3nec2//qvyG
sjdrQ0dQb8J4vFpwpScecwXDkqPZFmNABgS1YXuZ4ZavKSXN0ZMQKBf/vFp/YJH6
RduwIlNuA6zT17UMz8w09mcECUI/FVG4sYpBXh6qamZC4xz4OCdTDEqut8edPt0Y
a0smztsJFqbtAD4Gw8oaJSenxKl+eKsQPanp0SLDWxpqTJlQ5AygD6/oOQ14fk2b
r9JnfqUvr1GTP4Aue41XxP825jlYU3IzPs98iAGP31q6JZRM7lA2N/EVsjBSu+7S
ckO7tfa0bbVxuHwgMHeXkY4IRElNIRLsHKIKez/o6qLFir1hp1YFdn0V6i8phLQH
INy/PmgYBLrT0EuD9+VUs2BAQa0mdnMaKXzSbsKwhfJ4nfQ5ugFSJ8tt/iw59K80
X69fFp89SCvk7HbLhlXlFkwPYJmVjEIFWiED8Fx0Lbei4ezT5lg4GwvYa9fFnl33
uY/kMvwajO/B9HB3CViUiRWSWUsvd6ZnFo1q7dAiPj+qXmvxcfYsLZ2moz5DMj8m
+Sid/GSJfrXjrnGSRXfRpDQhz7+eCU0fwwpycauZR/9nidgoelOSErKGzJmLn3oh
h3q95QrOX4br1aIOYYNTFMOvUrIsaJ5M0LDbValxFxOB+yLph9U2fP2y9242U6Tq
Ef9v1ixtCk7yj02ZeicK+gsyE8LMzg/VylQrWuSLifLzrJYm7fghHMwtAWbu2ESg
OJFyG+ocAzKcveT4qYMlk4gCLgM1JwZFvjM1mJOE5IaZpdvwOkRpzOzFGdsZC3Nr
sfaMU1Ro+Ag26XM6No3zsEzKYB2s5pL42HeUEsIfzrtYt912u0pgdhJ3EujiWMLb
8OIF/LdTG9w7k4R1VNCFvsPwueCbxRAIXOH0neWu9NdG/21YQ4LoDdZ6GTvep9vc
BnFilO2Ss3U+zYnrwqPtuUi3X3UyQ3Q7nCKBvVZxqgPS43yicRfilrm0iZbssaND
DDpNFTxge6ok24RmxKpsqakeP8LSqC6Nv9DMRAQGqnrXbNlkRjizfGXZw1JridyR
rz5yYIEgGa9xfV2wNEhIQnGxZxUnwV1tJirr4qzf6pOcMZ0TvtvdYEQFfD2h7iFU
mDfEi8BE3+wUUzt/y0rwXL22jgMoeKW+VeYsotzkQO+3Lk/SQuMEP2rnvln//pR4
7p9mm3ueiqG/jElHwGB2BTd27CwwSsGlhgBFk2rA1Wc5rf6z3NhBNirbV/u0BoMK
CxsUODR4Up9s84yQU/aaesjc72oQnlSxPiAODKJJWR3UF9ksp4xWg0IW/9m+TjAv
GkWDymcyBUJ3dZb05E976PgKyvj0E7o/pVUi7czpnMBnKjV0dneAucF3WDhXtDS3
uxEWIFrVwkevzQVYNivxL+A2UG6LjG3yqb91BsNGKMSg6lMiy2ogfGu7totMDNIR
FDkeW9Ph6irxTEbgtD0LQgcLloADyoUGzOI+VMJQcN0WaDxFySqYnWJD/6mNokzw
ajvAW7ugQZiBkHEwkrSK8bb3pRMv4ArVkuYEyXClmCjnqlcs98Xdd01JJiuFKwzR
Mw9z1XW4L4atPIzRvIqjfh6aKIwp7dojyiOwgqpzcULao1H0h9ukoX24E6D0/vKc
BQdcnqkf9NfYYzslO6Ho/V7oWqbfiwnwYKoE2FeC2WOCQ6LegD680NC1dSoU95ku
7rCkHbLMDnMxyXjGL1ueAomwI6n6dz2VSfVcKNO7S5/4hVa/O1tLe6u8CF0bZsiF
J8GESoDTvkHEoRnGl0riIWhdoVTgJy6aMYTWec6sA41NW6yD0l3Ky+pexRBqA/az
/Cw5b2v0Fumhfn2QP4Jj/IT9GQ6XRe3CFvR6bnuW7p1pk0nh++IkjKSvUYf/NQKL
5tFYL6tRS4scKFc0+ldvRQ7tSAnWRaddDUzWqQJKlm3ujay4rgBUPx1aasHlgSPp
LuTITQR2umwPLkPNofUV9S2ZJVBa6dcdaGzBsnpxAva1zCzwWGSnO9ms9XbDYi9X
wi+YpOIax9LKTZWGbzUAobsHd/DmIuET07CpD8Jc5KEPMFC4H/VGkZmwQC4QOCvL
88KtM8TilIraaYpwbi2DNFtzV7F8Bo7WGoSXUTB5r2tyDVQG73DO6ct5/ovcFx2O
pf6AUp0he5du/xlYgkjhJibmKj6zmHQGT+WRBpEE7LzezojRrOYBQu0+JRQfV3ao
WadKamdqMP4oVaxAQw5YnpCoeih8Iz6R8YVm3YaGLAOGbwTbHZSm+BeyOOKjsa1z
cjGF3U3aqTtk4CX4R23NIYhJcGe7sBaTxZxdsmAhd++fsUg8jZzouJzc0jMDSFBR
nVdiqf6B+nxx3Y3ese7rJdHOHUt4nYbVLkyK67B9GUCIwLh7ILNYf0rq6AGVEV/X
Eka6L7Z1xt9fRMBMdmY8X5RyzulSvj3VzfgVhi7ucPIXrt7xFXYrLRxmUsLzNMt/
fZz95MTYaBki9p/YPI9bT9qmyoKwdaJxmwdxfxXBdtipiv8m93d7uWm+KoeyAWOA
L4VMgZQOz1OP15elOapE+cocy7XLNfGcgz6fAG5OPO/KQGCjynZN50OeQttDpSh/
1muIGFjtFXQjlTz7tjtPZ9t3Eny5jLbPVotshEnewkE3txMlSAsxfUR0UQ+Y9t06
hK9mX+v/+ebZrwyKeM4KKSIqJ9axTY3CSkYO/kpiCbP3ZcvhaMjhqC0VXbThghMZ
aEVQH8h/7loyyH/Ni+PNFo75u35jozahPKDnWzm7rSy96csTpnl8pgNk4dIZ00+U
KC59/Fa9KtujhXu3imSs02Gf9PT40iWzq4xeR205+B5paWkbLA1x0640sP7mOr70
yDYdlbjYnTrCw45EyuThaoYDg2q8y3YOJ8otSKCyJiWj04oymkIJocD1mg9cR1eL
iFfgrkB0A8gt1oVPJj2YKs+tiTNjjSZQLrf5owvqmFHeL4p5Ce90Fq+CgpAh4NaK
6V56lnlQVwUmMts4fGZmbNJMDAaOz3C9LkQMhxjzNXO3wDJnbGqhsu96PcG5BwJR
vdKKc/4J0o3Vq2juLeLNdqyFvTUaKnNZAkoDywyohMN+wrlXM2zhJnZkabgyr8sq
XjTWrHerOFKhBFO8hQOU+oXyVkKLFAKE2twYOiNK8Z2jWETvIiUtOXqD0d1uup5V
E6yf1WWxw/57uZvyF/MMy4sxoVkWydlAGXaa1lhTEtbyhO/RtMJ0nKxrEhT//LTy
oAaaWlrvE99TMmFaB1dUkBbHkMb2zlncPbvDljjdMRtWRV2TfCklpm/5f47RSERq
PWquf1ti3ZP8W8Bv2IgA7uz8GrMi0fXcVjnzB0xWleiFp5C9Rac97IaEefJAsSP1
GogqnUCAdRPZoQcBBHaAe9n2aq4vhmdz9vNnjlTj9xzjQEnftHDjfs8gMvMroyks
r8H7fqTJ8TN2nnpW10I5E0d9LxJyXlbZstyGD/wrCNIMOsXzUltSYIIJzjLS2Lay
qBrNJpquTHqdMJcC/GF6zLnvGHMncJ3fIxKPiR3B2/62Betk+7bsGyENre/GmUnM
rMZzBAKxK+Eiq5UiBubv3UlFpngmIDHLnsfzTEwpN+hs57FhKepgVwYUnkPsbYfy
Cv59IuBhteo8ftC6wlYTbKRqNpnDnus4qMa6YfNAA/ZwB3al0VkhIR/CU3GYz7lQ
yVNdwrfhsBJKKdaM4oH6WZ4N8/4Ge+wY85a8OvnXiqac4dZSxAWcJ9H7kAQXMNeA
qZlztWpj+kv/BX38OZk5jWBxOkGHHTu/XmzoJ1rG1mMwt3rMFhzoTiVZNcI0ubs9
j/Ea195hceGmLWiXdvs7w8djhhsqHYofccbswNCPrEQFAQUFirLuORGUwwVjGr8R
M2+Q1bJzAwNRJdvWopmrKE8SxM/nkrs9L1WEb2co4kLqwNcTFqBoUZC6qdzWepma
OYtkfysLTbOrbw0kFiC0t9X8YzATSYF9yALTUb/k8kLgCzodLpQHz11c+Wt/f4Vc
QP9TS05+/MqyYar4XgaKj7+96ksDNkb5ff1do24xPgA/k2fG43Bk3C3EIXguPwKF
dGYiCTYxnVaO95YwJ343RR5IVPGHWpPolla5TsBeowNyAHcO31ZjxwW+Ogqkfxm4
9iHFHN2o4hHIDucUCCbqD73S2uYYKZCAckDFfPo6GIR3bvqWoQixMl2l4WUIGzUH
N9+9X3wHvjXimBi4RSOxK/Sl3XFeFMHHL0lVnIBiirW0lnEJrUvMRRcRVoqb7lfa
sZnBtjePjLzp4Ik+KmtwJ4TIPPRw4Oe0B2bqrKW8OUd81E4D9TBSQiC9nnkA9PhA
6iYSAwBiJVGRwfOK32d1AohVRMHKVjyiYrzmtfGVMZbOwuz2LRh30zBElOcCd6tH
LUth5YpKTSP0ShnBu0cg6rQAM3IXXWCIBgPap88kv0yEfkLay546pf+sPtABwx+s
1jY9zJIi9IZfgds05g3O3nVhVQFNEumaHFFSR95B8Pj0xLj7uWAiaUCsFSnAu2GE
CzxRl6UdxjTSwmuHVnEjlZilAIKM36C3Sl95wAw+MhEOozGsWF4FIfV5Z91t1ZpG
3+vP0NOGgiSvILFQ4xDZBUNSFqmJPjvFjgQOKdvLHjZ2dpfkUQgFDeytTZHLrttK
JBKxjONTxC4R3ZYYcD+LcCiTSJQGNu108Lyw7L1v+X/cLhKk+JyngK5w9SpTHQX2
EGElSumWEU4TTH9thDjhWraaqyhtnRTY1drMdGQ2CF68RW/yq4uWqZsfDRd+f+Mx
Ej2PbAO+iEHb0SgTR+QfJzhu+ywooYEAmVNSj9tyqhtGMUmwiDvAC1emd9RGY3MQ
D1I7r0Yd3OoS0JrcAgss4uJXlHF7FdD4yGygYuc0LPo9nXB7aTC5JJY0ve090p4W
hFemJ0TS7QKyFUu4lGM5yKsgIVdliUqYjlnQ0hwvz7W65zItO6BnaxzUa7w6nwYj
GuTnJzY2FMdT66zPXywrXRGLEZeab0q2/D2RTRLRglRQXy9XT+105epqxH0h8kQM
tvCAu4qdLd9sTNqIbvUl2dGDhgI5w5jRos2rs9GEloJ/ZLtQqMubon7Xfk2zIFg6
YZ9eMZzwSLfOH/kPjhRfCVZw+obYz1HVYSZHczb36I0OQowLVjEjWENhnrxNoz5x
tx1whzchNk/AgNMrK5nAHaelKTiK1mIATmxt+nDHkGyHe/RBuJAxBpr+sIDlqgtb
yJuAmIFam3tdMqN2kmKwixE7S8IBaPflPA9FgCnqJPv6DCDT2yhbyDTbIpk4rca7
j2WzIUeuT9kXq79SArgQuGFEGBnG+BZZIcJ7VK9d0c8eJx9/0laQakSuTQLJ+JrA
mkKpkgkhEfKg75p7F/n8qAZ997/wGiV45y+qiz8HiI4oOFoalQDHr994kN1ZJBA7
+mZkj9T4UkClLT6Yp+0HYFa6XBP1WFJLhnsjlOJSp8Dnq1xDArwLXo8vK6u/0lVY
3yCNATZbYVeoB1AZ1YxID0b0zGrHmH+EeFYHyxZiDR8oC4HGOQpTafEwK/ME0W0Q
9jD+OgADiB31mmQ0EznjBAi/FsutXomvFjKbk7hz2Yk9x1Ikzyiwa4Wb6Ipvq5ph
zRYO5sBVmaIMsmrmhEaA8i8kViu1gn5I1HQiNhC5WaLxX/WqsMTzoUv8cjwCeUKo
Ma1aoVRAPXwDTA/zZq2t1plQ96njh+IMB4qH6WxsIVThJAfyPx2Jv8KoSqvdujwz
2Y3nPjnV0+y2PvZvAR+Mqkk6gLp5yLoYi4yuVh/XlitH9eCpyeQZuIzdHhWUdtRm
gJB7NjrU+kglv78He01Q5NmrEi0FxlfxuHK6M4KamafajPbOn7pi5ArNGwqkxFbD
6VeEsFMAWs5tvD7hrv/5aHCuGjAHRbHXuQbxQLeBYmP83mshK3uXY7q4Al1oSLhR
FFahCUXa+7Gzu9UwOpBY2TaKeWBlTNT6XK91Ve2UdklWCeaS+46Vv4OR9TxUNsV0
aRQXaJWkD61tig068F7Ek5N5+m2ReyXcsUYL05c8nbNHHABmYDaQTIMK1FvgFqh/
ji9XFQXRBg6Ee45S4vOeYuQ5AhJDzY5BkbkgNmRqsLrHJWWr4toMnCOew81g0zga
LyQ3HLhwMhBkYJLJES58EqUvtm3+XhRCA16n0mOsrAyzL2v/hn4XliKOA56M5Uw/
XV4e8HdrKLnVbd6Ki401uf7DDGpyTqAGLK7ariLYCYdYiPnCMV7v6fBEYYcBkXE9
phKs+xRhaa+RSmbuUBGxhK4aOVG1NDRstGdAB7lmM+QUE5FEQVcl7GBfKQKuMtoh
ohSDEA8BTpvOklwIkPHTuzW2Goypxt4I2UZJdqbMmh6W3/97EyQZ9GMkOI9fkhCq
bdukJWV3bO9tK2bYUPaEzMHtkmHSVolGLdrQ/Bw/4FEnMdvStZsH3JmLnYYH+WTW
ZoGQkh3o31Z5LO2qQsKb/NXlbQMXHJMtsmiYLPNATm9XqXcXaSZJNOdHzTzJzSRp
u9dMQz35syz1tgJxr7wNhLc4zDI2G4COwMZR378WqRxALbCcLumEk7qmK60Q9YPo
dnuJOE5vAZvy/n0GclsVYKWVgudy8wrzBeLt9obdFTPSMVhH0wRVytbq28CgVq+T
ATrwmhrGNGo0nwk827wtNGQXQsWQhukD5Yd0sB21L/Pp/WSxOsSIKwOpmHhfVPGF
ib/q9GYkma3wojaSB6df/HzchRGXbK9lDM9zgjIfhCqYAVX7ur+oZ89P4xBkzudL
b7QPvkrAYcxqbP96w5masdZCpJo9VNYn7n4EF+VMNfSuv2M//ERzXKI/PVAfX9Tu
dzRjzvjX6B+niwSvtsCUdC/WpPiEycirWEyxWws9rGqn+AxAc9ldMWOM09s6s56i
YKFEGkruEmnpeDNOFmavd0WgfOEN6RI7a5FxVKvekcF9rzyDcGXnAUM/QPqYOMP9
3SL8t3OEp/gGtHCmxGqymXtiyqASLLCy5nLD9tELGrbF8gbav+dFNT+I+sqT7urm
Ssl8zrkjLNDy6+JdxzGXsq4t0CUkNbe130XOIh2LCMyqxkLvug86XzkZE8UNF2GH
zDs7X0knGVjtfolBzepQfNGX7J293tVAQ8ab4UMQYUGCsxO0KDUMjJXiWuPPauJ+
1F03FIcbJgF16AzYQtCif5ehEbhI1V86v8f4s5zdGT4WREtcH1Vshj/c9mERb1Yl
Mh3YvTeRUzWi0UliOJ2wXXKt8GiDObwFubA9SOEha5EJwn7T8L5HPqW0YZlhrih4
VO1R30WYuceFHRgp2yCgagzyDSSuD5yCfjY87Xz3R5cRQoyXQJtF8gzI/ODN5BY7
+TjpnNG+u8DpGZeLv8724MlgmEqJ+oC9tvTbPnaAccsMpPl2AGqqh1kyAj0Ym0Gj
dkZhgzijAve6dIU7KUVpl8N9q7udiXdXvcO/Rkzrm4twM9WmEolhgQ7KGsXKwO7Z
YMpvHkC9ZNYqxdV0kMbVYuzsKX/hiQfaqiXnJRPqBNDzprOIkMkqZ+NAknlWvrjb
Nt+oL3Otua0OeayaGQC7/HWbcC01TNkOTpMigmZItvyvB9t/2apcJuUjdaygwCtV
AlOYnuWStFqrYLIX+z0nQe9StlOGgc9Qml5bBA3p1RLcf0V2/+q/ADc6omgaT2aU
c67kU3NwjLOp5nL1AQuk9s/XMwg+n5KpVjYGHNGucRbStTMiU6bicIf/C93h/qIn
d6V+dDeGKtX98gGQLvGEVyqYH5/VbT/6BoxVySxQsbOy/Da5XothGt3F+8340so2
aXh4bfz9sKHmHExudHshagFvLAF/ZzQsP4Jnp8LOv6g5psj7AYCTYxSw6QYK7MrN
XuQLiUFjDdmLTdb0GbZcnA5CjnscLClfkm47ABuLdwiCa0vL4p6oZDHsr9NkhdoA
RrGqNHKKom/azNQAOEXSdB9asnnnnGmAjqynd4QbIr5KhBYc6PUQWTd0rZHUZgwk
3kmOaxQy1nFEDLgwbcfrD0M6Ez1Hg9lp2XMiUPqX6NjJHzREJTU2ouWlKCVXEJ+k
VsAfYKRhBRg76tQ7BLAvZIS1hTazLvtksvlzChePTgIulL3M1SbulGQ5z4x/fPXy
4Rff7lF8YNENnBIR8LDGMzySXMAKPu63ATjYu87qGMWFwU9W+XFzxPpWpW91dMfb
u4edBvPWONPujhIswMhuDGS87xvGq6MPD0ddFyZyoTuMcrRo7omYkGMDHNiVvCbi
COfDS+bt1AloAsit8CfGxYw2qsb1CTnDfcvE2DmF/ZSZpf02Bt+LIpr13/9o6IQw
3zsmhJ6bB0cET8LZGNtlO8J8n3oplK+OiVe6qHXQMKA0oZsaMxI0wOMtQzglcAtm
8wlnwR6vq3TxcN7zzrhhET46IvZb3vTNn9soPkjFt4Qs78QWFgpC1UoFqZegawON
PKtl6aycsoPQQrWglLTWegb6sagIGFzdjcB/mOKjSvD1gDLuawL+zgZDC0Z7W7/6
t74xcEJtX34BJ92yE0khdJwzQx9WbSKMuHqoYP1NgBgvKtDLgoyRtiA12kGDoCVg
jOiu4SvurhXqhwS2fdChPfqIwfGsQXHyB6L9fYk2VnfUWtYIsbdT29Gc6eKQcXF5
SjusC7TaHrdRCxj++LCucTr9MUFwY0IS5NfQoT2Naeibg1Sl05mEF+ODb/olpPDX
5ObxswlL2us8wNeUb9BXxfKf7rupGADn99uuE1RycckIlQazMmYCkfRAHxilUwrF
/ZjoaiudiMRrwIoz07s/FM1OU+144NnfUkKh6Xh/Tglr8jFNGFEgOV6eMnPx8VFZ
XJMUiwV5Z8YGG3zp4Ejm/M4CEugJhJKpE0oJjD/ojlJ1eEkEzdcOo8jyUx5JOvzg
MeogcZFTMV49KJ+6Bx4aqmRR7DJ4+eE/6mGnOUVi5bxIeSqr0T6fI+Ts+IUttjhc
IWE6cMj7zL5gk+IJJOZevOkL6XGlt4IdD5WKYtvbQMF8sb/A2l2CkDyd/5+bWl9/
XpQYcD7L2Z8JOIo/zxtJuRTzK9DzdBd031mgmG7IMy0fxQmdpQDcLH1NieAoDcXe
IBtaggQnuNALo0/75rTmjwyQzJibAFBZ+9nKvNBdRjno2jSFr8S4YTjLYaUXaS5Z
j3tB/QxGiS/4bN/qpCqf6/Ccj4hUc5MBfczwATfZC9HyzjK2XjdMZM6JRj0wUv/U
oOdJJyOUlzKHXsWHA6VrCFPVa1eEUPZBvZ+momw57RY+cRc/SwDdTjubETu95aD7
emQpArdfqYsWLV9dE56yqc7V4az2l0nGT+G3lQg8sBTSFyS0Rx+moa2801S2BQdE
wiTchaunWGY19k0gkLFN0KBxMIVCsWHiMmB49AMkEPptnX2Ul7mLBtBYkH/1pZpZ
szeZRlKv5W88YEsJ3wjnLylZas8XBrhQK3zuHncy6VUZahVrvlDV8BMY0oZm4siy
vRNs1dDaeMfGawGVvw2ybzYXYHz/1nh+aq/eAW61o+2SySlJKa+5QwWhLACS/WyF
eokYlRCLy52MW6ht+F0svVbq9zMVDXvlmmVXJUDVvll17f8gE0gDRrhUqJ/iOhWZ
Ok6mFfoe70ZymQ8hmLAaS2TbEPRvd/xSco9tAb47ilD2W+YpqWDaLgvDAq6usnp0
2TQX4rHdPlPLP4QYzre1W73scoE9871YTWq+VNjXSOOX3Kx1E80D/Q7BRcUNE5nq
uY4yXUKqiVPLvy9znAp9lErh3HX4G/0TQ+1zBCyu11Ijiwri+truVqI+6c8k+ghE
rp/LOSjO0Zf3OETzj0mRRXD3Hve3kbs3n9bhD+RO78DRQ/M+oUzz8GDY7GrF5Dk/
iV5Lnraera+KCbnjulZfqdTB/EEyEA6GwtGxz68L0lRhzS3VLLhUy8vlVjndSNov
jSvVOku/08/gpExzCHpwsOmBgfekCbE1r4Dcekc+oUgejRf62ocp3dRWcIotenmA
1Iv9LIKt9fCWG5Hnvkh+huhUgLTEdNSDdJcKc2il8emXoWDFDxJlXFgmRKm8p+MQ
z83B8NFJPn91uZ2s159l1939jBj/Hs3wb/rnGK0546bGWj/kuWVsON5SzOu9tu6d
qk4o1Rngr/GzPY+NRXgzveOLkuHpUPYxxbjTAiHT00YPjqDZnj1ox7lSPYL/FvGs
IMnnDVpOdsV78TEhxx2re0NvXX9nqaOYxMY0fF5FTzWAU6++3mlFzZEZIb24un6i
ErUzAShFxPT9OcQ0+aEBHQ044uW6b5S2LECNgn7VDs8LmrZQnvtpOQiL0C1g7ESm
DSN3zd6Hfr2y5GkQXDqxE/v5Y3JU+0qfzczSG649HU5Qw166T/azgPH5hwz2I27m
83JfTtNY1XwdT0zQ+mVh3pNbHpByq8dVkEs1hoYg0W+7lMX8Tc5wIHV1n02kToMy
qDcAAPk5PDKDH8Kdw52ng9ifRaNAxcmu+V2hPGoarxnVKkniOwIN+r/AgM5tObCG
0H/qm5txh9f58OXmCCJpUwPRNhBagqNAS+Ko2eq8UknvN9kdSYoKb9i/9EYh8j3C
uLM3Nf4rcvZ9yg9jc1NJxvvMGBb/dAdU+t3dc1ex4bPGICK0Xw5p/u8feRyVtgrO
yQzAmUb8r5NP1u2VUVSY8c5VkCxJIuimcloRYIOZkdn+V8cN//m7LdQGh7P3MBJN
8r9yhKhmvkXkhn6GRdA9nlvsmP4bCClCPOkbsDwjVsACKwsdAq64afxcAEmW13We
zHLan739J8Ngl9cE/7soHyzNGIlbXmY4zKNIA4JrtWMunGMgix96cIzJMngXoaEd
68ArUTQHwGiSkNyuL7Kpgv1Xm7xnTnG1HI2lCY9CqN65aphqd5Mih+F6yVdS33Dw
swq9sXWw+dJzj1kF6Pq1kNqFwAgniMVOZIwgRedpoQo9+sJtVn2sqiBLSNzxhNv6
I0vckvvpK6zbZ9qREeXpQO+Hd2kFfiH7YuaJE4Ld4UKFtrJbF5R4ZSVBB/vPDmWC
ltUSgDffu4oXFXy+FvnUYqWh3SxaMlBZXmdf9RJqkL5S1rF0vjTBrZERindY4PX6
qiKK9iwMJ5CWY5oXcp8vQQYf5iSRGke/NlQ3SqwNqBRfobD4dIMMrduTj+N9Vuq3
xnpHa0pPVtq+oLkVjtFPQIjhVSquasTsHMEMZ2gbp/vYtW+mVMAC30Ctq5Pc100J
YrByg1D+6vSinwJcpoZ7rYlsYGpsVmnLm20Tf7FZZohx9hO4xvYXQXizqNuswm/7
X7Pdl68+LoO+FWHjj6TOcbNaQ5eQ2Ns/dq0RGzGeQazmUIPg+q6XtkI5TCJkatFa
euMvvDHNhGCy7DsdcOEI83ZVihYHqxHgBcMeOx7QwHrZnPWaq0g17DMhoh6t/sjj
OHSzxhmlsdoLX2vyDObnexFLk3owT/PRyroUFKvz1uN0F6ZPd/3QH5wqknQcqc+G
r4wqtINSUIazoQGSxsrx+9rgdIoX96D/x8vP+YCtX3er++yGRdWY1UcY2pH5TqAP
IUA8hl9IDQwFH8OyISIdl2sZW9ZMqCORyNOD+B+RlGUc5c8f1dmJ19kwttkqgmgn
N7J7cimmvFRgTBye/vFWahImNgMIquShPpN/Lhaai6M1Oi3e/rNKjuGf4DosUKGP
Inbj3kKIsRRSEE2wq+jS5N8Qxcr5xdRpKQCGRyyziRakRtYMkUX7yosY8m7q0NNy
tVhvPYrmXFfRa/5HqMU8rT+JsUeqwFLv7Uw7DV/hJQjq2hwKN473AvCTQCkxnJin
c10YIeETZbSIpEZHX8x3iZqcNvAYqRxVFyscc7XGZp1dnY4VYclqx5T79ARcv7/m
SkQQBZKbxfSGs1wKYWXhOUDD42EjaTKe1ekBAkN37dmcZfiIYRGRCJZP/4icdtWv
5ejO1+u1PbW5qMYjlYr24VzNQl+qENT1Fyf6bpZpipXHMsp+n3Mp6Z/rBz5in1Fs
uq73drt1q4lCIi9jkkvAxgXtBBE+gzGmFkGDkkELI/KGiPOh6b4HvgOdYgmkbUmk
qgapeAa8ux8tO1EtipHrQMRFfXE8j2WtTi9/lhPM04YwDLnThA6doYpGtF8oCd/C
ahklYNiwgjNoFVlgCtiIeDjasdiNmKPh4d3PxW8u7+vF+l3m2EM+Q4faO0YiTBbP
N0frCqnCFluOljP5UAH11PZonMsWpg7tLh2BWrYxIsYt84wjkFe/M4j9BXLOlBm4
Pz9wO2YIgHPm/4Ef8YcPfaLL96LUJQvkRbDAlQioQUyDKGqu8vg6fFB4fTJ70fkG
L2V8sR6W+YIrHZCsNtLAbsjX+7BUNFHsw/YHNzxHAFW94kTdsNp7sE5o4YViTP0o
G2bRLhLxfEpfD76qBUZMrOlI4Z0aD0pPMvVkl2pxloFHup2ie9GICH0xCSss+Gb1
CeHxvzB0qn3cyr75B2OJki0HLFxWEgQCWNHgLWSEbFI4IA+7ipY4C/oJLaXiD2HZ
/TMA3qY5Utcw5xsqogY3yXAz4zJJVhXp9adFMOiBZTyOSfQ0oTRfdu6+cCpUWuMZ
lKslJ+u3H8rVcJGj7rYoZKu8KZ/jzf/SE10VQ0s5WJvZ7X7RWySDfaul4EsrZrwY
KlA8uzR/vbHYk7CEpkhVYxQNjgrWUGWkz46yQ1XJgSxvn5ymjUZkctZ0mrlNJodm
3I4t1iF2O3PrJzg/AouXo/IrfZJ7k65NUfSQDu5RUfyXfZI5RcVsrCkF6TfO+f/k
swqPxEkvnFtQ6M7CirHZwClZEvw06jFH9GsoIS0QM7AKV+qNsku9aFYq1PgBZ7Ra
PeTgnvhCiMYvAuGOdUHHKDsnwbKIGlpyEygrkBl33VNpis517AVPR91F0FzS+v2U
7aZ9je8XptPTjZfCckmclWk0EkJfm5TjVT+IixXG836PYqhHdkYRzpDyzbwbPXbN
qiGCuataibHz9IDJeIS63F0XHPW0TRKXtifDaIHGvU07QKr0K7LxIxAaPPjYABVi
L3SBiKzpC4J4krN8/wP748UJ2Tm21dnl85aX74pF02MK82B+MdLtrOe1l2j3Jrx2
Cj9ZjP3FNPtZgK+VoDOezvPZgOYutDaL3HR3CnjnlUJbuXgzxUquJ3BxjnSKLdcx
IqZWWsAxc/QV9Cb9kQaPh/X4CENxVg272JSDcBmeSrVX9KCtYnCu6RUmTrEhsPQ7
wyuoaXGPKJSsNpAZCqPadzj5BpVIfipAzCSyboRp5qmr2ULmpd/Rfe90HEQsVLgL
xGwYfTUR6eyn3gt4aUbl2sTsqJ+AcTUD5Y1J4yYfUCbTms3wO98QJhqY2YQtCZEk
gjhvRdC/eEOGranLXfjzii4ydp/KTOIYmuzY59JLdCR84Sc2FBT1PbtgZ54InM2x
aSZNIJ6CwbIGD9wmG4J6t7wcj2ogzQhJcf237jLjWwBAFKtITihb8Cp9BzyE+OJm
ml3yqzErO0VW77iAtqMvgzUtIQkmPlsbwNghdX78nhwR4zupsxKfjQNQV8pG010c
iNiR3mRxfyRTec4/xMgBRHQH2ZNK8tqlZ1zZ+rvSG5imdjbEcXasGgNL0OR9vagX
koqXVFYOWYrHwucdST/1AFLnMw4w4hIqs4zs4siWAGlZSoNKHEvviqPboQscJDhQ
CqoVjtE3ookqkpdXFqSL8abBJjATWFGNBsL2kRkpvPfJw4eKESsWohpI60PmsScZ
5wAEY1lFyugPN1OWeFDm7KB0FC/XrwyPzQ9MmKG7pL8bFdGzRAeq3y+oTvOhw8ny
IpnFK3cFsmsW5YkgaUKZlrkUO2zGKD3WSKgcY50WkFgkLvT8pyHEvOd2sFCHIIm/
VZaFPN0sOd+ZRLCTlZaXtkT08n9BxnJM97/mHH95HSmi7URbtlsyJR/S0xrz8Y4K
upQKshB0KrJU6dTnWZDy7PsMyrYuihuk1U/otsG9Vsy14Y8IGg6OHDKwfP4WbFkz
6j0NuLTAf9Vek7pjowZaXocvOgo1ngdNuJ23TeRyZy76fV5DbXnMZ0Y1RX77wYfB
r6L3Syp4spDEJUNOr4PYx6v1lROMOP1B2ZjDP2sIoZSExaX+6o6ctxokJjpGJfvD
46BnWV3Nu5NipLFvrrd8OZjpc8hRMjQZa7B1tJZMD2507zwf9E5LfG7pEDqJziHp
hpoffyrh90cExsuhPuE8f834o0PDXmRFbn0am32e3n/PlSyDC0ynspSdqb8by2zh
dmfBdNYlrhb1xWUf8bJSv40DZJDav7ViC0MN3rSi0x81YrnAPRQCEGcPY2sjlCZ1
fcQehrRRsE3L6ffvLc0xPcqCKKlpPSXtziJD5v7uNwXimCOmGL2h77nstv1DSvm+
f1yepX1A8KLeicNK+PpEQ6r8eIq1iSNq8TER4+sXwdzbsaVpryOvtGz5RsYrFDNj
04Vm0NUz2lqdlvw5C9dUqXafBqnt4B1cUqPD8P6QbWkTZwQHGzLTLuTDCJ9PZpMa
PjL0vtZTP6Lp2T0dZNcB39qGjvGeBBPFfWERs7DKEJP9sRfYLeBtCPPjKge0lhqZ
GeUyzY03t+mIQWoN/OvJVvxlhFXGe7jNyCbKpfvA8rC+jBL5emWmhRUyjYY3hoHk
b7pIdiofELdgY3mx9h38ndjBcFVC2Zc3FIZ2Rsj6gf8nxAMb+b4rn6EER4L0khoL
MCtylp6T6k7CQI4FaMabaCCFcbe1bJRxQXUdH2noTt0w+cDUTTLOOXogT+so9w93
N5LWxjTz11x6aCzUAZsH3Cu4hCWenXInnIhrpGYp1zBL165Dz2Ip2CHfomALqXTs
1/wCx0Zo2FqsGg11y1LcAcXa6b2IBZKjU4Mp1apS7u2CGZ5273GuyhTKjzeJuTxx
/OmsDwbMrm3Bekwqe4aZ2nxfl0bVW9oyhv674prhy0CU5zvQUui7o5EBRxmgybni
DJnAFEUIQeqqezG8oEX8JvYsya8u66rNKy9lVgZ+mAWK31fEyUo/MJFj+RjNThTA
n4PNbeOwbG4bI86i6wWUw0GauL/4AHr0d4KOpD2FRcHcdrahZx5028SxZjrYeoqq
YlylbkbJ8PQ/c4s++BknF2Iqwtpzqm1J2A1X/xpRMPWmG6q9TX7QZOOCLBStQAfR
pMQweqV3ybbJfRvvbM0AeopLMyH3aZUaVdTGriotNVZucQdvPcnIFq+pmch4ssHw
9Bwj3HlJlKbzFE9aiSZx2zdBHKly9E1ubcMR0XFhmSK/SLvaXfg+3dDXss0w59V3
iwqB2NG0Ok3+wJLjQFmymFMCHJVX4EVl3gmnCthWkFD2IDClZQo3rRZNFTkBpGYf
pLN7b8IRnGt8hhy4M6AyYDJYSAPI/vuAx4BrPPGr+mlKkEj8xk61mjTZKi66e6Xy
xt9mHwoC7N7tX9t/N235q/UTdsc4V4sUuiX+rMoVJtaGMR84WGpEAsGN3tug6DDf
AiOnMzVOX+h3T/CVQtKW+AyIntyOS+pscZ6Kpu68+LJnmMvfC6RKruDNPeHn5bXL
aHJydUaFsxHIZr9O0gi4raz3IbYIuwNPpDv0NSTXB5kJwhHWSZU1yR7EAXbeYjG9
TglP5vWdxLB6VmtYqLy88b0wtFU3IefrZwnWT8qd7mNQJmybuTNueVugS5gGYKD3
dlY1+KspLhTnx10tsY3vCm0juox/Jp06m77C0gyeEv328DI/VeU+xFNMxDKneYpK
/fK0GkI8q8Y7UFbQvY+YAKx1/axjffN+RG3qH0STZAaYDB3TVBgaONH+GQQi+Kuh
zFNENeSt8Ygrfqx10k9z3cZgfWFUDdwccjyarngcuvVEaZWJrlBhoTT6Foqr621Z
ghh3a65WhFR//GSxQftlNLypZ1LUCcJaq+yDQK38UGC6OCRF1E5Bb+5cy4/ryvFK
EAEBdivPixeHE8RowMHVjw96doG5QhSf9Bb3/CJCIjKz4JqPnwZCt0TZYzdMzKDS
fYjuJZopsQaAXxKUTCFw180of6OjQDyH61Cxw4XS71APw9iiC0Pzuy4+8XMOJrQk
GxUfF8ivxiMmXTL4zVwW6+R1cg2AQ6ah2erq8g7RuDVFCuPuKERiCbGBOCob9U7H
yIV29xomDrKyj9GQqSUJR224QxE3729ctmkxxar9xNRJBzhv37Fuivo94yurnJQZ
ijkwQfp6eWG/VccyCLa4W4n2t5ZHEWQyX6Z4Bq1J84KJKYigVqujZ4yiWpVISQGc
C5bJl0O7+f1mCP8kfu2s5Z0ZWESht5HpbxRw2rJX8t1+Rnc72U9uLL8ZVkxbRviM
fZgonA+jBKNUb36drYn0l/f1w8Cd0lLiJUoUtuPPtU+29XJSB8Lz2teQTRLBxRt8
obMGRMg0Cnj+8bEQNnnxHGi+hDCBbyFSKxRoN/iRpAlgle1Wn38sNGUhZ1NLXN8i
OHpw/65m65SGyBKpCfWjFRqc2qcSZHk38beWNwXhTCzpvoxsX6M9wV12hKxnXwiZ
pcP8rQhq+JKgddpVgGOhzd0dl/xZys+klLz1IspCRpVQB78jF7QlaK4YQ4V5raf0
9eJsXAKDb3f7pGAva+KCOwOlLyqhVKGvuLzt3uoVcmIDqU5+jsnRg+A57eDSEh1h
esNCMKoX2EbVpqOzmlMWfqAkS3UI+eXO3BqYYGJpRr/TewDWt3p0Ilvqq9f4Nmz9
ALjUu1ZCDqMATg5SK2uY1QgbqJxFAsMZxUReLhDMXNzrfqbkmWdWbBwEsc6I3uue
rDXJ4GZMTwzRESn6yCJwR/6ZpTxn1HTltcLBlmPbVNqLgf7gB/kQdxCpep1qgkHs
wDrA1aOYs0JfLLA3X5hoQtoZ0ks7P2JGRf1okYQvQzOI56m/5fxAKB+TW/0VId0P
xuiqlGY3f8PuYrLB2UXAit2X3zLK1IYMqJYkx/rEamqAOBWNmWzOMA/GKZc6OtdZ
DiIS9T5P7Xvh4Zg5GPSfyIjut9Pg7v0JzY79cKIpWjUs2iozxw6dl98D2xLxWx4L
CUhavvI82P8QzKiuxkz7Wh/DgMGwg63JLx0amwyGyOuLowGeuW33JMzsmY0cEQRQ
AnG+Dp/rBCgNzpmafSZNEo9HHxZdzijbduma2wHeGTrW7dtxCFAZcTA3mtxyRQGh
rarRCbmALB28++u3/8SwNdprxDa5kqAAwi0TI1G9RMCmvCsGaxhQ7gB568BxD6db
QAsYTavHx6WrU+8XX8w83ujxPuPeYDx+VYdBQzc/0ObKS5v1vLQGtp9rmWiZUtM2
MFpuN1hNVWsn8idG3m51tlwZ+20/t4206sVj1Wy4D+0pThM4Iw3PoX64Jg+ghXDp
8STcZ9hLpS8DcP0t9QVe21A6ScrDvrqTH2L4kZiTDFAddVuYW1PtWGNsNZYRK7cR
8g9Rc5+uQC5UgRw6yOiDpKt3yRszgGrLueYSN9xx5q+UsdgED4PxolrHc3H4l81h
iJRk0KgDZ+4VlrJtQsSSHgTDogD6jiImsaGjGmOP97/vhxpEGjRMZ/WW77q81xPj
W0tgcXXSNvqiVtDCjnv4LXjejk7WX/ggYFukKVtsAHmmJofs3ZtIsxGbKmL+k/s6
udZIeHR/Jo5+RGZ4zdNHUguNPhRADqOI3uBze/Xa++iqkhL067Vpi5et2pf5RbpD
W7Z5XpnrN4VBOI27DGXzbgP+caZZ3AtYgfug3/w1XBPVpkAdSov7E7rr9+O6ABAk
See550Z2hXnyGf05hxaqHcmb0MB/u/D7Ef5eLEiPR+MslbC60Mv2NBTdCfEGWk/t
g/IxjRz/VnHkvN9XA5FFffA0FYujnLmND69dC0K6XxYBnXiqNO0n0trTGKOPWNAz
4pQpOmwkEsKt2lTqkufc+MEuZXVlDlGoiizL7DgtI6O84Vv4Yddx0T0LGFCB8OGE
Pzou3ssfjtOMhIjnBNNqsm4H5ltxaUUnfHbAsvtTwQWtkz5i+MnUy5pub1+mgx5R
3Dv87i17RqKeWMmCwxwZ2z1WRLNrpJ5/60gJTibYTBtEaj02RLrhkIVJPteQPIIJ
FUJxxOTeippIv0JTlH4YtY//y2iStGkrcJ5pM9/Sn1HCbtO5m9NZHR7cPWW/AKLP
ZA0VeySL5b90dQ2eV9sXguR1jV1eG2ZPLqhvcu1FdcTjNPPJaLwcUgmh8krucNWq
gVgIMb2GS3k1bixrsTaAx3MgOhsydvC+kA4FafMq7UHb5eomoQRr47SY5bXkyWrd
y+ThL4sDRNLMIOxOpbRocV4revhxdYo9yks9rzxW3lvW2Yjl2qz71/W3oHuiQR1B
7owxoGl6Rn3Ggg+TbhTZaC04T2wRXeHVqaZglQhKPMjhBmf9Z4YtWqQ5HWK35d8M
bV2dgbVelnnEzulRamvHXfCLnCKH+9S83U/iMRc7YYDNRlhxzOtuYJWzn5kucPQJ
j8LXCcndfic6ADtDp+ZDUt+hSYfiXO78v1C0iuvl5hQebft+7R1lGBeTtcefgkx0
24y3grj/wVRiwMBt8vJilO2YRrpkugnXTMt/wtKpw4HN4f4TuvwLcJVEFgwT8Ckx
c/cn7ozMcxqfA2Rb35Y5QXmwsY56458ZZlrXJH63H5QVbLf3QWuyOMofhBKDPw4W
aXvttKaCi5sVaRBNO1Viafhtj9mEhYokACAAI97iJuVXntEdooKa5VfQDYpK+vxo
znd/I65PkW24uD4KQfgexSWiFRCdkOM/PMrQewn9qotVcjyevZd6OAoUtkDNHhVN
l+0PT9wU8XYCT/Ss4mdtT23Py+7c6qNRudjQl5qE9Cz8RUcpQU9ER1rIF8sVu4QQ
P6alzstfD5HyK4jDa26OzCS83ZjAG+lg8a/xvW1fD+yncKCx+TwxwaTeA6A7DMbd
w3nRZoqU+yK5Cv4kCE3oQM7OBn2K9pk3BHpL6qO1acJfvqMhQnDuutApYxyhjvDZ
Xb4sE4W8KKSn3oqAicz3mgS9GyW/NVrd2K3cTzLN/JIZKS/CqcidsFcF9QA/t9cz
CzdeK4c6ldYsV6rgpVLN6ojFTbXqmHomTJUA/ES+tQOz0Mvjy61OOGQnxnubJbx6
Lg2/i9WPihjnFo3BJoLFs3EO0jk/z98AWoWokR3WOxy4goejpcdhVYlHpINm3JQ+
Acidtjvw7iFvL9+h8OjXy6NejXmrjW6Xer50dsbSFmF2jRwmxoLsirMopwzAKO6K
U0KpREObPvwqDVQMvaYux+F++X6PN1rq0OZP/CSe8k323Gr65NfnJYNK6bmPA+lQ
JKyom34nyIfhDQSfnA9NZN/nLmluhScA8YPr6AZFY+h6hWMl2dfPvd6Ifp3n4kwd
l1nEiZA4XfHufpBxU33VOU45H6rnxL0XYXtB0fkBHtTE4toByHg+t0VyoyGd+whB
qKa0xAkHwxcFzTw81B6RBBphVayc4lGmmn6r/DAiR0DC5V9oyVuRQ1SLIz4RZg2u
/QPcB5ZUcJVCGmNBAiMBxdJWX+b02uV31YmJxdC3hetX3i3c05kxWKIXeBE9XTcu
3Nfs88+TTd9eMoITmBTFa9T4i7wIis0f5KB7OrHeNSfUPNtQP/7ucB+VsfwVtcrn
qtvCSvnQ0XFOFnmPjLYNQI7Rao7wfD0qYR1JX9Rv10w7vS8Ujrwpr01mVTvErwAO
0uRIEy8dtjTvIYIdlpCoUqD4D5/OuPgWDyiBZtb3ciZVXyjZsTWrBGODXhRXkXOW
UiMUyrjEriTecb27Kfqx90AywzFvE2pG4imDrJxOfsgbBTVnXwDQVUxRl7jcMRtj
NePz53GdymSAFTKdIRgEskxdtsXWOrBRx7cY1f0pkdqf3mCirxWiH3Wk5/blFEHb
rmKyt8mlEKIIyd2hmeeuDeCuoHPcJp2BIiZj91sxWvFfBkXQL7RWEywRVkCD/oKm
PUZAnt68VvLhLw0mWAvbzXIFFl4ev4a2MGfaOw0kJFOCK1YnC5ELbml2kXjqE+Vn
qXJDF06JxyYzvWOfilHXZYjWnhgTxh3Y/5m/IjJ8P1SeS6gEGmCPcVgBBy3uinJu
ElrzfOvWu7B68gIy0iMNzs2sWa9O2pAbHwmQf7Of4GIwL1BIwnOObhmQPgpAhNNw
E1CCTUyewqAiB1xIlYQqUfvb3xq+dNHVkxVMLCAofHpVi+7q8wAg4eDlOZKPWBtL
/0iGXK/ZmOgtuKWi5nxxnmhlEnf7aztegXZh7HsAzlGsIg9Stz2f4bUdp3gVHXIe
7QGtXc53XMKxoQQPjzDPOpuCHC/ES20Hp671ODS+xoP0QmumRhEqBrWoc92Cw0TV
EV8Jy8RYZ4FuLRUqEw6GpNCpB1+lsNfuRBx4PMttCLIdKrT1W5TTfXREUr5KkU3T
v156udHOwwe6Wmkdj430I4VJ+V3+zLE/EwRiOWAzElc5UgBiYSfLIkmkMk/jziwA
WgBzD7QrNfumqJfwHYwk6HxXtDZr0wZgEw+o594FzwSZW1Bo0BZM2iO9ioaj+Ncr
DtZhdt315cfNPfh6DH/sVDd7hjPnECx4QEux1zjThzA6eAQB7bUr0jirTINbTJ6m
xcFdD6iLYsDW5FrrfdoL+vnpEB3TddRv+nTHxOeLDZcVyr4MdUo+Y1N4srYlXVkT
3hhld/bJJVjFdXiBiwDynhH9SDC5p37+PnXioF6i2/RCkWu6lkTYAE/sgb6DUA0w
7zJ74XQaUdKsol9wJ/J3v8Wn2dkZDjOL232BQ3P9rnW+B3vtrkE/JzRepk3CT60+
soGkM6gArjn6Hd/V5UQGsiw/dU/qr2eCUA8eRnauPvqc8g22f9ByML27OkFvwhiF
Lir6hRUg0qz3DKsNk0f5vpQGwHQNnpUT7blrO1BHxWevloLbKgx+mI14oRhGgeIn
j7djM6XztWt+FJCIM7Jp5wnIh967tzWuSUsA/DJHabbgQ6gQfYSvH7xwWKUqW0tw
1RM7znnlBLSCd0Km2zG6GpIdY60sF6x+RWIW/4OFaFzlSSYIKMpiZO6SwhTMZiMh
/OMPlqdi1y4ebFo6nYh6fhJ4SrCqdp9c6Q9oMgvZ2SWG+us6cQTwV8muzoz03K8z
0KzV5ZI84KC0cIaWD0N63IHbSczD1NTNUP9XNQMhnUiOOfvcYhagONLReOZ/OwcZ
2L6x0xyjsurv1n4yF4cmfXmeYz+dxFNUUk7PyNF2ALcwIitPLvCUH+SY+QGwLDjh
EGkjthEwnqHBrXJyljbo1+cSMDuKC25cBWDPg9dnTuzbq5WgWvIIwUVpi7I3ficL
hSAD7L2CvnAx9AmEiSdjiFUVDcXy5kTEsLHM25YOpDzp9wMRVU1SsLKZ/Ho5Bgjf
GkdeVxKRsaFQStWcIMqBRkkplJOh//KS5pzn0VqFt+eRVgk7Lnbg9tgNbLaHKmbg
MqKWH6PQ3TssgG/ze0XK51aFG6wY1Dnz64GZmCPMFCwK3YQBdzLlXdqxGhMyB+x3
LHclZA4OzH5TgBDslKC/FwRlpqfgh7iSyMeS7aIIB3xk0+wuqUPBWeDc76VCGSLP
LGoYUQ6kYILgpgxIuS416XbK/qJ/hrjOuajpeP5sxL7ozmgGW+mFho+cqEUuysZE
BtAN1wo/X6BdzDmsBHL7DDWI0w6qID0bBOGd24plRRUy0ClRfWtErX49UG3a4ySQ
xuqH0D0OUilAxhSb5owXoHSqHG+14z4x3+Mx1/pI5yXAkmMCbD1kX42DffzqlfL6
1UVqGEUSnx1dRSo/16yW9VOhdv4Z2DREBtVJwEnM2AnmimZPh9i6u4ayRYqNg7ZS
vGl15rWiETnw9tJovRNkbl9AVFMNWttpCq9akSECIVp6yTDAjA1MNR4TzsPWiiDc
xEaYGGckTPmG1787Hb5F+rhYY7Ce5Whtowx4fHEzBDv7qHSt+MZlB6YQB6/HobI8
vFZ1PSLwnlqEAZ5ONEoS7pE7DtXPlGOB0gyd+ifNVPWwVK1zgU5Kj0UMpJ0Qjq2d
0/uXe//y3aEKjqprjY8kC3sk3BFJ5lejFcTdD5T6j4yXwXnZDpZQPumXQRTLV7Kg
frhiR2sIWtvRinp6b4TlpkS9EBUXsrfVvkzJRBHtfqk4zG7kFBBjAAtxJ3aJpYzW
wJTr0dq/HEhvF/2di7kU/XpgXy9ucTDWRfmU0PTaBXkUnlQDk4jM/F5G7hKOhwob
qOPuZveOOQtsOoYKB/CuVAmpa12Qadog3grHjQ2JxpQ0jwv3dN7x+FXMJ2/7GQtt
wFu+drs7TEHwIi4G4qh2K+aHNpv7jb+6yn4qROJWPNprd34J37hlFy9szWLZJNNV
qL9PmDHbPfpyXniNeaDAaJfCyjqVq/0ke5DrLh711rHIYvbUJW+9xzVbLHJe6xfR
WZXoo9EL/VdCkiB3JdWhUqqKaQ0As5anzHrihBDaMC5dvsjNyhtuKW0H2DkbhaY7
Wib+HX8rLmozqSYG8BgEpx3Bvo1MHObMNGBhYriU6Xz2Y4bsybU4bKUV9NbXKvc6
DefHiGjChKVGcK6VnesXGUBxT+kHNjP04Ga/isijWErhEb6GA8ey6H7dqk5De2rt
BMN+rEZeUu9LKlmxets3ZAkPzyixaiAOgJPSHQC3Rd6FRy8oTolAbR5P+4i7qEOW
XuQlx4kV0J8muXAy0qvnNnvqBt+HY/BzXVBHzoq8Pyg8xBXCjB7FPT+jZyyFxbLX
0BfqMYbqCKH0pf3wKpD5OuVAXwtOehE77oV4+SOl+Wp7oci4vZyFy/KBEwg6jqMj
NYkqbNcrxcjkeL+KJBbhP1bCyAHpxcfIkty4E1uVXTp+9thl+y/z4UXZO6R/zTeI
MxDQ0IbPazALSMPx6tptoo6tvvxPGUUjChygnYKxcXW/bz3f3fib+VRp9A0L1ZPO
BEkpcXmiXdk38Z6yPLL05gw4YwzkZrhSiBjC11yFv5or7loepCgYzLJTQAUMj5E/

`pragma protect end_protected

��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���X��f;��on�# ���5"0 �T�PL7T�0����Ǿ*�Յ�'x���!�����*��w���0`>���M�I��M���M�At�YY?��w�/��
��D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��Ěכ_�fK[��Q�AU[�MQ���;�g0t��=#b�ػ���p"�敘�n�����o���{�N��E�lW��f����
]���+>w�d
�KY�7Y#0	
+��ʩ����=��#�r$Ȍ��!��s�U��oW!����JE����zd۳«�F���,��%%��
��[�9��{Jw���܃ҏ	�~�-���'��,��Y�&��T�T���Paf�Ox�v"G���S���2�@�}��&m.���$��ꎖ$Cݧ�z��!�XnUf�(�0
�_O�Z���y�n��7WG�Y1[���Qe�]p��u�1�(��9������S���`+��F�/vu7)4G�\Dj��R��ȴ��{���'=&J,�n-�L|ċX�(9�_��*/�{KYП[�,K�9��W���o�H0��Em�����o;z��u�\�d�Ou�����{4��r�j�Y���.6s�0�i=���o ������:?(c#�L��s]C�UA3q�e�����o�%.�^���T7�An��. a���m��D8���9�j��B�5��mѨ���i���dcD�`�Z[,�"x��m%��5�6�l3�-y]�� TqX�m��摪����>�Ub2�w{YW�(|�}���(H`o�}������*'ڑ�8_�f��e�ڦ�`����C�d�4��+������xG�h�k�1��� k=N�q'[�U�ɒ��5x��H�るQ|_��|W�#�^1Ӊt��׈�a�ݘ�[᷾��W�e
a�9ٜ3�`l5ګ
^���ϓ{��L|l
���H����%k��L~�_�6-W)&�h�[���i�F�X��b*��{�9;۷�p�x�R�,��<`1��^FU]6���[;)]E�F	 �)�Y_;@��)���3�s��~sL��yf4t �_o,G����Kh���k�Tc�ص���W�ϕ���N������]�5C��-�Cšd�� ߗ�x�<;�ڪR',>��k~�A�ұn�Ǆ-��S�������+���M��>�Ԁ
���	�B�K�_��j��Pʘ�v�E
�W���z2AO�rq�HT߯�F�Yv��ZP�9�����+b����^�a��.��,l&Y����G�vn�o �R��wvu��$���Q�O�rqO���t�DNP��fU�Ϣ�m��ȁ�@O�빠N	n'rr-�bL�+*t9Tx���hV9�N����5d�^��Rf�D��[�O�p��L��f���AՑ٩C-���:�#�e�H��'BP�^�m�1�i��g�=-�otx�e��]s��ԩU�RP+n_�r_�FG� �b)Zn����Y������e�n�1����\��fT�sE�ͬ繳�O��Rya�s�m*^޺��L���}�1��������4�o�>-�J���t�����H��۫�q�{*�K���ų�YZC�Z_[/�K6�AQ���Ϯ;aM������g]ޠÚ�B���͆�x��C�D�~����iUr�a:�.�<�%D�ٵB�%Z�-�
�BI�8T��u[;��i?�t.���A'$T�];"og�ǻ�eN�G�(vYA��B�*�%`8��q7���i�ۛ#�]�.J��^���dK��j#$U�����쓋���*$ȥq��cDB湛+���f���
g<P�Wg��C�HĠ���ܞ�]�O΍X$�5]�<!'�Hq�R�� v Wn�4G��#B=�cƟ{:��⣙Xg�+��ڵ2��x�W�V�(��Bpz���[��r�d���9V�ّ��:~�Q�w`^8Ҋ�F,I^ٴH� )�E������A�I ��4u*dQ��>_�CB�	yU�G���N�n��aSx�6��3�be Ǯ���-&��2| �
D(�\E2zq ����ɸ�*�'
Ċh�;h��d�ѰsH0��%W�8��/y���T�d�
���q�)���>?!�241�\�D��^A�V^ε�Nj��Og�
o&��J�]��MlX/#.�^�b�x���4e��x5�/���3�x�^�w������������=�E������Mv��8G��!̯�?
]/331C��_i�$m4<��=,#�Xv���O��h�
��TO>A�o.�p�6P��޴\�j�il�08��'�3ހڢ�(͟�V౼����IS����[nW�	���W~��V5J-:��'�*s�:8�
�԰�?4(&�<��4B���b�[&��M�(�Q����WU�E|��;� $14+eɻI�πJ��m�9XU���Z�)dm\>Aj������c�EE�+���vm��ڝ�P��+�uǆ5}r͋�#�y��.T%�=�8G	�C�<�ΉNK��c�3����n{M�uH�5?7��Nob�k��,������M�G����c�\����l(6p�fR06����-���v����k0�{����E7��jn��)�0��?�i�,k�U�Տ�d����G��9�,k�IB/�A�HH��{[!*���x��ty0b:)��ft�(�*wQ�*�c�30Q�1���^+�f�h3Է�P+�)]K��b�jTZ
�
��KF�1����p�zƨߞ��
�)@a1��͇���S_�/��m�S������)<����
8����o�����c�E�IH �����zO��.0\�8 ��^`̫�64���N�d_��z|�;�m9��/�E���8@	�D ����6�dinA��Q�a,%��	��X*���[���w:5�A��1�n�L_Y�f㿑[�q��9� �9�
��r[�'N��d<t�D:ܟy��i϶�I2��l�R������ �� �(��,B`��m���*�h�tb�f2u�T�=c����`�P�\(����+�I'��+y�nK�������%���0b�a
WUWU�s�'�[^H��R�<�Ӗ�WC��Q�� �΁AVcª��~���3Ri�6W��eH�*�y��,q9����RN�T�m�ɅS�T��oN{�L@�x��ӓp>"߄�OXW�^��C�g���d^�)��Dǹ�]~���_�[\	ֆ�o��c��@�NM7= &~\#Z��U�c�y��ܗ3:�y<�fN$�k���'W��� H2�@~���P| �k��ȋ�6�#�[��)׎�!�M�(o�.�˷�CbD���J�,���9�u���
_��*B&D�X�P������ nO=�7��a��T�3)bc�֋7��������7]����X7[<wD'c1�35N�P�y]��?���H�� �i��p(J�ԏ��X���5�;�Gs���4��&�f	��a�l�,�������$��ߠ�#	�M?8w�Kh�B�Y�б��(�(b_Qj��x��&s�1�ܐu����K�r�{��̓L�9�/=L=O�h� �^���s���.ǣRhh�i� ^�;7��ː�|œx����ÛX-�����^Ʌ(��1JQ��+��ȏ�q~��ĽD�ue��C�����%z���V�ڃ���c*�> P�&�
6�ƥ/a�s��L����'TC�R�͌�C8��V����P{/�v&o�"�j�@.Ƞ��]�*�m���"�)�!ڃ<)a����EپݛH��Ut�sqa��-��pr�7�w;��K���Q�P�o8n&R�2�������J!��܁��G��D_�Mځ���F6�$r�\���6���� %�mܖ�X+T�����ħ��W���C�d�	��4���I1YJ��8!�?yQ%��E�3�;������K,g$6�B��Ե�Qv�+�F�Y�n;�-nu�j]��ê>�sy	L�d�s5b��1�������:{��8/\�Y0�O^�M�)��>nw�� ݰӧ	�-/}E�k��Ӫ���Xo�������W=9a��T���e�N��MH�m�Q�������Q=��Lu����A􈇥����� ��Q/����H��G�%�f�U�WblO=�KPD�t&<M�V(eȡ4��<״��>�(��%\0���W�F�h��l`X_�byh�jP�I)�ߴ���rf�tK
=*9��e%1�d2C���V�9S�,��o-_��_$E��������V7%�?h|Ŭ�Ə�;��.ZvTi6izf��D%O�⤫���p�n����ݳ��@�?_>�Ox1�w����H
>��;x���tn6��8�\����;P����t9�����f/F8�?yh��nt.6U8������	��(f��DH<�]�3�������w����Wh��1::�� D,��\2I�3���:ߧ�ވ���ݴ�p(��@����X��!�~P�[h) j�U��k����`/lٮ�A�1��+���
ȗX�(�v�%����,R��f���X\�O>�g��|��J2�aYM�ND߉ySJM�M�����$4�_�-T#19Sb���)��j�`�5���ctH�����B�S�����]��x�H���w�!�جF\�a�7 2���9�:<�7����B�m�8 �0�{���L�TLՑV߰M�zו�������s��e'��8�B�Ӛ|��'nn5EY���B*\I@���S����Ԩb��U��^�G����$��=H)2f�ȥ�!��ս̗��1���y���l�(-�~���>զ���H�mI��AȜ���}^JƦf�hr�k �]@�O�VWv����v��ל�C�<6��7�d�Q
��i�Z�/�6>�O7N�m�����r�˿]�&��������T��	֫��;�)M���VuC.�g9��@5s*E��Vj g��w����I�o��:�2Bz��y��R�mZ�cEB�*}F٘������]ݪe(�� E	2ǲ�Ҟ�	���v@g�w${ׇ岼��+�O�ⷥ�!�����G���B��B�sl�&i���B��04�/���I�P�	6����[°a6�fQ�n���e�n3��դ���H�p�J���G�)V|:�NGnC��S�:�!N��	�Sŋ��vD��x��:��Nn�'Fq�>�h�d�<+����$)s?NG��-?+m9K�W����D��6C{�w�M��w�JB�udV���I�گ(1슩��6��|�4�Iz%������/�P��?�C=�u
�4V*C��!oD*���W�?ܖ�����mԅ+ܦ�m�C{%�dB�>v�8{��^5
wudR}a�����͠1᥇T"|�NWQCe7A����K�����B~A%#�
�gRhQ3�	d�I�M�Ub��DG��ފ��ЛX��!�e��b���i��LZD.�f�w������|
�@�hB�C8�{��-{�{l�]��
@�w�(��N�;�������U4� ��Ba���
�i̽W�����3\5��@dMd5��L�D�Jh�_j[��C���e$Ĕ��Lh1nn������-��|Mݴl����Q��/o�ď7���LG�S�k��+)p�X�Wt�³	�I��>�A���	lS�}����P�m�ٞ�˪l_Mi���A�~��ûK> -D���T��2���.f�W �O���B�`CS�I/�nȡp����>s{1.��9&%�囨]<���{+ʖ�����9+�!��p�O7^|�r��/���(���Q�ïI&Z+�ܪ�E �������[Wk��I��M�6��1�n��G���b� >c�̟ܖN��ޏ!�i2�u�*�L�Rym*|I�0���;�����6C��~W�/g�^�2��v��]�Hѽ���ퟸh�\�dѺ��Vq�9�Q�/ 	V�C:,.�;@I=%S�_U�x�`),{�K�f�@|h,j|}7�zU4��$�P�F7�.���l���CR���>�ݞ��;��t�N,���<�Q@�ZOS�l��_�$4i�L愖וې���ES��`7����PQf�� �|�)��5���]^U&8�4�AM�VE;��U���i�e�0�����`/aC,#�k�����e��K�x
xa.��O�7ox֠"�N�`��7SF�%�]ޝ����nT��7<�vۈAJ��l1u �_����'0[����E��D�n��5W8�c�Y?`�J�܃�K��aP�"�:���|�����'k�X���B������@���K��V�^A͉�� t4�]Y�?Fѵ��k�	~��㑶��?IC�h�TT�#��D���[�y:�m-(�;AkA0Ŗ����A�b��&�^>x����0���յy�.8y�f�@�)E�.t>���W�Z��2�sI���?
6���b��:�cM���%��IX���F����q�QLiUJq�@:�ھ*j\����!���遀qD�YhJ*���$����5X�MY,�z� 9�У�>f���C��
@��oc,��iׁ�k$ܰ�Y�\�\��Р���1#�CkC��
r��|����q�y���gQ� cr��w7�N�b�i�z���ۺfe b�KI�t�����?7_> �L�<&\X�2��LÀ�1{7c��L�.�W8l8��BY��s�6����B;>�)�@�8�q�Q q!%QČ����;�;�|8�a?4 ��1��NMI���z� ���U��(�9C9^��β㻤/�ԍ_c>v^�I���:8�2���Oj�y�+�ƛ�c綥���0��(��opڕ�#���� bJ����#��	��.>/�=�����~.\f�N3�ba0��ÿ<l�=<���*�T�\�W�A{��c�o�W]ba�h#�@b�-� ���/�y{D��ă�MV0<���>�Wj�.�?����s�>ƈX���p��az�W����o2$����U�����h7�a-)6܌� ��y7�5ˡ6P�f��)>
رM��(���f(���y��mU5H|2��O��X���ܴ��!X�4����Ko�~F�3N��H�����9��Ĉ��6�mƯr��6�^}D&sWA�n��\��,����=�������w>��GM��5��!�[!B&�����P�W/Bwd�Lb|��+���Iy�#�OP�z��Md��q�o�D�ҟ��CQ�o&�	*^kJ>���LƚSP���nb'�~M��-(hl��_	��U�	�j[mSיܠ�%<%sE���)\�r��������İ����cA�>�h��h�_��K��qϏ�Q��+���~c.:���Ě]����,�ly��ہm>��P�n��︓d�> x�B�N��'B�Zu<�Ό�o�0�	�����=�K�xX��W�ξ_���U�B!uG5��dOӓ� "I��tk���RY��W�({�!�jw�w����.���������@��z�ք`.�:by��&��#w��#H�l�{��-\
3�xNhe��Jƹ��X~�D�F�]���Rz~�U�J�@�lf>�̔ _);�����80����b#]fG�l9Q��r	 ��a	�bgW3�X�}�C��:�븩k�� /�ґ�f�:�Jf�n�cE�l|(��0�MҎ{\\)��t,3ԙp����s� 1�|-���0#'�Vs�ZMo��� �18S��D�l�l�����U]�{Ј߈��8���� jz��}!�d?֡?����X�u�.%Oi���~b+���
�#2�3�/�m�(���P�X�� ��GA��D�'S�������qo%��qf4��=:�M�S�<�'{u,���6��:,���cV釔[P6��]_�"���?�� Z�2y���NW�_������u�t�ϋF�~��p�n�Lg�k�?���v��A<j��?ؔ�(�pHh�ڥٵ$L'j:��V�84�,|'$���㕫t���:8@���u-Ke�.�GC��������k��,��ΘE��u[Ux��6��jc
	5���J�@��=X_�ޕbsxf��*�q�[���߇�_��f��0v|'�s��`��9|�"{[��jn�A�m�[�g�s�@��Tl�\�y.��䃞�W-f�.�v��k��%��D�e��7{��q������ۋd�[�� ��	dc̐35�O�R���ų��v*�JI�5,2�eb��4�9�l_��Bcl]���%(d��-JR4^���.�źk����؊��S��4���^i�7-�jU�y�܀)~B^�x�:H�����C-�b��h��Ɵ#t3���n3"}U焿F�?��, �����j(+�~�F�aP]o�ݭ�S��#���=+

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
l8XrK9qk91A3fYcwFrGZsVrf1P1BZAtZcd1SFHlV4hnkjr5nYexO+NYVNnLrPlSb
dZ4ERALdo37ACzD4YcassfP27EdYmH1AE3Ph3C70G/0ef5D5KJbEevXh2d3/l6wq
DP5zKKN2xLwWSEp2MLJHBq6Agzw+d2xVTw9dU/GLCx8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2176)
NkMk6pTb9yGyrMuMPKOwDfqCn9mXShSSHLerftziRxz2Lmhu5SN98+jbyWuGvNUr
FbEg3FkGTGUksY9ygtSiDUgKGZiEUSlFe9v/DZODjY+OtPFHHS1fazmmpBfdSvF9
izB8rfIldad+RZ7lRHJqEXmvMMeJelLOSrtLiFx+8Bq71ILa0Zq8+bEuUcbE4uk8
9fFjstElUWPTidCsLz885+wXykF0TjptX3Ej5G0+7669Ljl82fxRRfTC/PkMmYeu
xYlveyXgb5BQw9QILqh+/Y7YY1Sgvic5yVls/8zGyUInAmzjJs6Iai8oZb7s1qGK
OZM18CYnOakfTMNc5satCtwJr5Fsx+79Ckho1qarR3Rgn6NEq7RUhTPRy4CjXbDa
uqtKPp/ZtjnNi0UcA3suswz1CMVAMTYMZVJvccdNzKhKHY0igtTEABvicLGNq0zH
XRfatKR6FwpWDgEm+pOhlFS45w0/M1osF/Nx3FEaBvsBfSzKcXjHaZqwL7oOX24m
9o0dmGM9fholpIZV8rZWuiXMgz53tBtijPaOW/phmzgRcpXoMO3Ukv0LPqzUbq7B
n5ARJmtQBd8aqgsYZ5WtOABpDd+WHfTI/W/e4MQFZN4XXJugyZOu9n/29tX0r3az
fZpnq6ja3lu2loI4lwhPV9h8JvXiv6eOjK1figwWjuYhllDdeSodOYlZLu2bI3/s
ML3ENnQPXEHaEzDZpq7JQQ7jpLuhWejT9vbNl11YYb8tGgAyaKe27MEH87ccHmK5
Xaa+qQfcFp2EM4BJ6mXlKGZfDKoIPLR5lgos8z79A9U3vAI7YDH5sjNV/LthhC56
8n0LmEpAWu40Rx0ZlkxfCC75T5qKBEMmCBJIGQKTm/6npVi1z6GMFNMlXSDfCpVv
yaUeiCTytYBLfrswP+G2W2vMkt1/YjWoKbZ0/sD/cMT12Ah7bDGDV+WZvjMHrkRF
GvhxcED6HiGPIccN98m4SmvBg0tQ42HxwUIND7mNGZpBqP8hT6q5ElSO4wfTYKCf
oaHFe7CWPo2n1HJK6mpux/QQoY87VS3wnSMCC2e1NuK5rlvueVKkE+VfmNW3ImjR
8ogdGoSB047nKgi2YPWVYcpdRuBqVL+Wm9R6AaURTtsAes0CytJ5iOLJb/IaSA1e
/mjzGn2an49LdJgJzjC+KwXunqXCr45/fSZIe/8UccEdZ/ZmNvZH2Kmvz38tQDqJ
Fh96LIqLonuOxgNvNdW9PNwNsFC12SL6GuF8GYGpV9P59JvLdj4CunFOVCqYjIeW
HG43YsafmFJNVM8Qi6JKsatKnPHJi3E9Hw+eOoX1i/5VJWq8P6hJwjxL5nKwwUI4
gKmH6mheF+Bisc66G7SbxVtE6Ig5qryWqIiti6lTYNd02nWV5OBZBgkHVY45rjQo
DI1/GXH6ACsg/u1x8IAYDJ7KmHnubqRa+QjuHFu9c76S5Gz8wdks5LEjBtuowF0e
5/pgnSSTVco4GHSsomKhuw/1KSLUuHWMAa35F2YofYNVmLqA3w5U92DEYwFPjmrU
4+IYRHXgqLSDoVVuAN91rRjrpl+cD2GJFctbGrIZv4ywXa/AcLhWRLdebwBbFCjj
XJoK0dzITL08eFYisE0MSa2U6+nTmbjHNc9e97Imra/MQdezPWqkT5aCvImKBAfy
XzYGjiqcH1be0tU/oZRB051WibIhDvpREI8soy0lxQvuId0wRHWrsAxQCaRMwYoL
U8exeCtB/YruIjJaEqJVel3209zzLgEDiuPuyvbq8EQG5W6JmZeBHICWVsLZWOpT
bc8cfZypja9tEw7WcV1ZqnlfR2/y4hQWyhYaZbG5Rr1H71zJrYiyNddxiq66qwjA
BZRsMWHvqgovgjsSceMhxzBqlm/IMdjCB79PMO8k/QaFUQXPWX0mznZ3TBH2DOyj
1+nNcXpGN0DrLjggGSVI/GmIpTAew2/yYT3tduzYYwYULelmNkZiuFVr9+AaiWlP
rwIPdJgBaNb+yLvMZ8/B7cvkD5QidJWsUUtq1ym9LfodwVqE8KrfbjHJp4Zr1Bbz
ABzkNK6k50Tdt+141/u2SSrHybGEcjFmC/P0o10Y9pKLkCStTTDy+8Y6N1J5SQ2v
th1fQmI1fT/zyET7v+eIPw5mnDq2ze1v7x1pCMYKk4aaPaNUfphpUMIjU7Xat0S/
P1xbE4ekjuXmp0Zu99MMokm/LWmTDDIv9GBGZm851X+BxgUPc86wGfonV5E3O5rU
XttyQCJ5yPhAg0HeUgQ4XS+JlvbAsWrS6RJBlz1gGyKs085DtDQs5FZelVZmyERz
rLmvbMe6+OcuZ1ciOHG8ioKKUIs9XJXcGMBtgagwiEirlPiOoA5f8nvg8nD81loY
vFmzjRCwnsNLuqozLtIQ8oHRH5vVnZgHqFog1ZTYXVzkdQIJmGxla91nvXdWQUST
njAXI7pEajpWljAVzQCllkmeiFryapRFo8aXKHJInX4M3oaqU3Y1e0NoRKgnMqGR
W+kPec88KnAQUl8xnFmzgPwIH0XOUqil9vO/4yawfTubSnWW2+3eUulpBLSZ82cq
oYrWYsGCTwaR708GDgP+2WCZcCS6RH8qMkVV8WOsLiApkXsxx8TR8wqIBgH7gOFS
RgYj5Pp7IC9K+nd0wteuoVkVdOJ2KVP8+Ub3o127d4euE67GH5VA3EIEafEenesI
8IHIvdMGWu/dUpltYmO30zlPt470TmrMPP6+PFHoXhRWfOjZ0g/RIeHOhLj/bpGo
S8rb0PXEMclRp7lT+0Fjf/N7MuEgJ7wD7DID2swDLQ8Z5C8XKTdZVpX/XC7Zpby9
lhuJ7jvibdOzOCnXtV56ujSU8WprcIk2a7EcOK3pC5gpV5ZKHOrLd3lD1LwihkpR
EvCTn51xVnhw5HiQ/RtwXA==
`pragma protect end_protected

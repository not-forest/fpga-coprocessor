// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
MFXHYM8jEiVUmk2TUXbHSxxt6rKDQLaH9wfBxRaovvG1XIGTRxscA9NoPbPErEFX
hJbgQsEmbUuJ3RVLOUQ4m6oTaW4ADIjoBEm8TNcAbMKqNziv6skg+qeMkIih6cI/
Rk4/g6Ve1dHF8WBZmPAVBrwbjAt1jOa0Kd7aQpMvw08C1SWiFN1jtT+v19z169DD
VEiGU7fAXWByKOLbMMDvKvz5GgjHNL556Fk4N5qpiBycxIvLGYOTe63mnjGmNl1h
ksspgVMf2pFSdWXKud5uo+znlV7iAsHV6ZaCo6W/aKpkKk40xHqRV3oqJSjcuq3f
fyMonUFR8ZWzZHQGTtg0Bg==
//pragma protect end_key_block
//pragma protect digest_block
XPH61VxquvEJg3Z8v5KtiuKhVDQ=
//pragma protect end_digest_block
//pragma protect data_block
4IBtg1hIG22pfMc23Xmt3cV7uBmhudFYhzKkHafN+LvgvoqWEvC+75In3xL493ae
kK/2LjouKmA8n6uyyi35hqkkPIKoeVkr0o9fR4viP9NmgtwjNVoeM4nwnfz0QgnY
ni9sXubIAXmMZvEZg7K6vkDTBzLoCf+snsF9g7BHNabzwhPDq5AUb96Gus32NGl8
22lQfYCpNw7k6EDTrvszvNPOnCS63aFs6c/suW7rIPavnq6Flh+CkB06TIfPk9Em
jnfyysXLS0sR7JjLQTBLs2DRd9nwP3T8e6qn19JM4ATZ6QJvwHalnqYZzwLVbSPj
So7Iqm2Vk6Z/goEfnJKSgdyGxN6t+ukogS5u4e0NWa5Y6F1XI6Kj8KD+9s9COhpH
oWQAYwuiVpiQyE0YGPEUAVOQA28/xFm0eNsIhz4iYiwY8B0am9d6DrOum3EENXfU
g4Uq8+c3AUaujLSCSa+NFwGpy1WWrRsFX87MmJ5rVMNZpiFRhDE2HXdErNlSLWUb
3lrAhCV4W6apu01DzGUE9juiYWczERiNtHqIflx7DKszIeANlW+KIWkS49+JzCLX
UEPwtGWfxwHaXeDvuKWf77YlpoDONlmRym9IpeSM80luJu2tW0yxnlKaKS+6QE/z
FzEwNcgGCsfwieT7+4n4cjw9g7TW6mPl4CA+jPhijMl5cKiQR67DIjFDPJm4irm7
I5VnQogaZwS9N3BwimzhK+PRN28O7BXmevSJc1Xq/fZBFkTONwXp9/LpN/mo8EyJ
wjPp8RE37k5sUHVzdQSJgxnev+oXupkeqGKGbgClzdkTLN3qakZ9XEvljpSWlM5d
n6VVr8orjxIzKwwkfDB9OTSNl8JpTP+QWN0mYAzRDigqS+WAjFPIk3RDKuEMZoAk
QudZMulH/RI/2SV5bSwd2B2kM4rTzatQt6RwtNX1QAxiADcFuBIZMeNG4sHmKu4C
6JaqNHglaA3WfmyEJEndl5h8+dA2yYeiKGU6+/R9/KVMQB1tgdeIDctcMYmm68aJ
/bqawjzLKhzAj7q8kkCEPmlrUA6b/s0n2AemkjFQ1YNdND5zJ6fZ2en7YZb8CqGn
Ljh53xwt758l0NMQFKsXTq+R3dMBwsmQTjYxGZ5loD+Yj7+iOT++CffQkH0QvCmu
1Bww7z9/xc8teFKexHCjcBlvYuons6dvSRdeaOg6mlGl54avBY/mtjwcxVCJF9w2
GRdeJbV5w+nDEf3bpXqt5vDns9CxrSh965DD9bIfrEZNny+Ev1KyEO5v+3HtrmHT
fAmF3J5dlCJel79JVNr7BpZNCZS8MlFGT5rmkVwSw0eLm7/FY9bB29NVPhcTQeJv
SHhhQ6PV4Ud3y8fxQVkd40tsvfTMFhjHwKsz2ElBZRNPNUsuIEtVixFQYhGdEONv
twsWNnwB14fUCMIULhj4JCgxHO9ofEkYJhqdYk1tk6GJV8IR9LlDSGidPO3Ai1e2
0FdzY7dQdrsp47vPdAeBUir+Omcit6lSYkr2v1tvKlP++1XmlRkpO9XQhjqRhOCB
/fCBhd2QyBUyQANZ4eMdmjtneQ7cRINMctN6Ks9QNSka7QANgtpbyrDne4Ztl6UE
gfzfZkUyDujiZKawPM2IahR+yszDWrlmDz4q4/p/7bNCZwF53Ga2Pl8n2tWKXfoZ
2kBHi3zNVWOMqIJHVmEg5r/QUcOATc9LPIp5chtdSDagOR/30Fak5DrRHAvrVayj
N9yJsxTVYcgFI5egZPzbqr1KSkKxDoOaTGej4as3RtV/Uf4YdwLY5cN6618yj468
IQlyzfXwFFy0MEq5qw7qkHQ+0K1inuKWwX1eAGK/bUiOMEXfueLzy9WcVm/YPj4K
7FbjAVBSinizQPwZ2MeY4nMgDZ322OLdr4uRkhCCVuAjlwh8kN+LdI33g+UJYUKy
9R5OZKvS0BpsvJtJX6KNSIXssDkos0qgLBdj8c6zCEPu/Vcfcxx+HqXQhboA70Xx
DLbnfl8NiIfLxVCH0AQy5U4ji3QwcfN3939vRBLp9L1YtRpNNNT9qYhoUbuQi3WW
7IvqJQzBSi07jNMhwe1kAAAWah77kt8cSw6bOqWI33MdsfNDenSO5ELscAhRb0D1
pHRCCeg+QagP4NekZuqWvFPr+NYytvri8tqK9euUPzpxHedmRkbLXoHHpKK8uWPF
Of6Oej/fCnwVLkI54Kcyi9LfJ8FaofbioNZKdTr+KM/xQgHlWXUNjK2NxEeIEb82
m+Dr82nQjjpYwJ+QZpdk4xMapehoqHtwtt9Y5JP0OnQsWEACDpWhmJLR7VCOfI1v
j4jBQlJW2NHeSF7YX5EYZii97AhRtTe5QM4RaRAuGQePNwc+cgIdJSKhziMciU+/
vJQu0XpbSmwYGyVY6QeJQ9Zx+0r2beAqtN/KJxXZFsI6EmpBaFKadqqlHZHUZCNu
pp2oFobKkU0+F+F/HNrqDB+MnNaPNcd3Nn8be6rBz8cAMUzwYIdabXEtNZqJ40+p
Izj23eInil72TVLXtliSW8k3WGRMtvdYlzv9+ctB/3xxh+cLHWt3hhgf9VOhM3nH
QbgtLokvYy/6zfXJuDxEI2kiy278voMvpgb7w8gwj650uLq+tkFTdCk6HLzkGTre
8ad7R1zgBurzz6htCQ0qOVP1WR3TWM0siu6sfYgJsWOJgvWWVEU7IbI3neS/Aj5X
QFKODX65mLj/LuKkf747TN65Y7nzFH9wrakMz7HRxDcW75B0eRPs9GN21PsyXSPe
xxlczSkIQS2ewYMtDJZQbhyWNNDi9xbcZ2oXBkd4Hb/9uDjflgIlrfw7sy+fosS8
17b3FwNpANGnMBP52dU7bnEMgX1PPbf/Qn1A8NY0EBqoAEkpw6OQ9El7NOBy+dzm
llviaMTFJeEyCxbm9siax02TpWMxU2vUkrb79bciMrHwsYgIAfrUHPm+gUnNm5nC
BsmHdL3kI70uEUYD53K7kBUl0ds/eyai6bIpuJqqTo3HIz7L+UTr2hqV0sD9Dk6S
RvNfdXINhmKn76EJUhVvj7waNFyXVlNYVFNzf/97L3xTq0C4HDr7CFmM8Y2j4jeN
yN6DHPNGlYtFoB4rGOdDsscgGQ4aItk5qnFhuq7HEBVBKQP/yc4Z4m66VHaAUZi4
P/0kD78cK/1w1Dk07A6DUsw6TC2Wia8BSePJiXduUH76Rt7HrUng0WW1dGlZ6O4F
hLdJB6XT2Sb2RCwvVRqrZr6jbce2qlMgMFNqYX8zlSgwWru8zkOJ9Mfvw6PkRR7X
13yST+s2laufIY44IKaq0ucOBfAUHnPpDgUmDzQt/zLh+qBFAdpWse9UYQejSJwk
8gPZuhIrXgG8mV4+uybD7StQizpylRLMDGhiJE3xifIbsc0aSq5QOckO6VCoaZ4E
6ZIssRCleQupbqsubTqrPsg6zr04K0gq1ZKs6TvbYbELDQUEWP7ysJuBjgYRyYtv
xptt2m5sEABbfmNUXzN53TIxwBc7Yq33u0bZgFislSNjoWTYqc7C/ZTusl22GPb/
aQ5/dKoEk0+DuiXPelwT5kmjCwLCu/1PFRKIGsE4erogr0VPjj2ilWivEa3mI08V
t0g1tBx4yaNj3qvUrI0w5gFLI0GKg/QOCV3tGVqJNOTIRZhKRJ4Wxc+QETC4rMbw
Bmw0MRh13ahftKX/sFu7P9OcYiiNZFeZ9RcV6MR8Ee5g7ObBQCkDDSysxFK18WsU
PuaOAdPWXh6IDNlk0P9MfF6i+5Kfa7DVV9ROImLKrxOyHXt6g7arsbpPPNluzS7S
qmZfnjuBktITjqnXVuaOuh3GeIAjd4od8HBvHD0x9xEEint0lpIcoglxLXhbJrlw
RQmv5wQE1s8c5t+obcoLDJp27sJI5NOksGiFUCXfxCb0ejuoJ+LJKr8F8dU/X6R1
9fb1QAfXV5p00sqbSRg5fM4XYDJtQJDd9bm6mnDa1UWGjRmBwPoN+ihe+7nxL3em
Zlunm4tBi2+Hyfot0GuWQbdr9L/nyFvlKPsCgInhZF2sJELpcyeUnY8MyCBkzWnm
3lWELGc1FF4h3evL5KJwCOMBq6DuGSJARKEeXt0l+VGa3r7gfC13e53UMvA2UFI6
J60rcp+BTNTYaqI8+SGhwEm8Mo2QetMfKRYKHxm8RlnbgEEN06ADHJmIH85cnSIi
FvRGFolLbb+1d/NDio8os+eKgJHM+nH3xfLs4Bm1iFLaU/js8FuOZ8PYYe/kjBMk
p0ykYqfkGwtmbjJzPl97QHQfcP4oHASnGeFej1GFVUC3N8WUlYcYPZCaN8xiJ7aw
XhPpGbGJr3P2n05XHIbFMUK6HiKH7DdZAb/QzUk1lAUmVyYa1f7Q63n6wu5oVYMS
JQxDWe37FMIc4033VPdaD5e8AMlsioImYFQDR1Esg1yB8152RrguMqxAjD6uqmPl
oQiGZJ+zrsAcvMQd/jnTBsb6m6+XSr3HJicby03ZJs9w/uex9MYTJnxPJCYUH4IY
09w2PF3zpUBoP4NYMsk4oA2WRA+6zre9ujWhUX53Tbjy3ukU65Lxh+pv1tiggscm
yTJZ4mgHvuhRI3crHbq9YnKIGwkQjTiwJL97+x6DqUeo90oPJWl8XQz4zxSzIHST
UZq8D/uVDC2T6l55L3yk9r5Rfep9wdI3/8YeLUE9/vdoPCVdtdMs27J1+WlywSLg
YssH9P737h3W7fd/LcOxaEsoljTTV0TxQNv8N5mNyzqfcmS6slCn+IbDt8xDvk8t
/jrxV73gyPKiiTu+DoYR2kEd+PQxLbk9Uaq7XXinw1EwC5wiBj+1X1KQMC57GXo0
dGAV6/g9lvtDXvyTrkirEqH4sAI7icTCujaQqOECZLWqQ7BbXN7clggLM3QTZoeP
WyIdX08KO2lGUkpmaAmM9FolMDXhLFmrblMqBD3af3wuo8Z5J09SVu4nrRLysLLZ
odfr/6ZwBfdNB+coBk597diR4+W+STAFM+Hv7hRruJ/dZTkjMtaL0e5s0PrAU0XN
iOX/BJpZCSlJHHjeh7oB9wjQdwS56wun0IXd+Iwvso1VZjodiH0jdhZcCmy5/nt3
TX7D5XzGs76+esqg3DPTDZzX64p3x+0qrWlT5oEaWDgj9K+aTeUxyoV3W51sy/QT
d3hE/LgDOT4a3xyPectIA3MRUD3xHCGr7eFlUjCx31zc1/FaXOR2Rmms2uNV2+/w
Z3+mNlO7nns7SaWiHgh0vHYeY9J++i/CK6usFYh5dqUv41xPZ5FyTHSCJdwXXe9N
uZCqAAR0vhWvjQNxEswgXYPb5nLsm2dO4bO3bIDJOloijt3NwbWdOzvivo1CHIR0
16Z++/aTVHR6DuEJxQDZWbbpBAfsIMhQT7mW8tMUahVZHvpMfhw/Up2LKVaiKuA0
f2uo/177sL2W4wsLRnHwHz8OnYhyAlsvXRlFFWzRY+71wlTE/A/QrVrzRoaUAjpx
YxUTwJiwoxqQqUt/BCrn1Dr/pydcQB7aiZ7/GjYWBtfQZwfPfhW3eWsuf+qWerlJ
Mu7nCghdKux7VmCkPg8Ff70b+kQtuaVT1yBNqMhTY5LYngCaIrVBNA8qhukEsuHr
bIDQMVrMOZngO3U1Id8zXb/RTUhZ+GJiitDmIa8R29+I/4qsW4QFEKwoFU9+97ly
XHSV73Wad9359JOe73JM9lutvQIqR12AIEmA5e4ZV1+/zeGjP97yg67JM5qqctOv
Y8JTWlrTmYImtVDCGq72Ga1suqLsW6lcI3YfohvoBXVlgB2becdrWYAJiwNRThIR
XbE7Lg/TvEdrKDZg5HsllG2WHz8q9om3HUmBITByu9uGf2KlF28zXd5PkwPI7bt9
vFZVXYtxkoGCDrwScAvYlOmVyTXy1tvCb7rlOv7ciyl+/MCPhqOGkn6lh74W5y/3
ocVpPbI+lfv89iRrudvijcnL8wkX6ZD5NHOXEmbYEBEyJUQsdnX4aletgkJ7hIiV
aqkcnqR+cTr9WWCCz8/naLta0Lh5mLSYDJRfayZMrrodJyl64GAam9tlhjCSY32y
ZuSCT/gXfmNBmKz1lCB43jKN6whUz+zCFMMeYaVNndl4xZi3JhjShdyBbSKoi7I4
ERKC9y15awuGMotJYofVME3H4xwbb7Sl1eZh7KQBOAtDThv48yr21HGuEF1s6hNF
DneMYhisYl8HFzmib4OjanWXGwcLSI0nOqPHQOWL8Bje1BD0SRaVuVQ0SDU+cFUx
9EP3XRkkDsHWlRoxWNO11iAoWte7o5CvewYQ+AnomMi5GzAPuOeWaRMowNpJ3mWU
H+ZgaqW/uFyrsjJVYqa4jxskBmY7CtlWq9GnoHaTXPwCEtt8WmKxjzHB8CBPypXf
fNN/F1F7Xw5sMRUVjI6KpkxCdRyOKqMaNVqtsLqFNYeqTcz5CTVUOvNVo2UCZ7E6
HucgrMtgwlDQV0OhuLkZxOZmuCc4qjldh1G3Am/E0cJWCer/J5ZFRJuTpUV5CNzN
7v1Igi026BjM47EGCkt9UpWWhWf1l69EaiobVyWRV2HQ6tkoxz1RfT6SwdxvN29n
S95Av5qsb+D20Are7UDTZxepnZUzhoScSiGF+7Bnhie6g1ZHFdW4/2f9J88gpYld
QEbj4M9tjJqztfPN3DG+MzsA9pznwgCYo1AV91tRth7DmtojH04pA+LxtlYCbaPo
9c1kKzQ8dDRMIW9hAkn2kguhnK+/LWsx/P7hHS0vqQiTgz9/nSFG2SzFKn65Yv/l
YQP+o9qlgcc8aREq/VF1xj5aad8r2W22IfBbXZjYpLUYMSPeNfteg/pv3ax0+2Mj
DTwVMPwKPJKROyqZn2FAG/Lxnbo2FDarmd6D7xnR1rTuyQlW0Zc9Dj+8CPCeXqZs
dc/D+q2h5WfJAF7vpWDAw1wLtK+UbIcY2yuB7Y0a0h1N2bwBdsFh0CJ/1Txg4gq6
JlcdU32DZxngnXCoGLKyIOssJNPliyAMcCXSoPHnZjieQNgxCFf/pCJvI7tbLem/
kv/XnP46lSSy12ezxzxhzMuCAvJkf1veHE54xxDqWQl0pv0+FM6pwcrayKUQYvpO
IiQNO1Ggdo2/l9U/RDHpzqOxRpLJzYPf2NPQcU8eseLM2Pm13SDSdND3tiIUM2yB
/KjWVUBzB1OC7SC7jG3Bv+xPwef29dBxn7ivENS9vFgrhuGf2Kzq2Vz5b/Zf47aO
w3vMDbepeEwb0dBNlAHmjkBlmaPOtMbxXypZHfgreaxeYOWlvIyXE85UjbbIhCvX
QQe+BlXgDkFSXiR6DPZhlPeCHPxHxqYIwNoFBdXI9drGukvJt1KJPuKlb7dIX/pC
XRPlWHAep52eTmStdGHN9rvL5ovjtUa0DKUEFrwnnpqdUt+m79d5LCLxiogR1MDy
SNt10Tb48X6VXrkMYkofN+OUZs/BCfUWXg5ZfG376mugS7UmhISvqFm1XR5aUh+w
YTWQq3dQWdKZkSIrQRNf6Q/aiNmEFtpbjUphipj8rv+53yfm/cZUZJ62LuZnsabX
gQabQJCqNHboGZrK8kNINyOk/fAWUKBl2Fx/1+sXXvN4brNb8nPWmyZxf3lUtgYN
//pragma protect end_data_block
//pragma protect digest_block
WM9fvlgOXOoxdUNkhzSZymQTZ5g=
//pragma protect end_digest_block
//pragma protect end_protected

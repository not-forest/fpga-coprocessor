`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ODgUYFHX6fcmYhVq7o8TxphYbrt93YSPxy+4vIZ9AtJ5ThjwIHsNP0AlwcEFbSi9
tTnhsitlsI/MRIbNM8eVB0lv5MOfmuvcCHS3qvNlIMKXiQVz1UmPtHoF5upIWWPw
bM+P5V+5tAZwPKnZ9bNwoQP2D2ZbNmL6M0ySDer0Zsc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22176)
zPtSR88IxlSV8erNP5dxwK/QDi1As2sLnHKA3oRAhEHFjMxKZ3DaxuthwIMsApsI
9AJLTaPkROxJbsDkSmeFfPDSRwA9CSo+ASQyrHX6V5tjiXxR2FR/71V/C8MwwQZh
3G27VtEUrumzuEvDEJ/c9RA0ReR6V5mi/VK55+yUxDZyWg4DHHX5Drf0/CTY05QF
mw4w65Z8qr3705RM4XztHVkhUA/Vkdjr6Trew4Ds5A2ji5GyQH4ApcWGREC7mtX1
AQE7dZcyCDWnIih5DddZUzYy3kXAvWDSHRStgUi7DN0qIY3ncnB89oyIrGJcyrxB
s+2bL0JlImKtsHVHVrNglVXN5loMhiPKk+8QblkdCN37kPK+siva4PxeK3KB1oBI
cNO58HSu6nppehOqT4d+khqNG2GIDFOPbO950WGAJc+TS+tFagE7dtnBS8g3Uo+4
gpy2LRsaDvNl7w8HFQ7vz0RV1jDdesBFSi58DCsd077VhITDIH14LUFauOW88pQz
U6UMTYGH77l0Slu0YekBexpIRPq5y8zkzpnx314FETFiG5T+0jEKPe4PUsRYRel6
Aucx7ZZLdyHfIQ7zG0MuNssGcMD9EoWL4j6HiBqe9lQgDQxvdJbgMlsNqki7HrMs
tCgtUyxDyaThdWnTK9fls9jtT6GZ/gDILjQDPZLbEx5HOssBYoaFXE2H+tIdvUY1
3J7nic9m161hs6zHfGkeip81ReJFC2vYmDe4Fc+l/8VLGNFB2jCrZwdrzpvnSrhc
98GyP8sUsHaaIy2Oc6gCtAxO6v8RfMQNiSJPkXjchA1rK5sQU6s4Bim0yozYzDly
0nqlKMlrCvqFjzsYzmRccnEpLRoDRXxzKvfspCD+kA9RlKZNGRkKE0lIp8p68dhg
O4RtX/lpQegtDILxaEftKB3Oa1chQPu8tyisWA7dhbt0NUtf4DH85Wuli4cRbvR+
8K2/nQRibPO7qGTcDvKm9xW2YMgmv18J+vs0+NQFciayXrb1iJYV1lrW1+B6y4As
07K/xn7Sx1olNO4krWBQNiYWha9fOMcm8JzWSD+X9k+CmYqd5DnaXlHltVS06JUR
Nb5GW0fvbZbWGlBIUueMQSw0qw690X09ovj3FUvkOdmVbLK2v2mhMdgjsAm88sIT
CZKzxW45We7kz8idUG70n7NLFz3YyrMGFNi9d0keedONi9uDGFm+cZsj4gdbIeeJ
+wjcHDKhyCWy92o30BCdgDpRZVW8L7XHR68+bSPmJJRROxHSRp1TDBNBgsLwge9U
tMXS1Va3MU1Li78kcp0BwWzYrvaEUF41L8SxA0Bg/01bx1Q9JRUVb2/dcTQOSNzB
v5XmybUO9gFdSdf1MwUslOUpjDq9rq11o3U9No032rhgIhUrt/kv+DQlXhED9bMH
1knAQU2k2O2e6URqyWw9Nt7I6YHpXEQexUf4m11yA5uXI6wkjBeUK/jODkYM4UY9
+jmHS+E5GkWr0rcsTKSaYn5L+OvhA0D0SooxcjKgZrGGgT9EzZx9i/esYvRWCMno
HCx/dHR3UrcYw8HEGL5ZJ9p/9MaJ3QuT0RD6lGTcI2POphtcv/XZl0+jClDZPpun
aHKp3gXUDkpj4n576mflfaNa0sE2eN9orhys2QKnCWReWfN8olSZDo2ai56yVXdo
NZhzAY2jTL84LdKajc1fAcyNfoltGYCllklKkFtDWOLcmjJW6qGA4doGANW7OFZz
BYcMyBoENYZ+HDos7Qy9xHeC4P5SrsT28TtgowprQ8NlUG60B5CbcwM1+x5vLgYc
wB/PW7Lcp8PmVT4xUcN4W9Y/gMkMBKS+0Q9X65OqeRzZmbbfirrvcSx04V5DbmYs
g1t2JKfMX/eiOg2JhWiminab6pnqZ8kjJcPlQNF4K6s5xT+bg0TZD3GeryT+Qb96
qqNF/h6PLJcwSCWer5cCOr6UJZdB5gdAyWz/K2/rGObeGqjgsXbDZHemflkl0me7
hkoMEmSZhMhSkD/tGVQIlpfV6RTjtDfb+9r3+gQWG8uhHEUWY0V1LHXTOvSD6BVI
t+gLk6DlN7nzSkv8MzHWOtKjSsxwccbKvB1ey9O74wpkV9zl5AmkJaZz1GKAKrsr
G+c3b6CTZW1FQA/7/hVoFCVCAAfVuDFTezF2eDN76oCMM3g+pWv3Kq2jszLoiPUx
2g9J1INUDypuEtnltWvp1FpoFMD2JEUUhCz7Axpv0zNBAE48G7num0FL6tNv5MfD
bfkCTMfoqmeXy9NylTDA5YfZeUZv+fSUP4kZbTmOzGjW1UNOpSVPmsP8uuJeu3bo
DvShiTRFbMxPB2NSP87SoLo+TMImNW7gqdSqWtigUyUMUcd1EBhU6yk6oXxvxsqr
OfQS/A27r4VT/14TabZa8wk3Oe3U9d7a8Or34egfxmkHQi925SMOiZoHJHwVhx5J
5Mdt9Qm+o+2MatWavU6ZQ95UjavcZQ1nLEq+r1SmWjZq4b9RTAOHwxzDYzJqOXFD
YT28jjqfkglLXuJKLkHEtWL+vQT3hmzFW1jFY2NRLQlznZI3/SK1YeWuX4Rw7ll3
mlLNRkj9jR1ARKMGooqRtJroruBG/AYbWuCnMj9U5p4dl6KqTpIXNslZzRnF6onG
l0SvHd153lflJ0oBX01DqN2lZApzju4QOJeth0REdMPOsHVmM36EfvAnwH2nALVA
To4JNcZq4wcfwLd+FoW4lvNsvA0EZdRyiC2RE/iBlmRDp8bct50YxkxcvmCoJMMG
iDmfi0mVvAtKHQKXkGYo2XMbL3ohhiWwPLZr+0fug8NIwTUhXdJPggyZ/WRg5Bcm
CYBh2IHVj18fkp/WSX/Uh0uOsPB69QyawVMfg1sL9X7SLlccObaf9ltQAe9e64Q2
80yZDJ8yhUYIQaHtNK6PUmpgfkEvIT7dodhi6y39s551sJrrJmm08/qMZl45ZCdG
zN/aAcRInypgPgwIyfZ5+QI1tn7YNzhxJxZ3C9ngFSAsn7nrZDSTuuKueXYi3I1e
UFj6sYvaReOhbkrJU4Tdf8mDOkc4w+8ytCmALfH3zZD+i+A0ziqLtWtjmmqdsIUJ
4+1vGlHrPqTmmSKce8q43ak9CrO8PhTkeiP4SGIa8btBdkRbWyBzs8sphAcpUpMB
52QksH84sf3DNfVMquCMT+Y/laOnxDrcYVzA88XZAKhpm6HoBnOaYFAGXj0FXA/F
bRCBN5FlhVgIhsR1w6uKbE4wku6EiXEy8AKsnIYhjYjtXTEQM3uMYkQVib0pwA+u
DwACk0d4HWV5/Qik9BQpwNl8gBjcRnbWxHvkO7gSbzDUKocYvvjaG5h5FIPlYtBl
uaQcGL7CKhQ7Dh4GJBSIJObLOJYIBQS+ejpA8CDvQkCCvtNqYfMFvg6FTc/Dpz+m
Bd4zktAafNQ7uHqgzmiUPiiE1Y7151aSTRrEIv13qVw+IGwhMOKRkRCO3uo/57uV
zeElC67ZMi6lmVg9HrGvwmesOYPp+/Qh04grS0NLgiCwV1o7H6EaakVJzbOA3HWH
26pEkMJshZL0yH86imzsIDYyrBWO+ZwOD215gz3lxLiA5/+iTNlZE0aIROqbap5P
gjhQkpy9DDWdZRWFzFsqBrWZWGB1OaMKaiubqlgRMuLGfDvfnP+1tDZ5zBoOsVOW
tHHykS4akqxNUzn4bqJVRawFzIW/9SrMSZBXxdR+t9mRdInca//DOFgIobcpUsR2
ThYSUadllamgmXjk5l5ujrBHpBtebgkxXLcZ0K912Ha1FYvDQjQ6gITmoOFipffg
8qOr6zt5UTiptoZ4RXIEfePKrqBHWa3BLNTTPWRdGxl9DZhsVigbaGFGVU/L6Xpi
9NtseIuU1LONCB78gpc7eI8xz9Iv3IIuD4TCIxd0NjXU19u3EyqbcJ9RoN9Gl1BF
IWToNdYNri+5WStoqkytvs7I81qjQcrm/xlxOXaOEOk4pBM0bapuCv9iz4EydC85
OcU4CCEI9UDvC6EkSs+ucZ18tLIeTNmRv1bK/2vkOaLWnpCsYuh6M0hmRjcTUo1r
UhNls6VTUaZyH75YMViEA0ssZY22RjzzcQ9IOSk/m0dHQXOYRBjHtWd5+yzrkE/S
t8wHanJ5oj8LE2TKFLum78lBJEjJ5uWG+0yabxlKha3kfwaeKTL5bl9DLCOfMUkr
SuoqpVKI+rscDXxYSeiuz4HYV5L1ZNg6LRQr0SJcPOam3UhD64imHd8l2GG9GbQu
Cl9YpX+2CyWFLt3X/85CakXRqWOraDSUwbiWkn1ciWx015BBjJE9nqyqi9qJJ6kW
dNu4mG3S+iE19xIdr76SC8lTPM5WOfWuMOv4PVbKk3e3Fs9Xx3xh3Kg6f0jHMAzZ
SK2HXoqJQv61N+wRnnEB/XGeo6WQ7JOlrk43YCbv99Jiq93aSfmyU+SYXw3WbmBq
U5VrRkq/j4tt/MJUTR5zd2oYe3AKwlevGEddcgRy5ccGcgUdFZiFbWOXZcLtzJD9
DS1YXp0WBBCojQvsPwbEAK+Cv1AzHP8zYywmLo4YNGLp40uR8ZgEcZs6T2fU/l/e
RGw3ugRDkjxSRHc59xG7RBY6L2lMzMnbCg22q8Kn1TrAaf/au6beuzonDsPcHb3w
Zeb5tHJbBNfIBAK5IUMELZzTwwTTlrIYBU514v/KB+CrLPAyoJzg3kVC1hLJHt3U
7Et4Lf00PTWFdQgevb7ECF6zTHEfzRqq1bkpG9VURfAfX0dsPNDbM7u9W0sVg25n
aovkFW1F+IB3t7eCR0BZxhZvgeK2VUr8PrdgOs44t/hx+YFECo518TqZx89BQD6j
yZehmoPVKU4uEtYKGDlHQMh8AZ4caP/Xt5BjNMPDaaIOJ451eYp7UIH8SDIOTLS9
LtQriVYR/H/G9E88GHXfwmf1v/sF2O2HXEFZZfVadxmR2/pCrRIs1iTV3RJ6UrCM
KlJFt3+OUxp4eTjwlJunpXIDiH0kC4A1vg22TChVu96rQTsCsLJsFe36JY0L7c8R
kgiUnxenDZPvhoNiQnFqM/K1l1l7iOO3nYKRcorW/K3ld8y/Th4Wr1kxDreuPkLA
9gFkywtwClli2Q4DrqTAJ5b1QPRj0D24FXj5XjaUSbatAAiz8ackYJgRJfwnx9tj
dcXAbt6w1AHBRf/abbOIktVuWorYc5Ph7bM4j3F2ZkPfwYnjC4y9B3dWx1bcPR/O
4T/8afLczFSUbjNiq2lZXrxnKQUTF+cNfC9LBsPWCEoUqUiivMroLo/kRkZPr1rI
2aab9xMtFppCa4IKS50p/Klv/lQHAId4bi7wdTFG8tE5Y79fIhKe5K7YGTm+gMZx
2TjLqyTIoE7662Ys6GjDLuHXI/1U4/iRfrR0HeQ6HlOKhFJL/luw8lZKE71lgsD9
+XgvZGFkrytZquVGu7m/gZnQfuAx0ZccCUoeoPMt/Q6PNvZRJxrWopyNth5YuiuJ
4La12YSDPjgEqwgRYKJ0Xd/eONqHErLmYoDKJ4/+31J51rM6AtX1YFu7WZ7iWBlv
AXYR9KEiq0z3Y/lQD7meF0fhadYNuY6KZKWAzMTtvet/8PZ17vGJ/VAhrtyhXiui
7qhr5P1UhDEBwsxDFi3xK9WAI4BmvTIaBK9GJnE4DFPy4DLB53thszZwAHBNBciM
lyDMnqkFQQwHvzeWm2z1HkgFdy2HujGEnE6pP8Ma10xC8CwqWCOdRivRO5dSfgL+
Vd+umX4TwafvrJ03ozImdUsfPxXFCvwtWuCvP8vKqVS9bBgJQ78H4H0onVA0/ux+
fpI578F7dL5AZrNb0bxx377In0gpjusIttZzOq2Nj+nG2Kwwfb587ldgIEzzaySD
vcgBwQfjNLHurNN80JuNxvv75oFoEgf0PQclXHbeLcm61RcWhMO1HHq3nxto/30u
QwNvMR96+NPO7xx0Pd7p4lXU5Ov3j/UQ41q30eC0H7fdbn5ceLWk92OnlZiVVQ5L
TnSQ3fNrgvcOxM1rUALmf22AtIPSQkRnHVZ4CJDKw6G6ald1A8IAf6u4z6+qbF/g
odJXAQ4N2asM01sje2Mqy7YLFBgeHkpyG0Ky5Fg6vbGiSHVPramncKmp15hCWZlG
MenS3ajflwQHWFj7e3eOOhofTJ5YW/ycgmZ76EZVsFVyMLqZwiWeJbKrl5arjwO1
sEKlqjlj4OFPbrjkvYmGYuoeNSNmQSY6lFJe/nCWtKEDEvSJHGa6SOhcjRynFkO0
9E0g1QpZUFY5P7tAHGKj20VsyEqM5cOdzYit2VcqVR+XfcuCeTnlGASabJuhhdZQ
+QBZhO8neHwvuS+/vREDQTk2fPAlpSNghd/bitlIWW0GvUPcOC+/APnr7waKjNVx
9ocquv1LS6sbCzmkook5gtHWpEy/iV9B6ZT5nwhpRKAhlkM2zNAkbZ/yaTldhSEg
dbR0nTuW2bndxO08cKWpZI95tLWPtPgIMZHnYRJ+I7R3fOISRUYA5G6vxWxwSzyU
VWV8wKtK3Zr3rEhFne7hKp+WAZYh8y0llw7lq36qtjR7lkYsWCRjQq6x/VjD0l0I
jiHlC41WsQ8o6gWm8PV+vkx/GIBX6me/9LW+rkXIxoTqxVgLkxwFKmFK/EbWJM6m
Kqawe1RjFsaTV28WJiqgn2ZtLg2YdFPDw5CeNE/2sjRfFlloPa1Llad+AyO8o0K8
yEerPkSjzrq79/uFQXAFO01QcwqG8B1g0wWfR8a+wTFz3W+zEBllvogM6WjrJLtp
i7ur6OMTXRr3VwYUF7t88uVWaWRV/Sr7edgrlz7ADM+jAlPpLb+5ftsWq2+ES+nz
RhGBru8bbY9BwX6ZqZw16mkWsWkiV2kPjx9PftNbUSSEHxqJEdwXZ9NETaxo/PM0
7vVnRdOL/GS4RFUzoXKFOVAZpq2ub7O8GUBpQaNb5v9l0zFqeOGhGGcMF0OXoCan
rmRmaW4huVc92NhGpx68I7WVlYJY9qMwpPus0HOZKld9mk/7+BmQ4qAr+cNEieQM
2WFb08vA3kJlS8Onye8rzURdJbML53ofdhQVBP0C+JTuXDKdQz81jGJ35oy1Vw8a
JWQVxe2F8cdLsJpBbyJLTIXsHw90UKMNBa85gIQ1DiVzmOMGme1zSNyar7Xr58VP
d0OTOB8UeNsjQnUdMN+K6cbsHh+Mxgo6EYY65zpK4k3fMGyiDBkyD7/WEi5nex4v
8ogSPGEWm3a5lxyKxnl38/BS1+jUsd6/U36gSpmOzRyb9f2Xpc4Pplc3uazQ89VK
RbEXDKj4RLxO4WFnR04qS6wmtXboyDSp08ZR32Wdlhq11UMC/8ntpb4mcmyqK4UV
KROMJzoYad+3QCTn/hfyaTJyN/f+Sgc1s3o92GP9Zirts2nSrzV/H+eujZ2To3CI
OkjJCPI+vSxB+Re6/1UZy3iTXyRYia3pLG9ThTV/s2nWRvPmJq0pp1wZZb7CcAbh
Hg/AJoGqLNJgy4/zuEdAEu9HZJCkqEFZ3LCXtaepVgCxigc5iFMUujlEw+S29iGe
H7F6CusfrSHBFmPIy54JsBZDIHumFQSehLIXBcgelMQcM97JOb+U9NaeDdY9RCv1
ZmpfsF5y717olsUj2O9TyM/cfBEwddXGC8tR04kkUItIH59ZGhjqe5UwS8O99SJq
ZruuJZO7CR8/lJBQ+81NR/xFxWsJIqpQBhdJCAIzSotD9I7Dbuo3qAA9qYJNqEua
CBVUpM7pRko/PhYWy+/zvWiXzIcYzXsCOhN0pneLqvXFiiDjzTjKUHQ8A7X34Q0j
2rNI5Wo9yvM0cQMbKDIiMXIWfjvZwhLATUYfpQU+NFj71aG8ok5S1duAPUfZeiv/
UAfVgNLi6GOsf1tcdNx57yJC+i87FoMJwNAt1MEo0LsDTn9rwktorgX/3lTsiqsV
Vft8iw7tXEd6r5j4/VaEb/abM61d8fRFGzpxWn+Yyt3iDG0VRww1xbU+U1H8E8+8
O98GdlJv9FkxhBeGrsZhq+GmCUqEm4KAlOI36q3aAqiqOLUQ9fqL2KjQFA7DwPZ0
TbhT582AYHLgL6mjrT9Xv+ANXfUjDxPi8zU/zxcBkQqU8mvo24Zjb3p6wAF6mEYJ
FuHrgbSiErPnWiJLEZCFjQlxNSNH0EzPqGJ4vM2NUfci0eItU23v8NYSo+k4mZf7
aCwNBbAfi7WhbeXGsI81k2yQdLz7lUlUXC6oQ7HpKk54Xm+L5eUoyZCcpBgJAB+Q
sV5KO5y7EOoOS0aPC5V4+AdsBDhmIFO/L8yLUbmLUp2rlKea26pKgRvvVCWtSQwL
PBFL3J2cwP03pdsBfkJ0NTOfS4gmIFegVvLTykR12VrvqlH8EMqonbsyXGc4UJBz
+Mkpm7e+EKKl32DvGChGpSPxT12/ZKFJd3uBmkj6ZykYhzmsOF0QM5AfR75kogcB
rq94AoRf9nIWlGaimeTHHT1di7IIezzZPXw+mzal+dIpiCHdhiR2n+G60KyDQ9IE
Tb2qs2UoqLL4WbMsFxBM8VZm5/UmN8IrNZ2h0VqxDZPN/VXTGm3F5Jl3KJJM2b7+
soMV86DU1nSpzi4ojNiPc8V5WoS4tIOONqnH+kJd5imxa7pogdRRG+h96tA/l+p7
dO82ncGTkm4lQZIZBuSXrEgnxtR/XJPF0Dmu6oeS9EllYOfGXqhXJaiB5zEObyhT
LYsWSiIbuEU0F5m+h30vPiP7Ryh47KBVpWNd/y7QcBGwjpWTa53sjYB2vhzz37K3
BD7QDLUtRwtbHzCAM5xBF6WWhSYiDngUe4VZoxkjRPB9zeZtiEPb57EuSj5AQMWS
H+F9uag+9Qw/fnT4WcEtQeLpg3fKKWNtMLEoFIKXdt7N88Tx0SpfqAFfHqeb94i5
xbKh/G5iRcm57of0Ist/JISD9J2APMaSmi9d3dbM86TBwBXDGf0JQsTVzeJGaU/5
VBGzMKa+ElWtvN1D+bsh+zZXHVSLxJeMT7RWaIhAZIIpwli2M4Up68h6a9/oO8pI
x8Z1tBZVl5ucK5c9v6LMmNTkTG7NJMHzksuXJKKEUHktZH4+VqBI832vkjYwkfo+
jS1mQ5tItcdSEO2PcCs1lkkph/pWaQZYhsyR9jycFgZpgo1oa92d8xfaMes6em8c
e4BtkmFID/R1+PxnJ2jvZ5gQum+PAY5shDtxU59rFuDrhlcmEOXdmNKPQcJ2a8aj
qL45Dt4f6v1PxwKAWfA9Oz9OG5eKZscQmyU+Xu98AJaWMQqdEJbZvG60UhCiZwBe
fiEIyMzWY+yvDLC4TRM/n2dr/qiTdUoUUw1KU17BbzK9Dcr1adYQmW4eXrgdnV6x
9GX/2Ns0uGl8409SiqH6dBVashGPsuzj1ryE+nC50dcTwpq4VR5yo9WuZbalfLmn
8FxCW4I4QdefMbiJmejdBbypqmLXO5B2XobRGB2uIeZC4f59V+RRAP72bDuAUEOZ
l3VP0mHeYyUGcqR9MV7KCOEnL9WqhQsYltQrX1cYX1/RGkc1xL3XcB1fzQCQ3Rfa
Kw8XSYO3fye7CTPcvsDRbQCrS8f9cPGA3i8+pXYKOu3xAPoU6tvpNUbuBTxCP4An
aenGIgKrhSVPG7keOq8NN8BL1kCd1ICBE6uvM708j/Ce/+w+A6elP3pcgoLxsyQ7
tZZXEpCE7GBn4EGpmQrE/7+F7vRwEXYStmHBM0vRDxhDqM1WKbQe4hCXpZ/rX0+1
/7GeW4IGZta0IJjsgGww6FZs1smfp2VG8tSS9wYbo3QvXCFkaUVjYS6CJ/QXABP6
4YbAbqS1dho4s5IDXqPFjFLa3ZIAHhdyIwkHP0QtA0GSE0i2/Z+6+PRaFlGOndgi
aFgGgDN2t9V3GLU7WGXUOsUfL4KMFUvnsuhgQlPmGENOr+VXhdGTENnJNKi9BtzS
XTGiKRwmNhfHmAK0p9LjIf+kar5dPWClvkCqYVFdnJZRFBkAxjcyVhRydkA0jHKJ
6tE8jm3f20JFH/wMXN19u1wvwfWQFr/YO2YOF9QSRufcbHN1WUDrIjcS220pOhPz
P/rHJIBEJlhsagy38MVsYVjbw/l4/0IUEcCWUHvfegMz5+24YPEFXr8V6vtDkbHQ
EI08s9POR0GA7zy8Dr/qAyQHpAFco9NTOQ43vk/gl/Ay+/Wyc0PMwW30QAvE3C0s
2fX/cToOAxf6r4jL0q/Mhqxfg4C9RC16UagHec1KaEOSGM2CD8VLB/ve/hGzvwIy
Avodc++lbrV0KzZU2gOk3rTEsMy+aVLoCAVsqTakw6TQAzKg61zG6N9BBD9fLfUE
QZHDpwyPGy6CGt+KdgjLIzLJC+ix+zuznfaHuw8eQ3o8ynRvGPSjOcJM5wF9m6Kn
IdkqHmuEmYc4orewpdcx1Lczp+aNKRxOejMZv7S+4quJeAGtMB4VmU9AMJdsSVBA
YDZ1Zl3RZT++suszfKnM+P1kSXzVynDeW6vqQh+mI4dnIoVbm/TbWOprixNsmSWy
kuSBKmIDBQF5DGw1k38+YzOhffX+HAJWyj7lK3VzJbz/HEcU0weJ99b395q3EdiM
JRCE59OYsrbEBm9NhiK5eVBcYcqGZwrJ2wZqLCDALXUxYJ4g9iEYx7cBukqK3Ln4
dajPusjWTmIDVxeosahh0gp+cbWrP5i3kCpWDKIv4oUiz4qc4j0GSyn1nruvcNW7
B5l1K2WtNCVUZiNl5CFINJ2H8vxGrzktpjajYD75UhRNBK2fvVPdArFC/WnMKI2f
nLEl6KuDA5A/lh3AgtLb6ChvZ7FAbTiECiQlHmqEkHBlpJICaNc+62W+jo7KVif4
63FaCl1ng+gKlx/8+ceSaKkU5nDbQXlnwbrzzc3qZ8lVwnvE+gYJnU7xUNPaK3zz
E5GPyEbR+0fMhoCl2bBxQ1CVZaaK1NSRRMo5mbSIypXjHLRn9evEj38/dtZ4yK7B
qqOmZg4tiJB2gzafXdD8zP9SkrMchzsH2L8+E3CAtVpVoppTvhdCoSdC+FgqaupE
Q+fdNAGFQiCkXfLly3F6d/cs3ypiCQjI1RzTVr5o3ZCmSEEXfQ9HJ3kXtdqD05Vl
1NB/lU3+ZC1JdKEepLDDqdNDsVWTIoWf0N7FJ8dTo2Fd3EvNo7dq/qj57COyGeH3
9ZSp63ywJ1pJ3qVfXseQQKC0Oe4lTLpU22HdjA5qIgyZDSX8N+8rFai+sGuoXtk8
qgz6rdi/4JJOQXZWERGXojL/Oce4NNoGbIphLgS7JUolBegN4pmczc9oxmNA1JvI
iDzSgMfAaCf9Wnst7ZKyHtw5pBp3i4806YR6tudULrngRgAI9Fqppl2wRIro8p/v
y6gj+r8U9//2s0tQO5SMiZMVeky7DQJS9drxPWQ5LDntSQm1cYvWsFsI43zRg2Pq
sM4INIUMppo6iyCQi+tw0nNOg4g4b7P1kk/4jjND4TIjgyVHhH9wQcMxbUpjerzn
gg3K7x/t5fOX0gA+wdMn5gzVkOzCv5f8LIBc9F0vZSopGYiASyU6mFK1TmXjNmGi
F2hbukSEvpzpLRA6TjTzigSF8FsEW/Z4GfbEKu+kVIzIPi6PQY3rrHDJPVR64kZK
T6v+5OEbsUJHG7UufjLXAcxIT1rqR4DHKsWRqv2P01ofOl/2e5hWjL3g6O1vLdeT
ry0nNH9rOhGbHRy0YXoRWK5AxjDhFYKILtAfbecU1DJEKYDoaj7hQFuZEDLhrTek
rraGSsGbDnsfTMYOpBapOyTEXURWP576AKbrm3DZ3MpJkCKcRSFxMCkwlnDFIYrF
vxUBQcE/uvKI8lMOfv8SezeSka1mGBMqJuAJx3UclTvVgIvT0fuZGiSG9MLeYhrI
+FCY3zzrGDQPOU1hO3Ah/O24rveMzCSOIz05NnoHjXeVUUVB1DC70noTzE0qMcdP
bFsJjaoyVxXBOcQE7hDzaMFxcBgKC08Zw0Z5DBcIrWbaoA1GZ9bvlGOCW7nhZpWT
dy6nhHwuhZuxR2K1SLIvHboH8/xm8XYUD2LFG1Me9XakXvXAmtBGIDyG4ddwAebE
/EqgrapU1w7qFswTH8vxVILZILigrCM5nqW4idUpzQBKmffdkwg+MT5m0byFq0cr
UIlb/nUUHy7yJNZunRJvJlR2UnASwAK8JaObXk/Tt/2HcJpn8v6fVjwjQUdis/lQ
/wpYABBOM378QbkgBd3WNVo3NkTapnXWWtmbFkDDTnFYfjEcyJKxu6O5sgfmxuI8
aa429bOkIZPd3VuOl7juCntPaRhIe2OR3HnD508d4v7HmexSng+FaH6XewppYRQS
R7RCWibVnC8bpjhUgIztJLovhfaU+iNruF6JvgyLBCM/iqvQWn2FHf2I6hgbuzag
ZoszgdSAq/WHGMrIeDVuq9eBwARxSSciwR/SCLibq3Hynoivmx2hPp7iad/7kfeU
v0YrQDWUEuC7V/fu4XJABQd39PlSIlHeQo8snmfS5wWvoszqoaYiJVLYbQ0SvXJH
Y70m1iw1LyaRkrifyQic5juxj0qBRaSgpT9tL5mjL0X/MS92NupXxGeUF8gjms9q
aAmguQ8jwRhfncrcQXMx9Y0DsJnVlfOpFIY+J3UrBIIIQIuxNp60fbvEggEzzTac
ZVOT6fWt5oiUcr18KvNB0PKLPhGrXdmZmQ5LZJHtaReWIMx7KDJD/28yRodbNGfW
bDDaYqOi+vxpeBs30NEpZxbgW/kBO1WDTEnu0ap53gzSa4fFBa5bgVysIVYIu0+V
Xc+UCb5JbFuaNKn6hmY7hfzHWhKrr2KxgegKOiDkqDjdcVBCSEip4cweszvU1txo
Ho0idMDQZ8B+UtlUj39DfKJ6j7tlINlo6DjRsQ1vogy/xRqlw/0y0NmbLGB3Lgl4
teUsJ4bx7/d2Ybwx/SemupQKftGdPsBTnx7KWamj8y6kbRFQsgqJLmibAJMq2Z68
c/+rni8C0dNqk1yc6Vkf1ne7Um/QKQ9He/AybddTnjjlcVjIzHxOtetHZtgLfYM0
a8XggqKtZTQ+OPD0tYyhd46NpgDzEPrdHisM+ACj4d0EaM0snyvVvXbC8YDNIiXu
7WNz9mfAM2oHfWB59oL9TRwxmFWLGgBjJZMvbuaaN6kLvmXcHaj6QMhs4ZXL/9kH
sePqLFU1GaQeenrDhI9VL5m3IzY0P/29KEaQR9ORwhQey4/ukYebvDKobmgE7VMj
t9B4GlvZsI7COSA3YDOlZRzvTx8GOzsybSyrflSMrFhiQTsBQjUL02GmHfrmDNoU
ZW5jNcjDkvr2HjjOckHuJ3BuvJTVN64cVlnPvOoVnNbVRwGdqnMNBEq+qgBi5vIv
fG/4CU72fvbpQoI1yP+DpDYqS8ZqpAdphShsG3jDJE2UvHKckDGHGV4Gpr+MLfxg
8MfN9xOu6/l8SB/P8Z4j64C4Ao/KcSvILNbEUi54/hqKnYProEtpGgHJIXH2MxQ4
xWG6VO7j01YbqSfjME+SKn2RMYSsEgAiWapJb3f9YW+xJwRE4cekpvCcEv6aDEcX
Q3RlpyLVEGMtKAk1sEh6znohFMxLOK98VfiFjIiWaPoo4IgYjGZbHZBieYQg0opy
j4jg+OrI8Den26ABsSFdj/kXvIM+ShkhPtBoLTfIystaK518MaEif6crKsaCkssP
4Ye+ou9SKtdSITP7qwnLK3qwJG0O8DoAl/wbMWb+Ll8NmkF1Nt+9M1K2SStqBEED
MD8GaWY6rJLcIwMqKrVy+nd2W5sCJB4VDl6gJ28j5RAS05d/3n46qwd4nM6xptLq
qQpzffm1yVlFIbHisTl+pnbKHa84As9iEldaIqzRzFnRD8uRcIIMhXhS4ARHizOI
X+nS8SVcbQZiR6CFs8exuJo8Cu689W8b5G769h8xZDfgpm4Dw9KHLswCestTc7lZ
6SKgoYpcJweT+IGhDRWVyfGicpcPM72VGQYD0cthJw1YBEiKXmphbq8MHoRAzfBX
v0Di8dRNbxxNV5kvYY7kGKkof79S+07QLY1FO0H1wqCwDczm36NvFaX3NalQzJ0y
whMSgb19z+WepTR68zAQczozH/W7EhEPiUOGRLB9RKzsroa978jiuTMCtQnsViN0
pUVDVpLbgH7NoX4itRp89JXfgF7bFjbwFaJkbB1aATQ+Kzz3dKXgaHMyiLcI8mWA
9ou44jQK8l5HcjHcpAi/gffkDj70yhUCta9P0wZqsrnBBdnOzVgsXR4nJhViq1c6
/JM37KP8SMZppPaPRax1gLjDUPId//FMqPQtCqRvabM18JagJ/o0BKTV/XRFpyRa
w1u+lX/420oRcNIxbyDATiXsRsh0r90R/jdb6SovINufStws4TCpqW9AMTg5qdAX
W8E15d+WcrqIya7RBTJnyxp2gppkuG1S/woOTSLcsa+RLEfBjiMzFVq4MNpSGq9d
bsWR16Hlk4+OaoVxBjwfizrrjddvZmVrzoYV8TIk00gBCjvz30ky/m4CtL1cvkJs
5x9Yzg+lHB/o4LIczXqXkX2kBUvNjsCA07TA4ZCtVwXNbRlNGdYNP2MB/LAQHycZ
KB6LOSpZJ8DBwrWpq1xowrm6wTGGUhGUs9C+Tfz4muP35zaEgpb2RC1WBUhsZ1xJ
s2BZmGFqipXjYG9wHEUWRpoHnsSSFAaa/3vpwxkvoFjrSFAmEep1AIwJYDsRxFia
PkELr+KxFbwc7AHmMTcHfF1pUnHRhwfwGq4Q6AZzFNb3Yyia+/hbWWF4n35oHQrs
0cKg8sDZ80UswbFGwmAiZvajlhGNR1X6XgVeBzd/hAV2kTWeeNA7VN4R4//U4QJu
SGfDKXaLj71eooD8uN+jVmM8TchoK+/rh6kFQV4Gk8QTr8ZYdkmFHPz0WfGlTR4y
yQA815MxctLyLRzPjgdLLpyTHuIvQCM9VWAa/iz7I3YpSEIIQIRNlNAQPMq6A82o
NSDbnc89samtstmUiUQeNvbvgHdxFL/xGedcpU8G2zoavSB2P776TVML9KnDtyMp
XARiTHHEmpWLqFfIyIUtSTNYuaRYvxBMXNXGrwRR+tMzbRu0VJC58t1xYIvDXPGB
shTrhXzvwxtXv7QX2tzdKeHNGtRLQEO92LnBe2VFtHioonCRz73GSVtzyqTmgZr8
am8Ha3cL5EKKVlZhkTwOMgQeMJtvIEBB1BeoTCG/+M2nq8YFkN1YXyjHrCfxQobc
J7qoWd5b3xbavsrrdoJK1PWV+QT0twSghe9EpFtfUoxvs3L89P2kP9ugrmVYs65T
3AB4IAwUDG5XAUJOBQMWYe7tkNBSGW6pJGaOefEWgpLfxt2tyri78T+mVlOGnLrI
pvYp047ks/W2SwRYP1BGo9+JqyRQpFDN/D0kD8NEkajHyTyCi7pfubkHzhrcZpJ2
bUyi65gYJPv13Bm+ftlxntJNmXScpgXtdxYjBDyWdanHJVbt45eIcnPAkX+W9LnR
llJ7+UJT6CWvb6U/hubKtiYr9zWNver+Ri0jHgXQzIJaksKWFIWcufgiNspZc5Qh
89kb8Haubj6KFdugci7SRtbYt9/zMnhItJeU3GdMThQgLfJbQGEQsZEXiniC14FV
WSqZJGrqdYZjo0wmrqAGVANfcPZwAf3lDhK6MiGzefKXR1UVM3Aguzb/5p7xO277
R7wVPp/P2S58fV3JlS6736NEjhMr7HCvFBq9ZkJ+UDV10rPHWb1lWB+saFLXUR3P
6YwtIwhSHxj6dIsLDCxZX75Z8+ie3Hfln4Kylqgb1UBzu1gbNcXoVvWErPsT0tmc
omdMyU0km92zCAy5Oht6tWLH2wW2hmNN43TH99rfSikK30eJO3JYI5W3ujxPHzqJ
12/eqn/VfjxRZ8Of7Op7No1oQ6twsZscU9KECwCIGCcmwjk8pqKg7Xs5xH97CB5g
nAMssohq03BuxsbNCNKYZW3E6qMMI0TVEtNkcLU+a38e1DXpnOC2XjFD8IA8C1v+
y3r8PvKuLL+8aXSjdrFS4PeRIIiz08uaJoLgxW/K1stmGHqyk4eJkA0N/3LkLRvc
oveu4IMqFX0UPG5ztYFRlYYO+AQTEwprVOHh2SyAB675rqxs1v4aCHCq8AXydYnS
ZuVCdsgUUytloV3FzMQ6sPWgsgjrvOGVv99xgJbiZFzAwEgYJ+sgaaFSV0b01IJA
GDukV+W0vbHpe/LiZyRMPk/kx/rtBKqAmsjVVNfYk6tTgnY1kjdTWKnZZGgbavhY
a+gwb+MFpyXgqr8+lrWsbZAo8qTJX59f6AC7gW2hEp0RXv+HI5Yap6mL7nJAnpe1
mBY1dsO9GO4ABh7HGy1jbFZPdx0S5f3WXl0wojIrdbb573HZl3FzTKP36UidYajV
KsuPHuTl9s9cWeGhWKE9Y+Cmwn0Ob2f7NUuobaGQ/EnHLaakwFhrjR99CoS2mJU8
IBtZnqdct3jluQAWbFyyROCnSS9NAu3GjTxYv7ALCwW6E43mIaAJEWuTEx4Veb91
ZRp6AAo809YyzF2Jh7uz/YvsSerg4qsobDO5JlJnURh59vcaD+gJnDhDbGaZvf3+
f7ep6UmWy4Rn3LahDPz1CqdLNuutyc+rEFDHw6IvqIZ0rTBHFKcZEaZXljbi63JE
WYGvYgImrt6WWDZQJzT9IFogins/tbQXwrl8fnmD72ylbjcxzly9s38a8kXoc+Fa
W5zL+6wTbbi44gBtC0HnrOwzAIDDVFXr9SoO9JWjjxMD7BM9j4LaUwSNFbMUZru0
bqkMF/5OFbE/JNW6iOcb61QMBKfo048w/yX/IMYfXaFFwQGqunuBZQ2FYDmxqOhj
C1ba7oz7+QTFfxUndcNxtdv/MJBmQknIbL+Z+QmAf4WJGivWG9d9Pnjn3mUcFI7w
sFLOvQi9HfaIwd0S0wCm/XQJfIFsA3c8AFLK+GXau61Zm75lE8o1ECyUTzNNDd2d
gHcQVMZclagYfbjgOqDsVadpwmd0PU9Eh3llrZTojtT61AesuYWW0Fo4uy+NQnO6
xvUb54qIsqjiaCZRj5ka/Oj80fDsgZ2Xvl78Oe4DmllvQvXr7255+rRxGczRJNA5
7h6kvuGzDwOnJbvn1XRbZFYJ/6FwnXHCwJ/+680pCFDO+bcBgSzoWD3zcdowyl8B
kFwoOVgqAb+gZugiRsksABzFZEhilkxA68NAec0sn/WesyfUPn60zkAVrLggDul4
bK8MVEbhNEWuh04v6DvQM4BA66P5IZJJ7bnVN4x/8y9Td60PCETzFdNtsC4StPdH
qnXyKkeMmCipSUiU5q7neqmzAW+njS9abtaTconV6SEdeNDLM/V8zxYC/ZAKHBLJ
+HphfPTYVjJhHPL18EsM/x6gWwp0aA/aoxA5zKWWX1pageeQwU1wKCMN7GzHNok9
7SgL8lKuVKAkyfO5rwAgZtAD5kI1qJWmzaKDCuca4WR/55QQtDDuS9rCAvZ2KXM5
hOf+Bm0EVUCWVk0KcRfrzK3vP/QE5XzgS4MGdk0YRAoV1V1/ZJfBjZKYHZUfLesB
WEwfYskxf/nNwGGR0biPy7Nrpmnz3VZFdsZ6UU+2X50ufMBU0Z/8iZdnIQkFWWwy
C/sNqH6GfWpiWSv4ykpfizWkByhz9Xizt/NOmRzqs3vRzoT3xMFW9na3mYmaxTQA
7GNkxJn6+QgOT43j6zX1XxyejKQ0P21+Jh36z4hnEBggPySo28hH67zMl/qPGcTR
tJqZ9C2LuyaKHH8EDqmN27xt1nnbpZ0QyN3gtf0W6Qf7EJ2HrWBeCWehcmpVapk4
1tNKquFeT5FD0AY+X/JScbxi16YeqWD/P2oaGTtmiJ5lL61+HiUEddWWqg3bLW6v
na0IlyUxS1xLzTlBXUNAkmF5DslsbZlhuRPc6mAelr5SI/WM6JpivfJye/oM/iHy
pU0pVkJFdUIQEa+1s2WAq3KwI+FEdkdmdQLycjlsWoS/xKNre9KbPRo7SLuve2Nb
ivE2CtC/Ackg7deM69wrB8P+NuggfFcyh24+2ZVfbYebUJHTSrDeT/hxFa3CyM5d
KJSZ8ERd0aMW7RpyHPPVC3DsjbZWdn5GSHmxyvJmBLb8hUWAstXqRC5VPh3zWILh
AlNc+YJs11DKiS/oUaC3AhWiI4lANU5EHGwldvqdWTPrvJqACfBQpDcfiT5nBbYw
aQ9goLn7vQTDpopLfzhMAxJmukZCPJa5bQq2WHYcJRvwdX3l55vRbc3bheg14GXt
NKagLMzC2AC+8B5AhOqnQM+bWmgswqgoFhzgmVR/13dF3bAMS4OVRPpQ1kO3gv2S
bR1tPOZh7THyGuF/RvySW5pwtMP7aiEBHmmRaRMw5wpInhcb9KU53JjumNYx2D35
QtzNiopu2cPEKfZKXdSJtYW+S2VydGyclASIYPVZj4TxVhQ5fx6BS/3j0COCOnnY
7MKOH1U43E9wGz/pU86yBHQnP/UvI7MnwjSLcDrhIp7oLeLGqVi+fsXsITMFfqhP
y9OmC2s902ofkddYh5aThfbjCeDm+4VNPFTsC8AClzNT4kMKMgMZf73qOByuxQIx
0VpuZYH+hW3Eq/EB6D7ZVyjuvS4SbKyaQmsbTQrP5iKZUPsNwwQYiilZwBrWsDXH
Px3WJdnPAJlUsN9FnQuq6M+8zQRnix0fUtafw3RD31C+xwepvaawFFhyQ+JHGIlX
PAtJhetSdaSm7OmnNQMGnp67apbJ/o1lBt8Vh5EsGif9iDxZVGoZRtDGa3c+7TGD
AzAmlCxEX6czbMVyqrbh4zQr98FL7fgSJCMK1vYK5hTC+Rfa3CL0m4+pUBgdJXuW
sqm+FAsI9HELTT5aYvyCAf/Mp0f7Vh3ceV//hUisPv7q/If6yy0Oio01Q1c4IFrM
hr+IOCA2Qgk4FP+AjO7759EzFeUfyzYeNLBvTCXiE2sl/Zr9Y1FpKuP/UgVHI7h+
Fx2ehRJ6SRNuhoZR8yeTKBCO94waHcj1wefhM01ZQAIMyl21Ts3+GZFtRMHMFbfv
QFSrmhPXIdi3O+Lop5PKVaos8dbQn+Uwoipj44zbLjKQHc822Bo98sQyQlhl0gle
PQpsfCbyNDOFJPLN/samdT9dW0dFCYBZzZzQfTAKe6oSPg/FGvmCB26oHOh5ElcE
thb0zeh5fuypjgyFAC1nEJbqTLkAkG+gH+//A1Ln9jLBHJO5in8Ggbi6JFuhsAFK
97RW9ecMbsRKrKgmHZAyZfl3SUSz+sWP8IkVFmUG5YaqIJDgquFik3BkPPaWPUj/
B97jKa0aGXUnV++3ADbBqs7G49mu/H9oho0KpOn4t+8QsKrRcmY1f2w5llkYpE6x
fgo8u6Po08EzDZlnSTpjIUIXYmYGhXbHatVVxz4+wHB+QwdjrJ+gq3SDSzCb98su
7v4JL8IDQ9LiOi9nL10YTOS4VHz1nQHpuCyGvz2SKa7sha+9p9ebXuZwM3Q0kXoz
L4a+dYyZJ6rxIG6WV3Hr8bCoSO3zSaYk884z5ah4/iShHBSkQdLoxbG6i9TSxz0t
KeSM5JO0FnuQ8z2wnyrA/MnGnjbXRXeVzn0mo8YAXjhmmQKdWTNf9vux+/35QdoN
fxHcv6RMVH4b9CxwiltGIVFu+lP6zXO6ZQ4PbG9Pyd8ab8Mt2OOnePqhBUsUL97n
KPxdHoeZmylqBRKnfHXNCbF+xFd7437iiHtcTQSbopHjzO5Nwa9UUWGFjDXOLQ3P
/9nSOb5NdG/Rlv2LOnBMEwJhxc59/lgo05/FdJbA7rW2zsEJ+WvZTrHIBuntYfAM
tTIMHa3ItUhyGrmIHH2j62BSBXYm2WMBIo4tYwIg10UuoYfTwX+A63J/tVEAhSR2
Xtf/I9v4NOkBD87GmWm6NcZYrXFUm4GU7SvlaPByg3sy8JPzMlG2TRpPwPwTZzb0
mRFVOcE6mqVJi9IbUNwU9xuSCulJUXsEaMyHr1rToL41XVoRsb6jp6w8MA3RLe5U
k/JFMWhqojEg1L602GzWUbcvAI1ZJnskPRjEuvyI1QKzxjNluVE8bHu39gi/l+W0
UsgDcaHNUnRBlv0o51WUhkXoxXOg3LxTUVEcWQdcUg/MUeRrTwoC1SmThg7/r1kP
H0nKJd+Vbut9MEqg6Jk1ZlsSzJrs3AZ+j9lUZJabU67i4PTpXkwlyxQ6BdAwPRo3
Zl1FPNUdLGHGNM+w/16FqeXid+Rlux1fG+/TAVQUFml5xHwAGDVnwaKGQCoQxPt6
ism3CafEeLRKWrtuP1lUr0sMNOA/MUBRm0JltivTj4Iw2JvvskScNDRPSB8auLWV
vklbX3oANi544xNH3Fz3Q/gdcNrSIt5WjxGj0cYFuwwheoFd1oV9r2hlGF7LqZCd
4G13qzhcMYA05jYoYKDUmG4isnox5gkyypXuLDmMFWgQFl9ONVU5Lmi5wiEwfJwW
rPYjGU/KdRtMb5fpbPAnpxnwWNo1ejDuT0Iq7GKLAE/ngF7SbUGa2t1p6X/D78IN
yc7dWY21vTlX/c/CHT9ITRsHMhzpyTqTeCoR5Rc167qeRDirx6lLL0J7pKRIADql
qVCjYSnw68nOvwRv6bYjod5OF5ArgenGj7OrOhg6XfEpVQEzMxiBzSFfXdAXjr/p
0RmhMUGesGE9AQ4+D8Y01KW3MHTxDX8hzM4g+8f7kdzjulkSMyjCcvLumFqXSHaV
icAJ4TDYRDkCPm19oU0XH/vPOUxpuEFas1+d10vh5qh5TqUduS374b4+k9+pmj+m
S3aWLWmFLrwczVSvMUInKiQ5iED92bRB1klHLGAh/D10vhcEwJ66ckPSpIUKbLHl
GUSOtkwoutKTvkGT3OMQkDF0whGIzfCQGlvuA6pYRw5AEYZr/PtfahzS3LPN9aVq
BNQUhSHrlIOV6vK4ThXoCBU2KO01rdyL+EdpYWGovCv7o2HvWjEFfZ0iFqV4Uiwm
nszYN2R6XA4wElRNzPbigqg4wUFjlGV4kzyzkEGLI4FCSvuuNDeLA3lOGGMWqWEL
QOxOLdbMfMPP/7WDeIJDL1CVuUQlwFpiVwnVOLqy6b9newXSj+I4Qk/RmIEoS10n
ApxztBYcUiCHFg9xb8C9mpggEjKNwwh51KMBEiRZIaFRxnrmCEuuVI/FaLqothrx
74Qp0yYcprCcLER7GWs8TonHq9OZRWv26LR1S9IoM3QPpcn2CovQlYJjPYL3rzxf
W/RJRHVPaS5AvaCH9leXpdPHq6MJIpMfB2xOF5IKmaz7eERQX0GURBn1PQTIDEqa
eym4+c1UQ57aqBPJ3hoKYY8P01cC8XwJvQc4KfJTOdODbO1N1CaJLgbxBbzPmUf3
ePdRsqsHXKA7zbOedlLxMzOHYVRpol488veiW80nSoUs0ZCukncx3W15T/qQ2Q/W
EnKLocbA7waCtzyCb0383SdkoEXkjEZtLSuisZnldQOWE55xPvPoWc7VFYkWyD/u
MOmT0Mec24JlNqxSxjO3ApLWmoJLaUZUHy9Qgrlm94kPfJ7AzW41uh0iUqbAxrt7
VRkE5RrKc+PthJ07//wlLAjGXhhJW/mDlFbOUWdbrVGawWdAemzVYSy8Y2MnwM2S
MQMbY9aWqEaoFBKOLHcQsy6JtxWtnc5r2s3umn622GjzH8Yc5vt1ZvkBqyfkH9BY
BAG2OOcEmay6nlYKrxtCWpqVfMcfcg8kupI9Dg8ZOSUhUNBuuYS3TCeRyAwO7nMr
mTT2LQa3z69mc8OYhebpP3mlIeCVMWVxHC3Hj0sf8WxszEdSSR/ibR7EuhwErtco
4rWsL72aWrmNGu6PlYeYPQPVGj0DmsQ4RAZ7t1hyHo6ezsnpyLu2DcYn0EDJX9P7
muDepzqohmDXX1fk1vmnUkVRsiuPYiqSzwpUUCevrG4Y/oSg/bHuD6D/FkLaccQs
5vzHObg6kQmjY9etDkDqH680bVH/oACbQmegnQjHAIeOKTIfPe8XvgM1tgEf/qMP
HTT/8u/q+CO1iBJImEnelABPq0lcssNA0ztbTh9L2fDaNCGTtsk+53z/1d4FbQoU
GQDHlsCGk1NrA0LwRaiYpRHGfWpo1cCfnp0od36C5j67X93eCu4dypI+7HoLhqgX
R1rOIBAmyOP0W2KDcALAdwxfiOOvvxX0KyNbknRaOmp6dP4WkuH2rVx8gDDmrFK9
jAEy0hEUYqSiJXn3CLkM0W/gyrq06YIj1n9HtzSk6uyZDnf51pjveuRWKGpYv40Y
cnVudn16Cl1byZgYqb4sB015MoeV0apD8KJS71EwaLO88cWu2zEs/9fXAM1OZhwu
TT4HFcPunn2ejGcqZsBy1wdmL6fLUdrjcZ1yjk++XaW6MPLo3UrHZ7FF3MVRjcRP
mxXuP7DcMzAos1YMLwlKkRTAHS1PMMgPWBKI5glugDWc8HS3wU5JNaybYOWWXed7
R08u1kONjamIVk1Oz/a5KzIEQZyp+iL9FPXN9j8wHulhTzqU3twGGdJCKeNs48J7
qV95mgSLbSEGyB6slpHlPpGFJ39UwfbLp4AVcGik73mOhioSo18MJlH2Xtcle2mk
Dn5Zzck/VpKR+tkBDjJco36wkkM8mlhh4kw1BFITW6ZmZ1ed8878MYqcdPn7rV3w
ZES9+ZU8W4tOa4XXhZaw6J4Lddkm1Srw6EmGwaDCC8yBuZV3QZKFTSOavg/mOlGN
vU4ouh+U+Wq1lqqQ9rrHkfHLPgQxqBpdP5YPNQFw2EE1qEbDenL0ysFg04QQ/tq3
ToNEENWNr9ATbY6eCeTKcZAIOYNpZwjjDWw8z+1i5AJLpJ+4r949R09oSO6ZOMaD
ZDEr0NPPs5k+9WyVhSs9uUaXDigytIzjaAZDTN65eOVQVHhfCWv71hsEa/tSRLc/
gugmhceP9inaJ9i5I6r1vxUkyyVTTC/C6AwwMSCNzIzVYdDpJ4qJkhne7amKFoO1
cXxOLXNXx1q4Ai/X9jVNgdHsO+ZW3SF1vuCauUwfP7yTYHv3rGFza1tIsMAPyCmd
DGcSw04L4Rn5K9jaSgzdncd5yoGH1oswVjlQXbqJjPTWsZN0acVj8omnGGbWgkkd
drhf/svB8/OXVRHcKnPeeKBAc10UNkjzJID1rbPPg/golIG+Cgf06bnJsI9B8oiT
nGHfsgdQhF3gfM4DMIPHBZYCIknqrC0OK6+I8AShSY+9q5HYIDCye0/Ctkz52toE
h1/iGL8leiZbLpO0NZIypJ6/ug8CyZar002KNZALepVn51kSmu7w+0zHGDpkC8/U
k0CynWTlR/E7KuV79DAxtxt1nfcJ7Q6npo12T2L8dGbWPorkvjZ1L/5TkmYoJfX8
1SLqdoaodGugfT1O+95EHjt7FFAy9VX0IuqenUNjbq6pZT88S8GfQiwzKcX3GcBs
BP9pq3gi1Wv95fNDCg4kkf2AvRu3UMxhi9osm/8ewfhAm37uZsFV2bt3OR/c30Ah
wadte28JyumYnKYOpNbQeCF/P+wEufrwcAguHmPzOFfb4FQyOWuZ80Qs7PhNYFnt
ULaeu9155qHGEOsmwut769mvrriNu6rjSEdOVktMqLtoSv5Sux1D75NgyFsguBUk
X5H2kz3K3l5WN4rZaaoAoUnpx89IQDhsEwlco9HgaP+cumgX+7SuB8nFnE6ykmem
rl77DruGDV6xKjFvMlh53S0G1sA2KOikwZe1mH9uChtciqZI+0ZuzSiytGdLljS1
z2S+4t3Cr8WnUzL8dgUNMnkEiXWcxPhz6pI8xun6l14xIU0IDkBbF3rTbf8p+kuu
3gQEU8CtYwVBjCK5+fE2TdPrj8O5qekDQo5pY6VoslwI09y+ppGFfeP60Sq3Y5B5
1sovFNzV2xgMhv+svaIB5awgwHeMXuhjzN6OIib7JxRZ1WlpEk2RLNsYNKnq1u+N
bYWOsX4w/nHFxVYWgXZ2L7iIACtQTcgQgkZI7mVO71DfujGC4L2UCyY/qZ0cJO/o
BfppGzWTWE/5vk2BAfdMDpgw1Avvz2hlYO7rYF+G9WL70m2ml09RdFno1UzYuXPp
V3r41KCVWa2vWe6OdNGj8ghlqE/9yFGsLEreBRoaADDqggWk/XT5qXF4m7dgXIRG
jeqceWGHiYkj5C6XREllCEsuAukBaee2bNx1ueayOrkxhBfrTB+Smc/yu7CHS9/n
VEx/nBtWwzHoIW+0DXp+je8/iZfDAbo9PcdLh7W1mEIRMOt3/0MzLmNCjBNwTcBs
oTM+yiW+5uEf171u91t4s8Kh0eQ70r4IazXaXP7dQWws13XNk7F+uDi83+iN5ldN
VV2hhSotxbefWbMZRJ1xliZRT2RNO7ApmKcDf6RtD371hpDLX3Ju/YH8U3KgiKiT
j6W0U0n2YNAajjzlE4Uc7ZIEHFiEZIyB0huoInxBuFhjvsZhktf26m6sCX8J+0AK
DRshogOKscbIXhqTekzZwI0tRSamkdZaIox0FGwYQnwfSc5Q6Nb+5QZoRvYOZdte
jclKim63WCXCAmAn3o24qFTLj8fJDYO89RFCwFqRkp9Fs3ZTTRrhxqQ8VDGlPuXG
lXmORn58Jnv9l1Fj4Rj2L7aEXW59xLz8wkc/yzf352e2Cyy+z9NrCDt3SnWetVGY
c5pjENkOtLuZMXQMNyeBB2xX3RtgbQz9pYs0mECX9tVKaZ2pPWHQ1Cq9TxKAFhmm
VKbmkSTxZQ3KUyPE7Yz/rQTP2mfjEwhTw6BoCUukylWR2tP99h2Yy/z4dmMmetvn
n2eHO7EKqq176phAREeRnmyPoZVXgMBduNYCagbgc7gORNhJj7nqs/OgBv0MkrBF
FKa8LQ2QxFjn9HvzZA2VLxvnfmNfZqJxLQWAsQhuDaamhFQaRSXww1HEyPXM2ah2
I/iuiehMxdsNEVkHXTieTF6zgDNseaJT1XCxhRrKZpDN3WtSgELGxymEKUbidVdP
7UwO7jVUDCTxBXysQpA8RGpDJZ4ZPglzZclFthgRa7QY8sRuYqHC6y2IOI8fTnV4
N5aAUvjvLFF3fq5eHhAFY88DzRstNn47+rrR8SSSHfZReCH2NgtggvoKHtFAUhe/
T5aWe1As7ru5hmfSSm71vCjlK2KHp1h1/dyOoJu1C3rRMDJE7aaAjR9b1LCAtOt3
gLz8woBaryK11xA+Kci6wzp6kLigeZJocdYBBAdM5D/4Vbvk5IPSStjaItOSOasB
uMW4rsEinglTkCcqnNWw1okRN47Fe8NuFfBZC6sEHj/WI++d+Xlu9RjsYZnihgP/
ecguh3FZs333DOtOjFYw+2qezMF1RuMNfYeVT2kKQGGd5R22Jh6feBEk6bMtEqDz
l15p+SSH8qVscoSnoM0bkVLH1VuT3eX5pVNsJ/nu/lpFFrkSsfNZTnvO/B5EUPY7
0YD3JuY6tkhvWuO8EGy3A3YvlM44RWkAzcTj2sGOZsOGGKSCFcMyqioSb+jYs3q0
z8glUHj6A1WF1r/ixjpLdgW4q+3Xe2/WYXiYot2BTdIfov+KxB2aoqufj2U/Z/i5
0I71MLu6udhp7UX6MefFWyr3r1gjaYp6pkB5XH7rsYCXzOS/t1eGh7XpnKN2lMFx
nzKiVtzITLE4bKwFRCRIcWQeC/anoJZ7SjYJJP5SBVUvCsgO0qw2J/NEhNH83H26
kuZwv/GB6SqcxtkagJS4BBJQ4MQjSFZjNQLQdj1DfVbPhbkj6PWXPu9QesAJl2lZ
uLNxkEjtlYzMwVv7gbY2G+MJOAY02CO9tA+R7g60k7AMX6Qhd4FCoaQd1TpFIKP/
8Jw8hlskD5STg28m0OHF1fIonIiZY7F5UdELuhHVNdAZ6281Kug4O9FT0g88/AdJ
CBxtityAyNxoOkUxKgFBfyh73JAvZ5Ak+IRqinT1a4JFku8ageof5by+mtHxSEIW
R+xU+w6gUZ2AzjLoD/2LUHNQlSBKS81Lq5l5hPOyeewODZeubscWD2OtROlh6/uC
D3e8QpCxWlO7OB/N1IRQB4XHeGsNr3gsVPyaqciid4lWzzKd0oeK/ZmnvQ71uZjD
2s4H2jw0jOfO615LkxYqFi94XKxD2tt5/toBu5OQoMoT7xBUsUM1kRnaXZ8bgxzz
QRpgUTR+pxQnyDCJ7ifyJSjbj9mJHmob4Wby2p4LjwzY/jSOZeNu9S4gqPruAh3r
HAjHRgae4uy/XsHutqH7IaD3p753qv7VN8DXSm6vwB4PC/P+GNQX0xouVJSIqJlY
v1GjbeFI1mzdcCWQ1PSusQctH2TdNt+qPcX8ED3foSGxlC8+ARfIlMUxNAqOGL/5
0gvsdvo7cVUlpjhaA7MqQFAYUQQjHnMC/UUf7apJWwhAHSNixPi83VfqvCs/wKc9
B8KBXw05PzS94o+nE3xQo0vdDxye8JEgZ5/CCUXw7TOyP6wrNYvH028eKguFkgOf
fGBtkG89p0N0JJU9boSPd0SqIV2F3++Y1+/ichDxo19+Wcelon/ptryXmVf0Zy+B
nZH1uNVtWrEEBXXJvPLdtdqinpYs7l+RCmNPk3vhtuf3DwAG+R86FFEbNGYBU71e
PrfFM+HU5wFet31qwesZzRr6Oj715Kvi+BvwLbeCDr2mxFu+Dln3l4lH7/YHtg32
S3A5J+NnadnIqz+sYdOKCLRf1BOj+T4TODZYPKTf+V8fKd0A9gCLUo8GHfEXh/9z
qwk3PT/8Xz5r31U3Dy3/mEUF+Z/vwsGndVWsx3t50leHvxMnAL0Vevy/1OGJe7ze
/qHe9J+5iAdsHXCPEgQlU0m5g63ujyvO2VpErOHsGOsGXaE+S3m/2nXpJdry5kuM
Jm8kAAOH+mhqs3dphTJEyYvMDi5MgZyOAYxt8Szuzblfbwz8gaT821ZCBpWvgh/Q
46jiCFPfOcCjwDdTIY/sYAfqcrxq3iy5qarHgYnizFM+BEJuwBZjW8eonr69Ke3W
ZP594ca0+TyPHZH0+/Ggm7ckcz8nqzZYcFXJkVjHgp/7i3VgtEUBVy5lkWs4Jhu1
teyXm4d9EwbD4meaOwbT264aei+SX3kOklghOtWz+ScHwradMKsbMrqWuleV7SOr
BX88/7yjyfE4lVUCHDQ4G53VpYKIHEeOOe1aEmV48of98XlkMxRqK3u+cS49zJY1
WM2yFAKupzwBg2BXdoNN9KEvsmrYv3lY/BGb7MqSV/tls/G2T6/l8XUc15/INMfj
JkC8Oz0E+FmJGEZEOA5l3jIH3HJs19A2FMLXRB1VynZ7yMmHITL6ot8qcMMgS425
9jbyNld1PWAIJv74yEuui+INAdB3B5Y7A0lq+TpNocTsKuOwgvZqu5B9cfW6aqpm
9fE2FOMAKY9VEQEdYLoTpNgBpTRpZbS6GQxvis/QC6xSQaQsJwXTARGiFEfqfSAs
Zlb9ZPI3Hy1qDNkHDTYapfj4i8h0XGASKA0V3kNJkT2JaSg64xFyeVdde47ZFOLr
Kuuc2tmyoYgb/qQ9feXxxydPibnzGnqjc2MkG8V2rSfBHjNVXTw41GhgNZG+820V
rKFDTzGLiKkAPMg7l3tKjpvRxFEm/uoUFG4jMtQ4M/sThLzbJ67pmWPQ1m+F60+A
pdz5JVuRzdx17+04qhGOlRfvWuvUMnlQLydS8coBJmyQ6EzmLoWfqnXSqaqhj0N0
3uqzfi9DjNQatHGf46OVPFXsbpQyqlQgtlN5xU9Tukfotsce6VVqobI33jCh9yVv
m8NJu28Ibfd4C8A6Pc4+LqRvSlThap6wh9uZNYfKxuylb/DthJzqQn5W1kbOwGg+
kCTuuWYKwB19Ly6KdbT9AoFMolhSAXC10UrCVDpWrocpOgmDfTfOZZtConJBIBg+
o4yC6jIwVp4pJh7oC2ii+FjMB0wONQRliX7yIAbVWpdPtyW3GypMv6usj/RwMrx2
LDcQT2hzsTEqIJ4Ot1GAdd5D0AOeqxa1Xu9FTceE3/3UJS18NXH0mgnNi/b/pboz
vJEgjsiqRnMIdVGKHJ9Xt/SyVL4Pxgiclj461ZIlnlzEis0XZiW+JbiN0szY0e0y
+kmwa4mDL1g8IaSThYu/564YxdTekDeGJ/emMavDgBS5QjZAzvd8LTtkxrPQM+nu
Z6YUagWOXzU2WIuRK6QUGa7EV14U2C/cUGR4J5+3u+290EvYT2diAbo5F5ac1O7I
/I4dizr+WiuCLjr5PtWNamjJt9/EWeNYHyPRDNtlGi1mJMaPK688Dyttxa9X421F
gjWXKgpbrHPoTKu0QpnDHCQc4z9sA/dTHEpM+yYuZSflrpLiixtbVUbikbijZxc3
yBSvcnPmRjwKg4FMKz4iM9PMzkT9kSpxvnvUvdZ9xm1CsE5TGhBScxYMOS0PU9jx
P16vhR4Z2Qw54iABSHvwKuLZjT2VK59JYl4CSe/OeheRXZkF+YuqfwFd6kp12rvD
LbA3Qr0iyQaqmqiRnQPztC+qj09RzUBosiE95bgm8mq+Dc85P1Ryq9ob/luk8CLB
+tZr3nY4/owxzUmqhQCg4Ron7qIoYRL10tKoJ4BX7nvMZSXOZmPk9Gu7tnPw/YNO
K0Xd1/pim5M9l3rS+qXWbfedQSUBQjKww7wcdxvYCWgiODBjeuXjDQMpzfUjrT1O
X4ihcUrbG9LjRiMBjecikdPoqKwsrEozD9VVrx8XTw8oKhBlEyHK+bEirGG2aLSg
8/a5b7CCnImWKe/PnKoeomRvWcenc840JbazfxdWb/mxZwqQ4iB2YxGE3f/p0dSy
l/9jUXjS4HUjcqBWZhUhvOSp1eDEGUFMRag1JISQH3WQ2sFglkd/jifTxToBOpKP
w3FdJd3q8wv0mdK76yHxecXzLsGy+MN5X1r14EgfoR2ryXv0CMuhFj44Wp5s3dnl
vXwFty3bahEsiq8Nrd+bzr1r6JGef/EMdr5G88K/dpG7mup+3EYGGzXf2yk/ZpJi
lSSI+P0X1CzTv39SyZPoABldrN+jiD9ZMRZ/X8dgdpyPZBeeUW8iTM7x1vdCBpf1
cOLF7cBLZYkZuYLdtYyM4xWFUsum268Fx9w/hdCWiol9s4f+RCjdVaMIhHz6Ox7f
xrzICtaDm+ygc568zSXfGsA2oulGoEQ93BGKsZQRRyWqI/Lkjg0OPJ4v9Kcazri/
jYekuIM5yxYCXs9kZtd8EhtfqyfW3xRrG3wCFqaozXCGBjC/3sMq1z03mZnnNHIH
eQF1j7Pkagsw0ykskI/aT5Dz+Ucco50lml3SeEyBvo8SXdsHzCZ5Vro32N6fLNiI
joSoQhSnR6ZWgrm+mzgvpg4RSgh0MnHNCqqgNJEqqj3BgxplolggcKhaCHZED24e
MSayPbsKE9DU7r30zy1DapXMnm1Nmu04xLN9ymy+PEIqZcOutEbR3LYl8MEmm1cN
Mxxix7dB1YfO4MIC73reQEJ2CQI1K2bG49eRzbLRfhNiAajSFV80CCk3dQ03F/MA
dFt9fQbL3Cz4ssp7Lx0cttzo8ylSB/64GXfknnUOn56Z2KAiP3kAoQkwjr0v417t
7+pzGPLj1rI6NectmPgXEiH5MQ54ZCmfoUW9XpVJqn5ziwZ8i8fZjhBj2Zgdzlfs
GJFv60s4PXkgMjAgmRS2R+jxsFYQjLSzqPsN+d7xCcjLJpCCVtiqqTogSF5r9x2S
3FA/Q6jSdAqP0k6pob+KBSUViDGXv1Ra1NOuBCn4DIn1a8ZgZajJRyaQ5oJKkkBb
yjzAI/f0PwD6M57l8oHWOfEBTpJB56yzRVjELJobTIX3K0g+XJkItln9ddeIcmfZ
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
LJWcmhFqrZ5PsFhvncnftoQLSM8QOKtGvA/WAAVw09uQQOOmxeINctCRRBDE2/Zm
JWEcdz54N8pKphlpqW+tDFLzcBIY7+83T18Q7mNI6Uvd9L49wOUunIDWBjyTssIS
WOr8Ct9irm8ggB9pqhDLLGSdyW+1UacRdW3Nyq86qCU=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 2320 )
`pragma protect data_block
iuLFsLwmzvuuVcUDrpOSb1IfRspMHcDlC0+KQKaMwVJYyDujn+F3k2nJADqzXlcW
ToHe+ZS0M2CFheebAge/W9+i5tD1VpsOABkXzKcdNwoei1iuJME3t75dE1/7/hqk
oYiAy6m1J2ZI7GD2q7wyieGmuDrU1waLanLlmoFlkb9193Dj0j4J/rY6reXX15t7
dvOzIHhoE6nXFRKZEWd4Aoz4E357WcEj5j63TgybYn0TZ9yNDytZt9P2vgYYvKyJ
lOX1r8Qparohu2IgO+jXnHMev1eYZKXMv/CWyL2dg555Grh+kc0I4pfdr2IrOsfn
4LSgpx8xj0ALqScycGMM+kz7MdvECzJgC7Mea4okK62XlOVxYBKT+TgjuJrN54ca
e0h9w5FnLphCwABEfpM2CUXMgI4Q0VE0wkyM9bGmXhmm7NuI2NNuhBLFhNtum/mg
Fg5a9jJg7FaTAcDqGsSUIOkXYNbBx9hqDnQA6mUEvNIZFKMVZ8fyjfaqH7fOqqcY
kSTgnCrY7bzHt9xepG2Kpx9GbiQ7gnt81mm37wQLsLzHt2rHat/JjPub837bmUji
lxf5DQj5c3pMXxi4FcRYC57ewaXYZ1KaHhmN+rlyFhNstD8PtdlG2KGpvpaGATzd
orXjI66huxzpjy2qOsAMcSz5sBi0M7485Ih25oCX4dKlX2WFwkGm8B7Pl72dQDix
En6bkdt5PSz/k4bB+Tz5RnyJARVWkbiQ8Qov+J55Zfzgcr4Isp+lCO6IPEvDzwm8
cvxYmmsPu4qZsImPPyAUwQnfoWaObo/RLb5dsPeomKLkBnZoRXb9ISogxfnvSBOQ
DHYEZYnlVuDNwvOiOHz8U5hECNw+7LA49JyB+akS1/k2lUjkVjVj0wD1eQdTxu34
sdHhWa6by8ImoDYEwL9sO0noMHQP89KEHFq5wp8D01OpYRASEX1Sn3Nd5zC+LUjh
nr6sM4Btw3P0caN+URtK2IDpsV9uMyWWsDH32UajnxfVZ5hpizTdEkOzGwwJWlI8
Z41YB30y6Lu0mL6i6IX/Kwoi7/EpOURu/KWtNUAgoQ4HUfSh0595IeegCuXpPjfO
+0PAOCbjpgsKuh4Wi5e/CqlbEbpUL6NuAkMHQwuFiJTVs4ka8x3LTPkLs26Fm6sZ
4T9PHaZocyx7DCHDL9fpA9+rirWysDbtP5wNadVBDUzdEZTJ3ppI/jEIBtdK8CXg
xLWCq4tDekLAicV1vF5PzYdAr5ftrtzVfqr5BxjkjYeXrasryOc9XWeKpUojmLb9
YMc5HoTu0OGcDgbB4CEOTL/frnGVcpqNEuwB9IjqUDs31+8+Cv09D/RQKb5bq+Vi
Qe30GPIL4RWb9NSweP19bDuKj1smqlUgnW/Ja0xHipD1qGmGAYrNsHpPLhv1+WYb
H1oBa3qfZE0za5dKbVdbh93e1CpuFY5mC85S0B0OTsC/HpcFXVcilG5fJMM0cfjk
BwKbjpjvq48omjN9/0vTZbE1CQBHXmxZoOKWT5dWTXGNrL84MGkBCjJNhN/eF8nz
+2zCx6ujy7WV7ckPXTfLtYqdfeH65+NC48EhGa/Tvy8mENKiL4eO6/5Pdr8c7X6j
As9QtlXDSal9V0N6mQSU1bSFCJOwzxH96pAnQkgegBqUw73KSMnzIjWrOq0I7FwH
YnbYe/XVRTZM4UniADKUbtCJrhYPtAGFBfPjMsEBgZ1NdqTSl1uYm+7l45na5/Wr
RPEvFRbiADyrBKaNJY3OZlzVH5bDLvPxzY80VRbf2gqX6RAinRKbHDpJSZ89KkBc
3E6ArxVCVbNQB7LfRHJ9EdJPFlVWmIRb3v/80eUkwp0GOKWTF1kCJDyJ5cYxdc3i
yKadi2Bnf96SRYmnCGAmvMfBdK6PiX7WbLL4EohWblONEQZ3ELAzNCD9snWI+X7A
0O7TDnaJSs0jCL6mbTMcuCzBgmnm9L+HWq/KukltMH1iEj9gkE0mYFzwsev3JpND
2IuWpia+6xSe1uAW/eXgrPFXuzBVUNeqg/084Iye043qqfcnz50PNLLXF8nMR0ap
klOrsIWz5K263+9WlzMDIf4WnFpiDe4Y1GqaBQhOAGqGtFUudUWvk3cBKOKol3q7
VNJjgMuYwK5a0s7hql1nEfMdsegPN0ltX/LMKqvOAAjYdTEhLOkDATqrZ2yyq0Y4
SVb/BaCVQHKxtP1uzoQCGoCI/Bt3GSCCyHS2zpk2cz63YokZBsKNlfMdVYgNZXWa
A10HPZVWaUex6dPh7Z896edQGtvvwy/xN/FW7OrkvBKlagzHykOrzCmq2OsV2TUz
cLoSD8CFhj7FLBZg3mGkqqTR0mt836x22PgwVTlNlLE9pbg2y6KYgq8o+5rSqVaT
JIBguCZBXy/ftGrAKW3AUYAwXZk4LCshbr5kMrxXzI4Ff58bx2/iaBW5RdJoqYgM
VoLJP9YcHuOXRp0MIYFYUaFmobuqk/vLNFTAxiq2Gi//GiTdAntwvgG8IDpX/PWu
UYEi5PcgtxLzmF7k5ySssrMBLqNpvOz/rIGxcCp8zQzhP8tA7kUKbvaXFo2ExKGY
LmSJ2R36f+Yf3ygMFub8bypYGB4Ls+KlA4KcvWCnHH83hJNMqcrX/bBILntWHr2l
C1rii/zqoRNvQsJKTausfkj5mOI+qn8yTVLWQe+HbP3FZ/mRChMA5HuYXHIu8ddx
gFGXn65deJDopJ2+KPc43WEPEzlTGc3TNuWFK0UZqfH+airnA6Kvm4EfCPTTZaEV
aV0/iJOU+7FaWXtOfU5c8eWpM+evBKeteLer4iC9dOf4AOFCk0TX/FWVbEW9OsmF
huQ2+Cdc2Z+4syZC1oL73ZjkVwLdVmqSVZEFCpQHhXJLR6az8emg+wQOhoG4uabE
jw86YoyQT7EgbbrLD8XEzCb2L96iLIHi5BvmrqZ5wnSzFGVvG0msYG8MUqmTLiib
SPqiEPiBDXxs7xuqCYSpNsgbVH69Pg3CCsOMikOaK1OBZfErk8QZmrio2wW/vPsX
bw+DtKOIQNtH3iLi9m+6u3mn3khvEyPJMtXCWdh+Hx2YrxmrMUhIlvzz5Y6L6eki
p7MavjGF0ULgcoYyFy8C8w==

`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
agEydCaadGuzHA+gyAnof8LgEaQ1l9AsvlYdZpLsoxOFsSjRDMofjIbl6ZzFzq5r
yUPTaayQUH7OhsFcOhIUHmaM1+a2Ufx+hXgQwamX91jVrmqPCWmbvCCHXtXq2iji
3Z1Qq86HVxUUOoms39KEhWVGWh/WEkscdSL8gTQcXKI=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 7472 )
`pragma protect data_block
uAlCxa7nej9B9BryeDtJHqHn1nhzMkEO23qDocmHJn5GWK31R6TZ3pTdF1/IjMmN
sEQdthSxF/kkaaMBejdID0Ht4r3Uk2Y9mUComerjek2WkrIfCS3pFn4r90kKLNu6
1AyYXTd21uSFoNMMRderTHfpxgX7WT3Z8gNml8jHl+7vm9t8XtsecF3k3ivJ3whi
4GFHvoZqaCz1n1VCVQdCieUOXPsK7W9amTr3v355sBhtC+oOuZilcCJJzzjEuRso
I+QFVlWzhoxuuDcCJ+o8yykUgC5uZQGMH+pgqXHzzLTs//4KeHysrSyrMFp2qJE/
ZSV67ySXRmYkGeIt+huaRj49T7eruClxqwCiq2E+ZcHZiVoPgZI8ZYR5TR4cIuYk
zAzhm7aRPA2yppPgezoPBYnsonWD73AS9UK+pXZOpkp4IUOAoDwZO+tV3E9hzdEi
UnG2L8frqRv+kIBGdAlq9zAxsC71TwxxUFu1t/BPhrduPWUk/nsMjCHxs7UgqFpK
v0ed599ZSr7HhLfotlyz0n0KB/42ZWgGX2nPQgzBMrLHslZ5iopJ7PPs/Z3dBYJG
aMWQt4whWp/CK8ywrBAZsrLW8+Nww276VupNS0cs2zwouPStrO2/9q0YMLVwwTZY
W2C4+l5Iimwe9Be5Zvn0k2s8wLZ9sEUVjXVQPUC5Ee5+Jdl2sJ4GNrvFVW9eKguH
RmZ0Ga2OpvOK/wmB4yMcPYGJEuTOy6Hu99b1ZAfTsLO7jZfrZ6wsSfO+hTkSxjHw
HZPa2i5vv6LsOM97f/umb6JXuuaOV2nJYhLYlhQdQB6BUI98g/HL+JiXCOAkBfED
ELz/4ZBR5yxGq4C2Aw+h/jezBPIlbcDVEH8huKi2+AMkGKvaE3PIZkIkrb+CPwSq
WPSfSa9z/g10273SP8yxcLVygL6JOa7HZ4/fksSNl55x82hwysIW+2UnwaqYNrkZ
f70jpd43T+YX/up2CB8OzV2XXgviwVgex1WqAwR6SLyzfcf49UOeelWOKu7v9NUV
DlxtvtVEntDekkGYub47FN4EsHsN0vQG2x/Xb7jGaoMWmvgm5QrAGJGErJouJLgO
Ke1jabb9lEKhK5iAFmv6EjGP6JJ7BC70GYjvH5uGxn59rL62zzE+tanu7YcqSBih
64u+i9Ua28oUi9SCsQQiuvZ3VMv6tIKT96DZA2u6T/c7hvU31jT5sYUPOdz4N+8S
CyvEdgOkjkGAiI5Ywse1s0ggPXj2uhR5zPVPJ8DijUavVGxQbioWHM1zWNnjHwXJ
ZQEl4zrohGapIfbltAu+X/yrN/fMoJ8E3DTYDXa/ymd0tzzR575qd7KD1pPSc5D2
xZ600hUYeSyqEFgaQ26N9zBu07QRn6eav37Ty9QDGDvRbebLOZ+lP4xR5cTbuOeD
PhqfrwCCH3pTAzJf7IsKDEvGOLUbj49dyesSA47/cJtjv2XNxidkpNvHPQ2C449E
LfRGVfmu+YJbcSt5l4s2FvF0ote0yWizW4LaSWfpAA0XGWNkn63L5NVI3LGokhRM
dESTKjF+aSSwtMbjUtVSLVHDpxeQerP+hHu2sC/9I13XVK7d/AN64MVb8SGS3zQv
/5H1DjFRhljlB4tsP49uQGAiG+rLmpd7B3x/KCPxTxNV5dWQ74nYgg6yxwNWBdte
OCPxcY04uYeXAc5f720LjouT96b/WjiY4ap3YeGG0Z+Eyo+VvoBhDaEpmZOh9MbL
qi38xoj0sJUXB2mPVQZp4vX2vmnBrYuiL6g393D2bHtO1HPlMgaNHcSXPuMNUvkW
3JbgVe8hf4eo7RARguGtDS9NFviX1AsB6aDQOYYFxaR2Kx8p9aiDj3r+5SiGORFx
dL7jXX8b5ViRp5mZWl+VU4f7NBYtJQApDs29MLcEAE/IIpuklMmIt0DeUjjOjBGY
f4E/3GUOUgZpAMSBvI744GxcLlgTQK4dJE4MZCD09VOYubUTwz7Ehcz+3oBCDiTJ
y2aSdqqEnx+XOmrCvsdfAqjlBNH6h/vekIzDRKxMVswP/z+G8uccTc/GXgsCBf0Q
exXsZm4h+kupV1jBrEFhvmE/qNSGCPMQPZZtMZMh3rE+E6fK+eTes/yUhGNf+9SH
NFPuDxF6Wx0Hgmtw6Ggd8qEa7c5zxPHpHhp/oXB2vVsGGCkqBz0QDHGc+Nn2FfY0
4I3zfAiXEVCjMTThcZxq6K/I0KbUTLsf3sjmnJmxXFYMn/HFxHH/duuHOjjvMjiH
NbhjD7hzWN9SGLkRrLBA0yDXtS0knfSYXrCkGro5TUASknd6/u/lB5jpxuSlA/AX
I9qUUpp28u31gutnd7V+9D9JnpUMtihduKl7IwRurJJHbQ0EenNMPRl105UCnaIE
Zig9+jzQn4cXPDZzJtWYYpxP1zsumWvnY7ncXBHJfGLhGI+MZgEWi6m6oTqAqXRa
guZzy0TJR5spNiWRldt4F8NLLTsQ5EQnyUakIjfnnFcKvfZ8ywJTxJqbLpKH0jph
VPc+H2bP7Y15x3IHAFI/7zBpgFi1gGdNSz4+KugnQxj6pQCKQzy5yQc4HpyZ93/+
p7iHXWA8blsk7X7rCQMp4Nt6araaXrr3Bkn9P9EXIpk1GIf0sqU1o/a1QJfV1DiZ
yxumqsbJe+k5pmIBX9fkIEIbLCOa7KHjK/aWNZH6cYTofH3yBNEiY3DaA+X/apDS
L7HUtDf5tFgX2btW1Qv+vVEEEsigHZOhWPgVFVBGNeDNrIQlmx58hD5pkqmbfPo1
dlU2NpsCTBtCjE1EuX5nK65QHLIRxPe2kdPfvO08JiSvYT4/YKl//pxzRROmMziQ
+SloEhJLMGgYf8Fvt3X/+KFXa5zcNlaAwhU/twvgz4N50dwrSM24Raer2OEUWcu1
mSccC07n5KIrzJFVCki/+M5es8rx59GvAz60JKTfZ1ZCwvf0fTtP+g2MzpfAeiHX
GdLSOE+Yt4JeqsKJzYgbUTO5mjXZC4w2XoQI2BKZSCssakGKYrPef2Q3vmUaRzqw
lmQpxPOMvILOHrWbYVnMAtR45AjXGzcrhLqJ35EPGvTWO0k2rLoZ5MVXHHdWKoIY
BB7TINtuoDmCDl0PegoyEMNYacrW6ubg1oClmGFs/H3MfakvrmMrhdTAhiZ2xTYy
S3Wpa+jg6iM7i3VrL0DJ5jEEz5s6SAwqQc3K6hBvfh3GUq+BnUhpNvICN09ZiDlp
74StPfKAAl5qBpg/YHEkNcJcCweoEMNn3vVYWLpOneYnR3SjY78j7SfB4ZJLcWjd
rVHM+1P3wPZYQLbEVzU3mKBhWkIdJ29kS25F3BYPB2h8vhjOX/K/kLG9eQcdpBie
LxvDuYHL2rlQIz9nLotBDy4QZ4dV7TvdDmmsSWjUSJNogSIA5xPmDnWwr0zUSNEB
uLVHgiaFol0njHiLWhWSgtXCb6wHKI3Us09zhChv8KnDrWkGQa13BAXH2DTTWYAa
k9Pv0NCXuK87/7pvVfrVd2qrbL6hQm2HxJtEJ72lkrmtoeYyCJrn3Af/IJjQc1fi
gsUHXmRzP0f2LGifQ7cj4EeVvCZXyta0lh5wSMI+3AD0UTDClg7+GAqiVNYQMkXb
va4UIK+byLVtSTa3s36zR1bUAY5LXcrthBvnII1EC5Lgo5J7TELq1pWlYomuBO4P
1aL/Y9Xk9eKJAymOuzIS72HauUnGs8vxssF4tS4LpspLt868+Ju+zo5U7cw5PA7E
dObhwAoHAUbSpiW8594VFxAeiJvr45/3aIIu1AivwvkKRfqzgv9NtVDXb1I5rJ3F
xE4oxkF4OZFzYobAL6R524LSVx10VbT3oj4QBU7ODYMI/UzXJ1RKPnPghmgYlaRh
9o+W82UBCbZ743nyHlnzEFiTARIvXriCkXPOd9PH294+OEX3UbyK7a91fZqpklWi
lDkdSZZsuYbjfNIjQkZR4f/rCvu67Jfsw6oRi2nrk6hqeOd1CcLId3UUO11Xzhyk
GCeyK5iOOb3h33txzOLT+L7Yn6MVlYbcycGhtNvl8MUsiYJJq74EAKEDD8q17lQL
7AlzhaDuCK8thv+F2MLElGCSSykRKvRwV9x6eZgHrgnokhbufaxoqGbOtolaBeRP
OjWai10katrh8OqwkRWuB9P5A9ZFppE8QKyo9aW2LqUVSdM366shkvZAQsnduNJC
OvIDGl9QPqOC8Ej480tSfRU8k9Eb/YwhYbMCnsBUOlRdu80M8skmrKDPaa7CoaSc
xwOMGEzjrcKRKHwLf/OaHmbZJ+jxPx6b5q9XmdBcqUYfeHXlQw0o80kdaq/AB1Wk
LO7e29G9onwI3xoHSbHemG7C0vE3yJBI+Ys5WScVjZinW9NnC5Ege06s7K0mvQ2J
ONdKvnDseJGVg92Re7RY5rruWGU+0Hoqd4Zl8UcqAX4/Lf4VEFPau2CFqqEMRg6c
te0c9K/jNRa9sRFSTPmh5E0WWeUnm0i/+/QzHoJEN/NAUpiCxkcsX5luAYkH5E+2
JrQMAkgXIbgtVcVFA8dVWUnxZm8PVwEO+feH2ewnQgI2Dcxq1YFU4BharMzHMDjI
moY47CL0hyvExm6y9CmUP30h+qR9FiaQiYulDrEoCkf+5qfseFofWbUNiS4IHh1U
pypypJ84UWeGThMMONf8XskhviyFhfwpi4YzoUvqm4jH6tCXvX3JTx/MgoqLBfCS
BBk7kVMg7mmZuJHk2/U9Vg/esnNRPK037NdozNQ17NjftlX1wqb0ikeCy7GMZdRG
Q11/zHaXNmVnZZqHNdkJQ68YXu6C+8wcYMSrf9MrnPxfzWFxmt/WTiVWafEQ7bYu
7K7AjB39hJGsHjmJoFtHn4ZnxrDQjVuZeDF//xCrAi8yWvA3/OY0IzmOhhDDNOEb
KVXMEIV13OZHknfvzXyX75YBUsCcQ2JhLlRH3pTIXnSd8yEzqzM3UAMrYBduuc1m
En24SeEtUNMUOR+2w5hHNQYLh5wACMOy2COHAyB2PiuvjHVxOZYkqqIv973+UT5k
htexxkAJ+ov+k8dCqKRX7LYpRBVVOL16ZRDsl26SoD0EmAaBnADPbG6EqXQKwJsy
mrvlC4C8my5ZlnUBEnmSRycF6Mmo1XnsqMfNC3/i3HezzfxN9w9NH3/TzTFDtnzK
yZEH11Owl32dH22FlCBS1+iApuNPxcVIhM3V4ocMQvEcEVqFWuWT8/Wrsy43syyj
LJqLH8hC57tbmDwxsj9t9hrw04W0fNrTiItnUv3EOMM855LK1d6URX/rcUL6PyRw
r9ZKkqWvII/6PMdZyokJv+GDdOBfJ4tOoTz4zFXHMyO66OoMHFaQia93pCv9vL4B
cYx1fD2cElldpXFH300bc9F/0dlL3rQkLrmBIA2eSkjMMQPWe2zOYPhm2Uw36pQS
0U7Wmky4Kp9Cg2nZPucOxM6XRsqktyH8O/TYF7SE1B83ne0bHn0M76C9k2Mb7YyD
T8MaT/HWZYSLrz8sbD/jtUpbjhfZUtr2MYCodt6NAJiAfWk1SlXuPSDO6r0bUwFS
n7sWEu6TRBzamYlNi5YCdkWGtYL1BGyf1Qwe2lsxeNWYBxn57jQVZNpX2zghZjP4
K0zWr38Mq1sA1mVLxV5vXrsStAz/WVgyVTFd7DZfd5BNhAPYW8JSz+6Fx1KH5jZb
IPlv5oEd1lwEH7ln/tLAbLQGtCt/6bxw9t763dDKju/y6Bq4PLlMyt6Ww2xHyPk9
MJ4VZP9FhPWJUQ399shmkPNDXLaobFyWdQO1ZmwYBzX79p05YWdSIY4wSK+FPmzH
/QfOOavIWBbOoBRZlAO4WLp1Pm1o40/oCBMJHveufM3tCi5WU8Fb5g9dbVWhpJno
euUZOmmdyz62f0TuJYIUeSp1Cr7tSWd4XZN7a6s6WZJmbZQpML8scKpnBanx+2oh
nQ030219+e/f05kNlmxU+ZzAExHJ7Dd79GCGT+GijOcgbPKqRsqR6ZITFLqMBlxg
oJfQgkEWDZXVQWBdwhQs19pCEuE8jKUPTdRKGWqEs7H1sVa7ma7yVzKnCStbHKhz
XBHZWbYa04zhJ/nnoGRdpLZvF5Hq3S2KbLclVXgcV8OUVShTRc0KeEHHWUVI5Fm3
FkG9SBgBjw2O1YQLdoeJ1LypF2cb8QT4x7u17WXJUdKLk17Z/S4hRcNY42O9lAZs
/JH9C1fbJxTeq0wWGxyHeWkjFi9lH3qmfAt1nWZsC/JPbwBLPys9/7Z0mkvQHhu1
WVtnaOWo4itZHzeELlpUdqVhXqA4AWFCfOiHVCKjFCe2jS/UHK5/gThnJ2MIFQw1
gIINO9lT8duIGG/CKgycRoUUbw3rkoUSsjs3SjpCeBWSjlSVT10klFX2y1pvwCP7
eC+lkqeKD24cT+eU6H1sczfxbOLK2NdfoLXxAjtQhwjv8Y7ky1XzCpMiLPrk82Vy
Wtyc9NKYZnr4IN244C6WEaFH9/i67etb3X2AW++sZlunv1TGRt+tkdRm9tfE3dW2
cLE7eWQqJmSV0no5X65p5i4TqRya2VZdr4nJy97YXjaK9dGWph4oGD1SJuUX7ScP
1rwyxAI3lQn/y33UEjnRl1BXoUYB+XiRjZJmCVxovhTvO+460vFLZ77GQFku3j0J
Wr9fqIlpowk5ckT5QEfVi8tbl1KlBBrCjwqlxWYOFvJI0LXl9u6OQxFX/mGvbKed
6PDZ+A6kKJb27OfwAQAXZmT2jYkoIwtYd31ELWCl+bd5uugXWZe69atP/+kyCLnf
8Kv2OHqYIqO5j6UJGQOH9LP05Pr7+6rmgTOJGMpBNwedRWY73HL1zYc3Y+pebfsS
ij9GYMoXnZfxQHSB6J4mZuebFqovcTFD40CdBnE75P1eeQhc90mNeP3rwMAc/3yG
+nQ4qzU7Ate9Jz0KRkM2Ti+XIpULktHjAsOpcoYtx9oJqvPDflLpkcz104EBafg0
tCvKSFAflUYWNzypo+Y7QPuyeSIj1x5IkbCYUOdL0iKDs1esDunRTrsKmuQCbd7q
gr9W+o0cxMQxkfwCGvg87G+RllybAAi4sb/snVDY0/aL4EOyeecdqPOdgVPW7m5D
4NSVYxmhW3K/hiw0WEMeCAmOnUdC1oEbnpxdeneLiRuuVT7WTKMoWlUBYjnrHOog
R9vft3NrrDk+pRnXA65p83NSpB9usf1/8u0nUT+aPCtEH1fHJLz7sY7+LSDtOoPy
KWR3v/wosACXT1UbAPtpU3e1IXX4EdD4jF7fP6HadgTVkkyh82pF92q7roJqx7i/
PTWU0q7L1slvp5SSJNE4gzBFphe5LFWQWvkIBHyIH1MfGRbRATk2Oc0RTfIsi7D+
ShRx6B2UCKQiGSp4vwYh+3CoSEH3XaafELX6WmNHHlwdNd0PH7SW6fBPVwLGlsTv
Yc8NSzb4L7+SuuQQt4IUjxezoUdqIblNh0R3Xmp5Qy5vBQPi1g3COpY+KFwqOixQ
J1u8emDPRBkA4bM7iJLrW+EAy3YPLm1RSYxqhDy5A8RRXSpCy3DarnB2ssjmOUtn
sEu+5F+uO99qj6HFySnJL5BGs14mQmYt+mxkFzuf34Rz/3QuU2ZAUANEOG0W2YRa
RM/7XWtChdJ/utWveWnw/I4t4pDtzECR3XxGMBgJ+DLZKBb4qJHJetX/f3ky1JKm
C9LQp+H6cQ125VlTm/nuw7n65BywxDrVSMkbJxI1p4eOrgILihSrmDK9IBSGihB1
fOTPbtpM/fSnrx1mEbQHQEJKUXeofr9Qsku9L41w/dayQ+7IDHPB0xI8L0qfZeLt
VP9ZTjGQE2e5xJPxGrLNxqnySJ75SbXDd6jpvF9+ifGc5FulRFHCgkgst3WdJukh
L235pM9vIErFxWv1GLImiJEFGJjAYb79qHokX9uzz8oM17YxUDnAE5KEdu/JVsv/
Oqo97W1bFJrDbfaVjNG9MxoZnXeQ0MAkSiwpaoITJxUqOdAmyylS/yP6KgZwkzNM
sunGXg5bWzDjlXPWqN/ilXqwQlpMb/x84no2f3eJZyotbVQKV7TJSC6j7S9XZNsb
jf1K1GnFwWougRohKJral/mUG9jkMsJxbF8I5JbJGgY/nInLpf9EYbldGcF/9h1y
A08tmS4WMECWNijYx7jVbb8AuvwuTg5bTozP6DMdHAO1n2nJhFKexmWLqgkRpCr0
maSeobPcrmNjoDod//eWcVSnLjJcK03aEl9vQKbW1kspYVSYXKuVlxXEhvu87dyf
/BRpkfqyMNYdBHAPpY5hcyDmBZxMs1A8EkvNs+6If5o5Kag48lC5cpXq5kDgXGXt
UWyWb0HXDPIB6s/21F6x/gDjlAxuJ1P+kT+5nKcs8pvlxGDES4IXfxNYjXv50oJf
7vMSQHPsHm/REfpP7I3FEiQYMtwuwR+T8gU0UzTnL2gjKzyRIX5081ipEizM1mMD
BMmXsXT9RjRuwvYCh2v1AQR4SDQ3K+VifpoWeB1nJxGz31fZXCK2rkiKU8IXt3vr
ajkapzC6FkMORQUQgz5rZFoGQbe6iIlLmJDsYrtxYWes+JDqYrCvekx8y4Ogd0Q4
heDEcieHNXf8Y6HxF7Ey2puWAAHYmipRvvk4e9HVNBcwfVafwhjn61w07SJ0Xgnw
0p32wwkSZvwGBsQ6Z06cFo+p4w/NlKrRNIyl2mgher1HbGv8aMYriKgHkUD/crbO
BmWj1K2ZLz7DP8OfL7HnYdsd1oh8hBiFk9l9Ib2gEIAzaKc+muGNXXglcfJ8LuDb
FvZWYQpCtsfY4kqvQwaRJFfqNHIkGtDcEpRN0jQjBl1Jvda6UqMPtrjDR0oxMDzE
SxxsgzqsJ4qZ+8gqDOUesZ8YP4I6Ut5z2WwJHOOn3B+O+JB/LTFNvt30j28S9jNU
wJgnT58vK7OCuCszBrYMJfZNBxgOFS0bhTzkDLNyFFv07O6++dVV1Fzp1L1IUtOL
pxD+y3mWu70+aWQ+j4IUQzdWXvCkzwUB81YNm71WFhRMXlM2urA656m5VW8EOCZr
pecCTw14t45/OAc427aMktZv83sm3PwqwUWxbdBg9oQGws/m0bb8OmCaS6RZLGAE
RXvIHNjIgWIu3Smut7OCbnP30bUb0MItbQVtARwwe050KoGplK+vBOZ+2s2tVzVM
Z2yxWVQx8HVRuBBz3bcnVquNBtx053AKcGnrWp5Xiv8vmEhwSfo3rlPYr1/qSLot
lbsUMjROMYdwQ6N6v9Bq4viFy/AR/xMMYHkqw+AYuRaelbbDeINtgy8FhGHYZCxc
MhwgaFLq/9Is23ekMbZPkYhLtliXMRa/6Hkf4PsJR2x/BfBCr0yKwv00IyZuuGQc
O8gAh2Spx6aGgcN7xPIPNissmt8yDJa3OlymJEc37gZEVFz6dp9+wnT+RqbH9MmE
7dnUugrQQ1WjcZo9xNHSPqlAsovOYQxi446ii0z4uEpZYuSSbbllYYmt6dO0UiUM
CBzA5mJYdth4c4glfY0gTAaGN8LuK0Pkiz7U5Rw2kFPi3P/eiAmft2jKePTkAMgU
s7bi7e/ke+5tcId2Qe6Xlufh37zE2MqLzGo/a4BpYwUgtP+vLgrehLUC2OSTZqjz
D0wLS0p9o04BFFUzOJX5sqz+3RltAIwHUOrV9mGJJq5RUWi9pmCEL/tvrogxOcJ+
4crmdCAmOjvyn1PzVVcBQ7PfNO70KWjbYJkVtuC81EAAKTJDXNWilFLyX0Zvr77z
6T6/7RFgyyf3ZA0a7Ue6K7g4GJgROnsSJs5FN3M+XePS9bPmuMfFZV1vdwX+6G+k
VLOqKNAeSaDlfLF4Uwyfu/45fuebkk+slyYW5MeFlkNIMS/utvxORMixmTyuuqwY
7xvkzHbEC9RMTUqWQJm0uFCyUqZFIxAMYN4T8r6ZXYhPE6QcRUPsKY8MwbCCbDOH
IS6ShET1DMHlbxjfTuG9YPu45mfn9Cplnyqmgbmkysy2CZKI3dCeg78qW1MFpxMe
oHEypJqFjeqegTkYT0knJnj5gMXsTeVQwO5ur1hNme4=

`pragma protect end_protected

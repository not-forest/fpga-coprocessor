// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
UT8bLlthZVKfCbDCSZ6tMWJccdWvxJ8TO73DTs3jzSSiCW85r1z4ppfPFLwc+lqy
Kvr5KnTng3f/rrzCaQdZRuFjbsNjm6UoJYKncN/Udu9RzhtZVnzokMdCYTxwRtYE
J3IjonWIWUHYiZedKwkVsgH+jwervyMQVHBd3xiiPpg=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 2080 )
`pragma protect data_block
9JLfqDE51QNdmKVQkvdvso9/ohEShqrvqLbELbZ1a481Lb5/HIqEHKoo8jSNnBNS
ob9kHayxwAnjsbEtgL+tcG0weXY0gRTmohlszCmPnwr0i2zHThV/gcaN4LFFLhuW
D5mTlqDoI+MSx2XRXjII+/xOiJmUG71ISUMQAAqTXNq+cwkpHu/CcmzmoAKlXiZk
qPh284LciGxrLOAEIa3khW12f6M/NXx2o3UJvT8XIF8m5R1H9v93qm5KNrbM+UL+
MVI+DqdW0Ba0A+i/f8N2ET96DPPUcfoJFb62KHLkFpVBy6aJOSYZZ4JmMNWQqrox
G2dixGnokm2K3K+9qJZQDa3kCwpjU7CxQwvHGJxZNbdl0td/isIYvd3oqi4vdynD
dIVtFD6ZTaxjC7F+iZc1+65ojaMt7Asd8kvimxF4No9Jlsv9E0vJACEi4hWsJlC4
Z4SOsaG+E9Q6ypdO4NlvOH/Ukb3mVFifov+WVles3xcWZ2nGZmu9HyStrYAfTZbv
voE3CsBW4KMoSfI9vq70zy3AvRfIAEmAjbnPc9L6JkHBgmRXMxtyL0GxnC2SKQoJ
ZJczgUPzGOuaxUYngb5AeT2Su7kYMsWFpkwhJ8DO0ZfMgW9ofYsJ6RFm0/W0MhXU
8owENVIepPiL9mgc/maFpJECuA/WL+va8TLlQJkERUwnEPcAfg6zYDmByFOzeVW8
rKFCYQK6HulWr9aFdy+jbqyQguMvc2AMseTniL2Bqx+hd/h0PJ3IMuiTLyB6sZ3D
zswbBbOaMD4Ap93BeygT9WLPRqJ28PzT2sr0JLUSMH5VZivxcYqiDOi1f4rI+Yvg
z1VxMxUF54ZkHR2Ihic0Jb99rwvVUORQQ/EBWOe+9ZwIUSVW2y560oz4aR3t4cXY
6AhGK6I0KyXdoxTixbxtC4PadiBs/pLxWpdMd2yyOkumJV6CT/qfLXaWaJzbrWVE
MghCcU9RHgTsQm1Murn7JOwrQGWTYW32Jq85p2nqWBc8pj0rOJdam4KAKtfvY1H6
qhIUCDDXmYMP5u+uGrVPPu7bMO3qUh/muTi0itgBYZuwsd64yufK0wyAGd+vSdja
+w+/7rBnat3ihGdtijdjnV88Bg0SlFi3sl9ddYu4Az8doqqfKgdOWD3qHZhph4pb
go4CksY5B17wqzMAnDaX8zkFypOLaYvPtF8GOPAUf4gFcTAI7qBC+1sCwaTvdB1N
lUNuLaXc7E4ZTpYHTsLDJ2LbJTPkWaqrk5NoR+IU+7+e7epsiHh4ES0vFWZQSsgD
Jukvjwzc4VLhFNYLNN4pkVMLqekOGaknc9+DPNHnhZRNcFLXWifrBSjv256emzYc
OhE1f3iVY1/lh/XcE1fUbmzoTdpUPaNY/g7ozrjz7DyR3U3lQk5sumkt7TOGFjM2
TEA8DVX9ZOZKaN+iUEmuS99JBPozSLya+FUZJx5R8Xp5z6R15nMoLPQWTFbB7nUj
mTnfEIGdomZkG6k4RFU1yFaXngs14N7d4i1o/MIjHIQDvcdn3L7wrnhNO79haD5v
gDkvfclEdOyEyeCU+PI4Co1hloXVhYldakN/VRuFPdyI4wypEBnNsLiHrTBp0WAE
6v3zyjix14yF7VAo2fZ7ObmkfDsw976ahCaw3YCuBPQE+qBYUUnq5nkahmnhgDDr
kif8Nd0Xvz9/TL+3HAM7QvM9Xm1H46yKthJenq+m9vYlyNZgGIF2O1DaoDSxzgtZ
G5a0ikpEiinkViQSasCz1FjwSy5y7KJYCLtlit9B18ZS36rn803k+rm5mTd6oTwa
9SZIeZHkPzOA5TJ59yfZxLhmBB2A5GowWma+OKW1+GcVzCl29Aue+d7hiKaT5uwz
4/ia7fjABEPtB7Se/76cctxb6/7sJTEOtSie0H5N8VthP/Z0V0x5mnNk12jAnsLK
AfucvLkdOw1D6hlhq1tfwMT+clzz13WjfQfqDQz5PBb9xBLux8dW9zJ3oufLq3A2
5/NUppXlCKYDjuqf2bC5eUVyklduwE3vqStBH/4S/D403ZRGu/rG78O4rZIDVpzn
/EY6ZL5/Wa6N1+MBB+VZ6GwnK1fIQJ19IHEwR/3A7hCYdDcN3LyuPmKabL9+5ZJK
seMcvss8eKgw8PjVQPDZ3M5Te39ecFTZMoxe9ue137buFfw7bIzGpfuup6CZtOES
50wEOxe59OYAQPVFGh2zfZo9lifNnVa27OvPgn5840CY02+K165xzGCk/aD4pgaG
rjSspxncuRxf3KTS2Igd2+PY6Nfii0SPM7DXm7n8nrxQQtpaJsDyohi9rhuGELbG
rN4aB1XZVFGeF3HL9wrhPcxvE9Ows95rhfmJEectJ++Q9JMjZBUeWV71MIjK5HHW
dOpzp1eDU3+m4Oj/wQ9UVPgEw5U8LtyYImfG+4AGpOJ2NbapEO8YeQacBmxfuFqM
MJh9wf6hzAyefmLAMo+LOBmfaRZ/o7YRxTI8zEXa0r7ZVWjw9bAQASyyZh0giApd
jpc6XTrw6JAbwXvdJERMrdQOgGRg6G/Cp1rY7Qi4JCrdVynUaYikuVXoPeTLWGQJ
HE+jtr/B5Y/xKSlQEJppUtG8MrdGC+fTEe9MEImISgFEMA2oZBfpB8lfS6mbYXGy
Xxa5u8rSBpDJcvyhQOISrRzU2mPENGXmKKfbFm54tJ1MoinetjjRXiGP1yfb4cr+
irXXrAQxcEM1naAb7hcqemdmCR7yvlt72/TDfs/yvPwU+nyFGptfRg4KWMG2SWhk
SVMIbyLJYtLrcCPx19dm2Q==

`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
kP+lBftnpndTS8qfn2Yhz2mKJKwplolYl9Wwrkqau4AAyHFbi/TPTMWlzbMe4UMO
Wpo8MGduxm/HKAJ15oV3n0P0yUI+jW8CHGtuGyPIj1NJBOoFGCz28Fl1Z6pUTC3g
4vqyY0qkLIZt6PSRhA9rO06B34HoBUaerk9tkhJGN0I=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 36736 )
`pragma protect data_block
8Nyc11aAg1r4MIWWcWQulVQlEB4Alwg5OoQInx9GZny2v/v3PmzCNYBNUg3Ktg1Y
IMwnP2CE/FMDLYCU8hblY153z0yO5ciABiMz/xLaSkvxcGtmEloDc4Rvd84YVWot
EDwz+zlk6ej++zXRQ+5BbimuikShiwuY9fWCPpra1Tz1IH1IpVIAEY5li/DEHURO
aWsIKMQAh0QsbjH98ikseFt6Y+jBd9u24ZhnERtwljBYr78euUcbKfHppDYqNdUC
7a5XI3u45ontrXEkQC/xZCo1BHH50X+qGMD911HHSxkRFKzIxjXEyoxhGfyCJWj/
cMLHPP42Kb8MEa+6iUkH90Itu7JBJrXjJVVtKx/c/FdH/zsoklcKUjoz2PPqJbRC
bHrZAkranS1Nweo+kk0JVYof1ScW8BOB+r9RsaxiEqRUb0S18H9g9SuDtQ9ndtG2
zcWE4jj8t5y43oDscBDNoGYh7aHYynyQe85QtQEZ3fmeUChxloewMIVOn45Iq0vc
mMCSZlthUcFKRwiwLPDg+42OyYFU/jLXoYQboucdn8C4T0Xl4FTTh+JtoHv+dU+X
xTqvDWLWScOp+io5xqUwdKj2LuTB5F1O0NY2Mp/qRdxeSA/FNQ87HEiV1cToqgze
jLud8nHI/abRzDK/CeS7iLZuxYrPcu3o79d2vXqnwV9kSDbKUbjJOBm58pC7ZIwo
nReuvubyy5bqxbGanK3aubdS/Rb3jhpqq9Hslyg/i5GMibCBXQFLU7OdDfWf0Fpg
xPhY8pZQK9PYxq+kcU+IYR62soeMHZrBVqGKhML5GLJejG00yJxRiJucQmj52PG5
Ea5Ez5HdMHLudw5x1VHdx9dRhj1zgLurHcnOZHW1RbRFIPE9LX83va1X6Z6zWSRl
55yMEnZfWLTR9tCHSaaSAnuvkqEcHKotYfY19VrNmKX58gFbTXFzCfPNMn0hqdYP
lXW2vkztRoMU2rSkNq4smmQGNC4mZozEiGD+sFRxFe82WYSeIjSJETCMsNftyYnj
BHY7xWrWZJ5rLSj8dvCTajv/vRQggEp2ngjOCq6flAIVjpzlzEdHPu0zg5bo8IZJ
5Z5smT4aFQyJlbF/XpBR4cb0qIBDgSPVCUpAnTmLRgIo3n2nOZnB9n6K02o5M6QD
LPc1wePO/TyizNpsPVVs4tIswfkVsayPgcGFtNrW6RK6RiCrx492Yk0DMQ1Y4oQp
g9oDSygyJ8t4gIUIVHFeMpyCVYaQmJPs188Tu+/xFeznmJ0Knk/8eFWz3eVV4yi+
3or6gPKzC/cM4B2YXTPXtsPr9Qba/+AKBkqWf4xFpbf6jluc8MBgBkrWbTGJh9rK
YhyaRPZgzMpZDlooEueAIpzcZH2OjmkMAHbLX1Pgoy+gdpJp+hcMW6mY7bXaggWx
HNEht3V6s3ExGnOCUw7SvpUEKOXKtp5kcHjulTB2sFtq/vGFBYJrtOkjTKPk+fvz
AGZtYEjT7fozh9hY0IYNT2Kb8tpibXx4+V3qDPOoqzOzeiqvxMWEmNrqBBCK73oL
MSUIsALrPbXnqG7j8IJNzkVBgNHP8ICUTYI3XXyqBHLeFKhBsx3jSUZ8Y5LUDG00
+2FvQ+qTpk4iccKYNJCK6zmXd4Vii80n2P/f/3r9QGsAYZWzN2Nliv+an9olFCzQ
RbIDXbagrh86FqOUICvgmbZxs35nL+U9iDHm6L1xxe9uMTvc+1pod+XF/r2MQe82
E4mCDpjl1BjrieZ7X3Zwbn6D8zJzxjc+uXIFVfwhzzvl9gQ8zNbztDPxS7Bs3Ie7
sdXXK5zRW5fF3uLoQ6d3KKfHWpaiQcTHTJTMcNYjosNE1wIuClJUfdekPDfMJb82
20uZxT+SP89hk5QEPQSQKlOSkH6acP2cMxrfx7Zko02hkH9UTd/uV+l8oHxMiOlx
x3TIJW+a3mpwXjPSF8/BTsVFrLMicng2SfkldH1m31QTYpHTt7lNsnS9Z63GdfqY
/bVDhoBF9/ubc3M9zBih/xjz8ZYNbde1lt11t3pS4FaVNgIL5yJ7WcNM9ZfGpegI
6QLl2rRBjoo1xJL+4CQUySD7s6XNRSsbeV7YVmC7TJ41wIJ8wdh0sUGBk3HImI/N
9wkZWIwbvKkabRpAO+q/8sILhpBchYdcx9GgE0Lnf4WTUC3srgAIkznHfxIecgZj
rEf77SA8rUxtU3dVrQATs8rosc1w5ltZ5pZSZ7Biqx9cQd0l7jMopBIMZJcut0Yp
o5Y6fOgawEXH+2sdaIak6UxO1ykmSadR6vnBQ5ev/N6+4shfEy3O/CrFfVdYUWle
GQBSLhOc/6CLlzIp0dBOiqEKAb7cVGn9zMy593cqFoxJ5Ipr4KrTdBHF2Wi7T7U0
irLpBHo88XcR7vWGw/FUNZQ/qnMH8B/S6Q4bswcc7ZMZuCTAfvRSid0Ase/CcK6C
E7iliGW0lqnmDUUtAlYoVWYaac8e3LqaO2gQGa/x9qz2boz4uYOro3KgPh/nDdWL
IXItr1/ctnkCA4O/Fof2goHHWn9S4rOfTwDk8V4h8ES4wL0hvlfYmDkBbMOoEcWV
rcThriDhE87PDv5yktMZAGVNciVcb2FocaPXkwN0ALF1JlpJlCFsM4cHl5ddyvtB
s5sJaicfWm6Ovv8LdI1O/4NKQ+4sIrET8gXniM9jnPqj8eMYRJ0lr6oIIASS2oaX
KFJY4hkKMhKY1mV9CQIIQ3bch91UuMf1PIHoVTEFjQStIPhURCC7YlD9VmwsWN1W
Hfz4Xa9QCt0D+6tp+NNH2FFPbHYMPH6NiDBIn+Yh5M9W5NvkKAnPAVVhB4tr/s4Q
y1EoHRYmQ5+pHSaUleGCKPqvL2IAq2wKL2whjYb4ljU00I0wQ3YcOMcewhmjld8b
VJp0GPIHWgAReykc7HJLJ2SYW78nyTRrscegkw4FpQ6spuU5f9tpnTQO787kHYz8
koTjnBdTCMGddgBiedjuRUs/CaDPsrYbIm0ywX2g82fDQxKmCg6TlBAS4+49L0XR
m5MGlJaTmjEaTW7/myTMojhtN9VBFapG0rLcEB+E7vn3VSv8bdPo+ZZs/1NoeDHm
6MH+DOJybt7KOQmq2Nhj2nkek06txMQS07mSTPIeJOI5zW+IpznjUEBsTbMgTFFP
2fOuyNP2EvXKgVPwRyYqU5Iqvm9pVv8voG5YJbqLsNeSbEdtMurF/SMsPA/ZJ1xK
T8Rr6r5pymczAKnWzlnDsozSH4irV8ISL93kGxC5r064BvwgQDvvtyonik3NAYZC
jBYgUm6P1n0oflBEyKZyFA+XFG+snCxC6x/gQZorveRbNsht7sOCJnmA9WgzBnrb
+VPnPv4ZbZ5uGYp542KIRX/lIW0VS0txfUM6TE/va2HnV9wbLaNoWjouKn5VCAzb
5jH/2GT5z1af2xW8PatBBd+YVJoFa5EOED7w6VhTZA+PbwjAPYanZAUHCeGSc8i/
m0s2+SM40qFmr4CGRxHNfgO9Fvi17ngoN3q0OfsezqkvtaeHrTuoSzBMNP5XJHyg
vBcx2revR3LbY/YF81a9vqbaMe7NwvpIXUhjf3ipZuugLJ0Q/NVNsxNAOd9oJTKH
q2w7zR5LH9W1nCeMjs6B/kpBvs5cOrY0VDisD6ETdJ0NPQGdNjiVThzGa32Pfcfd
L3dY4EuwbABlrGFukPZtAzcLTuArJOXeG5aHbY5Uk+kPKPQL2PpNIthsImzYfcua
t8xMETmSz4gW/SkbYIoFI8pVDKCNP1H3VDuWcZPPR6vKMiRiWj9AlA3JRAj8Z4lu
k7xyzZwtK7YO9ZFNkXNd73nkcsrG5qI6Ynt7G8dTDofMyo8n4fFknzhbUXukmLmt
lbMOhyQp7JCUlFHLbetNtNtPsU7N5daLey9DaC+Lu/l2HddbTsjjt2RwzLxALNvc
xR1Dlf4eIyhPlIVykZH14tZfRy2CRt4Q3sBe8A8tVjLT/8XODmU7XYojhkvXz+vc
UZvq8AG5dNuHJDwpTfTGoRKEGdmNUgRuje6RmAYKNg8afJoS97xPJBGaS7coNNXd
P21MOcklafLSwKFrG+b+3nC2fx+1zMbLxQHMLw8A5VfgXHGzhzaUI2TGPkRN+zRH
lm5cR69ro9e68MdNu/h1LFv4n0FHdLFdTwlqNIKXvCL1zOrLvUsYCIE5SROszOi4
iuOv5WWKiWt3OUiHTATh6Z4T+IghR8/NQolchm1iLe0kcUoe4qTwrLWgnPDMV+Kc
OD8Q0FUFfpB9Z3Fl72KKF/AdUR1FjgoQW+PVG8pNK/XXDZjpSQ9POPaiq7M4aXw2
pBwbbNbc3rcBwGJw3VpGk4BZpj3LjmSv/W7oS6et3MW7/pcrG4/G+Fdg9MO4OIq9
bTqUf+ZDO27z9aBkR868XFuSe5qRJI8a3O4A89C5+2tlveqYOcfBugyKTgIFkBwV
ANgmbZTBDiBsiUz6+JaTgqH/OJtBYAmiDVTCdOPPNwtT3CDWcDgVte73Bo2/ma76
YLWuppzas0XC3vMtwfhiJMsG4Uoitk+rr0mhYZkG0z3SF3ErREinBOkMsHmrSMb3
lb5bqLLbyXt65xzgGM6xWa+RY5/R8QhPtTsi9JpHqDwbFCB5s0q5tWsvP5QhIuq4
Q6tidqmGpnZepvnn53JLUC/ZEk8Jd49lizXR6pvaVFztZPnQKrMqd9qjleh7XiEe
mm4Bf+5nlgBzqIunjXTZa7tFafZLWt4b9KoGZ1+ayt7wmPqhI67mFmtbXnhmT7VA
tEAIVsl2XB6iBNueyMtPu7ZmYtvc0/wHq6wWReKTIKa53DBFnU/h6LTod+by2Nki
+TOk5Ef6ZRdA7pmqKr9fPhtc2H5GBjTZWEFPXZBmlOL7aa6UJHEWlf49Ae5apoDl
EDMXPyITyROYAGoaGeQsdqavRj4YLDOTC4S1JV4iwn+hjyFzbT8+ovNuorF+7e5q
27I/5MPF2R1yenvFWPHZvSORedlyaP2H8hmRMjc+xKYPM7hwjIFVPgOsMn1t9VlI
ymHydBv7QjQQeF1wJgmA4+HNKBnJ/eaXGIt4TZZCX8iznVAUrgWc8bSWuRc2DW3D
xFEmDiNNw9b3GoMIcPGTvOgNzjR3eKBJArwl0yvYyhB6nref6yTJwzujoxu+WedA
WKYQsDx3ODcaKHrU3A2bDhkc/l9PwVEXRjKfAvQFcMF324pVX0ye2i2sM67++c2y
4n61WRsScHdhk6GBA/QijNpOkNpcjvO9YEW/xjS/hZfLnSmvS0KAp33dsJ7N1RxW
zGnjhDnuUs7WWq6vQ+F9fiufi827x8qxcL9YVBncvKlq37tiy1kfLHAiYepA3ESS
nFxkTs+mESkJNsARtviJIDPlvOhmqH1QwlNzQKr2JRxHjxjgQ2ZSOCo3f+IZg4CQ
kpkThpE2tBWvb2ck5jEG2yfkWeMudo+Wx7n3NRCnqOo3FmYvRtzl8mfeMT7LZhCf
WijSM/2x2UsI0TYABbEtBw69qbaq40ehAjHOVdJpQya2/Z7Xo0md+yRuHCXW9gOu
GU0ouSBI1tHcRuxiEwoNsN020Nd755n1tIfidbR7L71SAWngpX7nGK4cTCQdJl7X
aCUsHmrtJDNa56DlCojGDgXGYozKgWOM7dKPxW4814gLwP09NCOvusaBLaHvybfb
00ER1vURuZ3SHy4eJiTfmkKMO62le/llarVNHQvX6m5Ii2ujWvkIelvFarsTWiSI
QHe8HwNXQPN49VJWyLws4NThWVy8eRIV4pF/XS/XVlArwIJi9ozgVd77RbpKn5V/
pBAUWMjLfCcaR82kWKXQ2/moykiPw89oJGRVf8fNxZxxKFaf65EXieEra8pn1egM
s606JkUq/Ubjkhy5vMk3q0SLB+mqzfFQowyCOwJTJpn9oOyyaf8wdkSJsWzgr0MR
yEoLLxvvWV9zI/daEDcWStXcYUeiWsQZl+Fg5SjWLXQiAjQMLZFqNekGe4Bdmv8K
rjLwIjFmLlJN4iN6V9GI9Jn7etES8TxVtxbtoaPFcrPPVAvdZIY4eaeP1cUtu63H
Ybmiy5j+YArwVpZzLLHwchOyc0oughbokW/8tUyIWu5xvGgbjibuscSH3lYtrlA3
WMI73bniOyfBxH4CFrGZ7bFqcPlOB1x6DOc8QeybsCDZ13Y6I3KfrsZIzzYns1Bg
i+/RC0+WW/Scw+kffvJm/432jqghW2H0Pfg+ZCS2nCkOB7N96mdl3v683CvMVSgp
zh3fqdeemz3Su+pWIcx9MIOJFTW+eKUUXCjA9a6QlQpbbZA1pNxiNAtDuJhm7alW
Ut+uxq/wD5zCi32HJF5MEJJmsPN9Ph/IbuwWNUKG9RBLbjsBOFCmDpGmU0+lDF5X
s+eM5q2t2m/MDi8ObuyknTTLG0pfQ4KUEwxSspyuy75FoH9bU8cTDofFo0Uwmdl8
0vBEkrzP2m26DuzDxAAnzcwRWV7nx8BQl5ju8rdMK/xAi9RMyOAzqQUzGl6yQobD
zqwPQPimmJpQ11qC3n4SrmqGXfJBMoIs0k6/wGXRHo5Agj0j+lls85sRFgX9ZkNB
uiY//SbzvNH436ppvwIkVArrowzNIS8tZXO75kmZFSzsf3QuYEuKkoxtTrDn2ylQ
txr36gM2ylRuG/gGRQgTsb3rjm+t3h07kYDt1hErpCSlTuKfoDDUSa54wmfB1KZB
/xisi8s+ouLZuVi1xLWrJXDUMTfzTuQIsc6iCF+14lzdLFHKsOsPXNPK4AGEE8Y0
KY+GOlz4/G4jHokPno1o930q4qqIEiHyfJyBScmY+6ZsgVxDlfnNggv9bThWnclO
ROzuXwQ7caimt1BJf+ZhIv0NYPVQ8kHuGUSFZondh9RClgef6RR4iFb90vACgJJQ
NzAtCUJP3nHUPvkSKJGcu2OBeO5Qs3ttZbp0PBdWCuE5Tq4GbW+TEk3xicEMX6fN
0GztQ4fKQPCFsraQ6yOaeb2kndcO70x2BS5tmaUVO2eh+TxroCVMMfHr0yrEj2sD
xyySXk+taQ6Z+ffcE5hucu0FmhnfIduxG9Fk3WujlfAKpGC27pejpCKs7+ghGfRz
hA9d/GZxKi8QhxfYcjzaGoYr6vOHlu8R1iI/Wm3jq/i/TtcyqtpCyUjguHgA1Q7g
wclpdxOR2MqfBEJA+9Y0kVpqa6QLFKtBAcd0BeBzY5SgLFlI2W5NKj53wkFbKzFx
zWODTioQCi/CfRWrBoGE3IIPOu98Vi5h9XMXIrrB5SQ/fava8aBOCTMwa5dYoWuG
zjrv8uKNg6mm+TVqAbSXWcyF/TPayIZb38iE0aIe3me1FwSKWRHHywJmIhjpt++4
vdSQ6g87uG7PAaXTo6FvMqyI0eEh/8/07greVbbly+0OWuHa7IpNpnvIFmDoZJy/
0DQWCzJhDOjMVTbejEYZ4BR0lNgSpJX4agYFu/Sp2evP8gpwI/T5rles6CguFM32
rTv44lNbhNg8kW9JNKvZNlGjOHJHMBu3cx0cZEwW6PGYS42K0C5MytsGgeQ9Lkf0
0smA3hv62zz9OOQV6I3f89KIbZhJHoHBP2NbIeoup0JObv6oLcbqsXEhHWyoGsjN
6+Y3bCfIqNh97N0EB1rErBrbCL8l7xSqX815eZTyIt6caSuKNp8YHY1F+8bQ/I0g
TkcVJTz3u5axjrtOxBOU9B57pg+irT7SccaRxhUOA5LwbF1Yy0Owo3p1xrTOGWfJ
Vo3wa7+2B/X3Xf655Ohh+zrtj1qhaxBkEGBGF/o5P/2I6Z7DLBaGYn5Io7FCujAM
SLdKoztm9NVVRQJzj0qJvxfvqa5oBaoW9GlvgXxr68TX4QZ1InUIr9SAtYOO6p8j
bEnCgdVC7r2bz7uF7wL2NR2AFEtmQZf0Zt71NFgXgdi4Pf+XjKayImuTu2sqCmnr
o9v4dcHeGFddiIHRHKsJiBjJTkYCdYqxoK+y/cHkbyYIMNKlRvfH5CSxG+1cHCNO
PAYVv0oOdBkxLUrJWTTv20UX4dd8NbKDQxlFqeUvEosvdjZeIyQFllDiMkiFbTjw
EjgU/v8/MpxLeeobY/2sFIcXS/fDLROaOqwZ+8mGmfL/OhAaiM9smW1mo5TbHMzT
gp2JHncbV4hwWQNbG3SZ6x53B4Jzr4j41QoFi+33pnu1etjmGUPRGpFpxgdVTtYZ
GPS6SV/CtidCJPzU/OPjVBEo5ykuH95vv0wHJ4mtJMyhUcuoHpXqR2viH4sI0aNa
nBdf2I81qIKFB6b6Y12df7r2BqHcHv4zhxfj1qTzIAOTsVVPLj6u1wqRGDpSL9XY
+TZTlGgUSuMABj/cny65PnayFUisuJW0vkNklowUV5QkxpPQ57ShNNvCHPm62qKj
EfoBmnCnrZEuZ6dN+zuRSIU5CLEh63IJqu7xbosTRjMs4m10NfBoqPXuO0tFA7kB
2r0Nh+mCnYsIuyEk2MF+52lStAMB/igds5FgnWg34v8ngCYRE0EYRowH95C6h1kG
tdkhJMXETmgTzMRHO/fxSVQtHi0nIpkv3itcJQEvvkJgXa9kdr8ir5FtBgjdb15h
yE43XBIJDuqOhnun+0ulHct9u0uyOe7hU3X7jxm2QWi9iTLr7BnbLV49sCl0gG9a
6F710yAZvpJVCH6chSKs5ShOXTjb3Jrs7fwXqscIh4dN43Rq7foNJqbB++XHIVaF
wwYsUHxqL7lj2nrqHTnvJN0PzeDYsv7xE7CpwBGj8/XjFfVqbeJjWgoE1ZqWSjQ/
JTKr5nfkiP/d466YvaK//bG8z1yxEbRB1qRwQ3GKIsjVAXP5THP9IHQC838mg12S
MaG6O5Ujlo85Fc14BP/RFM7wGw8ioC0498mrnLu8zcEOtzGsQYN/68rd9FLm6KNG
d6ju/XNhdmW3O5l2kOf7ICV6DrHGptF64/9s9gI8LWnaGU157VqQP81FlBIBc85I
fTwitfUem0p4sXorC59WzEzhCnDTj6iIgTcmF9qLi6wgb/zKEsJcjCXH00QLFgsV
NRS2dsE3yRCLR9p014ZwQcbnnhw22w4E+cyk56DqI+GmRGF9DTTHUvC/t1dn69Py
xV0CMdIy8W90RcE+lUQSgnqkAXb+oBvazG0GQvvh+V2C/zt4AKdIWrfCBUUPazMX
FOfC9KDMx2Rd5yMYMI3PNQ8Or9cxPQ51u2FZfW7su11OaM4YUVbH2J46hULhld6y
MbkBIntCaxFgubacwoZvQ7Vlrt+QxNxEHY+eO/GT53l6N7u4ptd4uoyWxW90Z15V
uUWuP1OEyJaK74kaN0dKlkXPthVfP6wT/0MSvULNly3T7r3R0FRFQjd78+H7JxK/
kyzkMvI3QGyFKl6pz+45BCNXLJuaql08cwj8mtcwrB7ZgbsqVR8OY4WOAPDF5Mwq
wKK9/VDNZg0sZ2HUwo0UxFvW0f6dvF1OGtKz0qmUyFFnbcY5f5tVyFXeR5mDtbIh
5i5gm7P/l6jWafwqxO3BUEnXjf7Xu1a/iSJI35pgOgTyyL4nolAjGqTEQe+EIV7T
FUbjnj2C5O+ZnVw016rvbtmhWlh1eWQb2Ots1vMpXH3F2jbCjN6woG6+MfJLMtrb
PBb/0AS43yI9vr7mXqjdPOkmvjRDVZ8E2Me6BJz0Xh3k7lY6U+uUt9Cds6YbMANE
3Qay5OT0kCc5F8yNHTT6QNeB6/xjCT7Kz/LpxK4B2udfr+qsx94I5iLlybXvszlO
fCqAIfFAg2A2BOpc9M8HulDphbrFz0CojIM2BekTlQ9lnUKEsrlYVeo9pcYFzXgd
rYWvsvudLiZXPIhc/7vdzKey1C47gc0/WDG5CyFNrkUK30GStfRIvlZGwz0ouByS
Xhfr5QSbejyYbWASFZm5k8YRO97ySy6ZSUFCBL+OjXzUAOvFyC8CQ+hD89wMuPjx
O1H9P0rgXkgniFROd56RdLQu6zibZJTpthQG5PRHnE3XZP4Hp6v5UsYP2r4foN2R
hmXBXLEbSUGd3J/VLzcQCwjZ8KYw6agCS3rJILgGl658JZY5757ThjwuCb/iBtdj
qeaF97lg0qZ1V9Bq3wjhCF21ZMA/+/pXYYkE99rThakU8LCyesujqmV8ceY4RPji
ySLzI53cDhFFYu/ZcYq6jDW8MKaxR24txztDZF8miOrNDHGOA7OMghIPQHfHNzrE
DXheN9aUasgMPUPTxSZoK9tyM+f6Kvg64YOPz51vDZbPLmt5OFHfZFu8wXEpEQ9E
QIfeDNCMRuIAx7mwvObCnQijZrfpXVqdQOcUUrHzfO9jwaaXZAuYUFb4FJrqJX+A
H1AXUtHzM/81HvERPqHhinsS3MTavb978/LeOyeZRHrWNlQjMqwjbYFKY7yyW9+I
TpwtjF5YrRP5ClBoHfBqJpAq/lsVk1nQDUJW+de9V6yJ4vNn71+hexHsKE/q84Fu
50LtYKmqYhL5xfR8Iv5FsunJ3x7liN6i+VMZJc97XUkQ7VHctY7r17eKNs7bSo98
Noc4T2OBEdYgoz1dbU1Akb0ZRw85xJMhXdT0G40xgEr5IHown7gcm0uXTJdp2jLR
Fv/N/a70zs4MXrQQLip7DWjTOej3JGFxBl7UcS2U09xojL3hUVkzwFSJTJYEiVRO
pX2BU4Y4lVpp87jBMLiejxAtxokGOwcL8Qy9k8juZ8RGLv+ieFChP2576+taWikR
IyWhLQR4zIsexJfqiy79Hwjcm2fc5DAoSh7ngYO79dG/2maTAi+ku36O6vtTKjUg
fF+yVYsYrHZVwzwLHfUgVUJtqKEP91XbKnfY2veC+z7oGHaCpsTobFABlJqfCVV9
lWSKUdoeXAgxa0RxSEWcJruQaMbM9LESdfS6ppa3N5m7JWyin8byWAAGmI2eUBUX
/FQMLdFAF7JDjCdyc5gmSW1VHxRlzWdMddoycS6cUdAiPK0vjNDkAEmdryUnp1Sw
pCtryz6HYiG1IW1GbleQslvl0l9v8RhBWvchgrfGvTrBLO0T6gEjVeJfk7J26OWy
sgwVALybqVSdw6pwxlleWCGLquZxATslZ4ciNvpIKlgT2Orek5hdcDPC+bQOCRdu
Bxi/ew1ePAyU8gxSj7EwhXhp0vgoEL5wq868+ocT5J5LQjb6+KLUEMCUP0l6R23C
ZMxhTJAYlnOge5uoIK56DtNzJakypFkp8Ftl5ekzUfa49uGygkxUgRwoGrA7Mu0z
6cNaRLtlaBXDgsLix3Jy8e3R0gjnKPVAugnKPvBahBf08VOaAQ7ULOI+zKKIWSU5
+wLbBAXNLLj0qoz3S+BhUvTP60InKNuWsx75+RyIXOWVV0exL1Jrgjgb3w7HqL00
JlWEJ83dJo2AnuDt7e72KG1RHGGUjDQF6/BVzCJSTFHB7krgWZqaJsZuXE97+/wf
bRtkw2yJdu7MVjIWnloFJ1el8YSvhRv7miHk0uCG7omfekJRJIdzwBEg+8xeY79j
DpCDlVdGEXXuTA354aeRfoatzU6s4hDxHXGmqdXNT6rpyhqj7iTTWI5y+cwFqZxp
fbhctvJr1dk4fLxmFk7CKHdzGYm8r6tdE1H8ziCO3FF7d/InMZOQDEllhHWtkBXT
PGrq5Y599XyLSjGtmwcABKczL4xhmwskm02wz7AHG5dSNLorMx81Fi1xhHpRRtp2
fXL0I9e+8vIEV00qEeaHYWJ/dS0lwJRoTFPby+e5csenfPHF6OW6xZwoGWjtpk/a
5ImLFK4ceYlXpdqX/A3Yr6UBQ9/tHQ7JGA8GwRSPdCrWNqFdih8gy6a/uY3a2C3o
Up6TA0BsOJxPLZ0ifSBfhAiv4ERSjr5cyySHbYv68EoDMIESEzCp3ZAw5xJ0OWbk
4TcvXu6B6q6K6otpqGRCvwUQm1vscHcscE/v13caDETGzPLkvvWoAp9UqpxnctHp
BQSU251iwOU/MlP8AHTR0l9pJp601PCW+qSe+C64suf07muhJVxBpE3M5bRcj8He
Ng/jPqVW81nleKFdQCsnaM3VV3rr8HnzpEAx/Je+hrIxTZeDhtjhR+Q4fmO1OZp+
DZw30iq6RPxBWqg12MJklyjdlCtZNAqevaUZKEDIUE7Y5p9tOnGeQqpl5lfqBTVQ
29mdzXHLOzsknMYwZBtKd95ocenRxOiwWlIfq+bPU/T6U3xFf9cqnkR/n3ISCNM6
QwpX1LcpWbchmPMZQ+kLvEWvjulF80l+LlA10P1nSsSqgAfviDb86cNx12fVUx/E
av7QVS4c6eBT3Y7evp6kR7eHsRlXBMxKczqNZlzdZjKVFeKDhCOvQ3l3uTllIHlY
+aSPucZyI9ZiCtm95ej4wMoQ+21IzlhNO9xmwYs8qn9Co+qbnOTJf6X1E0o3Cryv
IKMhms+62b+ypVT+hoyxdqe7xHzgUnPNzg+YmVLyRxUMGPqLsIgVGGvjljDlX2SX
8BjvuIwTYTLvcSfyGTey1cKOqZzUaG1r2BqM+0vRWgfCwohuARc+1E7uRPvpWCnI
GVsO2Zv5k/0Qt/0MjKXgLILgVJLwYzPo3/3PatfNeUkWdmN20O98/JIw9meoa/JJ
lOg8IP9anRInVBYrK7pOoSp4eArR3gWK/Ui9fIxp5sFi0R3rKo/Ow+tdCPdl9QaC
IpZ1aAYvMfRQaexXIEu4KTEkcaJuJa5d0Tqh2Eykz0fMT4wV/xe/JND/wMr2NBKm
yikMGz9zBq52n/OAPFDj44VYoYRkhJUrlqcI9Rk7Qq6ku1V9+SRiY6FeTGso85PA
MQGbqiDTDKAZPND4FgqAEQ5LJKF5hJ6VgrGo2sgH/i2pFYEKiYplm7qezobokHzA
IJ5BbYq+unpHWnKPDzN1cGpk9tfDlZJJEr070PFEma/bJrJzS0VKLZ90q346W1s9
FC4cm3M3S+J/f1yFSOZos4aKccE78T56HwrCO/o0Uik37pq5gcImv6pJNNW9KDaT
2vu0aYlunbvh175EFLoYGNP+9haIaBqQqZpYf0GGE0RA4gfNWs4Cy6jRTQEbK9Bt
HrfxbsaHEtoFofZJrBctNqMN1hQ1uJLaddgH/cq9HMODCPblHghbh31yfBi0WVMV
USvxU7/kON/Xsdo6Xvv+tBusTLMfv+zcrdcnpxF853bhzT14PTyZ5v3HQEoCQ/FF
FMWsoD0XiRRpL1KxRH8ACwvOa5nN6UPOeU1OMDrUe/n/X8fnisJUOetr/Nge833Q
TUYbC55G5ZvIclSN5TZwz9XEjpxggLipBlAha/RKPgT7EHoebMWP3eGUNg5d1Cz/
V0MYZoqbpo7SHwpgNGz9HYkuqy7B3zUmQissIpNn8zR0JiIXColYeIxwv7MSiCgr
jo6tkQWLnV8CL8f7QadkC3iVkyRWbGCPXeJwUewMC34tdZhM5FzkIZS7iUxND0Fk
BEeSIOouIBrFLqk3RDGGqfZcHOQPcvWsxWozn3pvqLT21fAYNH99rmxdeM+4MT2f
8TOI+BYR7axA/rT83INcF/h5NsINXxlH2dE4Ax7A5HSYKCkx37CIun6BZKSAbMgz
95ngKE++mD02CW/HbGRCtd0mCvFn0/va0ImQIR3qoYYkAaRdTjMXoeQh69AljjzZ
OhrtKHW75JRy/FbKjGSNaOqLSRVpKqhMEe+Mcda8/zwIp/X9RrEThe935vj5Tphk
m3q1n0EKcKid1SLBMs83CW/8+rDDgS8552GSwvx8lUVn/d4pdjC0XyDF4lg3gJR+
Sn/0kiBv11LG+uIbQSqfyLQ21Qw4euUdC8ED1DYGw8/S/xwjQbMFMQ/uA7Q9KScQ
ZXuvAtYcXrnz+e5uROaECMqMbJo2Qn6CAP6/yE/jCCLYe+e5Efuj13q0r12ebbE2
UwXHeEBQsPKHSE0sLu22O8bmfX6QbYIt4GRxSzPYUaWEM1HFBDsTfqyX6Ur8KL8t
EpEQX4WYtWtGTHlNRUT+8IZ5uMJHFbde9N7nhndi/IoCnNvPlntXaMhwgVCa4KF2
FBbDmVlCBKoCuyl8skonYBktUBCwttVCLtWZO4arihCbpmeR7iSMIPHaCyfjtFqj
/2OvWu/5c/00qlHeMie9T2VIAa0xU6DrqE/gxldOc7ymIcRD+B5Q50xfWpPXwZah
5srWZZ71+RjFHqzfznzzq4FLlraEGaoKfB2oskN9tt6Eyfz174UrOuLoQ9wYJu+8
hD5clpL9Poc2HJMarmamepGzQXFQsfPSoWVHzin4KkxH+fJXQLbDT7XguCiRDB4O
5MDziOoO/S9E2RB4Me3UtXiU7II/ApEmMjqfjEtqf5Lzeiex/0y+FjNhFqv4NI/w
n8dVDPFlMdJPyZh2NAtt94JccUHRzbq9rBGs8E5vJwVft0EMhqMemd6kV3nPRH9I
gdoWFsbuTWz65GYEkhe9kSNMI71UVEFWmBlgxe8+LDdMh4xzH/AlcTgv/jKc43k/
uGZ+WfT2s80gq8d0ucQ+QvLleobDms3RmpSPoJm1R0l4dSmBVGj3D21h3QxP0iq3
NCe3ZGqzO3FD2j6X/s38Bk+Ex+wuHhCMC/OziYNaLae9imVmk669GJUdL000Ufrz
zKLSjQX8bGP0XURuBVbSKicppji5Mr7C72IfwDdsQXEwOPCWOtJ9C7uQojsK3xpW
CJ2bVJoQLbLDK2Dc8ufKG5i+L2ZNhNBARjz0W8939lvfg/K8F8VGdihI08fcC22R
s3gNUtV3KxISVpvxx8T8wzkY3GyBpjMOps2QRb41thzoNjmURkzL14pnDzZo8nJk
vVUUpH/EOMMHtL02S+RYtE7t7Ij3UzEqegpsDlRYP9esA6EPX7xQvnseeTlcw1t2
szaKY8UiBr1TUlGJwLlxoZ4vzSkyTYMA8wtu0+NfPNa5xfCYUuRUuocYpqPzK0K8
iZPiLIGA1XTjYGlOj6YjNiLp2kIHoW+OZv2makQ5Qn6O6OPCUWSdTwnVOm+UIf5t
4P+xFMFBlNwFTJRIgDsPxgWU9PgBzcmPrK2xy01ncmMsSh5V3oqKLm4ipzVoAyd0
75C0hUW9bLiQ8VV8QDBG7Xqadb+Au4PbzOHH3lQTzSlPw3cwadh+3q6Cg84HvQGg
wi4C0TkbbG62RbPc1F/Rx0Vo32wJtV7RZf8BwoZcZpwzXvDYIB7Bopt51HRyklsf
CsqnAMMviKVMaqE1MpYwOBvvzjCu3HW5FurrtXYtQQ+xRQeAw9pvht5x75ecWjRC
NpgxU5ICzAWiCiVzQIsVKny8BFkWHwWDrADmHWFtB+MSbbS/yY0+CzGsUpF7Te9w
lI/yH74p1tXRqpSamb/SzD/RfdJYlv87oS6Ikv4JLFot3ZhPKKu5ackxDKH65nry
JRXTZllTsFC47Zx2SL6L7Wx9fxv2jNhI4Zn86mTafas4ogmh2+LCRTzpNyf5lGTZ
epev90FMVwFSa+1O/4Vz+HunTGdc22MaeoaMQU4eI8V+lG63fOWFSObryeaYL2ws
Rfiy86LUuRioDT7sx3M0bRB6Cn/vOfpJ3UZLQtGnbAeiss7+3E3oNnxdmfwVmncV
bnY9Bq5Ul7wbrKLQ4WxZICvQI+7CrtwP1VaGRn8B0GdxnBiPtWFgkUpifBM4z4qJ
5DK2jnjYWVN++JGHyp5BYhQlFrEut1a/EizQiYmjHAffnGGV/c/UU0ES45JJnRXu
7MIQiT3qLZ/A6/odK5c4x6NBRfTB0H4Eu8tfEGtYcgIPFyhzahqTm+Pj1O51JYSJ
AVgo6g3p04NjbKxXKacFH5uFQIWC2RHf2ZpcRQcSEPWd92pitlDZxdpArDJDXzgT
aUzvnQLLqZxVzHeJe8yA0Ye098qqEAPVR2rKCkOOPa1AWU6D3lWDdyxY+SEI1689
YSHmLQ640xAGtmqjL8oCFPkQkV2pVJpzMUb7I34OiTohEwilP2l471C5WOJ2Ev2N
nE9TQwIYUUjZ2SNczZEbFfqM6rYXg85djfbFzdq22HVxnuqgO1rmf1iD/X3Q8Bi0
EamrbfTX3T91I5SM0DWWGlz4RChIzd2HytapZH9T8F9DVf9v+dWxBsAPGrBNEh9N
iIKHC8TqsAXJktWKaB7e82/vRKlh24002MFVKA4AxxDxH5urW0k4afu2eAgu5jDO
lP6NJfVLfX3kG0GroSyX5sW+QTid4HwRRFE0hJw21g40htG7uKFIhMXAC21pILfm
tuWynSf0d3qj3eOXRcDreklFFG5cxkrf3+lUvhl+0hiPdUqDWoGtFppngeBB1BP6
4cdOIcWax37U1V9rq9MbSTRt5N9kFK6tQg1a6AvrgzGh+Q26a8VSWpECxx6fFXzC
SMP43KPnojkBAAn+Ot8LkNhuQLJ1vKfrWQsWS6N1mS1Pnys5gp8MNuLAX5LB0MYw
4LFZNBKRY23QQ8jjWZnulfuEvOMIK3hZPmmzvwQiIg5ao+e6BNjJ+B/73gdyndIO
fgfwsWWeZWbx4+xvmVPcpldEerg0WLmd3ogKiYdtc1Pt0jZdCrAf1yvBfYEWmVNL
S69bE66vBI/WqzFjA4b14cuYfhmdLdntE3RTf+KlyRPgeAZ8V4JLUczo/ziYiW9Q
rbV3IouZR5UA8WEe+SMGOX7FSef6jYpugmpIVds53fltVlu0nXpycoarLgMQMel7
7xkg82MdneSPxZR4AIn/5SY9xVZqdUJWEt2x8/XNeWA1dCtRpSPnMPGUa0v9WU28
Bzg+6f26eT813VsMvttMrywM8bPWw/TBP5g6N6YU2AeHSYA26L95EJscyX4gzFYD
XkbcKHv9gfuVkMW/iwmCuzeNaNh1y4+W41Fy6Mj0+JyvchEY6GgqVukCLl0dTJWy
98VVI7P+2tQRmJKokftHeXvpz72X9IKEvg+qU4NFIco8CpreCTuhhc9L7HVMgPVa
ehR22ooWdDkvpz4A1wmlWkfo+YBgeoHTmbPXw8M0XnzOJ1mcMdYjej3CfswZflsA
YP53tGaTWQbDcASw/17oGHcngUeKDACu+MifwQcrFRQsr1h7Qo1mXzNPKz7L2c/8
UmOeA+jYjaUqNnesQc5BzimoqJAKdDjv665T6HANKnelJ5yL0ojR+D99vrv/5CmO
X9SX2YYMuXRDoWPVlbreWTHXApKQfTM6D2gBNQPhxdKD05huJEcDzEvXyRrNjLre
wU7p75CDyhCPfYglVOLJHXMN5pEn9HB8xXbXNh/0CwdN+y+FSjY7p+M1Okcy087p
5FV+YN/1EF1xHVj6eAnLgJLw5H/z3lODl+WGx8DGELRj3J2QXbCashpAm+exEkOe
0eirTCd/qTR6SaqFNakIamm64IWLF3pNbWk61zBiuD6+PG/fKbWv6D80Y+v4Ahq4
0SkE64OwzW277XFvqwMzAV/qV9tv0wpmThh7SpHqSBGWyhMZejTFmTZjN0wgQIdr
v1L1qjipiyg9UGgYwcNKVDxjrsOPOAryQ7YxzHv9RFe+DjrPmE8OW6CaDf3dBqSR
o9I7ueHuaQOO0F1gR0IX6WUHbHhZBRlelzTTmq55udRCFhXGkj0s+PhrTZza5s9u
R7tfBD8bsVUCojMyv7CgaKjKxde7WC80VQnpO1IgeGaB+ORIfYYofw25eZlGmP0b
r70ggRdG1jk3aLKHV90yd+SfEbRJLz7f1zLagbrr9OHN8W0TCwa9pfosAi/Qrfm7
wN+PMKgNuTtblQJS7KL1NJWu3s15db8PbW2m+76LkvAZvIorLYdDjgaKSxBbAiiY
JeTlpjWurxerulVzJp1BSya1UoRABygI1K9QNFfWVE4fxqLVXVczi3FidsggZqJE
BU6Nanv2mY0o7XtC+hrfLhwg8M+ypvBreQtg7WlNF+x+F8fmn6alWWJGaCpCiPJF
4x8oEmra0wmvnNtprqw8kCbhVr6pWrU9TyLpqCYlFhlqfSS4B3X5L+KRkDheSJwv
PVoT7d3/0CW88nE8DFHiXGMx8VR/fqHcBJrxLIiMrl2s77i3QuaoGyhS/eMQNjyt
FVd5YFfn6RcFR6aAEGzkrOEoxwTnLeVnzSvYEGJFIpkksi7b03IkISRn+zJjgyyB
L2HAbWyMgqV0BGlSGqImcM9l553QodKIrkbYUOpwBlgSACLlGscJtlUCNqmGsqBV
8f6grmhBwaDSD8RU8VWO104I/+Zuc35TZLsQjuru9jvLPksU+a3Zaibyk9myMb32
ni/zSY62K42mwgGnV6SyWzEXU9n5sYdrlC8oGEk+UMjQQoNewhA90MxzlrnrWCjL
QpuBWx8pU380l8QJNZh3JmLoRFwrmoT5Nwm5qdmWSF1w8OgLM8Kid0kanPw3DsL9
otyRjYcSWfiNgKsTHU06DuKl2kdPNf8yzTivNKBUaorTgxFy+ouJYsAHPPTEjwFF
ZqaToo/Vr5LNeWD+6yZPMc0IzYqfdQ6fRR53z6o427wQjwckBbGK56dx/u3vMHpx
WJNQVLGcouNcbsKMHGgLnWGk6giOvMgB+lg8gHTvfNpcPVTwY8jD5S1QkRtTFBj4
bxH9b6MueH2RklIM6LgAM9lN9MQ64SF6A9BeUKha/XfbN9VSTTIwLk3ZrHAvUJbY
OsnzXw8PTydHccLjEqEY6xdjD4l8jxBD7MKa1+G14K/X+kkccOfqim7TYffFcOwe
qTF0yu0w7aQyKNN3ivKnYJo/3zLho52Wvl7V5xIek8br+WdhtlnR9U/X9bxYvebT
t7f4RRs0xZiDelsw27OPsJfengUXNA+sFDY1VwL9h6YNHjB0dAhLpfBl31rVlpYL
ylcVO/e2/d3Lt0sxoRP5BsUJ3SVJHRCu6KQ5vFEJWl9mSJ31UYRLpcH075/0jxci
dDzLkDZUClK6jgFrPjkK1iikA4CtdP3m40045tykG0Pmdd/ZJCD+d9V3BM7mGv9z
BBDEriPIJevcWLYhz7Hxq/w0/lN95WlTK0xR8h93UW5drBjIwJ6ia2RsKwK2ZIde
NtQaFcy+r5gjHzbsPqYDy17635W+1uCpxyeqmF4oTBHgwVP6Mi5u/GKdgul9Y45L
PrRCBIK9IRDx8r1irNPqb80P1/7flqJN64tXoUSzBrznmYVkumzvm8cqmBXrOtss
c2vHjy+wmGhbYEF0lEv+3JKPHSKZ3XXFgqAKkiXqyNTpN7LNZK3I20uhwM+XghXm
u5hcmLbL6jrG+tBH9XzRUcj6Fa18jJo3XKVTgkOuwcBtApH20Chq6f7jtuAUw99/
0Gd7icl0Q/fdhuGb6B/cg4ywaO87FWvObgkZGN2EVhkb5bpY+U1C9PoU7oohrqvG
FruqFALLOB2bjw/LHtLNrmXpjQ1tVj3EnyXgkUD2rdSFpdvVrqFPNv0VHzet3YxP
MctBjSGAhAg8dirv4meHYqMCtx+AzBy2ws51TAmnIwvdS6AhfCfzRgpjmp4XfU7z
rg2db8P8Rx6Su9cuzuOEvShkbj7DS0txHKAgIBsMPgYfRkfdD2Y7L72nAZ91ZaJZ
P4hfuauRYtUmXzmbhB4B+eu/8+e3dEgyYweAnzBIZ8lI0kboxtPhv4EM1DPejKqE
cVdI5H64DPzDYVt0W/WqX3L0u7MTOIqNxc6RfNk0oFfTJCbyA/S0wKmPpn3VffI7
oIn0BTWoVIn5YbSlfQ2UPXt9ZjInHsjtnPYu0rk3uG3JVFqLUb99KRzP7uQKqsyl
osJvn9oy6+yMbTbFcn9Yaer4Q7AedaFO0x/0QbRsXvGiAS+v+i45BXR6RTXmQRcy
rHANw1MWTfXcCge7+juqKJGt24vr56E516Tg3olz6L70DJ/2XOJewy4BLySveJiD
oDV8qcqmoLUYCiEUurIle0+xzgHWLoeMgCMLF7RchLrWcEugaAE8mxI25Yetd0u5
Vld8fn6SXcu5Ca2bIBjcnrsVSj2wZtFWkyE/M9sQRkSLulMW8VCFsL7nv2NHMRrs
rIsMpGKI8g8M99I245u20rhiJq9s6LpJ67TA1Kk3SRAC3OiX9nGNSxfydkplkBjj
bn/678NdX/JoEr7yrjBPEGo95WY/NXIry3/hQf8PXA8vpxqDgjzMUFRV7n2YKQ0T
8FsQFGMWZInjeMXuJ+l3ULTFBpBMf3/3tc7yhPh1uZ1POPtbWmKMX+9PLxKTzzom
IQLNNq4oN3Jfzcw218QFPyxpDnhF9yu7+AyLED32Trz2RbM3XxjQBtfm+e4PdLfq
dW9GGmSYrAFdHnsfhrAhhRWPsbRjdAqrT6YZwXghUvckDZfn5lSbP01UvEYp9KCk
5JZrSgnwvNkuvykXM8HdMg34iKqmpQePUzxIVtsuQVQZfTrURikWIIqF6jHkXkdX
i0M1DG92gZnWspovt8+La+TSH5ZQXO8SrQXmfbUif+GSFVkvM6vLT2PB4xwE3i+C
Zx34aoKPPx3OoVNvqA10AvCZOVWT+Bvkyf7fikNpqdSx9g6swatM0lrIM6qVtomF
1sW1Hy2tAaQ4BCOXiQTiUnih7/1hqqSl3talVIB5RFkX4lk0R/HZv6zkC2ZQ6d+Y
ZCOx8nKyS669C8HTS0pAnA8NymEE7ITWl9ZP8/Gzn5rook7wARivLM+5IZCdpj8m
LgbzQNni5H6y40L2qCS/9bCWSqOvWJN5P/Bpeqpz/gahI6RvqX81UG6Bh0VWmlwL
0d9+DiZ7NXy3W9slDy9wkGVmo9OSUL5pMRBGRCfVf/eCkahR8znERJZo7GeIBVA8
FPNaPnuhvho7MF+5JOKyAYe8kN7wUiCuFREcF8NqXerR30fmH45W84b9KOjLgWym
MVQwzvLR5fKsDI7y/Zp8ytuaJ6TkqAnRZL1uTXO/Jn6tbtJxZ6DEf8Sd57OCJHRy
izJ8C4uxu6EFzdoHkAxSLS942yIEM3ExDLufziyMz3NVTUQnQYhxQmNfk2VgSISd
e0zz3pYeBX9gcSGn7kKAakm7zPmyE//pLUMM6dJDw6EtcHBNUG9QKpFHVaImj+u1
DhIEc89wPjPBB55QSKD/BrH9p1qzmPySdVG0D2IOxg5Ikv1LEKK1t1x/9koriXi/
JEs6FLEnWNHUia4Tt8EHXtl6pdhbtYVhnZkik0NpBjDGjDF7npwFLx51YkmLJxAQ
fdidh64VmdOTAlU183o0cD0U+dCr2YLXJJJPinLEDvyT99E6pOEIOJpejnqvN9cV
7IXmVwy0NZOSdDHrODU7BaWj2rC6zyuJ08WHoMispJKN5tSLm4QCOFvFwb/u+F59
d23a+nAllxBy2wN9+tYXGqW6XO61/9gS9gvHiBP/SwEd117UOfXsrEU+nXjRaueK
tGzpCufbx8IH3IzT6QGuDI5mAJHtNHN9CnKFyIFE8QvPeL7YytBXo/C7IAAlhybJ
AURDGdRJH+tVCRzOT37NtAA3WsMmOpx3WPduGtv8ZRq4KEWOUUYDMF1BS9GxdU/A
KhgfHvC8nruETb7JnMO8rIHOmlW1Onra3lnSXgFpV5uKRobQkYP7QVaVGSuKAdLH
TDE6mu2x+m9jXVM8KDfytqcB4QOkEwNnU4eeaVIEKmJIA9UvUNtfXM/J0UDWh1PU
YshD8kT/5/CkqhVTS+0ZwgwOMKpReR6b4iaIusSefKuxT0bQ/cg2TQp14+5B9v6u
lJoGwlLF7ZurpMiYs+eTyBQFZU2fPisV9XR8xcF9J2OsYlOi2O6S6rS+aXdDa1vO
AX0mRli5e5BUK4gAQl7PxPcPEfPFzB/tguRA4fhhJemdTVM5gkQxXsU84s+HmbN7
fkCjH5dGr1AfvFA4lVQ6MNxyRYYUzHPLaBbL5ajYcDhKJW6hyT1whABZMfMSvPE6
3gjU8hE59YYoTSXUWRyeHmTS5hHQhBDgcUMrpWQQSZn9vhjkiH6+f8eLBtGJ6qzG
59pd59EdVpKxtpLA2RS1kzERXI7/+7YunySxx+c6f79gvIr9yxarHRcpRuAMv6nU
mNVOkDhHzn2cHmcviaXAsM4DpCqXCtzhPrYGFvGRlIU5tRjlHcjBB/ApgJwJ5DgB
2yv0BYPdbvaBISaPhy7KSRNpPwJKay0mF+jbl/n5Qf6ivNBj3+cUzMP1uEnDJuUz
JH1dC+8PbXF6/DZOpf1UvOGqGe/zoP4u9+et6rQza4ToVa87DBXNpPtpXqiXizbG
2Z/eYqI8IggVkOdkMOmWsGULrUR4ZYjNqWZvwW+1pjv9qrQmknbMfjQoG7XlQmR4
QACD2MRlEmjoURAqf4eGU6t/FwG5aiLa/WxbN2YRa8ShZUN3KUVdBKLu5HKvkLR2
nZXRVJ30UUkYHFzI/VgdrL3phJSHTrWGfEeAbZaoRukWRsr75OIuRSfg+BbGvwGZ
BG4HXAS/aG5ImINGnkNIGsaIi+YCzVg/Ibu7C3HK3MuBu/R3TEU+gTWDEWjxX/vy
663F3R2kkSWFGzwaX6qgmXlRCVRIrguEMozV/ACsTLOX2Zv0koeZ+B+KV5dfsq6V
BPlsG/3FqKtYX9bTsDAf44SoRxxKnRvpg6bSv66WWMeiCcgLnuItU40y+AJJPaIl
vMuuZMF3HYsm6I4mCKeoGZHPc5iY8eLDK/vHr+PMQOELKGxVbsAX+hDSVYGZRQZ6
myo0eGMCyXO9Czb/PXK+ZiLclBybgvoHInEJPK9t3KeuDWwR3G09uQ4rhWJ2gBeu
HWKkyWysQkn+TEGe7CLizIJ7rbHhTOuRsLW0dq2LIz1Wm8AcCO8ddHJwXBCR5Wog
SC9z9uylwldxZF5vOsmthixpMx/xeCq/w/2HDoUumH0CU78XsocZIkq+acTKvC/h
XhT3NyNxPgrhz6pKBRJ8YGacZdUDC+AxW6UYe9Mv7bbAV0jLIIKSOH6EJWCRXYwj
i/C6Dqa74SXFQ7DPRwpeOtPwn7h07/V7nd746IDMi2oFFM86AX4iGnrvGzxl05iV
5QF681Y3+GRbBjK002wnZ0lEuNKZso54TAl9HvWUWkGZoFNmncN4CM8n2Zx3zlWB
GzMxL61Muqcw8U8CMJQaxa5Yicle2oDEL1MSVogyniP5yKfS+dLyZ6s6qNe0RvoI
dv/9Yx5d+7deL3B6ycRbWFIAEcOmkYR4GPCPuz3+wpbj1/AKD3u1160tMMWeM6G6
UgsbBnBN6KJcPNjbGeUQSGz0IDuBrUdAHD84ma0JPKvpiIJpTS0CI6h2JB9oAeJQ
QZY8hxb4hfTPJmJ6gVKovC/8iiMRtqfqf5SZgpMtBHDbivKQ5jxYfR2gc8HxMclP
e7GVZxHvex/L3LPhI6yqSxwQVdjlxMxxVlVg2Qz0NPBa2wJKO+eFKnjacqdVedHT
emY9LjboKe870Rl2BTsluRQXik/eMhOf3DK/t/D8oVHVRmn5gcYxWHLGkHDEvfbH
JeheBpvRZWcKDfAddccaK0J/f+uccXPw6/jcQGCEjG8m6ZF5TsDz1bsxtoOpupz3
N0T1EjRGoTd5Qaayhe3e6rty+2sCxfYXHR42yH9rAxXIQZX7LYaPV2Hqf/JeNkUd
uctCMhz94zz4iZ67sfsXe0rvcj/LXnBGQN38usrwEfmNpTluCkykjsuTPL0MwQJM
vrTeZsFATznlpA8dYOfiafJtvuX7D9OtzR8MqAXtcrGj6dzSalHGLSeYB6fIuC7k
21T8UCc93b0hX2U1x7Ps5BY6fgGNRSOVEudOINtDiI3yZw3VAcMNeyrb0NWaWOSc
4F6MxfN+RwgQVyGGMy27MRFXmp9WpyyBJbIfPqKNPaw2BdghU/bOzisdHCMVKyr1
zv+dk44eBELBap7TKboJOwXwPgGVBnFKLFtf8yjEcx1300PzZ+7p/P4EVvMMwtza
FU54VIv9wK8PPvYXaoPdAHhJteMAudDkX3gXVQqfhob9zkFBQ10gP5C+/aPN2Qzy
R9UiSJAaAGiOoj5QMQtZsQDtRCIcdK2gSvhMwkR8C3JIUtvBw16oVe9ud1bPquQH
366JVmv6ob+bDjRSxj8XWpVvpKXcUG4Z4u/4UGlffszilgFY6GRbGr7AgUAxWqEc
VutEV4jubb6yTMwWrYBLarVnMbs+0RJX3EeDjTe+tXBGVmjmkhdBxCeEdWpQb0Jg
R9/hX6hqGXC2+aXQ23oRfK1/qGAMvmSWKbSjSEeNfoLlJFP0h9+tT+MzPMLAnopA
Ba1BIBOaekosNYKicZ7407sl2hL2lmCjVMze9AVthlAfWjZWSVEdH8vIQMMlLnsm
7Oj0LN07+aeywy9hwFEeLY19mpsA5BFPRRaRQ55XIu9M6JmI/hsz7kZFDe5E64JP
IHXTGU6il+c221llzZ5VH+vLZ5MArh3RSXBn2OKARA9K2QiWywTUTwT+P7J7oEvc
yzit8CjebQoDC/mCqY6Y1i3fu+2r7lQ1aHlsmlwZObBxU+NFV7PtsxHiBwcavDJ8
EbP2E7rs8Rhco4soCiWkEdQfmjL2JDWvaaRdlkmU5Rk9ls/9Z7umvZBzqSe1EdRK
m329LyFDjgZycj3MWHykFRWRteyheUyeG7iZKA9Xojxfr4TXIJ3/AdwuIfqtGU8M
ufemJdmD5dfRnBcRtY501mo6qAXRybmArHP2Cq+6eYZKJIa+3gf9TmWp4w1mr3k6
qqGwwCh9yr7DoO5HoNslYjstFNByu/NUK535iDuc8MD+AD1UvdhppwfgkQB//UI1
XJq8RtxeNpNmif9gbHZhzKOYCQxDfK96DNiyfBGSoBSDFM360DvLYmtZN/NYyvep
ar08ebPJGU4lRHphJyUZSbj/UxlNcy/q1SraQvuhlmyVITeVdm42iqiSTpLTr9o7
HIENzOm5SYBfYOnBZ87EP5nBnZbqJQXQrYW0iv1XsR1gWmYEmRsphmAytyS5Adop
JSrMft5AApYrUCJyvvRKmuju1TUbmPQV2nDRqwjkl1UpSxkNEWp7+pbKaRMo00ap
BzpM4KC58Vejb20PCn32ker1J+n8o+jRvIOgjDH9/6HeJNuKJHTCH3meDbdZl3gm
lklx2eaG5S93P2dKryGjFHrZAbnCpHZdMEP6CbqEnIu9TBDMmXQKN3NIAosq7wdf
4ZntTeBQAQzAI84Aa82Ra06ShanQqRcUrr+4seiEqCRB+kGzGrJSJxSa9uwP3gk3
kDcY8qRfbeZFls8BiYRjBqGGgD0CujJyA2Dnc+ljJuEvaPdHH4pM5YUSzZ9VyKCk
KmS2Tkymdk959hYfDdBfHOWK74YuQPSphBHglcBNTiUoLbI8+jwmoavZGe4phAXZ
g1ID8l5DOsrktwjsCYDuOzeG1otztX7PUa3Bg0UI6ebj3rP16vC6MS2S+HyIo4zB
miBE1qZ0b0kxKiD/ypGn6Pz7pFdsCh6WEQc2ICKxs8RjL1DJmlwJxIng5OFil1Dl
WWSZLJG2e250aAgdBMX4DguSIPBUJjvyf7HwSAghJo1zFamqkwlCDYFzAPK1Y+M6
QBOtjusKYntBR7RtXr4huL7hM+pOaOmWXl/YBPoyBB5n2UrJIy3B9HDwN+NhYs5c
hbcRV07YjUOuOCMgXqquqI469F29db3Wv9dcJbgFtUM+LDL1zlip1z3rqCPudfyT
3JvCMYZlKfAyqJPzzxPaT+R2CE5bZNHiZlWMF37hVlypBJ24qzZxiJ+gcA6CziDk
30XjOZPI3/siDo/pdHrGEZWNu3gqdcDSWw3fMjxh/aVVkMwIM5P2GLlD9HeZRnzN
/7HIALPmCvqTtG3nLXASxO74z94jE8Bu5xQYlMzvc+mCMff9883A/6FQXLoEhq+f
hmx+6LmE8Cr1m01tcw1q3y4sziOcVJ/r/FbXXrmxon7urRDWkjvY/OVopJvBs9tx
HIIt+m7M4WI08+Sg1z6MsYoVUEUF3fE/lKCMnbPmVHC6J3zGf9WqkWBy0IaYx3IC
tkQutld630bjg7Q+oeYTJFdjybcn0cnBHUfs7zbGUdniw+twcTXcRgqj0HKTNeZo
+VMjj1oCfkLrT0o5i11Pmt08ecG2hjjP/f65Hqr+zlK1zMEJcj9PI0ZbQ3L7ic9d
VCRdUFFylrjKeBYSizl1Z98mt7mxeHXc4W+/DqzJgH3HEIuxHaau+LwXf36DRnac
iKyORh5/FVjj33xByqOS9xyO0u2cOqbuR6oxoPwBOdnwYHTiVlXfTzC+EkfJDp8j
FSSPs6a2d0mIvRKu5MXH6aDLniEK83PUyAgtgHL94ihSxHfpkUxK0Hd0ZDywf9lG
+80o+aHTgxSP8kBgak7B8L/trCyQHfTlOMjwxUq4v70QIylUpRqs5U3yI1Hg3JaK
p7xTLimFlHItqbp7dC4cZX12pMW3KY2jFohqJLolMfE3E6j4rSHoRypyXgDNY1vG
M1afu9HR8UQSEN/RyUX5Xi6r6SLm7nSq6yDNrd+tm4trvgXZ3X4bDw9Zn6CLSwJx
MnpN/8o+1e+pn0K/NaIeFBtUvRwoTvFBlDsOm/X7YtfN6MGcpoVLQNjJNUcwx9jV
Q7EHsT2qD78/pIhVpcsc3TisJhuBvfWzQTLZwOQKUd0AVstTzfFmOouYw+JJwxL1
LVRJ65qOfo8PGbPxuyFH6zB3YRYua6gOZVscCYmwv6PiyUAC65mWupiFGdDSkcC8
t8wYqSaJLNVauLnMDrUlaA2vEiaWkrvbfRNPfe1QlfgwMD3ipPeAlhO+UmyhSIXm
BIfRCPvCw/J+i3gv/7/N395YUKMXoGrqxNzvfw34HmMgHkQWx79EROoWmgGA360Q
In5CF5ZqWX9QO8ZnGKbc11A7GXznw/2pVKtg3zRvC9+15O6OWs1MOErSL8uTQx6H
25iKxaVMgDBiQ6A4LLsqarHm0rd8kCLkZOwlKznW3457Q5tDXq433EwDnCWHVcgQ
6Vel3O9Jpq/dyzKKf8Vs0Fiibp4PFzQ7zN0tLK+gRIzLrV/gZRFc+w5FAhgljrdf
jN+vlzFXV7zauGSrS+GKZ0j1blXRc+t12Bv/p1ZDfTifwCjDSheotpEL4lzUYfP+
+Iz5zZ9BRtupMtMGNPaXPjqRdsrOENONv+WbTuwRW7n4kgsc7fxkUGUCEoYLrKSC
uG3wWyMw0VyBLHbZimVJKLcpT0vxqnHDt0Jtr3SXbmBGNHiR/rRANUHhKmAE+say
0ZHZrS1HHHQCdSxtOi+K/3foh5XDtv45kLn+3EczbFbZGxUtNcK1pq+G9w3BOcyO
AQbUlJ1JnDmsmx0c8awlCw1ncirD8hO8Iq/djqSlBsLO2H8wzfyKpnOHIx+oWu4V
fQA2Kmcjncy1OmY8ecKF4cimsDZZdx6+VDzSecAuqFAZtx+PoO9UMRJc8T9FuCHo
Poy4hsg4i9oHptwGyGyZqSf0arb7GIFa8sVeIYor0pm2x+Z7OdhxqxJx+OqBQ+lL
c+780aJXzYGXAcpQFE6QEHr+8xRMG8LQGc3Iw0uypnRzykRy8YMnRvG0L2c7Odp7
iuWq7w9BwqQ3DrcJRSK70iMCrZtJT4NlmGc0ZUr1Nj5aArpDIZQD28n4A6+jcxcA
PYrbtkj62Y9QkjWoATmaH5TsMgQPuuWl3c3psMvhwe+Li1UzA9zEQDEKSs1bGmQB
/d3AOeHnXauBbvP6fIE0XRMPy+SGZZZG8AB8PvV01FjSO/0dIZipBwJcjOJ9Ew+F
z/gT/s3W9uBzwja7iw2GljqOz6khmqV6Qq1MU5Jkj7aIh6bodlFxH4LG3JRSTrI6
HOK3GRQgjYBfuPjNDiV5+imGYSLwoZ2CaSp2bCHYEp9snSGYsOZD9Eo36MWbc5to
LowP49YjOqDsgzm6qtpkombCwI3u/1b0VRcM6GF3yDloXtUx6BzKDge1riBE41LR
Ue5J2bGap9RAODNrHdx7HnI0U7MCth8Z93AXmNUKFvl5XtQfLTVD2N4dlobO6SrL
WHj9yf+Z6MNwxC+tHMgPXBRdjrYa5NlirvxoJowEtagpB15TWI709LvDNzIYyPpG
5YyrmfQ4DZLqk9hM1ZxrVmRIp3fqynnAdkNDdrV18FBHzWEvQRsJXf0Pz8ADfjof
Hou3iqII40FL+wUrfOf02zS+6hBG4NBBeCgnESSKAgQdcJwhhvuHwU7tq+ZF4hcW
HiyosyM4BWOAZSGMIGxvckyb0UWqKle9fYO8kR122iVQWPIC6rd3JSVdkzzPwLZd
BEMmiYOUT2hs+c7wQ8MP2AtBjQXUJ1qUkYtVtCuqLlJG0X06/8iEAESvhAMeFBYi
pTYvvl1NGGsNHQfted6dxdt7/QbRDgjyqYCCEV9vqKUQJS7UgVRPSdBP1UHdKQVb
A+YCyBjDQ5zunPeYXKcUesObquN6letnlaSEP9SoRf0MLklZ0BS56yaAT0ksWkcd
8naZuce//YmX3IgiJ2zh//nH2mlymy8vlOOGPptRAUpZmYN2PnzI19TdGAE0wgX8
LkLGayBZ9Zg0iq0/OEOYM62faM/O7oROUwLwz+dY836QcF79dTU0JsROEWDOX9GJ
iabwG5S0vZ03I/b13LIMggy+WwhVsWaO9qfhsi8p52q6GO8CVuIhBsjbXedtd36B
rWhBYZl/wSETl+3U2zGDzzzDhgnLag2INkU3UHt6YtK5s0u/lq1i23iJoShk0/L5
Qz+4LInPz/qcn60ndjM/xMvio92PISZKrIQLMdQK6Z096kOHcpopK5oGPiBhcrxY
6x6A4jDTOdJtn/iNWoaW+O9BtpbS+eYSW9mXLk6G26M3p7f5UhLoadQXqMmRt17X
TNNzLvtVbnDBqLE70aztjCBuz6O8H5FuKIC0t8MfN+sl2CksrhZn4nlsWdkjVmtD
QMCiIaf+rWv2PaWH5cPlseaWfayWEVDCgl6TfhAh7XEkgi8dHjJzXjdF4i478EJb
B75AfSf+l4OuiCw7YqXTk/w+gJRemQZMpnmwHEfYiNwp6eDaHmkBfOrArG4BBoqz
q5BUTvFvy5VVpvrOIQ/b9P5nM55wzMf/ta5cTfh3rvYjO334OqnrlvrKtFM5NwEi
vpOqaLjvAAuLpyqbiwkNRA3Ki8Z5lTSnZq+2m5CPhnw9sGVyIjoYrcKIbwTaRwhu
7H7VOadDPD3Gd7dJY3aPsjq+kbClrue2yCQkFVh3rtwFAphoqrBs3ERqZNzW8sdX
cszr3znDGeIB/5LgWXr0fHhxXqSvXA0YZoiNDE1tzSCWLS52en2rRwLkjj/tHEMY
5zL97xmNqgW1z71g0ycLLmu3oud41db2m01vk8nY1ChGh4CrBOtb2BlmHlXAtqrN
oYL2F82BKBJgzCtlUklQV1jmKkexPazCl6sxa2ZOEc9uYOw+mNfWtHiqDzMJ5hRm
oILAaMGB2EfPROsd7SYfcD3q86Wm4E4a0dYPPmUdU9P2SjgicDuLn822VtKPEiMT
ybYn+E/gxDHsK7u6sRu1bw/5+F93LBPZOpkLf6r+W3pFsmdg59/lyiXUZ/c7lQsm
uaeax9kXBE3FLYjrZFWz4necxxetQfQvsEUmJ/J/J+nLLn4t/R+UzXNGd1j9PMYX
hnj9UAQt3oZbSCkFpW5ARwew2BjJFQJTL/unk0h+5cQDZQZxsOExKBhDjMuWhKeQ
g2gp4ptMfZFFysDJuaz2WwKTe+DeZtR7WB/3z9cKcWD2NAtdhyozgdgI9Shk2MPn
MZ15HEPK+Sm8RgmwoTpsTgZ0Hjal9baiKJpnEpDNroc/809o0TJ86cqA0WElE6RI
hATyRLeVvY/YpmjHtnTXFAuRJkISHGJbVipJgQO48EB6hftE7G422vOLXqZp+4U/
aDhN+m3ELKM2CkNU7cL+73sHdj+7nh0XRHD4Rz6bWMWErYEYvt3j5ctO6UnBI7DX
sg4MFrXergC1kKaj1mbZyO6Sk39tX+M77ArBUX51DSVu18MPp4AhazJ8UvaeWOdO
b0S4MNnxlIEVlEekwSQeW++ekVR3CQdsHE2SYXz9o0OCHiRzx4OJXTm3mpR/E5la
mAN6CLPa1B9UDelzABUg5Yawe7KZKvd6SQGzkUdXnZ+vkZQzOkI1vC9J/yAEYJdK
3SU/WRbzoWsWqi9uDDuvz5xvbjGHuhW8ZigHqBvKe2gDSA9HOQigjcIC+x56asyO
BOraD+e8jvcP9pUCcy0Sk96dBir0/uwPByZX1OgtTI7xeCK13R7oQCaMnNnQmtXb
0LRh2qfgOm4IHIj4UX+HKOwF9FBZZp4K6HqakQNvNUJY/HiT+94q8ejLlcb5snPo
BUhH+daYDl1Seae8+F4DmYLDRCqITfGRlLop8whvg/1UlSqVn2HYDCIX7tguPImR
O/87VKjzDPVE/6ev68eAGAbbbXbolkk5+JTTCAd5E2zPby2IomiEn8a3lTfzEw9E
supIPQYqrh3sbVlkcdrcVvwU082tfr6ULyVFbAaJSaJhbsE+BvYTX/nMSnIW7/fr
Cq0XfGbnJ7n2m8B0E1zhyCiFTGQ4sh8zGGRH62oeXHAkBDW4I1OIXeCmsT9MSVyY
/9nNoCHpdnv+o0uTVQ4OIQOm/NbQ/DNOVFe8SXz13rZEUaQcTbXMciRW8tl5hw0u
K9XKyNdX3Wv5FqnYIzl0xz2USafuikCBFIWCr36lp/zc6JxgzPGFvlzFF8lrmNxM
EpFSgkePzFXBZrtMGCF14NWDeP1nX/btzhvVHoT45SnZU9H8o+LonV5hGwCzga0k
JbB39G8i7jd+Ipp1cNSr0gsfYwov7b7Gw1qcySLOPJQM7ru6BAVQkosmY40+VwTh
ADAyrsKA1VK5YRPOhT/SPUyuKXGPYb+AdQNAPiwwy0v9DHJelRBXjTGluhwj/UCW
e0H4sbpnQPVU5nYjGVHqNsowfnwjDDyL5oPAY9S0kNRlYa3mDPBIEcxmzXodsL/6
luIovSl97+pJ4lAb+G0kd72SNuZsW8g39Y9yFN/DKigLlZfXzX9oJTkGNMsykBE2
nUFCHY07r5WdWxCZh1uBq0I0Vlt7rzxDK86ATNeWiWFADii8BtTyl0U7B2zezKGJ
YQAgvbgD4YUgc2ttoK+emXCxfR3/uVaGXXf7w+sUUq/dIc2JlCIMGZVSPR/68m79
bbpkx5pJnke5oS1fivi3FFNeLkVv/Fe0zg3TJ1SoPslJfRHxH3BIcm+FBZ2uitOk
Pj2kWkaSyPUE2z/2nSXp0c6x0cZ+aJ8iVgvKmqMHuWQSAs/pcTQamma/6G0SB4ha
kiBxl2y2rVDbT6bmQxnajn2RVqMYxgQ9R/GimZDYqzitG7HjUuoYpXorUur+eb9y
rTXXY8LWQyZJzC9Ka8vKDw019OwBAtdaGmvL4DlOIxWGANYmC7wpYYrxZZwHKzet
cAq7+FS47PW4P11kC9tTRXY2++NJ6HkKT5PnWDmYKGfkPhDAuFYr7cQOjK+XfaSg
fU+LwzM+DvZ3YjB8s31V4xJ0H+EXvCBukzKwNbbZp85dORGp1a8NdFMI0NQ5604k
QJ6eioCkn2TnVAO/zN3UlBSDaRPEqrwDsecfIk0F9Vq0sIaqPQFIxUwV2ZA5Ekvm
OVxKdX0who+I1UCBNtI2cTopCVouKaB2kgx7+bugHSBob0Dt1rlMRuhYNBcUJtdR
vxjvvsz72IAD62NjEsPEcbfo66ytt1eEjNtwCMe3MYvtJ3nwHUGAaOxNeOpOqeDh
dWQdnuEElmcUMBs8yrZ+jIrAWn0eCaxLn8ehnxzr4/JtKKBVKUzN/ElNrVTSy1Id
TgRTzj3r7eR68COiGoEA2cpzy5NG9x98EwOZG87iJ8D0yH/g8zp5Eg3u5aDqjnZQ
2uLEiOpgUaASRUaVh1ZxKtdpLW7V/PigmXiF1fLkDovbUwYcQE/zcGgFcKMvq7gN
nd6NhE+VghJ4+6UoKb/Li7bTESHOw7jgzLpWtQs/ZfLq/NC7SGsaZVD0k/TBClhr
tqOc417lDlfNoNJls8lILL7jdOXrdGJ2hXrotV75P0VetgJuSLyH5X8kQUMMJa0k
mGWhj6dVvKhs6tQDIROFSeVoCGbXQ3z34M2wcQ1Wx55WGxfyzFJFFw2RkKBhh0WT
2BBqW48dzwLWCwe5v3uAhajJZdOW1Rio2EUxxDa0dEUXA71N1byxJLIjYt6pYk2p
2ZmvsEDoTggsXGwvxhYRysgCIwsykD5otL9Eq2cNvJcw4DNR60RDn6USuoYTUTCK
beqtSF42pjfUfwHxmQYXL3P/zSM79pLzmuvXjm+JGIxoUISZdxuEZVyCfPs35cBO
GzStw+ZA23q55vfQSRfIW6mJfAAZrILbFVzFnOX76VBlCfEjnf4laQSC3EV73gxs
DUZ298M5TkMxKEKZaFYPxmlMAnZfmIGTpHNknQgXTOMGUy4jEqr1Yezym56S7+eQ
oDJycSBqbdQNX+9YvnIv1ecF6Sxwj07LQJmbuggQDPSNnVKDIL4cDIkdC1JdPwCy
Ys1G3ANZmud/vcHgKsQC7bXM6ftt/g9KzaD9djy/I8T/hy/ZTY81A2H1J/st5DpJ
2biWM9g0BHdUBt06nzxq3FMmoZSPArXpmrwq/hmzw81Oc/pitBZPSehrhrGAor9X
Ihp8ll1wZIzutb1C631TaSYHegQOAUHCjl5Dc03QRB1P9YPqZXiPcuHpmuCyFZzu
K7Sblt8byJUs+eVC4yehMVfmT4kKuFwC+E6PQHy23NWBrarTlqBrcozgdmN+PhPf
16Y0YZQrOMMisSZhJNSm1t/L7WQ/zNgPO0YnWRWi0pdjlsg4012/pLuL1O25+jkL
aLckjZaehmhy77+gLMEr6Aq+TvPjl5u+FatfxQnsZSrTMsbm3qYgug6F6MVbAvkT
gsBTuL0CJAdBOOcEfbdhNd8/pLRSjODWytIJtfBTMx/VqUzur3v7gNLCbLRcRUaR
2p9576SIMlWX5eGXcHJXAll23Ir1J7p3Pa8LSOutgSpDYuH10PoTU/cpFa8uySdw
ZkbK4m8RxBUVzX3fQRUqmps6L0pFCK/2B1ohjbnu7SmE8WNifLSTdDGoc2jWOTmq
zap/3CrK46CuitWePlWpP6O07S5TUswK5nRK4wYiJr0vDVSYgsJ/jK3UHOk9P35v
bkO9udXgM0IHJzkiFXe88TojeYukhgnpddDac8aWHafToe3wYbqpoKbn5MD1KwzF
+QwYB6z3sJdvhSv7J4wuJbjac+32K3OktwDnqUkGa4FBNaSkip2PxknSAaj0SzU+
/N/Kwqrtjq4zJOkePSi9hpn8HJpiiq4CN6PZtupIJP9dw2QRAPDNwwd6zm8oBLaN
RMjpjtuzOuMx6ZYIm5NvtU9dQCmiGpMgcdhAK2h+ZkPALHZSB+LyANDHFy165iYD
F+hsgxyN4DF5yWBgerrX1xDpgo52Jc1xrKIhT8qy6HmWN4fmYw3p4lOfwpCCPMNT
MxpYlhV6ZjkmB7X0F65Bq74azA4ptA01kQwsOoGtC8wTYUvpF0u/p/cGiL21eS6x
c0u2UDIsYQZOITO5A8xbg1v6c7VnNnSdaCxYjnUkeDu4EelmdGrufFQuBwvcgX4+
0yPxjdw8zU9QFQWxrbiq1u86/xKi/bWXyqf4N2kZacAAqdw3vBXLTzeLGIkxkjbu
umCCngIJKDTLCfoGnfT+RJFNRN1PGCxwV0WnTJFkGC3KxdlQ1+5KxeXOktCtNu7v
5dRooR2ttuQB3Y47dAskShuTvA9REkgpfo4V8kVoLOeS8kmPK6wgChuenEreOu0T
W+oAFtiy5BcH8F8bnGfhwDU2QJY7piNfGeQOXjZ6Lkuul8PrnThTFDTfhLFrqTRm
tesoSUwessFWCjsIhTC762iWp7sd+TQS6MII8fT9sOvNBTbEVOn63cE73GbyNTIV
rePRiyA1lTSkr7gmyVEQoTn72vyOXNg+mDHM2fP4lagTD8aidC5jxtT8du7ljwQ9
CG0qiHlEGoPlOD8Dc0GlGi6061rC/hsnZuommxNqjahKn04Z+Mi6dz0Q8IG+CqC9
6QTnSzO71uXXj6QQNrjvce0U3SqhwJB/o6y8OqgR0AO0RzJ/SfeZ36mQEt9Vh1BR
DmSzOhT8YQuSoLqGAdURSiABOqgle9z6Ddo/Z8ecQC4h4EK3UrirH7QJfVC8WImW
k+V4CAZJvqpqMWE0BD5RTFGvTsj6hvcGqikbnyDH9+4lcguvr6yEzj2/NHpiVms8
fl2ocLNy3QtrHnTYHPbY6KmbBVh3wrJdXTX5nxwSia+80YUtHbaPK0rPVUrh44VT
pske4rW/TX/HZxTf8o+OsySFzkRN+0l2ducfv/aSDNRuwslLVZicvmyKDlIKUO3X
T7edulpV/M5nG1/6hb5nc9fGrhgjIrRvSXXt+Gen4g06mSoKJDNMkqagzDEAbU94
GIkRODg2GLVavtwhOmz3XHq36/W0GUEC/ETakCf4lHoFgLHDVOvq8ni65bD2YsbA
KXhb25p2O7waFOd8HjodfZn5siDZ1+1vPgoWGYM3v9rN/GKakNMRa2LJ/x9i/Xug
XleLp+le6KhRjjJ75NlnHm5dhsFLRaN7GPgDjIZagE3YA3OibHeXOBvMqHlzpuLa
3YZSS/Oq8DnYlnuoYOhY7rrNFfjD/ErwfQP4d/b76enr7N86R6Y/bBobSZXeQacS
uryxZVGhpsnHDkyvVGuZzmgidInBcJcO/xr0QzKTpOn/zlSyPkSo5H4W+PkjDAxB
Hvkf19jeZdwLAIGO784ufYDhAx5uaBEHAlFQkucMdF4JM/RcJllR+vooTmnDXGWm
n/UF9J1QeUFrsfH9lEQSYYd27ADaBRXG6ZmALqAfxe3XM/h7KEYdt9CHIRFdWNVs
wVv0V8t+a/ChAkYP1z197TTGtavq9yXCYP6BWAw3Ve22ajy1Ks1OSurPwJV7vr2c
KVb8PR5rnzN2bNHU9MB9T7rXfJsuSBuXkVCVjMVaUC35S9TmwL4L2GIWAlLK4tnV
s7Y/x5GUcsvL4n5DVMMPnpckPVnOygeM3Ql9pKIIM6I77kxGWnOuDdtR2rpiomao
rAyboLWnISDeBslKxhs6u3SD5nVrHzNSfvOLJ4Gen6ZB4NZzas0p+H83WVO64sYF
ATARZdRpqFKUUtgYk6V7tzkbt+ZZSviWDiFKK5HnauaJBUCUxeJAdtRmPYv9HZ4G
jtoGi3aze0zXHZuKX/Lg/EVLUXUx5neycQSU4Au/X6btaZ+ZPphBSpiswWGQJCxJ
CKEcUP4M320egvfUC8QlxmcEuAiWutqQhlvRsOmty5yjM9O3X5lXMyCW9FnHJ2q5
jBENX6hFGZb4X9s7EiHbyfumihQpbo/anXKduR0YAKBhbpAJ1QcisT/0TO2UAUXC
Q6MVt2PM3Br1E0oHVlIDZmG4BhErUPayBpeQwSKiiB862QTLFPC3IWr4MMmYYGhW
E17vAkX/QRK8woebFbsYevqn8mOu9Bm6PR9EMhBqOVeUtaOzdEI8yHyR0kriD6ym
0uje/raJfaxyXL9+zjXkkPclnVW3+WTemR7S7H8sBItcIogu00c6ckKenGXLTGiN
/qIb/Nf7aSl+w+iVqEL0yYOh7Jw2Pow5vA9xRoFARlWVCDWfv54c14uAqWjxB9fZ
mzf+J2nojuNTOaR2mHbyihO6/rnP99HCDolrg53FNPttz3YfACuZPKThZGGgkZPr
GbQauKt38p3QTzZOYbHAo845MJAGmx3Y22pscluklNOPBPyKFyICng04NF7P1htA
EhR8k1fmee3bh/4v2D0iD4FAPUKt6/A7T6RyrEBQgcY/kaHaVdJcqWJIPDY/zzah
TWzQmTDcyr2RffdAXSUnnYlUrlikjbdDCTolIR766bHG5/5l+VWIW0ZP/RTnlfZH
7MxOf/nXKZLx6XMhCm0mxsrxnmMWV91nEfyzGMhdUPzMpaicY7c2ru/KsLbOhHMI
GEgICBDEEY58eVRO8vZFLJ4/C8igKjq93gLUxKPmoDERpBAylA/sCjAlwvM7iShH
hBvz1THAnnBpZQsX+fHB9TitXkTx+qBzvyjx+DaQXW1bCMxleX+q1Ff1m897++7b
mCUzG0Pos46AcI2aGOEA/4U+6jlAOACGhiU7etfwt4yeEBqMoT08PO70osYYuQc0
eUvKWM7ya5LB4HBT9ixoGmckFC+PHSGG14oue5cyE4LyEnNkRcS8HPYOxryphsZ1
EyyZumaDYfiT3V8wy7K0OxMhqBcUqWhIvjnb6KLDLeCkO04PVxtkCo35R/Ha5DE3
KqxYqG9Z51Yw8eLhl1UvqbmHZeBK56Q4JTOt0F/SRxbjQhPRa78I4OhaJKDkfNXO
FGbqWtej3Yfk8cT3XasBWozThABbe3ks5+z8LAa2DioXOm/Cz3qm7SJWqQpFkg92
QQm3XrEDDNcgcbaQrlXddEiRw39Cc6eipe2dC8Ts7XJ3zcI6qjP8MhPwT6nUzjzJ
xBQJuN+z5uVLQouBNvpxKWTobYj8vgLmww890rcZ51mqKJ5rubuKB8FsSbz1QWcZ
KBTuavGlKoF6qvG0PL5TNNor11P4wWYuPJBhrbK2Soa3RzbbZdQ4IrOI8cI7IGRD
wCYqqZnDDowsBLcScQ1N0DMfjhIHrF7JmmCgQgypct0uia4i1X/yqVUE5r4JFAHU
rs9v3Izyd0nHqUFwJ+fzxWv5UHWWH1VuOFb1pSL9yN8ZKjBqOfpMxMv/MCcKPYI+
hegg01F4bCjLaiMlkc+h6/uTZYeTl2hDUA2nsfRRbEA1jGHJe2ZXXvYCvIJVFT3z
wGO1sCFIQwYCfjmABLwIP2LzUEGbRjqMU3ekiiMqOjHE1WOIQSdHybPnq9GcybB+
BTs7YEv9hOLEgew+/OEuygIhHxTX0IxIi9GJtyguJFAIQyRGPkPjN7JAY9Fp50SW
WlGjx0AkF2B/46DWMwBalIi4Rjd00KgAIOOcVayoZzXsWixFBzVnk6qoOIlpwo9R
ZJ7blG7c+VxPDMhwa4gQHNLo1h3jrOZQQMEQQX86VwGAWgDy7Jp6yLIiJ4mIBdRF
NurN0wOjfz+j++8M4hbNEdhSiaa/1attND3XCbzy7c+KlP9QWsurPWZfdA1bsLou
p5EW7nygFpfccsn5xSFlxbi4MzDgj4sXnzVwc37dbVsvbeCdLgI7GBBHGpknM5Ks
/gLmkCxmJqqS5efCMAg4vo7+K0n1uv3ZIz/7cHDH61zd8I/LbxiXjQIuLsuz30aF
h0NyYlarurT10sa0KsBl6WMqXaQy8yFTW1ebdK6KBoQRogiF9kzv2gTr4dxepXU8
+v5vGjA8soMoSsNDkCCUXBM1vvL3YG5O41EGVqcLz2Rcsd9A1e2l5bUXcbW0km11
85ULX/HrWkP8WI8l4gS4TyCgW5thHUcNTZZBKWiaTAvhCFmLIjtxpy/f6qEZyvao
fUGsOyqDix1t6odAv3ijuXzV4w3/4CjXTzKmQCuYR8SUG1JWa5L79Ln+r77B5nB9
uB08PwZAtAw/V+1UWkfKwJcnqr+VT16TwW09zgHiIs5uaJ5DVGPXZimx2aKQaguV
W1U5cgcWVzGtuUvh0Me0uEdCDY4VnevcfATrmg1AotVYPsC+7F642S9KBRtyl+et
u33b/mQrq9/Ogy1jNnf0hA8ZCRskz4aJ/ufEmROosXoBYX26Ys+H76Y1zb1IqEBp
pf9A/TsqQ0F3OD1E4Bwi3YhQ67Lp9wUc2WI81P4n2YUSdGGgn0UHeujeVitMO4+I
yo/BuXE6IE1jep7bCd9VGK+Fsf97HfcomXu5tqUWvmpSIDhsxCf4/6Chdx7Ay7FG
EeHw94CMBbbZkcd7cAFutSy2I58qZoGAIMc4GAtxfZ47iZs9rANV9e20zzL5anCl
3p2vwxVBAlNtcQyfBDAIQjJSWFeA9Wka5opC1FI3HH7p09CjqYo/dBYlS7O07o9X
it0DvtZaKPagJZvtK1tgbOBPJbhlzbXxCvQ/y/SLXazG4eOYMsWdGfnbeGN8AWgB
2QGBeNxmuD73OBGZDCQ3SNL/wxRcVC1yCvQBmLZmDWWjndaGOYkFMEW9H0IC+hsB
h+LoHBuXvPVi9VSxMtYoUzQEE29SQRem9O2eJz906cYH+1Jg0udc/wVY+NkAvCzT
lzOPF9odbYdQ2qssctj4/P3QjQBYHCTyWbG1EpuwONbg2vU+nB3EpIkU4kPIIGZY
A5I4736Mo0+x8A+eznRsTAznpKjmGLqJ6ZTjkEACnxvndPAnTwrHnJbnjteDtRtf
AHZEibse9s6ts2lEC7mfdTCdsALubOZsBuZM29YUyz4sVduUN2VbQqxo1QNgLd/8
p25vyK87S90uQPIkaFn9z+nPobTAgT76/+GAN09tTbftThLpXjnibIyQxx/GxHYP
qSRVptkuMoTzy+dxeL4LtsHJ1izBhKijqyp0Ms55tKNWPRvH4VeGBQBlH0tvtUKH
IECJQtG7gWpnoicooHgbGfBScZmLAt+JGguRMNlSoEGU6E3unt0mxoyhxRamxJ9B
HMporeXPU7NHz+xmcQ7hmrthsCU7mzHmqVoi0yD/8dxtmt9H8bEQb1oKJRmHLgpH
nw012hnY8k1y/ebOshCRK0XhhfKn7HP+QwXVEixMVZpxhzyMkR5MUNvNc2/KKLWP
wmtIT73GxAtkND+XVjx6zbKDKe/MCZ+QD88xcy4BgJN8FNPswdWhuEgXHY2aUsre
7Q7t0zzr/4YKLvUe+vINsWhSrXKhNvW/XZX72dhOYkPOzhPfPX3JxTyQxGd+5L75
l22cWXgXw9Xe62ETOlwV6xWHdGeHk7QMnurFuuWqvyI/f0+jifgxpTcvG9XnA/U1
Vq7g+VJ4nHpwXmPYQtLkmHaTlC36edsUCyf9ELZTIl3pt9m9ABeRF8M/hsbG4clx
DVhTdc0Y/vrdB1mbc4198zxxiAxdnegmjlw0xDRtNxCdZ2FFBDkIY+IMKv+zcolK
/vMgguss7Di3r27TtwcPnvvrScF5kgUnymFZo7qgfSQjoC8DMsKQf/PHCG6oY1eU
5xS1vTvgd4gulbJUBwA+Cudk1+2KU6fcrPAYU9Dj7Y++8Rqv3906mdkjw1tghg2H
e+JhgMctn+Fi1d1F1drCH67+iODX77oYFAnYZW9LxsvmcgFWpoVBUdITiMWGi+Ut
chQ8iqvgZk7SrN5IHUiN/s8YBKqVtmtDobfnzrIdvIyxTNbQQQmFvNlkt3ibZtCj
83Cj2KST979LOtZH7k6s/Tgshr8dbiCPFAgEeJ6e+4S4Szmwj/5j3cILhLnvUHYE
s9x+CJq2pZciBXzqU66JBU6OhmXiISt0O+kFfKbA8+s1O1InKFFDh+Ic2AVaKJyk
WtfzB4i+b/+y5jOH8QsbB6ZFuNAE2JH3rrIIS+EXvN+zOeI43TsYMRnpiUFTQkug
Re6ioUeYcxwXGSKhzNEEbdL5LGodCfy+zMpu4hrsUUOyl8pNKjFDvsBLT4iC+Bqt
ak2AmP56jy5DqktY2sA2thtDB2ofOmxUm7UAQqDJGEIFsQfdx9gLRsCrNp4gBWdf
nPCyJuqCqYSREGpvSZvmSDmr7gOcCHo59G1TZWvjx7xSYXr93xfOEq71TN+y4O1+
2I3m/FGfe6S1i4znCkoQyPzWQWm1jr00IR7Oz1mJ2y2LY7xWl2dD6k5esCAUFz0V
nF+UTD/MfOscV3BLRiRIfnme9NDu7QjJYX7kB5eBaViSvL6JyRSqyixBvY9UD6nx
ctyQYuV2Khc32WfTSgK91unjidm+Y3BT6kVBkkrbcf7LuRHFbsQFlgKxbFVNTw9R
dmKxsp+tK2Vdp/v8K6AMsiX8Hj59214BHNmjBospoc+x0wXiFbvYTbbwo/CUbEez
Z/1SgR4GHMd10TmM9Ydwmnp9w7U/28Wh9r/jbNGinbCFgD+Q+QXBp5nXLAeG1Rxw
jJOI+pzGc/vZrObw9Am+rFsj1WmywNEaz+mT6J30b6mzdBokQM5SwvSbdxOuwEZu
+3dJEZgNqX7RbE61yPFX2mt7+scs0TC7JyyCeaFxRX3Pw+pJtE2ddDOlNUz9WtOG
ijNU6iFvJ8y+7CzF3+Tv1dFhADoRZYCVtRp8Hx5U76wNdAAuPkXi9GA3+ag5xp7C
hLXVf7qCZl0QHWHv/xmLgRkySbfgDNGzb0CWY1+TcvjqCJ8ILKg6WSEsyd4uMwI8
eEJoWvMi2zaqwxbK41eN++MjxJ2BIgzFVQmGp6zmk5kZ8DiourNxvR5H+XEp7K2+
e9BhoplTDzFtnvLd2tv4mJavTEOUmhY/KPVfHnu3+PPmytYCY/BeIhUZqeRYGHQS
2R5uPI8eCflDjsNZlXTD3R4jHJ+c19IX3bpMNE9s6Qzk2hNCJcmVzjJFrh+Zxg/I
5dIiiza5O9ukVZgS/lf53zR30wqQp0C9kLOmKo92dn2MnlhJdxxtGPMneGXfYAIP
MIA5JW9PXX+d8tOZnXc9sNqSfCe4UlffaXCBwKNKry8KDOtKSZJV3sKc4UZJDu4m
TLj2+CXLF0yp4sjTYLbpQQEgJhAIvYSz5kjbxvnIjxpajZ0LW4Cv+QJ56DUvDHGp
R0vh47FoRNRnE7fizKJ5a7bo6Dz8emi6qO9NtWorhSoo1Tw+dr7UAbTSInI+8XUp
MBHWZ8AYDkMWCis3Dg7255xuCCregsQb9hIxuNOBHx7gY5V3odMMjEzNoParmXU+
8JL0vH3N0g4S39+p+lj73Je5jGOZ/Y8VQpeUzpDEX4hb/WdXGyZmVpfCNU5LvqIR
Tlmt5oRVMUwpKJ76Lvx8H3A/82wH8TlIKEV6MKmksX9FBXOGPcIX3/STkq8BUAhg
Bvqca64LvVLIbhfwhoEXo/+sHN8iB7zkJ4CbmxgkrD3rLtcgFCPYXhTS6V865KOK
TAiUxrV7Vn9WX6/F1ZH4AZnoqiNGRAyTJZheEV42Ao/xBajjGS0fqJpp014RYPIt
P/CaLwVyVOkUoWKZw1KT1y5GTf2+MT+atRP9VkUS+PnHpQo8MPO/sk3D2fPE0X6D
05roFd3qrIdvtHEZAzVi3nXX/N7EK6RSu0jiLpa+6U3EwO9QSQx5SEWe6/MOzhqf
wMMiHIBWvRDH52WSgtxPjuao8Tjr3eeA4EyzcuGnnb7qIQpxpH6NtuRsQDYfeXTA
uL4cfRLtU8wX2HXxYP1Mm9h5pEV8CHd5W43II83t7+u3ZxoLrKtqblIeQf+afUGl
qcL4sTWGF84L/PSebwxFMRO/zNQNdW69m5xqGN7gsve9QVebeTqE31YqsZ7fNg2c
PelT13OpZH8SJ7uDMPwzJ4Gmmc+6W4ItjV2Npmho6m6UhGovq1fGfp1KCQCcR4Y4
YJdCLXIxAAwlJE4OqPf9l2119Z2XfrViP0m4qTv4YD0iRciYkDPpm3blUBifdFNu
fyKwsGGdHs7ShO+KRv2yAuMw//9p9BZWMZpypvrq6s3YBq8Z5Naz0Ypo1aX+cBbY
iMnLXp0nWt0oMdVXG3vrEA6AftAlIBTSwNKRB6IS+xJxigtUogV/T6/DgOeYjmzX
zGsHz+njytzKcHFVfQEAzp/XXC2tyoooF6hAhqW6Bg67zwHIIp0wz7/Y+yJZSqHd
+YxAUfmZhjdKQkZskE4JUEHF3Hs4WIYaxfEh15xVy2C5BM1FQbLQu3EPfh2z4RGg
PzTvJoSRglW0YAErdJGgcTfv+2+L3fxvPCiMwVD6hVIeQZst4RYHgzkLX4qva7y3
Zd12okZT5yT/wC4eWew6szo8jFyq9Bp5Jo2hnMVxnNfhNuJuBZljHqMk3W7CbTub
BT2ZuCevJR6W1TCP1cY2Ta1wzI+nlc+SENvIUe5YOnOGJRQeD0tpslBtahjuB8Lu
Iau/jUklTKt6U0ob0uyFtVXcv6hJAFiPba0eaT4dnZZbYs6kkvP6q7GIIZFyS1Kn
zgR7Rnb1FHcdP7qZM8DsTCKDU6J6NkPCHrCuTocvS3JK0aO+czYmxn9dExoeAlf8
N3elW2RebW5JtCRAmSqYqkYGewyFzgrjXDWt6V7pVtSJv60LQpgJanuDCHHZmnjv
0nrKjC1N9YDUbdZExQPjRrwVDAjukI7YUIzIHpnXztXUwKADM6cU4xk8iyA0M7Zh
3kg4a6TQWsc7bPtImlMLfoegliC2g7ExY9mqo4B3ac+yBd2zByeZrLwFyG6jnR8F
b9E/VhArtzQjsm7YPhdU385CqkDGSglZru3Kok/yGehM4FImH69xVH2cRvSJWTTk
uWXrLILIwr2DhGhpsPQgH6QC+TzgJe0KbPGI1hy9PZzmXXC2uKj0ReJ8JbpTA1A1
5GtvWVo90FUA7Y90dt3noMNbwur2Pzi2lW4w9Nb4MQ82yMlBA+CDDHJR/CLC9TCH
Y9YkVPjabc7FMA3VkNwl/11AFqDrWGR8eFKV3qAvkAv3bim30EXEpmsv7F0+IChQ
0vo7U5ye/9ylLopSDXKOCZcfoR0d/e3ADZ0pok/1ve2uhz+74hZjPDaVYQoIPnI9
aAolRZ05yGcl23APDZTff/klMJJeURKt7/zxxWLcTYgLdmVOkFp781b3mPyV0WRV
v4eIU2KwGqU9Fkubve/avSCuq8EpkMPIJTZYgjCXGWlUirxz8Q12d98g3AnINVl4
duY40nvi1GH4i6X2b3XqnjMbmqe1nm3ZBsRfKeO0x/4UPSbC+x+/1+PU2sur58HU
Z6Pk0iSogSxOn1RzSh7gK+zLNS6nD0oGTCjBysMvBpCRIxzELzw9V+qZWWou9ulj
C1kjWI7gqsxz8LCpyGNl1t4swmrf/gJ2lyiqPPgkMm4rnVdNbWf28sEIPK+Hq4JS
m1/BuqSRhsqNIkDPDif4fwtlrcBZiNPelRNpLJ19lVN8qVpzJojau2pTJy7RLKoq
pAcRSHUvUufDPXomli60TGOvc9BZrh1XmpJtGM6GaCGi5aRWAerj+YsQUwrVrwyF
VDiTz4zk3tq5IcoqfFM0HimpyCnZA1Mm95TUTH8CE2oFWxdUyiVvl5V4bXd7SD1g
K+Cb9+RvktWzUitzAqgQb11OxQF9iucXnMF5ZTaVXBu+0fUWBYlE7rsVly4Iirxs
wwRAwTidnTbVeXmpqfHf07RoxCbqZKxtmq0W5JhKk+CVHAja6RgNuMF4jLTjVxya
mN2Cmt7r535oWLRBgPbygrB0SFcMxRJfqqAtFvOn6JEJw5uEUAKjkmlg4Z+kxLZd
n6OrFAVTF2tat1DS5P0hylVfQtEikflwjxrJG+fiJfNJbwWCS5FB6iWSDyX3qKEe
1OZCRzLWHvSA8xslCNl5GPlft7vKTj4kVU/NofsY04djHzsaUpQV/mxVQpc2Q9sT
b5Yl1+05CuSSznl/jaE5FsufHhukt0STWKSLeG6yn1p6IFiTqvZNggNzpruzjprK
YLYCoso87rvmFTbfmuUx9ApdnHwNcq24Kp2x9ZqiZbzGgZfkcBRchsNieNSQEESH
sZlqCUY6d6TRcQcnSSp9LIg2h8cZfjjnYhssn5BVVn+yjY80XkY0s0DZVn4BKypT
Secio9gS9yqGU0Q7e0tJuJmn7OQKGhGz6g+ocN5gwaru4/tM94GKttQ7hYlESZtf
M3OsHEvuB0zH+mWIVRDejd+uwI1CoEuV4qW0dK+Aenhr/ZDmPKkG5y1TAa7AqkZd
si1ZJSjufK/e4Gn48HgIotQhKM8l/TEzwHwSU9rTsaUPjto5U2qb3llgguW/J6hq
aiMkI8dMiuYKMAzl6YOCYNd2jZmquq65zNdaN5MATjBdU75dfTLmSaj4axJd2puH
kT0sMQITAuRsYqJPEdtQAQx1r+/TqMSgGUBhxuzMStrytu3OJDS2g3iZvnK1SC3T
TzIL3DsCXErgEB8giDVTg72yLsJpVkHFVRaa/7RHtpZS4fMCzpzWzUIWUJ2B7dhW
ve1ph9i6plV3PqcDgJ1zhCzubbWoyyEbACzIY+VZW3lRrdFDcZSlpe87AU3AKZb0
kXTLNFfGpivOo1N0zbyW3FdXiknStsCAo0zQApaN8UURFltpPwybq/Vd3DCwjynH
FWGjMXs+fOGZDHV4AtgdlLVFiO/Wv9XFOniF9ljuvU1sow4L15nZe6PMfD28sJyE
pJN21EZiqQQq+A54L6R80YovXLavqhVfH1Bng5kISIGpvQxZcoZ7ilSIXdPZ2xBL
0wNQdDkwS0zy8JdUTEvUexGTPrOTQrLLgVLbmm+VJI2X/vcYhCmthuCbJYdIYgBo
ZPusnLogD3Y92TNJZyTy5pftrB/qTSvt5eQl1tnuQ4mVUGNqVu/dGu9aAP4BGRtF
/23GFjlOhRzRN5t/etHzGWutGnshtvpZ5K2uedAihOCNAswBL8sohtMHUCB91MrV
UH6G5LXJScj+5CT+jsluCy0fUEtTqwEG9VtwLX/bYqx4TLF1E/CJhyQIokIN9wU3
hKgJDHvtJoJeiGTRJMlwbsTeYYTBcuGb1BDQyHPLdlFqIKr1eUgEKmLMR2ER+Sh3
HqNw4WXh0qrM5jixQKtjMlwKeya9NlH8aAaJNoTtzrTkR0px5QTnBISp2NNRN9XT
lA5yCKsGO5tnr5N9s1U6MmtmfejdDWS7LD5IKgLZsMx+tdY/SlMXQXZZrr44T9Ew
3wCc4r1YdTNj2UYrtyYjYFwQxdzpCqnS8dPYA3MJ/UQXCU8lCi57HHD6UmR/kwkS
uuhoqLHXxWOVlg0gP7YACCHXuqJr/IN+i3pHmSmxsv8pZu6JO6EFt9JqerNgp/3l
iW8ssFVsXi3rBkxNR4sidtiW6PofPoob9n7pSul6vfzWW+Ne0Y7/ZeE8gcH6olk3
m5rQOFHd3MKnAPYnhxFPY5o6Be4Dfq5VD/7XsH/9F2BbkBj8QnHOTlD2Y9G3xeMv
04axB2hYkK51amFsxtHX6auEgmTM+51b6hp9XI5sEl/SYGcMyxGmLx2Z8bjgrEKf
nKm1sNIKZKazqPI1kL1KYwcfRGaMisgUFQ8sdvwKhP2iyhlMR2Z5i9M0F3vnLWHn
/ej/DWNeACztbzRHFtJouhy70HfO3czhVgFp5Fad93/QNSCiI+a+m2rihHVp/vI1
pL13GdKZeYkiiHTXSJnqrWodUpgUbbDdK/ZmHp51DeKl33P9vB6/yjwGY5ewY0zb
k8V8OXc6lWm/7IeqHXmgKcCro0QZRA7Br5+LgHxYqg8JxIaNUAPpjkFpdaf76vwo
AY0tTQ1ZsCVCLWjRjLoImO9q9yq8eo3NHckEvu3SqDcC4pVpa57eYI0+dVx8krpN
mecisS4QqFOaWNf4nhp47yWNOrODlvvvEy9DpSwA2fl+X5cDh65cNPyUxzMzmsQp
IFB6a0GNQTma5qhLgf7+7dh1y/Pb1ml7W5ugRJncRD/tdUX6paYaqZlJwFf1MIWE
ZmscEJdZxlOB0fOQs7WJYEUE+DcEyevLj4RLI+4OrU35mXEURrw0pOMR9bLUoOBd
gK9944ekuQFV93JRlDoX9oHeMOpO1VKBUQaTiqmsf9ni1TRanhYTq8R4gTnGjZ1V
UQ5SrVM3bTSWDzH+84mTT8WDWLrR+OnsBDNdnnLHcFB5FWrXuULrRslBv9ruYV0x
WEsojJpQF4hiYoWN9RSSh0FPSvLzZmYhqu1vhy9Y8gFSkm3aOwkqFIeCmAN1vHgC
MxTxr1bIktvAwTx1EGH+M+KhDtvoCAYBdmyb6kgKkMykEQGiEw0w9m9Z6gK5Sydt
tFrLM2hdfOZxM8LbmxPUGX8uyGJaR2SQ0P5+b/WnB3u3PMMopBu+dHfSm9RdbQxE
Er7N7uDF9b2Aknq0ibS48YwnSRJHIlQEgk2hvOXYVcKTkBqaKsLl51i5WHh60At8
OOc8B1nEwsrS+vcRNChQk/SrlNe1dV6DgmQYH6ugdYzbz00I9hC+8WHJVDfM0Ihd
ZEIMS6Q2ii4tcTrqVXx5pNRPG1Y0lyLefhezBva3gxkn568d4wYYXZN1d5dvdNbw
SprPNxSMivF/2QZfXtpm6wtKrAKtIxKI3lD51y/APlakpQnduVvQSIu1jQRb8F1D
y/sbVbvEHYecYWYMnpNsZnN2ERA6h9qVbCOgNptuAJNBfSlk5+TZDhAs3VKwf9Py
V3lu+2ZJ86EV5ybxOyC1pXe76iDReIEjCZkXMezWdr8Y/tP54vANzGbaqKdbQpEN
YMlqem+ED2npMxs9ykjoNaLWEbfUh9b4dI29fo6WY6uK7ukakOV16FnllK13x5M6
ldqNKxkUiDaI5HD6eGeZIhmKViyihK6Gh/RRJ9yOM0GxNK+ZYztdgbp+YfskNI1F
ZdCZFRGHo56qyhXUD9OYqBs2Wy5PWV9MwPn9UDmCPjv/6AVSQ6niVQJ3jyLhAVl3
7XXtLwOM4k/r6cUdr+MQjZJ6WRSzUCZ0jLYqogq98svLyRwHSljiIKilnkZA50bG
mU1IS3mg01XOG1lrMwc+yl8XMd6UKU42ERFOIDKiLECALRgH4bSRmSEJ4TcWUtTM
WQt4QSCMEh/4tjCSS2lRD48O/+cCqsNUjTetshHLBGse3j0nTDMqnMzfLsqn77lF
8fc4OvH9AstPDpTAdNJZZt+2oaWlXArjEJYvi3DXSjVFX6A/mmwEA0v5R1Wxr94d
fl9tkUtgSkorB/YAVGt2RWK2lkgnWd6wXMVrCNaDzG+2MuoGmIXuDo5aq8egt98V
Eb0CiQfM+Peh+E8JFsQHoWGAdJ2OKZkxj0JxMVW9dTW2VQJc01U6zo8cHTYFiUN+
Ea0Ke3iirSUTa+4LF5BveCZPqY2a9hD9zt6O1BrEURnRFsb/90XA8mAHvKimsNMc
zXigLHTMDAYlSTDmuiLdRco/9TkNROxj85oWjLnJR8XNZ6yhyc7wOvPHNfsKHRTu
CIXqdZYHBz5Lz2EU5BnyyK7LeL3Dp5GXLx9lRJ96dr3oa4EVwfSa/tgIuwCadlOL
zWK3bmahN+DtJUPq9yK+bigzMHxy90bpJe1Vs4nrTY9jClVgifpf2raxOYjOL7vF
AQMIKEzUNyNU8iB44v15kdOGk4jyIAiIC5ml+eyzVb8bffpofVIWrIqhZXbKVr/F
zMZge4A5QsshdSsUIoCJjq6gLCo/gVVi0hzG3kfwK+ekqiuPrWnZNMiMp+Jy33zR
KJ47uo2su8fV0OHsXzw44zrxp50urKQ3rYTbzwhUA6Q3xZy2n69LhOOHzqdkX16Y
bfJbydci3gIQni2QsWBekwZdx2MFDrqD6qq8wVEa5UyZlJwSk7dVGzbE41d/xYEA
aieCbKGsNeR9yq78AcLSBY5+S8uRnjWYGGVyumVnMF6wXMr+iA1/5CZbp5BpG1ld
JGlJwPfo9Larg0BnE04w5aOjIcduLX8PBDBXYeWZr8YTV+yO5o0S6LvdOXKPfmgS
H8ucRa1Oz6kNBaem7TF/d83rHOGq8zhC+mBGt/EnDw+89rJQbtJbiUtN6+i8bWSl
Ak1X/+kIhO20QC0xGJau/f0eZAZOf8CJoS88Y4iSElXPAeSWNPlQobBdePtjuC3w
AXKro3/jZ3XGPpqK3zlEZOXX/3VIFh7UpcFjT0WvjjIPWW3aaThUtHf2s98C4ajl
m/SWeB9yJ6E1IgfM2knZ9ZCVzbw2h/xv706AZmMnS+QxF+MIOBQTG1U8/rxM+ecC
QmYrdud6BqXws/AzYiDHKYm/+KRx2gfZlEnb1mzb/GMVmGTew+YKTSJKvO42aSJP
1bpVEuM6HROxLp5zE7Ltn8dUQcz6GjvG7NCqznufhL3Z84o9QZ5dGDI7NjZ7Nc7X
jAJuJC+BtYJHPJTfLhhSmx2k1kwwJU+dgb54iZvw5J+vyIf1ImHRdlYYDFsi4f7w
L+neo3mMms99DwmhLaRectjk0Lk1msTlc+RLNRjJOp2rGZNt7KvzmRJDVA1KB9V7
LHdlK48R8gqVRSno2hlmIuaZw0ZMsz16ZLu3dGlOOklkGFzAk7LG0de358iMfh2G
NuqZnloflTP52OfpPr0w6H7HkMIadi3Pb/Tl3CyqYDQPXVgFcTzJuGP0Y+EpARVh
XVHMUpljhi5LONBF0ODQmmHyvqOQffEn6lzPpfRLhgrd+whE0DpgPKCOvVzhMQAn
vGAk3q6DG2un1LQzcJM0tIpQLqCP8i/Cu7y/6cfO6FXtKfIAiMAxxa8gmG/yXW0U
31aC7yu9SzJaF5DTHVzYKWZgnLqmHrQ0c28Ajlu+GBDk4X98ej9wzsritCPO7aOY
wuscR3aeyr9CoPclJ1QZFbIqvuma8X1VFE9zTDwzfKwm/FUsKcFNYXx+LpNzdZs6
t3K3ENEiMJRYGFmN52eArig/R1EPZRQ4hHALw1OFYJyZ1d9XddTnMixSLvUV3iAv
9Wu9kdSSWieFVKgsKcM9QLS7viIUocHB77IHAXgGFOJUSwgm6RydJQL92euvOzb5
a79KCltnoiSxt+Aux1tb7HovhV3rFIsCWwMA5U4IonI9LnI9lG4kncuQXoXFw8sa
VPsyWtQl1ZfQt5jbpIsvrgQZ7wEznaPHNCq8R8eDVVVrroCLKc9HPG4K/WfX6jYe
okucU45pubQd1xA4K9lZfeNj6IoZHYQxzCazqYp+XwJY9JUa4zt+6X+RC3BbDPIt
U9Cws8eM7eB62qTaQgxj6a/jggqXpLRKa/+MG4B/VoPnZr6OfkLfIb0Fn2X5HNDw
6tYaAJHwKEky8gVR3/0VeDASd+3pxlMPbYijAOk+0Hu7KQZwxyCXMOIdpdrrs/W1
JaBV5i+ChMbFWpYRc6IFcHqplyzJURvfSQPDSPQ/Ptk8Ll+24uLe9RciBwQKf1o4
F5nDa/Q4Ms55U0z5/GZS9y7a0+LShwQoO0QIJVg8uuvpj3urIAh0QW6/+Hm63hU2
U6E/p/PQXAHYphXrCnsVM7ez1tlOL13JSqxv63JHHTknjJARwztV0BNumRjXceRQ
jg86yiv7pGOsbRMJGWxgu1t0Zk2Q9/BRxl68LaoculQYku2xiTvbZMCG7IXy0FQc
WAfcmcKV/HbS+FMDpxqko6PFJjleZ6mVsDKS1VNTBnGM/YYqF+ghbSar0KCEs4SG
TfZySOejzzaEj681/norB3GPkvBfDr6+8EUKAxct5K5JSAFJC5F65xTlcX8cIL0j
pCFmCeSrEWIdRz+MPt+Ez4J+bzePVjnip/VFnt5OfA+1zHl2XfMMm/CvIbiego5h
/HnP7kICPWyA5iWWhVmyw0TQ+7OWW2gy6NKOBvKtFcEtJbQn31BWVgqALcCGteQ4
P6P/TaxVqYyEM19zjr+kK2mMpgPwUC5edlPysF1yaDrJeyVgDtqU2LnoZfhvGJcE
tzNTT7xmfEieopTSdjnJ2Cy+aLYR6aBCnXbZgk21TzSoL8WY3p5RlsyxwoSrHotc
+lUDyp5fd8LGtEoNsb4W3A==

`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
YcSuXR863z5vZj84ZI2F5e7fFzJRkztX+ixojJ+m3bUQ3mxBIZk04GgVKLA7qgvLdVBX76gXBCLG
Sttm2IvRs6GiRna3VftuNURrA4UEkIWONmpg9lTc7wFzeKCrhehySwaO4PoU6WiiWQB/GIlaZ+vN
8rebFdL4rPBpq3IUNPyBne0MgjoCs+y4hqDVVJVO/fDs71QS8QmjwCUS2BDkmyetaiHTKCMJPR4m
XwXs66kCNmHnrxGm15X7NZa1fIbuCWCQZTiyBEGO9qqpFIl+pMJpK47b8rNmGYsxa6CK9NDRvaun
VTQMY5q1qDDWuloTASCS8OyoqIyrRYDpTsoeug==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 2080)
RULDgVd9tqjuHbQjlQH7NAuc1+Kfq0eYKDEhObpUOJInBlOhsdShvpYeRormi5Uc4uBUX7J2kfyJ
qsHr+Zn7vap7lUzlpiX3hvCOcIAV6/FGNDeemvLM2XCNslyZLPV+Y5JcfCi/dFn6J/Dg3bzyC1d2
YkVtGIe6gMUH+E5O668szzCPY2J/WuyE5ulPeGHPG0TUETRZtiW+SgRZsYY3Tx8EUjhxwGTQummc
thYQZXGRk+VlFrZlPt4a7ru/5QZaHXzpzPIonTlSma6hWgayw4uiwyTiUhqtzIUVBv+Kg/HUgymY
4ds2/mnGs+7Q+lQAvZPZmcAtxdt9XdC0nogCPfVCFQwBidspFXYzIu/9GZlAzGWOLBgM+RHPKlxa
MiChpsNBG/uvc+FDjII8E84XtPz+dvWXvYx5j54/dbic+Qwb7lvh5MqFml+xDr5qzUZQfFfPWi0E
wpj/XeN5llVomhXI3qAGlaN7Xo5VuiKOOQc3fFKQQbV9aEgSyCuWRsMUOv+To5XOjv5rRvnwR+Lv
Hg8G1M00kY3xyaCZ+bCf5+n9zqi4yjz8gC0pxJfh6m4DnumV2CwR1oAVBnpQBAu0MO9gRDpN/UfI
qPYyBBLZQi/SVphpsD5nzOjEsXpqJuMw3ommdRhBDPbvTTogBGsZ1OdsjxK3AwOR9pt1nvsESLSU
GtgeRsNEgLFbCaJz7WMsMveKYwPwHqeB8uCRqv+PQmpTgDv7EOCVasGcLm7h6Uf3gam9NA3SHBbm
KnIpTVJLv/oJCNq23BOP1qWtqbFJ56b8jTbN5+uCtxm3WrvqP7Cq/BKgv53Yl9C7qqHSnkMbQrNw
GJWW4NF5dSIVYTyJ5saGc/C3W0BkxuLFSuoyMwV9yukhj/KBeNx28OEvu698Pl76Eq/JW1foJCeg
DGIKYK2qX3BJzFsd8KTBF22sQWwnC2UF2O+ovmC0YQ7VEEsHtiYos6rWTaIUcN95y59uZ++SJJLi
IqKq8738bvJCba+H2tB0pC3ISUhU/DlrHnaZZHCNB7uVTQvscSp+uTXGoYUed9FsKDlWiGSEaZQx
wq46iARwwaE5N58PKsIDGS68XfkrWOxBs+mcfMXwWRr8arRgtBJ5YonB7/EbJvz4wm+Dg3y564J8
8SEm/hIe1zsfGGq1Wb/JNdqPRNW8kGiFjlyPoNwdCZqhnBepP0l2JItghtQwgEMVocagp1J/bWrE
facOAOiwpKY6leUkaN9q4xkt3YPF05mzMZoFNHOVafVSwK5022nyDhBhTVTZd+33htYZY3K/2d97
q6ZVfqp7sABFL90OYbEfzUF/UH2uZVzcFgtRQYYi3fCEkb2GnpoM5QYl17qimhqqQ9UvewyaWnNM
vPMrNjKBbTCsMf7mLQB4rbhumCAKsz6orj1DT76/gI2QzX9hHgMhWZltTd9h79v5eis8BdXNZodU
EO+4DbdReRR1aRfeIOqpDs30gMvOVYXcEKU0QyQrnFDs1dD+ymlmveVPhJ65elVi1rbfGuM/XYhv
ubA+jPyi5KtoiFufQMhShmh34WI8Y/gcVYVXnFf2YScPpoK8xQKAECYYYQRX/R9aCDaNAQv+tdlu
m8N0WShFufoqdD4EwudMIaE3YT7M1NY83KQld+cEIa5Zj1R8H1q128BAAeWbUgo1r0GsGk2KqDbS
141toTxUh1XNnsSpMsr5yYhHCTMD3nYNgMGKDBKMDKG8apY/EAzn3f3g4ImPb4uu6kpREEvS700l
FVgxvIL3jZx1bwcSYxzWYGDX8GofRyMVOc9nZM8mm9pDGJ2UEr4HxsypFRvHxq58y+8QBVQS+LmL
iQoNxQJtOePhXLaSYnjad9mjrNXEn7DZ9EL+WWm5rEkaetFnoCBJ9hTMDGTieIOBpmTchfRj2wqm
wvkopRZoKmPKFET13NYkC2/4lttxXJaOW8o7VQo82qg19XaNgUlam0XJ9Ay5iiTD+1Fjf9lid223
rT1uCP4mPqBR5SBS86USV5o8lmtKuigLFa9V/J6He+eDUjqKuPjIpMEcTXhbE8lxlSbSv5jf1nFZ
ZJ5yhScv6l/uRIsM4iswCADZ5UDDFM3Pg5J7yS9jon2VoLD8GYoLms1QyUq1FPpfthm8aKeAY1f0
Nn+Oxqm6y2WmcLMRISCr+xC0n3bQGNBcEHiTMh05rkon0AHYU4Dl2fIIormpnS9VYEDw8xe1jbAa
2S4AMBzjp9e3MQQ4DVLstjBO7rdknezADkdzh5b/TC233o3nMJLwFFAWOOTctMMAC5SVvKv18ooY
bPSQ5QMMVVNH6SAucykXdMy9QLblpMcntcnA9CLbJmmu6u7c1YpokSCQAU40mZjC3Jgk4E9zlYTQ
Rn6/wxp5ld1iwjo6nH3WNTld9V8/uG7UCz2nWkIUzxfBJiC3ksDFgSKOF9EnrOOyrAw1Hzwn/jQ3
KPMqUYucB2lMva83YkGPcy8igA8r5BqalbhtxWjw2t3E2krqUF5dQrpB+hdnMk7mgC8WJdt4rtYR
dEtDH5Nr15ijqlz91p98ByFq/r2O1cbsxrcHK6GzKF4iugq2cchtt3nJkh26g/LI0S/TSItlo6Fn
/0vP9byLGbxNMZgsIyIsJq6GSmzgIPeW5p1kWzj/7oWE4r3oMVtO8M6oTe0kRzdnZS0ilFLyxxeV
+/FdcgY9y/4j4IoLm91v1nz0A3DZ+DSjO1cNDEIFnC2cZMSNsN4eWTYwfnRONHag5aKXTGwVyhhr
JSs1d9H4S+KNfXmitRkjFNgBpmN91UJpb2rUcw==
`pragma protect end_protected

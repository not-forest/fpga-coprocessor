// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
M88c0rf3DC6pIQIvyAQ4UcTFmtZqUViVByP1MaAOaGp/H4iPiDkcmGzjgMVtG9lO
rlsExAjcxK90n0+FATTLNupF+GgqU49WAae4h6LmlkpmFM45DOmnsfbZfg6n9xGL
eqD8gBG5gVidOkcjJgQdlnprr1sBAOoabJQ+1l3mLvlvNgv6yX1Afpza/HNLcDan
Yf4HnXj/NgeA09kv2bGjtHwMw9kwk/zfQdDyibLjZ/C2aqrCBU+k4MeKSLnTjpid
2KRJMOitTMFvHFaaWz5LgF7LSHXzE/O8S2wvZqSFukHBXcPu55lRDrb5ldNUCYVs
MFuPivrVXus5KklLmnprFw==
//pragma protect end_key_block
//pragma protect digest_block
4npCh6uG5uhznsJuGTSB1PVlK0E=
//pragma protect end_digest_block
//pragma protect data_block
2ucj2vDNV976wbnk9KmDN5VI0BYb4efjNU7xjkyRQksy2yWvCU5YLh9b9qX0A3Pd
u9Y6TN8CuDaH3dXcT0PZvC6nqZ357kzdeGOBtbemb28gflHy9d/x8aI1VNsi5pvm
IJtTyIWYYiV0020X60RrQF+Aw3ACE5GjPnWGFZ5Dtk3slVuxzJmo90VcmLYcc/h3
Mb/S5gVR8KqrD8aFSbMcK+H7G9j7uyIybYSSJdLLatQDnam2kMb8/F3L+Vl2QCD1
cHKuBXwsxlXO8z5a6UHMIe5oAfqxS7iBvw7G60n781zym/4grmZioQUZ9FfoX8U5
ceDV9Uc2+71Nz4y6trZHu43mSDpOHLN5S3wiLmiRVtRvAcc+igiB7SkM/Wz3lnyf
BODSFEyijZR0qL0RAzYtV8bYv2py64EEzbqtxeX54XDGJTWUuk4k/YmcW+ks2JW9
Trp41Zn3P97JDMSpXu2zphuW+JY6H41GzKFOtpG8x6qtRWyLNPUM+wqEGKDFocjC
GGPBsGY0//E3Ef0riib0j9gIqSBlrmzFEV3ZhFJyW4GkDz6t+AN+/5zSYuiMPzpP
qBeMuQAQ98VBgv572FxZfoSgJKr/8iHZ+XDrjNCmXG44nu4NP4Qlwus8x67LYtu/
OWTVY5v7qP9jeMv39vHynm3apwWvs5LY0dQf/LCjpx+H4APRprLzN1q5dytqCWmW
51h6rJmv+RchijVhf7RyJRUCqD94UUWDGbC0puJWKX17KbBz4mgnoYkyX1fEndQt
hiM0XAceUCSQTGXXbF5oRzU+d3kyonmQJE9LvgUhpzWtA87zIdPnJOu3rjIsfvtX
rhsylTDstqytr4q/X5C97YxuU9MIrJ00BjiRe6OjwQzVKduIEpb3z5udq0Gl5QfX
eX9UA3VHHGQuV2xGS4w6VX8Bv23qxy/qqI6HM8vH/GNeOcLCx5hhWmIN2M9Vfjx3
RdO/bVk9SnQhugnV5rIscnAeSpwSJF67GT8J1rD8uRORM6RzAmiICP/qIolyM4tF
90632yO/QY17BK6HsM3gIvKSBsystChZyd4Sy58sJ/05jJXA6LvbxDTD0LzI2bv8
yQktlIyDoDgIOd1lHWA4RvAPpgfpV9aTDfd+EC7a3ApnLiAgSro6kA13hfw6trOv
iafE2feadz0OCEOBIoJ3eImZ49EhvkdH2W4kjbGIe/4vOcuQAUhwMAa4UMvH7jH7
7yj93g71FAImVAtJOckJ2mwKaI83zFxTzf11PElhGU4vMwI9Ie2o0PanyO7OH3Wu
CVz6cHW4aEeq9q682FqfX6ZjEFtf9bWDVBEToUfas3S7qtjfQ5WwFXQRokCYvUvL
6Y0cb5P7Zn5ZlIUd1ACDB/x/KM2RtBKNGI6RZKzr+jaFNwJ4r6vHFS0O+ArQFhaU
LNy54dhRhNfe6XMVI3F21Jv15NbVfjsVNxrMyoaUVY49bkX5eoCNNS4peLk3K9qc
j+WvG4OfNlfS90EOKOc+WPc7L9HAm8v/FMm/bKgnhzldeDL6KOvZhi+itIPE6XyX
v/tBVLKqPNrQLOG71prcWR1rwzmZGieohlyuvoT6NuoyX0g1qCSJ+1zeEPtHo/5h
5uQoWP/GCDPVCc3mWAqelbsPmu+U4sCQWabQpQiGCD2iQn7mJr2nOiYG6qkZchpH
n9jIGrLnImAzrU44Mu4TLckIOajBSsLp/FYLcxrvBDfRiVktBq4qWxm8BBVOMJsM
o7pue/OV9+E444FOfVOAqcKJkMyfzGsd+qY6fH9d8lXMu9D8PhJ/5PrEiE3Bv3VV
+VZRW66IpvtCPmSFbKqZwiZH467eUzHOXMyO47g/TG2BvtyPgnJk4/YAdOvFqPtu
GrhmFhWlz0fmfuUTdbTq2RFCPLgHOTezfk1WQ2PshFCVnC6Xh7n99BXtqHA9HmCT
i5QBm1gPw+/YoNGAqD6jd8rSx38cyONfOIuk5ArnRj/poqcOfGCVQm9PejL1ExYq
ZTRNrxTOeKzGqRxKMOm75Lirs1O7+EYjsyLDBPVzdYIXSYq+AO6xdWCCE53oLYcT
c1c+pqo8BgzjJVn5MBcnkdJT+vVxKudzfTwsb0CKqrW3nlm6Ky0ZRl01Ek3bcdla
ZkBwoHdT2i0lLbkLb1bc5R6XVnRViJFCZket64kZFy7krSVTZ3G9qGs+dajfxdYK
UHNruG788JdTttutpEh7fQ0GlzIN1wo0QVsBeOPUymEi6MtQZBVn0qnTnLeU29Qx
hQeIbGjjB5ogXiHovQW3zFdcDuzb2QFFzOaDKRqC83myAnBpdjzIYzptFHdLf8rI
sinhk2f+upJLR5XezXEPFS9ZiJ4VgsGYlmMt8l93YQJkpKVVoBv7CuvfPyq4Mvhp
Qfy31cTNwJ91aUP0T+eozDDF8H9trx9UXezF4lsxWcleYn4UE2dMStO9Vy09KYet
uXPWrQNnxSYTELzVVbqLUyGlwicFOUamob6WYMzpyESLvHEEvIuhkhvdF5D7R4F/
c9TcE3B0zhBixbrtBArQANjAEn77ZvMSeB8GeQT2mf9jt15qWjQBc1HGlD2Fq8Oy
8Q+YqfML3sE7JW2l1dq6N2t2OgqeankTpxpvG+HgT+k/PRjxTrUT3sSVc2FmGfjw
ZIXuW0EsE3bVGrtOWLkojD4DFSKD4tRNco6S1ytjjSAlkUYBEtNgl8Q2pLbWA3sG
92bzx0laE19PcZy8I38hedxZRiypkOh+8aoLMb0kBdlROEfYixW9q2tqZiPUyW63
RBZydMU3nb8dWLpBrcdFbFXQDRjj9rKMsw+fhtqAGR+wKXo92RT7VX15LcCFvqDo
6LVM/94yMC6MFd3bDBIZLtnyD/sqGvoa0DwPVBa/wEwUMTSNpE8i+LEiyp5anSpP
hl8M4vCKRx84rq+uQAkRfazn4bgl33aTQl1XRvG0d0bgYWL3ZmpJ5pnikere4Cd1
WIqcPJRwV+SsEb9wAPGoaisB9stMIHfXa/gr6nlEt0/SsQgSzlHgUS5nmwB33tLQ
E+0LBFrO03HnXYy1hJ1iIBgMEj7GGcjngRbmdUqJWiu43+dTDBKBIHlPnvwB4zVI
YEIYyouy2ePvEXLNw/l9C9zfC7/X2Ri9YWLhIJmKM4fMiFFXvefn5nWNwnGG9Q26
2zLpdxvVo5p1luTO+B5ltNIXw77KTLZlVLmkoyV6ndSX+qJF2JrctFbE6qiYuTZk
jLXdNCXAIEB3152BeNVyJBgMrJRVW72XDU6kAZCSYVHXylWV5WDuplHNVb3XoqL7
vus3bkP9LELg9piMZCnYNCt+bp3xLG6DDi3PoBJfrEpjwK9KMTTYMdeoVDR02J8g
j/wNNY42+pbJx4xYhQAUf0ZUerxAYN+LLPQ7IIwRyGpQqr6usdy0F7BiXZDZ5AYc
v9JcBr2oFH0LREqnKkoEDSaer9zwwhzFWKeKPO4s0JwRw5MfN2hmn4IxfYOOk2bp
MwuwFdysRAct3XzuzQSWpFIxdWpSsAo9A7P6ICmzdKt633wcFF3c3VJNd2bdjv38
rf0AkTkjebZts0i7XGTSmoGklBvjcYDux3u3j7Ncn8/Uvt/6zXQyvRsktr3vB8Tx
1wKl6DhXSqkNGqhQUxDzAZ0yGYx5VWOdY0AG/xb6bWJONZOrM8pwPe/C6UBrT1SO
0F42prXA/4QtemF1NTl1QQWYfV0fctnV1lZ/j8rvDu/YQOH9BCi6qN7oFBYcMrYY
guPdNMlmsCeZMYukOAWbXtRhSygiphWzTN1Bxj8lH250hfU/AoX8SSTPJtKsNaTq
2BeET0GifDTRIcz/79vgZtGoLMGM6yqrlr18ALvYgMi23t9+xsDet7+zZ0qfq7sv
1vv//bxGUKioSzGsDjQykRVdLel0C5efOYEmH1jGpCFvGuRsi/6ddREQx0Tmk9L6
hZbLMxaKPt2ONHiKLKfonch4VGSkCEvTamlLiAbRU1A3U1cr7QDFE8IBwA7KJ2Qw
zwjbrz6CWUn3ffbtLovUhG65h2XnqKBn6AVvkZUDRhkmJUcgOsTLoPtGorI+hV7p
EXwrjjPvaLCBdQ5++KHKW9UtkVBEJEdSguV/GqhoK62qLB/uiF+7iYDxHGjpC8yi
So3wAL363XWsttZCChMuJFpScMZ4amILy2c3RaD2W/241SVseerzglUSTnHiXblT
h6474IyiOYRX0DROIU7HWLfgL1P/nziGQOZlpQ1UMZmMEgY/w1HBjH/kh+08kZM4
RA8I4pWJBr8cdsMQLgv/CnJiUaV/G6zcO3ygF6LJaLbm/jrxdTdX4wdU7ykKw9/e
pS/PL6YOEhzhsDZVIYqC7DeXn9qVosR97N/c6McxdJfo3/B1aHOjnWblDvQSFh8X
+85fV6p8GUd81bBlQbhNHkUzqOO94nFCldjvobvFdsXKsM6Vp4JHHeTpZZ5pan3X
+xWItIEXS0ra81fPga6gAXcFt7LUHBlqJ2qSZz7JJDOmttLs7mqErx522vowWPak
875o7jiASyAdFIn6JrCD52y/uXg2YgWR+43lbNNjpePsMBa4BGnGWulZdMvh47RO
hdiKGDoqF/VGw0ZK3jvZ/CWgraeKKjA5lX2VhC0kdykiHdsKf0y2VYPvhh6xOv1w
FEyfq1lbnXEtIB7dxTnm3se2IJhN48QNmmaLK7VvmXY8fFV7gc/eOUMVZDz0wWh4
SaloXtizHUQtfvwW6wJD+S9KLCpMcoaFGt9xqxC9Cxuz2bxIrkVFaRrelfF7aaVx
qh+wNcCgrzrIb3LVOxKvH+ADM6cs/Op8Pc832D0vytO/8f67iKuIA+HqX9smmCVl
vXcmxAImhjXYotOz1LoAAz4tbciQHu8/H3oJhuONG1po7U2MERpIYBSmTpSEea0V
K0E1EVSEle9KSowlltccwSLAQ8YFtrq3yGCll9rvEFi47MEdEtD7W8FfvD+bED0m
mE6bC2etDLLUnDq6+ZPIIxRXsZxiM5o+SHVWD3ZHPh3CuUgyezTkQp0SeXsM6CwI
0zWwb3dtkQlHAi4l1WtylPZIWDVE13NyrDTNfRmBUM7mMhd7rt5XIQyT71dkv1Pn
HdqemzfGyf4b22IgshXXSpU1Q1FOMlNFYhR3LqJSQpHl/5jW6zI5Jd++sghsIZ+3
+Kgbs55Haq7gw8nD8K7Nm58zabmn4tI734daFBQarhZwwbSoG8eWfKFN0mFXR+sx
piPqZHmpnDFi64343P+AptfutzATCeCAfMQm8H18yryxqJQOG3cPjcGNJUcnLaWO
+c6DE+kJr/uwzf+y6SEVD0GOcpTAUzntt6n4jfv0PAxdOtoozugBwyOvdlOr4Rad
emq3g1mHKLIOxmfixtFOSHr5jdniklropJae+mEN/RLb5BsAqwx4LccS5aQ5Aj81
uaqNIV+LbmbMRxHdDawh7iJW4r1Um/PKexHzro30S/IaH0bfmn++/XGRTOSjqoKJ
j5ZCjHLHjWOKXnWvzam3RmaQmnjJQKFEINZ69hD8I03JIxiOOT0ljxGRmVmptTMJ
IdztUs8nRuS7auGy766SnL0AODng2xkr87yBjSkZb26veAAVbtTpDf/XTZMtnmrI
0jEVOjMlBVMcNT1peajWpJYE3JaCd1x+HZDUHOZ782kOyj6E6Jw/eVksQjc1gHbe
xjXNRKuC/BHkZGLm3qxfFUSMxE3fvR0VoCVFTzmE7tRyfJUTs7v5cbiSDl1Ase+h
YLN1WwPNN7HcDdU46QhKuZ3lt6S6YmyjMmHs0VgHQ1L33QvqO2CfZRtSGB7KpWx8
8cJ+yYDSYZN0T7GGufvPeQJm/Qzlh7LFXNDbZDYhgRgcC7zVvrG+kz5pQmk/9EkL
+tFg/v5/MvO3uR7UWfTFFBx+76bKbbxMoQbX1P8Um4Y7w0oQnlH2MoIjVFsKPwgM
ykc8ltFGrWBkZlUWYcbVgQQf8C5Jukzv92e9ENnzDtEw91J9X34NI26GADLqHmw5
k9ifWwgRxbjHCjnZ+kaMXOUuauS731UHzh+5HrjBuc8shayNFTujKpw1DbiaQwYD
+B7se14TuxjLzXvwP3pX1UkTXBY8HPaw5EmRufZ8qhsOR24/cTg6cA88WHUDmDox
pVqIyX3L923X0+AZO6MvoW+9KBVinagwId7rVlb7RBMCiutVvdiBz2AomnqoDp4v
hren8VwisAzeQMjuNq2+Bbi4dnrNY6Jp2B9fyGd0qzWddXrw7I8rEMt4Uo9r2CmA
fv8xGS3jlGz3xSdyp9bL9O38QeHNtquuyCGJWMbLabCsmCwbCMG6k3Dv753idgZI
/lIixDYGIBKslzfhrJb+P+f84mIkYXbDejYYIMi8OKnc+I97U+kyStCFKpt17IeI
uQvWfPXux2x5ctolb7WjBre1lrpmqmrcBapHzWZ5C8aFz5xlB6G68c8YSs3v8+DO
EMxSFrodz8Rk9CISBVVYBd3xe40vWR87owosUm7BDHy0ZhSrE8R/rdP0J3jtUDU8
XAywJ72BIDWAbsBJcqBzHkBJiRazKsRUsABQ4eZa4M+PkWdHVT8i0PcOzJBZ53W+
PeXL3PDB6R8Te192RoNrvM8zMHtZRA1antdHDyPK2tJjsdly34r67IrTeBB2P7x+
IiKJySg/84hP/nedTFd286D3jVGPy5GJ8YA97YWsPrK1axudGRQzKLHjh3mgq7OJ
DrVbLOZO/G+bpujcudu25sGwdXG04EuWMvXf/sarE+1wTOIh5oa78Qx4fW923JDy
gw8rTw8t5S6bPn3xlwoIRW3PLYapazkHWEt3lofuDE8c4+Aji5ab6BaG8oIDd7tX
dXk70G8c3lFBMZXh/1rNR3Yl40k3AGuXACcO1uwTLcRqlLGuf7iWRHNK08Ko0RsX
4l1+i5S8JvIcMnTbl0XJovO3071uAyg5aUd9QWHHdJB9tZoVtom8FdbufU2OqU+o
PI3tbth2uj4iGXT3szME1ywNQtOKv5fPBRFJbt2ZbNotMJPehE8TuEcACnY9VH0E
fQVtYV9tRfTFk9SC1xf4648kAk7baSCLc8J7bW6eXjyB5w9hST+jyjXRW6aCdH3z
X8ZPMzv+XQyETx6xAVpRiOS67zI9djoGBL0jvqchOxRxZNAyY6Bkry014tUsmD8F
PGFFlgnP2fKmNbeEZ9psAQ2hwLcYw5c6WXwFx5hb0kdtIUtGVJudEYn8Sija0RUy
ELhTs6KzenBFoQEFsUy30x6dquerncW8hUInHluLzfNnBQ2/o5T3VKRNhv71m0X+
nrVxaNTytj4rSe0IvCprbTnNWQWzi1BUZwV1dfRhgPQ7qX18h1SUtSeRKFtZ4QzP
89J4zvcaV80OA4w+gaQbt850r79FZvDrl6+K3lia7JP2HkSHbyOJRBH7iqx3yN/l
CzHLr1SWB6CYM14tPRedWZ9D8qZXYs8chJUznI6CG+3yvGQ5pim/Ht/EzPY55T+q
vo1hF7db4AlFgX0pxPwQGTCDR2/1orZ5HqpakNtvcoKHFHAyQpBmX9AVoZfdjYrX
omCHVSbceByE+VO+trTzCjLZIZBBSxecDSyluXsTtLw/CQLY7h5ovt3xgJHVnJj8
Mpy/q7/aWOnIsZCsTwy40wnod8fVA2oXoh+Qnwe7D8mdLUPPNjAOpy3Pfijja6Od
BRvVFYg6icAnyOSL8OUXHVVUSDOXSLTOzFH2QjdrXVeMw9lV+keBwOzdWBry+caQ
astlNK5CDt8oMt0eDGX+Stj1QynyqzKj8AMMp+CbBrkVsSl+MITpy95wAPaou91r
75InuDuCdNgEqGJbqLTmfUtBMuHBTPFEyb2pLt4yEm2kTUXz3r3qUDJKabY1MKFj
kR7V3QK8hl4fBoPJ4gdw1bPRC+z1K9uR92rQfkp3XwppLwuihqEQ5zSu6QXhk0HR
bnCwbalKL1UuijiPOxuOGYhx5PYwhTpcMcVierKAd+FDHqxEk/J5qDgb3umcC+gD
PdCeAQfLTq+wis4iQ5VYYdvRdeFxvueH5uoxkxwOiAAoEvh+LTzYhovRtdjb5RLe
np9CMe8tsCjf+VNxMc9AA5QEHm0gMB1taqS8JIQbzni1VV/C6h7skdI7qQdy6la8
gRjW9YQ3Vyx/YSgVa7GPWDy4NWG1Ene+xlrvo1nMUy9L2QyO73N74DFqGcxggxbi
M8SW5mSZ363FQVATWwb9hC0ZDXdqKOMbTxC8TNEiBvc78t2A0+DtDYML4RIZmK/+
aaHwyqETVsZc/rh8wV9WUuXYHk1ImcBh+KWxQTbP/24v2XdfRUPNSNw97Y2S4at8
uV1Ru97uy0xEq79K49gKG8bc/YmQGBOfDDoZJZkTrc1fAEV4Zyhewl3/xk2zkIwq
dGwjfdlwBFGgkVzzohfifzcFmxMyyfEQCU5gZJinMOc5ENgH1nHywxXwYtvEEhDF
7ngsyxvql8JegXVxFCNs6vC8KUpfQlbj9yXITqUXvJmOyCzZt7y7Bx8AjLVp2us/
eAYFBlTSVqI4hbZ9nKgsy2oPVe9dkKLoBq3rjVvQ7Qa6lAOGpd7sMPG6USwlz8On
MYYYVKpXgauT5Fx0wFu9wRjZjtLMrmKKjlN3fNsMH0b2Cz4dsgzfzvhz8Y0J4SM6
C2mIiQVQCUQ4axrIzSCAD5y2NeNCwz2Vk5N9mQKBvYc96omivPjd2v1DCsjyw7f0
iHLItOCdKvijAy+gQO6begyRCxLLF1CcVLT0WaEPs0eNhJJrlISW0MlAvFOpVRUD
J+GSzV+nqncUnXdPE7nSoWAYbB7ILoLQbb3psv1DgFU+e/3STH4Zdrkd4LXpucf0
+1ZbB8dHqAaRt45MKpNqtZ7g8LdEvYTXqI45Hv1N9r3q4eS4RaZmYF8yBET9E5UW
laqvwSebStwm935RxRKc3A==
//pragma protect end_data_block
//pragma protect digest_block
z9ZjwkzmUO5ANz1gt443DZhqUuE=
//pragma protect end_digest_block
//pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
S5uUalj1deuzxv62J1yNxR2s5PSOV58tYBqsLTnO8aQaBPAH7Nqo+fKlr0Ue+m9u
j1OGl2YYEarKWh0scuIGrSIExYYRMWd0EiTU0WcP5S5xLOSNz08DeVLZEBfbfE7k
jkbfwi/BKZd7qSN2Xd4O4WxTPuguWNpzgGu2Rgbbuws=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 22176)
a4VVeO9qTioN8vaxP/56LYlo9+F66gz4SH2RLJVgIpZ5BYX9qzLUY4LpaRYXURJ2
n5zEcEVx2pnlSSmAlgVdSsC0ypVPoZY/1IWkl21lbAPKN3PEfdEDcSismDh1iEih
oDgxUr1EYIpjwrAQg2Bsl1Qr8Rfnd6kvfqoYmIpshfWUh+eBso3aNjWQAIUzUTPY
8j+Pf0ni8j4s40XoAiq15R32SAqkQ4503icPxxvc2vkrMpDfdg1Hvt+NlCeXYM/w
9qv9wAYkfxNixnlY0rfclFC+ymuu9ufAitEKTXKY8ltM1GbmNJNmKVH+2rMK1Z06
+fqCNP/G8jgJpDlva7VsUj6j/KSFVwa377bvhXlRwBMV25DVrO2Qfy2n02D2Vdlt
aY35Hd8qc1dEPLxYjRlH2PL9JQNmOx5jbTNUAcI1jUx8rcY7FF3TY3HbZwMzOqwo
6yq5imF0FpiSihC9uZPXTnqMnkOd4SQIpDFvz3fu5zbT/dW8+4g6VF2lMOKIq1mv
tKxk0Idp8hmtaUuMAYzTO3YiR7szGZ865mfDZdt0tghrM736fSRw9TRkI2zVKKj+
fmQ1m348QG4TfsAqs5Y1rMt73NJEREHTkHtf99erNgKNCy4gntkVpVr50uhJ58do
h56V8cNqpnBxIo20SwlZ0V4DyyJ/Ockg5A3Hg3KERU/L4qO1dgwNcXyxhO2Pn+kK
bKohMhoJvXgdJipaOBdEGXt9dpyj7Z8dMcpuZ0z0GQjLoKueDG7iyGlL87UX/zn9
IupuiztgF3nuyjkxCjdY6Uem7ldzuj5vkIouc2wQMFaRFa6ha00AWvcJpEUz1aB/
LGwbKuhyNbjC0EtRJphYdgNVsvP2LRITXdVSkepNL/VnHmFr38YFmRYrHe4JosI0
zLHL39OBJbY0JtXhy/xfy6Waw9Jx1b1dtI8/XKnpWTrpRSOEj63z4hJNziwQ6eUN
T8qB2ZcUAek6OUTrktGaiXEOuiqTLNd3BIXhD/pFw0pvMtjcUkZw2QUPyp28Smon
kDIqiy7q/Bgi4gQ8f/7rp+0XLDlDnIeivVwnOxMGLTMcpS6u1xDknHvjv88hLkFy
Xs5+3SVz1NQazXwMerGPLBcE2F38B19VGBZctqwThS2HSrt+kBtfnwawanuRmGbf
3gviEdJCEJSj5BwRKmSGk/uxC2/RFlJ5txrG1d1Bc2Ftfh+UgOrrNpS3Fl/3FSAk
YwGMnU05C67ECXTp3a/IF29Ht0vwYzlQD3zmGaQzoWp6Z5wEKNJKrrxIzf2uHs0I
pdIT9DFs4WcQggVWoXlfAqgMmKePlSGHcTVEXOaZPg87ZAgrweD5tmqEuH13/2WV
v3FgrWRmYEObeT3oxhUfyFqntFDd0tBQpnUQhtNpM5azeD2sLzz20DTzkmAslJQ+
byB80Os5Yl7Icqjr8J2i9Z8XAY335sJJS7z2Snw5UnT+iNn43i+AQGq+jf/ubsgt
PtM93scyUgggIjDImqW086SJ5mVA7ixUMDNGUPMF3B6duINdC5zOvEvsu7iF++Wr
EiuECeJJjqc8buzwtqk1V/6imZKOmhe6CAPj6KCyEkiDG0zw7r8BKKMI5RIBYgQF
FS3rt8E4wdMGdUZPzWYTZL0eHkS3rwmIa3KCsImYs5rpa/h54TgTCl0zvIPe4PTb
lYEWCO6l/2nrCEcGcUlhvSkmpEWRWAO+s7PSq0ZtHQAavXqq/pdfNcK5C6C31U4Q
EXB1az7bMACkYhAW3jHvPNXZ7DLmCd0Hy49XyQJCzWxcCTQQgdZaPO73qlcZGK2r
3sLbLdsom3IPdMmi0gX/SUPi4htMT/S7146kXHUmnkRElvqS42c07TxXzqcBv2B9
fQaI5UenkvQ/8sNqgDu9nfjyvm1mtioqBtueoBihLqoxP1V4ZZQ+ro5tnVkofV89
Pn9d7mGU0v6ljgKopfLZHR0pB1ahx8ivbpa14Lyy6DKtjFX8M/BmuFbV/JQiXnc8
K+79QjISrNkLm0pvEhOMdVgRQhKcZFk9vzXC6ucXTOQHXvO7oj0QaU/zD2F+srRK
LL8TanDd96WOcDOhyAy4MsRJlQdgbj+NirZbu1tdlR43G4Sa5ZGDB0ICvW4Sk7XH
dUEWojY7u+fXmAIfXGnY/5fqE5ddQRhxJ5lCbEskdJR+rRFe4vVO2zKMWyFrVB7H
zH7JF1x1c8i/zXt8UXas6A46j5n1gvOsDu2OYsUQqhEciirfL0TWEscle3FKVrZ/
Z3u7RxtdkmvmQTEo4VfoWblcXlYPZSiwtVWxttXh+ljSuUEBDkMG/xTJFvc1M0fA
/YV61zEnwJv5hdqbVImyBrrBcAC+HcB4ghI/eeNdQIa4C9Rr8eY3U8dZAkj7/xU9
S2h+gZTOVqM+3m9LxqaZX+1cv0nJRO1iunXod9yBxvQMQCMsPEf/l/43asjZfRhc
wFWFGZ+6h6iwAmThsfghftak1HibRCvotIc5adp7UP2iMPGqiE94XVcX1omrkE/b
QxQSXrla8nDUcEHLcJmWW55USLLmUwQ7Kc61Uq691gLzFMUj81znnuo2hiZUGp98
83DqpgK1F+d+9/HtLLurcaJy/h0VoBe8XtLOLE1sOffkNiyM2e4mRX6Ts8Xoffrv
RUYGFsrdeTIJLYqft6Cv1XuIrwD+nbqUKgZzzEL/jfmTf4p7S0PmKg22Ej3fHEwy
Y1QileBeISeTyxOCWaUprpuaFHC6uDbpkMI3DUyiTY/2zZrvGLe3r092x3GA4CSu
adwLZnfNnM/5vEDZJhgqzpl/gLHrDvu1/mlcX44HX0yrqWrla/BCe4jxZUjhGdR3
BZP5GxZUv1nf8brxpWbnDVnOfRgRaTaSQQl4n7oLATvYCoAfaUR9UfyMl5cSEITY
hgWMY30BszeFWtjpC1JOnvuThGq1oR5tod3rFRFnSlyuyjw5kYkDoHm1HH+QPLv6
lc3OI68HWabYS6/Dm9ptADm1jlg10mAOZKSXQUsc23b7wXPjfysQSHEw7yj2fZnI
Hbz1u8qCFOwcvq8/cyC9psy66l6Cig4V+aF3V6WJ4RJIDXFAEvIlBnQeH+LJfuX4
WBO/3emekrg1LJmjePMOOqQIfIVGfGy0YkJQhyPMUGc/SACc+qJJHm+OwBw8ZEBX
hC+hiCgx2p7i2+ZZTBL72aLDIJYXNPVaLRmI0py3+YSIHM848r4K0B5q2zL6LW0w
0MaK91bmAJwF+jiHn8OUWU2BW4TDRg68nylq5XoVVZ8xDY7AISK+IaNYcR3KSPUe
iB6UTLArvN/AoqUyzgmPW+J84/IsFbQHxIiJbIm4fQgzYFpPQQr2U9RmdDvVAoHL
55zqGDraa4g08Tlj3CtQ99VsZNzo9INGGLnUuaunFsIue0vcVwbNa0Van0PpEJTu
ccBO5B8xrdAJujTYOX/fXrxFmrphK2aGll+PMn5w7aUWLYtQm5Z96uLXq3TOHC25
NuHraCDox0v7t7jQCW5VMUBFcuIlXoAulgoJQta3dQyv1fAIROi/iA/zu43JXBeG
0U5bJ7u4BL3CLTvS2ZzQe3d7sTcjB+8BXo15EYugdtHCKjn24JtXpKjddRO/sin7
YM/otWYHaVdFdfQZzeu01+rH/wCxZWKrHcS8TcxPK5L2Zt02AFO0QPLEJ4kIdQCz
Z9nW9c7mikDVnBiNLXG8aTlN5e43cmYKz7F1su71p6VPpAZMNcvSxJryrBTnVI5J
7MURMzJhcRUvma11KJCmlTplzpraDh+eOlnSnnI1/BLwtgaHLczK4mTI6vBBcDqX
HJoayAbIu320z8nlLMz1ZFe8EIRak92LmD5MiNpPzQ8Ifv9pTgKNryjvs/dCT70s
E2NNOXwzFJ6QIPu5+5aFLEhP3zNpxX2ByGH/p7WfGNPBIxRLEM76W6lL+vl+lvSe
mt0ozAJYO1xOPDBHIW6q5TCimBACqp5oNmi06wZ0DQzFglRVpr/LymMLN3XTWl/h
9Z/pDcqrAdgtVqpJRVJ1gApzkE8fQKjAhpmF5NHOqyEYZt8+5ur4nsWNGz1ytm51
ziKtaVqNXTi6gqdQLxHyoC7v+MChslJRj0EK+fGLW6AQKHMywvUihS2/B9/HpZNs
IXrZiDGLqXvIfjVz0aV0MSZGvgbQveXVyMFOAzmiFRaaKxpiHLwujIvqQPxjhBM6
PeY2/VWJ0vP7zdbmEJ/aPa/afw105PO8GBwYacphIFY1LrlriY8tkeyTcEwQXge+
+feMeu9Y17wjTI8jzBEG0jkAlcQ/FniRSLtIW3osEc4e5y5FEHubReeQih9+QDaS
5b9gOxQLYjuMC7llO7cX6WnRGbjuIaQaYyRE4q9+vD26Rvo9LtPtRO6kYYm17FaE
eclncOYVq6QyzYSy1ODZJaqUB5sLE8SYtXURvlw2QwJhSis1D7CmE+oJVeugd+jB
DoF8DAxwaiyjcFKz2QH+5blzTYH6eibzLUxgkMWZy3xC5sIDPJtUEMtdJQW4wpAx
t+0C5iiOxdApHkY/84QLqqrGsEpaAN0f6/8pxxtiB0VSu62ZmFVFvc+Bns7xVqVy
YtNsIRDQdYfBm7V7xZzjcRuwtnKOy6RrcbrgbBY9bot4YvAjUyWidZ58qKpkLh2W
QPjpmLmM+p0CFAvMrVEQkz0FoS9qQb1LXIkHjdbbjO+GpRD3zXUZAe6QinNN4YAG
zP9mJTM4aDo10aaQrgxtBfxZGLYizoxVsyLpzsASZ9tTM2FAebfHDs6wSFKGFXJ7
c8KR5AxVps77Y7k1cHo5eovKdSP+lh8QarXIieQTZxEbKXzus5ADKE7ddGJrIUWe
HcHgUOb5IqBXOw5RR0NaA9IppmBpcWoPfa1YW/bd9OJ3TW9MUn4Thpdqqw28EyGF
h7R2PDtRDDgSxfo4r2DfhGyVufP6Wmj3uH1mNqRrp7TIyqzY2eAuXQkIO7/1HuOf
rAAalD6jqlyaEPILrzodrP9Y33slE9+W4QJe3mbodBxgcc5ZE+LIi8A50KhtLDXY
KxH1e1gro9+gilPGjJLiqp9/65Hvso+OPidD829MVob3CaGjZzwc9NGs3Y7PO4LP
0Avn7PlKzDyeN9N7W8F38rXsqqFYzCDqQg/ZFIUs5bqx4lGEy+N0C4Bk86CGBBAR
5q1Wg7TU0RTd3CGNwr7FKF0OdgS+pIqNGJa5WRflPxqV25O+vBew9PYqyINHt8jP
vBqddxsiMDmvb1dVof8ii2/zcJ4Cwymk3wRgYyOGr8VMQzsraSr80JZ4ncTKq6y+
ytuOhFCnqr3szc9PsEJVLUo8Q6BcknL5YHFNQXNeblQZQqTfTOeciSNABB0C/Bxr
noOC7SkOQGr7qg6gEWSBebJCDocMwVNWAWFoTDejjH5gxuBIMjqVqAIct1JOWglQ
7n9e9bO8y1MvAB+/DrOv/sJgZynkE7O2b+G9RfAtY0qWByqvbgVLuxmQl4u6J1Ij
+7b9GDcdd4kXbQhQDQdbFaDiV3+WrHD50XegNlF852nwZEcyiHXnCu2zO2IIbm7z
Rfjg2oaxyYcBBhlhuvTX2uLrtn32vB4Ro/hc28yVOmulUpylUE/ZgQHkhIhI4D+B
NUoAmWl5/A2AMApqOXPBkNo9ObMGzJCoB23ydoOigdebdZMeX7BOwpAJcApt5EDl
IocpB0Z+EDa3ORL9AO2Fi38rTNOUd2WBNPT8PvneaSPUhyPRvfJURX3y0Gm38Tgp
+PEC4/S30j5ZSz/vCjX+QAjsgWDvMAbe628U63Z1coEJF2CkPMJ60t5+37pmzcLU
6fIozDOv1t9P2QKIAG8vocSy7cdMilTLUprD+jFq767oVPE0nBkKfkYEGyhTGL8S
xmeW75CpkdplVpHMNQiwQiG+J9aXDr2+roaPPztqZpXcgOW04FCcPM5yZ86WBeI4
5jtY3wPEwfQraccc6IdG6vGq+J2IfQgKnKQtsT9qTh/RCEuL8b/vvaephcIuhBNC
jsyYYQzpRB3Y7M2YuJiXXspkC1yZ3WFZG3kH/D7q7yWg+QlyIH2MPdhpJhEDGJFs
1cEr+TUjBCdtCZaH+oac9+Te1LfI9q0o/VKmdp4OSef/y8YzVlYTrLu9KGSOwug4
DMCdVNMB4ayb7+odQhnXZ7RlrnUucQNFxRCN00oZb+l1g2E7dnWJdXhcgI783yjG
e+M9ZUICVQVcOm2PLOGqjLnfnqYbzJw4H2LlGJ75Jqzu572NsxMgVWofLk3KLPkG
N/y4mkfPzwGks659jkMWqb4moZm5B7o+Xwd0fHlwkq2sX/OkG79YxZE+XZDptsVN
WNtod9kuZGDDOGBElZ8YC2AVcH2YAk0zZxE8jerrI/Y9tYYBPuDFPzK4knXXz1z8
8gqDZiXrVncEZGnE79BM8W4Z7s+/SiYdx0I94qE78JfeRR4sj5/Y8ElQjjPrHKbz
g2UGteizltT4tQPNmN9BgxZvhMWoyckvVDXYsUe4FZmrL8Y9aAxVJuuWwv+68awu
gNGWaSsHnRH1cATEwoO/cTdl0fHxR//Smr99XieXhBg8n0j3f40Tu81iPtus6JdF
mdbWQU6MJ0MOI+f4NFng0iTFEGPtsKNo+t1Tq6HcUrSpwjkfxy+dbazy0AXiVhoa
qe0m1awshUxdyVF34jFnrWEBZxqwtGeDAoxLTezaHdBbGrBtAnvQvp0O4dQIwCZs
P6RpT97dKZrVwjfsDnEEbIpMkv9IwgzmicCjvKgShur+/JnpVZC2WLVwMfvYll/i
yJLv4Y8LPU6Lx/XvStlrhXe/KQ4UoemvPO1OySUI4LU0bdrpSKZE2Ds75jKJ+TkL
ZvGV2O6fJUJcP9br6C+J2NuMsqsRbeUTsaqbJc7zH9gStsuxal57hfLXPMxwHhsT
+ff+hmtpsWN/LNSGnAgXnmAPukTBrYyuTdVGndrPzxFULkDuDtLhnKjsdt+IwCIa
tGiq1sN39msTCZAO/Yzb6GEn9rAOYbejGIhA96ve30zV3OitCMgf1Xv+WJJpAp60
aBAS8Bz6zAYYL7ywxIdz060HksD5mb/DATaoKyI5Tjp8jS+9Jt+oFI0/t6rPeiOF
2B489iRXziBt1i56aWVdF/PeV5pNcTdbgbAa/aq1phplgHHfparS9Wht/Y5GU/pX
xYXXTSivzTqsaSvz5JK6rM1DtYrxAlkKv16+OpAMUgqEsCB+644DdxlEBV5MHv8+
ZJmPlCzvoQSnezQMEc7ZkIBtBQIJvzANBX2DoU7BjevebkX8bXPjjTJuIL/UUnYN
1LGxEwAEWL3zp79/ylocoM3BNvElEjKF7DQBAmatWgD1c5eSokkWVoyW9AMYTiah
Lz+kZEZcRYc/FibOjUY1TKMmIKNFXePqNntseLCs2f1DGDBbhSlG9fANHIVkGVCs
dLW0yBABOssCKJ6rEHyJNQ4DBVhuOM5U9QpVBMbrkyWIpBIrcb0T9MDIv6Mutbj5
68tQs1cqeAP4vg5O1qx1oZVI5w/IhAjmLcqyM9ApgkP8cUAxgFYb0sDlNHAqkJpP
eeqmsugEhbuzDrvqpd4t80pVGkizu6VOLkEK/IQb1GC0VfzsXtjrcuoUfZjovg1w
v+48UQKGlywPjTQP4Wu54TAdG4FRkxM4uCrTOB6E+0vARZDVR4/6+RKgt5wlfcK9
JjB7stxaYVGFuXV/UmDG0SZLZ4ljGnBWQ/VZyN3o8ioL7XqLc9jJ/WaG/a8v2a60
Z6X6+MyZEIDCAPxj3Q9er9+Xbf3pEcHOMHN+ix7LueKVFFluBKWs2PzrFWvSv5r3
cnBLMpCEq5RIMxfW0JvbAfKP9va23hBHxSoVCFn5Mo2Ay8JfQ36TTO8k/QQNYZRR
SU/qF3YlI/gRkiHB9qevfkl6kV8y4oeBbTuIz1vzOUrP8ktPGiNmSzvfv7xSc+5D
xCpJf2slFLFM+0a6DhavECscWE5YqfEmSeVPcKEdxvRz6NrGIqL5gS++AQ/BQ1ee
5cIzSJNUZii/E7OXKsn8t4DcKbtPoE8C9Db7VEmRVGFQ7qngx0lyLe2/V6ixvO1Y
oT4vEDD68LC8t8TnaTr083oUCmbtzV3+wACarI1gGhTG8M2FjcSALlSUy/DgNUi9
JY0ZMv9d602TN61Y/mcDypFj4Ic7xDiOGEvhvF4whq6JmpQmHWpB3+tNykKmZGuM
z+mXk3zloG97Ak8nR5ZvgAvBDAi9hsDa1sxeSwO1rcsakFaaGGnHjDY5IXe0qWKr
i/mmiUJw1NPM2YI75BwhUe/mR6MUmJWj7nLuK84u8XvJPvDVsYI9BDh7tJ+akGSM
8D4bLQgY9zKHV3743iQNd7fm4gVhoIiLD23pnDXWqM0gxja33DHQa0djlr49Hi0l
RXgoQjx/kNY7oWQbgTkI7W5NElrSxTZVlq88twRm8+W0yvTeX7bNpkxodHw84H+X
Me0lDRcqBmJQCpdTEUBh2LC6aPk+oVqyPPDV+AEB6wQOg1ooN3k8/zlV3J+v2av+
DyeGHkdvK/ePqLSpQbM2A4dJLgytGSiZ83BInGNDr6/vF9Ux4XniKYO8BXNzUkAJ
RYW+o2c4FiE4Np3foNovejBoAvvEqWv1yF65JukZ6DFpTTzP0Cy/tpHsQycPVbp8
zYbrFULQh3SeRhdfyaok7DupjZmho28trvgAW5LiRcoZQquiZFlM0IzxbX3PIWrk
U3RUVvWc4mk9cXLEEtqvF6ROvosBiY5jx7XqGcgMxkjffH+UkrVpVPOypvSnAV9C
b6xvOyS7J7uU9qHww77jGGf1C2p06QonMBLn+RjHwHikZWbmeZQsbptFv18CQ2cC
n5wSYoEKVLQFlEQiGk+08bkfMrsuIe8T5hlNd4DU50SdD1c/LZPXk9R5yvO25UsD
2ivyTgiJ4UUnCKg64C49AJhIm2aKtg+bxJlVbkbhk4162oyZDVWoONfQBAZqliVQ
WlTQE3x2UUrqDyZzCtUr/m/YUBekVIlwamP39mRRrSNvvR4lZ+GVDWMudMT8MZbH
GHfTpOWXFBBOiNysxnHeutbq1JhRZgMRqVNf/GQE/MYdNdFsfExT2v2pOnF45UpE
TOtD7lsaP7v4j0ySF7Nq0iUDpx+qrLYuwmmm8rBeegs//c/pbxsSANUNeDJ4zGc1
DMMPhqgji9QlxpLOgUUdJreVUE1ylzJ8JKj3Sztxd/LcGUH4lsdwuFOcfLUXWzjC
hTtNhJEYggueJzpXTgze9mg4Z7RnnUCCuB6mXRlH3XwfamFDXvpHZRtfb5uSIxQj
7DwpOVUhNLR998Q8O8gV3LSmxRm0totVunccAYs5VLvK6QpqQ1UmmzxLtYcHAdvn
Sf4dx+tuCwBqVnCz1P0VP7ACRExubTOZRuUTFmT24Yn1x9WSKQWzP4u+lmj8d71K
93y/IYftEvjkpAy45BfKYGvNL9JRmkx0qcdg+PkDzbmCMFrMeel4q4NssMK2K8Ju
PKp9EwC/RCRSIlBuyb42dlCnsCMW39cHkO2flcN10iLFT2f3Qgr3w8r6EVA+HoUJ
Ni88nQImVKby9m9I84zinLAxBEqT7O9DG6NMA42R76F4d9yEbBbN7nuG0T6FDDtd
ujDSsu154afEOvarEa33dq+4zaFi5YSD1Osvlw2JAfL/O+sfiFad0AMFL/OD8P62
kwJnKNtgEKYiTGnK/G9CZLTQ3OoZy0DUCC27gMvDDbfdIJjp6gg5+uS4WetzL35G
B+IIM6Eh/gvck5DPIup+2VoiCnTBlHsf4oVe9cwHU+sf/7h/X1QKub0iFrCkkPss
tewcdOBlOltvB5cblTtPcPdGYhLrSctztmNi5FwIhIsBX0MzgU7KLlEsledjdy4r
PBDW66sO6a4XhHV/2kcgQqw2kXzlfcQtMX7dRq1yRn0rDYicQDXECK1l76Oewwcn
+aokyVubkR3X0UEFZ58uNhJhOAC21xT2Xn7y+2jTfSwmfLQCTG+eyf1F+5IikHt3
+1xMq79Csme2kOyhkvCt/z9O2vueHQiXSybuTj5vzG4gNTu7vqk+zz6ZFyDeh5Ps
ns1EYUn8rM1Clu7vxAtjr1kCmsJP/Muz7S2YImIplYYyMW+UxgvSbcKdhMlfAQ3k
2v3fhzgCtgV/G26jIoYzvNe1xKJBJMmGPXWYu5iz3+Wd4NHbDwV6dJOiIQQVmfp/
6ylutUdeVRtEPbS+t+8oQJG1joQqkH06Bnxq01MLzTSmGg8MGSMsEV0DHi4Q/688
YlL5tzCTn2vuOUl0oyILISC3k1dq5mRMWVgRU9+MH8inuBSg4zs7+YL+M4yxmXWw
RGnyb2ArIhNmcyCq/WBO7UEQoQDcNVMHswKTuUDal0HdT+u16LSLAriBQgoPfXbF
c4xK0ti9pTGlOVtgh6TtyTfL+OUdw95ZrTil4Nf+0Nzor01We7CfcjlIWcfY+f0X
ptaKy8Q6pzu22Y+7ZVlre3fwMm1Jf7Y3wX+8pAegrkXXpCamiH02KHOZY7eQLKI/
3ss2HKV9g4fuh9C+SsgeTgDcDnnULB/Ag22ItrPY/NueVDuisdGtkLgd3rIYy99f
HkigZzH98B/dx0SWcnwtaFy/Xu7aGteCUVS+6TaYO16XcAhoSrqs8pmXIA983HB9
mPgUewbmCulY4SlBnVkZ7IY03uIKcR/Z9Wz/3wjQzCS7wdHzUsVzNSJFGCX0XxPD
60WFxueoGl08WMkPycb7EucTzSMPXITWKW84lADYirzvy3/gQKol/IxdMTKKvpXm
nGQNxA41wBZft3RTJfAeGlor6i9sKneNe4+Sz3DoTvZm4sMtKJ2qjPbOmxP8b2Q1
9nmCE3yyMkP1Uf/CbzKYL3YZ3Fc8Hy6fHrUamCtUVjyiTo4AtbI/ew0KoN2vA66q
gIeIIVB1UK/l9yh3fzFgcwCt2OTwi72fThG8E3Ddnbx47MMOpwCsVxDLp0wRDatO
xtyZCc9Px0Hs88reE6ScM2xDqpziPOreQoshhY3yeIxnH05tHhWBa45+Fj8FhORW
ib3NWI48phkzdj7Uplj0PbShRcGt+1qPFmC3CzWh8sESQVuzr9QGQOGrQHX7xVZK
MkCmnnsKE8DPGGQAWYZiQWDaFlZrwDzIIvFJfj9KWKIl464jcAhCpdfe3UZTOMwg
yFEJmKDlu3yyobhNfIRfbr3oksm+L71hR9i1kirxC0EnO225PW19IAYtBUjrqT04
Eg6MUMD/BdemurTwfuL/HSLuL7xj72f3fIhdvmwrlWC4OdMWWfpRyvLW+Qbu7Pol
o5Bk/6ZsiHZqeKVbcZr4ZfVBtq4Ac7oZhraNXbuz8OgEjsEmbiINa5WoWc9ruaL3
mGl4Z6O81efdREw58Kfg7ZfTa/wiGYrbb4CQ9L/7DZYEiChFjLCGBVVrhjgXIuCy
xvIFkmFxXl9Z03bBja2CIj5CGblYgiXENEKJlvV8usRyhCla3IzUK0snJXIRGNZN
w/wtw7JMO5K1CqEw5Ma7oAHAZIwNfPhaJVQDtg3G11Lhv/mdYtTcwRoKuOHLl5Ir
ntvqA3cTya5Itq+9d+/LoyvYgYYHF/JtwlbSulpqcWNOkod6htH1RkgTsg9RAc0Y
Pz07G9A6hYq0mWrucWV0cJZQJIVmiPvj7lO3MbX8IIVy92LcPjio9PeXHsOK2cTw
E/1aCKdtylcHd1H/ZKEW0PD7geOTj/TzplqqoW/r5X4X8mwV4zgdZLEyRKaWA1Ax
fpwQU8JUVM09bgl5D2WE7hsjouFO0lhvGO2DtfPULt18EgMwbEqTdEI/TD002f0u
moH07jt7uNRISJb81KE+0x/MLEJdSPEPltakpJhvHysTCTD6n5ODoNOTqN2tblo1
xw7KVT2XNru7L2kSZ5lylAW61Kqo23P75lbld8BuPGfj8kPEBC9hBvWTDt3eNBqg
UIX9XYieT/GMpQdpQh22OaUfj/lvVsLm03FZrLNnRk7x1IFpky2NTOq4sjxVvl8C
oDlWd481G+NIdfPNcVr471dV+C+d5mlKsQRfx84i4/LhYwWnAh7zXfpJZdi2pCjy
XlY1h9XYQBnzyhuc1CF5P5KBaICj7MADO8EoKFAqR8ts9jqjBqY+sFMWiOOLzbNf
MwrILmWAtTz0EVy4HYE5k1n470HUD5+Gfd11W0Q4TobZTNslPxvYsBqMTrJJ6dAT
VwZN8J3qenHQIOFQV6LrrhHLPrxrUDW5WYKT1lSJeRTRdDGU6XL2ZX8lAatsVG4E
9WtO2Xzs5W7p8NCNGZCbOGe75BobTK6pIou6bPZyVmF7iUXal+qQhAXLHUsh8P8d
XPAfaj4CnuL+f8UOefmFVlrdzepPI2/h8k2TdMRdbf5byH3GkiCHJt1H3B8CFrIY
dQOI51yGHCNSKk8+x/FghBgMxoc1EfSxBTuBhvf312Rq1HoAz8U1BF4Nk9Nh95/b
bDImXXwuorDMj2K1fR3ho1tJ/1gLgSe7UmBDLHAHtra1NvXRv9N9FWV1KtQPcPuh
0uemJmllst+jjilU3NZx+Qwf/ZpnJSKO+qYQmcVDdsR3/GfBMu8QnvkuEy0DiLlP
+TZ2z9rsUpIVIVkv/MbrKQGkhz5WBq0Wty9UBEriOX/Q36iec0IF9H9yNrVkEo+s
kAAatdyUKu923hlYTekI7Pi+RihCd6ZrslPQ5NlmXV5vjvgXxhhkt0q/a1NmbbRv
AUnbuoWlz91qm/rcEaYVNdjlXZ/hMM9WYQjMw6K8oPjDbtFuSiSVWQ1+jGEInnZa
Eblh+Sm7zxZpuqMgD6468Vm22+il2MOjBwP+CucoPV9NFT2oj+2nk/MdQumruH1t
E8y1dA6WQOuNjVfwDKFhhDzpW8f2SK7Ys4z4LrtWxZrKwDuURwwDL9xQy1WDTGsy
Ewg25blnbDD1J3GK7298Pt/7i1SMW/AkTC9QFQMaxwHfAZG/ZEOJL6wCARzR1QY8
OkH5W+9gXMiK3XKdYZkTESm+eIJMx5w5JaH67P7dbnfQjmc2two2K1IVs9alsqEg
Nfp9yfuAm4/qh1Tlo7jvjuKVS3f4gqW0yjSLIeNMm8QiHTTNIf0Yh/iqhcyOVbVQ
RtNlMG8phxLBtAxckK+VErhNlYOS4d3TuoEf+NERMJfv/WwngHVFYQ9s9TwSo1zn
e3BC7dZS51w/16aXjkh7tOVwp79ZI3/5SJB5xTvJWISCAIdhVtu4aiYNv7HcmkDe
F6nnFfZQ5Ta33r92QGc0MslBJtuhWSMH0XMdVu4FrN78u7vp1L3q1KdEG1ON8Jpi
P6ni4xWnJrRjug8NcDSkggtSWa2bdVOHgglLoYZ7Bsx0DiOI7sBIBwKJzbAGv4jo
t9uGpprYpUSRtbjeVn8l/SCGlgU3JWiU/m6FAGVMEJBTMNXdIrgaeKhB270P6Rca
+ozdo09E00aZe2UZSzE9kN6CTK6lsRbNVnRlEJC2CWXHgs2IE2C8Ji6oouFx52L/
c3P7vpMGC2Sl0ZP0f7epQ+3X9P/PuJ/yrHJkVIiHUWjiJg8iMEJxfE+83nuGiB2p
tRSE2+FaCukBQ1tTbrjY45qOWj2JMQSuZutD39AA1GbQRVYY0hdzU0VdTK1OnOZW
1QDVLG8ExjGVbBtyec7op68uy6AX/Yo7drGlLr7WG7HbvMPJgTck7lHW1C3PT1z8
ga3ScQ3M29sPUZQHR2hNT1qUjeA8iLXXdLX57ytsCqXCTNuVWuRyBXyoE+ieOnHD
3Eizms2X6JJAjuw2uX4y9Aw91LDGoW+Xh5TCRSrx0psR5tTEuGne/9PEvkm8TwOO
N2KeeD8lz7c5XX5sAAGYALFQprB0m+8gAwUuJOQ8SXq2y8F1X6bIMVDrdnCl1gJn
6dAo078ltqpqRXd1tnDxG4ME2CAot3NZfaHkEm7JjgLbVtW0Iw56S2LOYXPdww+9
l729BNc0UtDLafFEtiFW0IWiK9rLMTj7sU1/BsizxU/mMV6Jb00xk5zuKica9ld+
70lvems9EdV5me0qAOw87vT6C700oqg9/J3/iQgoLEgqAi863RhO8MFuUIIQPuBm
Rf7W2AjXia0pvIG9KRx0BNShB3HLXVnCCoCZqpdMKJCQ2xDnBX6upqv45AdQ3S6y
yQrK59QGoL6n3yXIW9jhSJ/mQEoZtuHk2knehg2UtVwZoreftflZalpezyfAo3CF
SBVABi0nEqPSfbsM0n0XbdLa+kQgJvvzOBpWw1xhC29/K4o+vHBb+hgOf8VeCSzQ
0DfL3dGkaJhdAHxZuMFOLnEJCV2MeZf4VVbKN/cv834HIVWhB/RMJVeGLM4KW7mc
adCBCg2yg59JDLdrXw3tD3q9JbiRmGalNnH2fm6dGoSxEed1+bRh+voymwab8boq
J2eKOkeOnmpztAGe3MRxhdJUN3FGgf1vtahrmmm9UDVu0pzHvAPe8v0aGsqiqBj+
bo3ejzAy1b+bp7JG82o65buK4R1C4E2bVwZx13IZUEvoWoknrwbz67btN+GDN5+q
IX9luwl8ZPshMTWp/RwZsRmj/QK26WVe6J5jEKtJY4Duqa4wszQs8hc3CryfQ6KB
uSPYJH6WQdpj5bE4a71OnGu7pbRWiMRbuNDC1XF7s6o5861JLTQHHCANS4vJHrCT
T7xAgWNselz1Gn3Qz9HkGTN888k/3MJFMpHCjb2KTfbW9sOiOx7PinMXqj/+YTPC
eNjals//4LmVV0t7LgSgaUUT8jD4hUXt+lIfWxhtefdK7yIVj+63z/lT69pc2GjL
ef+jnplVRfsN+Zbpi46uNyHPzjQOZgfrtX1r0UOukgP/lZgUXh7sFwy6wPL8HXtO
KhvdGjIHjkuVmN9GRFzF8oTIlvLze5yjoOPcidKNrF5aL5O00JX1COWBrBtFhvoR
NBP0LO+0pR3JFZFo+SDeeNkiGk5gybsxb+gUnI+I8mMBcd7eJh72G46ZrSJ8Qeph
QdVc3x3FDzgk1P2Dktvedy6I0cvWd9GNjDWcUBs2sHLcrzZCQ0JkadiEZY82CctQ
f9zWH6dzqr+ivQQsTI9hA+I9VteXzyAmYLeJI8FIxxGuqnEgfSGW2G6zrIinmqcp
hmsvLXAetikqBeaEmGoz0PQOGNqLPMmFKPjt7+6W1YaQCqCjkPFu90EQEtoA1a+8
jI0JUAsh6fgIxE+JI7aJuOTNDoUOKw2HzlKyFYBEXF845G2RNzWoJjnSjmlRpwLr
hIP9hLyyktmYb+m+YpO3Y57tM4/7ZLKyMhckzLcs8q2lsJtkJQTbI/sz4gFYNpTO
A3+6psID+OiS/oSS6vnt1MrR/GGjNa7GTDF7mBh7irXUsq6ZtennkpbI0nSBA79O
ZLjo5S+vTacO5otsDAsysI7jqex7yZZHxLPBvH0niwNm8CO4U4/G9J5GlIOVOyfo
bdHV1k1orbpcmRGe3yirEgjkOfdSRIv2uXslaU4q+3V9es5QordW3Sh2x3+4YIz+
efQx6e1wP6+1l3oeZ7He7UUgEeUdBI2dG4RISZCzjREUj3Y7h/mqFK18/+gb9jNu
wJXlwjUmzpk5LoPrsIjnjnALQet119J2rt8/ZLO/1vc9GeVBsCel3HjcfPJOmFjc
dXZHJjHDfklhZrntInwpXk9t6iUXlHUz8XbpkSM2VPG8tLanWjpvkz66yDOQih40
k+9BM6aixEeGN0Y9LeYj/eUG5Y/fvUm9WKO8Q/cURvqCWq8E/d1QJNLL4J4yNii6
sZPs36YKgFBTZz62U1q9jtRLFavQ9RjFrRjykHsuXd0WR9RAJGjVpUrzyjOpyyEO
0+HunHINB6N9jqPAHJXR9i5jew8toqB8nH6czJFE44MGpEj8lrmAmOkEG5iZFzV/
9vL1eDzp7f3CJp83Km/yGkFn6xFCgY0qXeKh65djq+D2rUrZ65M2cyspdPst2xY1
fwjPxi53W+XsiQ1HbFqIbDFdTzKOXGjXDC1IZr9CKYKwpfjLiKRWU45GyPFRX6mf
maCc7GKKO/BeZKruYVq1Lqpn3Jgn7unvyK1MLas8mNhDQGOXn583wG9rKpHLuonF
26gkAU0wy+UogREvPKTlwmNNULJI0k1wUwGkzPjoJi0wL96X64ifyj9ewLxHQlun
dcrx+JbcrnrjUMrM5GCxP4NT9gl9cMOSPgNxZpEdjjYazJhf+Hls2GwS2zRGzBmn
xkQwVvND1bKYRrBH+fpjEiUMrbYM8m9pbMDY6NuYIv7FJJFpXIKFEctT6ERVOGWC
h+6BnA5FhTOa+WHOKRTR8vgwmr44bJ20wsvi0Qz7NodLtiK6hi7phknNNbhhGCJk
7lif3GTLE7+hw6ZMIO4YEwTF/8o/dVQkC+m5FbUwyci2roFwE+fe+EWtPU6JG/Ou
DLYNN4MJW/WiJEOvpL0yNNH62elGqJNY2GmKBYPQXg/Lul18QDipCfn6X8/7Tpbj
HN40uk9VYKiux8jFu9qJ/Ksvymdj56KNH4sEIVVbLtQbBL1eUjy0pCL/Z/qh867U
rCDgkX7SdF9WnJKL4HOAtQceczItaL57hox3FuwqoHRVyrfJ9Q+t1X2RH/FA0uWf
YVM1Z6vtTFhjE3czlyKISvGE4UsNO/83Xx36rbrPrbPhvX2KvpikmbYCZfDb4BID
9J9PnSDtkfCmjfO70rh7z8H1TkIYkUvmA7OTXSiv49MoodK/dR1XlMPFM11NPTFd
c6PsvUSiatHgQMC0hIsYsP3V4AXDA+fGo4LDOeiilJPbf27ppixIyCuabSidnn1v
q9ZFlR9hBHvS+1nSeJQr/t0YlDRbcpvEvsT93oMV8MMNi8KVi03fgxSfMT7+Cmqi
A2uxKpw0wX23DPObhOm6ixDcHWdnc8e9g1UqOd+2ui41ZJpx5i8AoYUBJfnB0dyv
SM0DWc7keEywIAfGNg2cWbZypNQdvzUKi4r3r8twHFNOZSagMuoln1jXOrhqd+fg
SNPaC1HEfHgM6SWxmFcIxM66UJvZ0+y225ER9z8hUJAwLDKr5I1dUSE5FPlNto2E
l0rQi6mYXm3856p/Ul2NqqHPWNVtYG6Go4H6Wo5juCEJjiuWwlHZlBrSxNsep8P9
rmfIDCFcBcaAHZl0/NvSUhhd4W7lS8rGxGr5SpUnK8yw/QaT2gXaOqbIuiCnK2Eu
uKxVN2u44Y6CQuHiXdN+miYndZ4MAQgis7PnZxyg7nM1VwyQV7F9SeFy8VYyt6CU
09qMCFqni0kXtpkBquGXjrA/0fDn4wlogNyCh4Pr/uEGMa4mLvagfx3X27Gk4SIL
Of+RwfMVRDPoRxko+Vk2WHwfea+jD1QjADiu5cScwvZ18HS/VfaePb+0Bc7ibVHn
4LFU1u6+ZmaFBWBW7fC1CnAEA/mA2MQpZ6eK1g1d6eOVStg3h4+jnKxaDbddxeDD
bahEngxA05+rxtxMwDzdO7i4Hruo0f1cQmAe0ElYr19SbHtd3ezapTjEifxbTBSe
pXxe45cKPq4yit0Rpoq3Jy1d4uSqadJa4T5MG131zYrGWM/wWuAWXVm0uwnnwkZs
nV612qzsllUhNi0ja3sentX4llmQK3TAu3ajz8kR8TMd4wIY6oo/1kaolTTx4pzn
bX44VJU7UuxWpCv79Sf/Ane3CFChl8V0CZRM1f/1+kSdUSJerbJF0ihLZAAY3V0t
WywzhDxsc972RtVohCva0MlXW+fQJz9AVbmw5v4ltmUlER8zmVZ9QVHyyZ4r+Y7Y
XtZIW7gSxy8yLs4OaZxC5eGDBVSC0j6En0K4bDJ4eQ8E8tLMSOVllz6HokZNv214
uT+7pwHQV0IyIQti60j3jbuiKbKtPD/j526pVBwF8j++PK4DGG5QKt54745ughBJ
cosvBWY5J7OhvZ7wiL0BvZZR0eIs8U7Z8g6NODvr/707L3p0bkH1AzHStUlxUrMo
jtSPUIBPGFLlD3E5bz4nURw6O6Yu9ph19i9tfHdA409sbPaETUNjsT5QDBKmy6+Z
IE+1iAv+iIrz/gjQl707HY35mNkGkVE40OeM9rgyIZ0dv0HtM4wmSkhja7w3r+SS
4++/nvwJQ+5luIqp+6Bb+vRgX5dqQR4tTqIbMXekyE2bNoxMMgfdocRhXE5LKzsh
wVdX7hzctb6TQcodQBv2mXdWv3vwByl7D3/M8bCAMkjVuCo0OLKWUYUoJgMDG7Al
9OsBbrt6MyhMLMDtoaa2QwN8vXRqfbAMtWAoIf8GktWknTgF0boZ8L9Y1hc/THT5
rodu1TFpnr/DXxWhtwXqPdGo865VVurQ1Q2V+6HH6vMP9Viyb4dp5u2bPpupoUrF
xW+nhqvrDixDyLFV8+jFcoqrspgJd7OYAswVRZtN9XPD+EGB7xOAfxLUC2C1+eNF
WqipLgvCIPl4fCauwxnrzDc0A1kF2MILGdpewXXT6jJ66LSbQzIoqDj4J6VkbG+H
j9OkgEdxiFEN9IAuTllbiFI9GLgcwDwZOEcU0A6+SiLWbl/9B38raoXFP/Jf57fm
g3FKt4GiaiYeNc3yJ6aBpkFmUFr8ZdNzU50g05Ys7V9KJerCp+3hFbK5PXiRyJOl
ci7MvnncSR0HD/WqFOyQqP60X2iul9Xgv74xwSz7E04apiB/qxp3u5lGbPrTQarW
UHbxakDu0IjcepREWVO/fyUO9znWZA8S2UAj9JgdMEvPOBrmkPChnt0A4P605pa5
fP7PnRXX7Hb4pvhFZwy1irtM+opitHZPdZqIYoFs5w68LAx7TUcbq9S7M9yMcyTt
FqHcOIPR337LVQ1lfZL+HVC0t2dGUVTiZ/8bnZffosy09K8ZrZvhl+JGtmy7e9K+
Fzy5A9L3BIAR+VfI4E7Q6o35bhKGVs9HX63bsb6TBTAhptGk3j+o4vgTVGCfLsCr
aK/m8OkLNo5q8yl1inPVzTnQkxN17tbhFkL1Rg3ey3VjM5UCb4Vtt6BYZvaxYNiw
dEHcE31BIcCXeF1ZqmjUosMA216BN55OICAmgytiv59FJQZvfV52kvXqT3E0G6GQ
TCM3CkdJ7WFn3+6+skM0QlsR5a7No4ASc4FF+waNeza7cNxIRy3adNIgNeYXiUr8
pV44x6xTsFyrioJFlxnAjZ6Mh8vlxMdIzCIvSek98mWaWBJadUtEWhcoH1KB82mf
ChqJyxa9O8ddqV2BQ2v3Rs+XL6zHyXoiIcGGZOnk7NvXIeJfnfjRtdYm85gueLTY
3sk26+/jrkPzlosva8ikLGCxhv01fzIrBQDCeyUdu2oks4tyZXkmxCQGYRGNkObj
Mkxg94FnqhSaU0qhGHjrFXLFu1pdfMEpx+B5TCeD93TGg+6UuWr5oMAkXIgPFLzC
wWtTpy/k9yu2Tc/PB6Oro0riaFxYLSpXInyWdEXLjLT9R7k8SRX82iKjvDTxGfNT
jvlTmN7Xezb5NLuCksuHbpiNHaHX0n8MwlW2M/QFvDzeh7hsiEgieP0QL8cph2j9
BM3Pj8pq4dCiCow20HrkxwYtAhCY1uFeYQuqqhFEYfiJKh64sjRhKxehmxCEhvQV
N8qmZH6nudHJJWVxyxrww6lXqBoRs8+V84YVihEnU1w8j1I1x9U/aNZq44r48PSV
e+lB+ldiyUjQvGgC1GtSFKdS/s4D37PQBDSH/sSuHcrETTNs+LYv+wdkDJEVBFUz
T2dkiN2Sho0uIR1ZJ+8mCp2c+Z1QduK6jWVpXyE4+jPeO2gyU3Z32JtNjQG9oD7q
9vy6fl6g1r/Xfgb368ptLv7b2mgVnLPFp0HnwKD2EuQ0uSPhl4LaiREpv0CTrcFt
meINXsaFFNVl70rAisd5iVeusAbZoBtkkJDag+DKz9+qd3+gJdd4c2mgxZQmdyN2
NL6mJrICti5ZxIJ7BTsI4MRu/GcYjrR2kUcf7YdhFcur53/58w7Tf+zLcxP0nq0W
wgtIaNfC2bpBXiWRnIWpMt4fu3QL8Ug5SVdHf7keQmFekpAszred3j9+lj4P6Gmc
ID/eKc7i58MPlnA+SpA7OufrxHGwNekl6Wdz4liePHsZP+2xfzYbkVdVz6UCyAOG
iNElkaap0gSsK3aufCuUGABzDFI2oRj4tmlAcocPhuPWcKBsWaX22UJsUehUkwsj
q0521GCbV16ka1llar2XfLQUOUu+G6jKXRXmFdDsAsn/QOrRIEI8U1RqvsdUgLUz
m9hgWUI5ir6dvRWw8GJJh61W0HEcWIk9MOmrNJwxc/T90qyLwgIH6HcpgVNUOl9Y
U0kks9Fp0X8UvI7hIbt/QZsNYmjqb0c0DK4j+fZbEdKavW0LkcruEpVk6eG+kthe
KEhaaWyzDnYnQX6h7cTERWZVw1rVSka5a1j5aY90agjBetK+e1JbZ7fK5omV+mdp
7kuSZ/gHVk3lcvwX4fLJDzY2PdvE+HGHh8PO26K/Bo6SLk0FzfAIswubrKRLBpws
NRhJiKRKYjiwR0OjmLMUGMhJmAQrtDOSYBB+Te8bhHK+7JGbYLIoaLs5UEtjlLNT
1gRT4DfGOf88vWGFc+Gw9Nb4Yfnwqszi8pQX/ne3uJ2dNTkmDizDYrHL+Tmfk7sr
WCM24MgNq1GugeBOCddYVFNjgTcxJqbANOQoV1vL2cA5BmwOBPLfW4Uf21nsZWgh
50RGyOEFTWvtaLgPNsR+4Hv8eu4r71iy/Cbw+5zIkYVSTLfCwGWj43ePsJDd8sBb
kJvQnRwoJbJWHb3tcZrBW32Q/hU8Fz4URjIHTbwhkeVkutt/txMam/WQ/AityKot
3G11mKkagz7slxTngcQTkubIYX5pwi/LNpT5L+A8yFNiCKDjHU/jI2mjrIBa/Hun
JC3CjsrnDlI/U+LFzaY7IJo9IsFGfAOsSLIEkpupaTRjvetp8iEPncHvJHxxcjAI
NQ2X0DuPQ0WzDwseeSVsl0KRGGIKlH3JFGNP1JL5Vk+EKMSIKJ6CR0Tr6dhrN33R
RJWuKbhjlvq2gPLnJ5IYSelorYJdpSNmZqGWQuoDIRcO9yC/PKuzzq39rPilwpjH
/XrRxkIrxB9S1Qr5wyMuOBmg5c2Z2Ua8pqqEgjuYBiVVPyVAVUKgL5wf9CRydK/M
BUh33yyBeRDh8jXNnhF4K7RuBSPnSzwBkuPXDw+38onrF2I7N4ykjOGi+yq+LCj3
/LyCC5crn5l/9V7vRvdXQ6+2tLKcxNqJDvXSs3AvyMd3c7fB1vKIHuWiBBW/doEA
gIAkmmApuL6WPTdOPaWuXXC0RUisDuqkLYMIpXcb9o5oBUGgZc2+cZ7xat/P5rhw
U0yC7bdPNJc0EeJXglBwZDHdciqio6ytCasSXB5Ae+s9U6LAWhDsOxi49+wTrB+X
yMxI4lh9gY2lIZ6F7VvrJM52vROiBLqX4SQ/eHG4ttvy5a9z3fLcc2GzwJLU7/oB
vs9uEIFIlX+Lc0GwyM06AScvYE3kvcJkqPhUcbwuNXKqSR1GKjaa0XA6P9wHNcbN
3FtG2SHSuZX7007PKbUuDmxVKH9IoLPAANDip/TX+xHGoubBVNj8ycy+w9YJ0Dnh
XG0ULK+sWwloRU1Nwywkokgbd1X32XG+JO6NelnZePA3vrCjdQcJxmqYm8yjEzPa
Xk6GEOVZYljRIyIqWuk2kfaKqU8oniWFE60pKLIX+LeagsFYJ8rgjON/8bIwIbTc
ovEjdhD+d3etrsU97X33XYZubLrOZ85AiqH9OqqZWl8b0QRTlpHo0QnxVTG+4K6b
9ls2DF6YROeJmkN12GR1KGr2gLlWfkeS7k7Dlzb3oHy7wwRA0KQaroNFZPrHZDia
GHw5P7tnUWvggIsxjC588Y53r9xfsGMTTUGBf8v3PBABMUBm06vayxPprCQccozB
D+cEZQHLOckSummxfNh7NPjkV+34ztHKrsnOO4bVrrblXnpZKe1HKq0rVKduRMVJ
UsezTV10AFdvm8mDgKbfHU9iZ5gLWH8zSu8+QtczsKIFyFBXx/JPSbKRBkD6dGu+
CW78m2a2gj9kqh3qq6Fz5KaxjPlunZcTqPGbOCU8eVsyZ5ijj8nudAC8xBzYh9ud
qmkg6DvMnKa8/18S3wRX0qn82u6vTIvPFozDV1U7VHSL3zsxggMS4yMnWXWzh1yw
Jb8VmW3UCiaUxc6D1rD+Pc6Ww1rpC6iD/YbRaiehiBjUdDA6aLgCBiYCeKd9uU9p
Aw6I6RezG3axiGYU9yeT2EGPsvC1FuK7MC/OXiz3REfHmxE5WoXNnetF5y7fRIRi
ruHzoyB+AjmsjvMf9NLBegTMTux8HObOHjUrkX8kYXKolu4XeeXihGGCJgFi5QSZ
RBg3F2hV1FzwDBZfvE9wm+29pZaTPe3wwn6Iw2ppjJnJQBNjWe4tJw/fKiUQZjAJ
iMt3tU3eiC2kCZhg5VkCUaCtr0ad+UMUhokJbXglrEbtew5Yz9FwuoId8i8CmB0X
lPo7NLc8rI8ajcD9Xc7YcnAO/QLI5TVMvfe3ItTFplI2yNt5xPiB/MkAunnMy/CG
/HHoU270ZKGv4T8Q18BB2BN6ee17yMYoMSFPzPwiEGtatchmtVoq0gaM0tUoA5VN
kg7qgZUGPqHeKIDJnjV90VWiSgjAtlnV1OwMpaH+Am7+GFY0lvK5hzwzZt8R0DhN
QP8ik81/X5S6YaKHsh3K0kTjqvdO+AIwoIWOuCylluFBVFRb3g9dH8X6VUgvj5WP
Vthiy++hWWrYuBBEpoxhrHSpc/frnJQHfkJl4c7wLtcA4+vJur92B/84sb0wceLL
QXMKOz2fnrfND6BirfWz4x8rK/hSEYTua0i7ok/WZflGW6xJJFY9xg9wve7OIMY+
ztG3doEVjy2df9rqGcl72sFXIVrFP9EgAYlrqqe1BxB/vGet7ZTENcuXCFWwaZA3
XDVaK9HwV9ZO0/Go3YuKOwcOnMQwxaFHiJjeI0O7v/5LRa/4a3DC1BCE6ADWPulN
6qiaUWpb1J+gg4zgzeWflnhs/OoKBWGgq9y79tMaS7ChFwLk7h5cElQ2Qj/KjB/g
dXwRYS2PneEx8Pu64JymTgKUJX6usgOSl7I4ZKp8kGS53BsIyP/aJkXgTDeuvMa/
MF0/bHt34BP4Z7dDBtpSfzCnvIehM/FvjYyh9vppiReWqoZdhDxd/NAyBlEzg1GD
XmHoTOg32okJGuLYBfR62A4BWKWUzxRbqki/q6OKmklH/mKJtNzAK9RBN+mj3vyH
0Jb38nbvx0/QX63tyNcO4tC9Ue126D3mEeU0VwKdr0OxtSeqpSV4C/+B0/Lctywl
64KLlxa+krVv59dA0xQOU8UiI4KGZv06OB3txGZNYIk2vScOtuaViJk/ju4eSIRx
o0PGyLLbW0R2CvXjfD46WLzgQ9ZFtt+j/cWjphXPeHcUTsHff2WGb/mXMM8r1bqu
ppOC4F1dxg95nIB+nxsP4zwV2XH8BkZuyiyLQg79AUxsE0mxZjsf7sdkETc35wM5
n2HsrEj3vDbAKC6CrKuj54TXRLfMmLiCrHYDr9VvFABxvcLtdUvbnMNk1LHSQoBW
p3PpkYZmQcWo9ikyUfuvyJhXvOAzdSQ+whG05ZCttkaYnwXQfkgmzDMgIbf1gSBp
a5TFVaACPGHNMXzAIUs27D0P+J9oz2M+lrn13g5ItOhs8u4yXVlsKaoiEtYmHDpo
Ze3nGjG/PUMi/1demNbFjVa9s0rAKa4GqXHApXenyZiG7qtlRgoa0nAUARNLQGd0
u2ZTbiNClYYk0rdqNvHjTxRTTb0uaOZ04+qtkqomDLHINQS/gfUWLRz2Z6HSRhEQ
QWP+g5ZHsCjLaVAT/28WL+NB5JJEcc2nLwVNYYI60LAtydglNoXIsDLbcIHqaEQj
p5kUHS4XeAqAz13QQ2UdrmGJ6mue5VH4nqMVpnJ3Q9M5VvjugyMOWgJg+clWb3dP
XKgqd/5vVeQAVaINF+K1IoJb+CKM7Oj0d9+3/YKAjgb1SUSF7RSWX1w0A2ZsiCMi
gd8XW/J0v2vshV/14ZUEdVEBKWpE4sRb1iU0XnUJ8sJsB4g12FL3SQfT9xqGOXdu
vLUGq8DWsclie61MQRO1oRth2KnODmIern91fvg9MpF02IcIgaooHbm7g7Lpgl2T
2ZlF58JbRrwarwVKB2PIKGnxPuWf12SRKv7ULAaMBuvcAUb7iP1sVPt0UEhG6p5v
ZMqLEY2ZuKM257LMmVhMBprzBmxCx5r110nhYV+QeMp+ekvE2yD3RBzadGOU3xR0
bRg11QyE56sSeJbEiYXM+CCDdz5yyyyRafscljIVJUDJt1QRMvkM/xN6xwrTZovW
ScUzFYwE8df1E+DyxaICwIkhm2vhi2bRx7vR1aaRo2sg5R/J4m6oCP1QUlvuf38Z
1thivwDQqTiMgJ27xkFqpKbA+c0CBxFZFohRf3xH4/WGZWY5shtm9kG1MBTk3gDk
yiRzd5abzNMtTgPJQ8UAVLf8gk91Q/PG0ERXLAUOgWKScivpOz1ScN4f7ocEmCwy
vGz/xxz6scTwY8OtOkjPPwqjbSPjRsLiwRQmkR2oNnBWGc+4CeMN1uUn3vK710IE
fZRSyY7/064oHixZjoSt4+WnVSPt7ZrORYs1xE1gjzlH4SBUnF9fh8ld2FcUTfBn
VO9koLkp9qjV1fTqM6rnakm4KrxXkmGQb9RE/hs+o5sDvKt/sBZt2JyGGVk2wFM/
u8j2pmGnJKEYT69yzP7yAOdXpZACRPz1rYNfmOx5SNKO5hJLK4ywJOIFsv71QAA8
bfnkpJZ6lPNaVr/rqkBYpLwRw1i75HKl23n1RO6Rx0QNH/P/hKf6yuF4Pmh7F9nt
0/g3LFPUR1kWC9wTVCtMU57z/3H0rz3n8ndkbNtocSWJHkbDpBL3aUEoZBnGXUT9
ZXFRvEtcgtMlC23uAJgmFBk//7vDYHOownAoDUdIhlQdZGsYCl422mLG4WgZgMwF
TvJ/IKHKoMlFgbxrJlQM5hMNfuQ7Zu5J+3QHi0K6g386hz/ftf8j7mlt/047mXQN
UVZmxg4Xzds/a4doOquzlyxILViXqugwD2JX5heC7PYUBOU1pLm2QNZfPhM5213R
MXc45Jijl8/Zxx0TEa3KXzc9qS0LggQ6icE4z0sb6byj4IKDq8kCqfBLvQef3ZEi
nh5b96vmyB9R+mycuuWiVIRzniXIxcRq15HsRUpaqB7K3BzLeMR5vPgV2BvvUqIS
qDlxrYTnoCUtSm80MOxFuE/xbmO8yRsb3HnoCJ8Mege9HcGKUX4uxzYPoUQSbO+K
oYHfBF9XNrTR5Q079AaeMD/yIePZnNwWFAQu+3NxYvlJBqeuPwQBacntf4mmjRDk
TTtZ5VEad4FzWkXwIBL1WmjxXmMumbA/H9gsu6TwmlJDic7BigkGU08YNkck8SdR
l7nhcjO7Ebf12DxX8BARbzMqVeabuSlUh/U3nJfiZ4s/93OtFBh+s2WjCynJfFTl
69fN9a4th3lUI1j58Dl3hLK8nfMLXq5t3cLw9GBpNHIW5lrGS+Rwv+a8G2jFYNOx
VSssZiZoyq1LpMofafrD9JyNIJ3tzZcH51jfqoZRIyJSQ3/danf/RzPvEfMELFTu
Go9W04MKL0TEAcmSetcoW7qOw90oJg1i8NgJeQsCnmbqy8adeeVxYNssJNgoQGiN
/puJiXaE4vd9iRRZLEfV0hrWjD8wFD0opfaNP5B1pCEXP0A7jaKULEcOOhyTO9T1
f92CmmjiXH4N2q4cxumUm9b/8kYCSZ0DbffXtTvWZhumYSk6OKePi3LGGGZizREH
ajhSC2xaAKxPh1vG7VbabxbQsxgTdE5NIlqS5vBsXFzlvawpigUUbFw7QMj6JDNl
8q/6QH+zCYgB+OBaiA6JdLaQ96jaBzfjWIkGPxgjAiQqv3mzaxu+EVaVaoVcjGKg
qLb9T7Q53hXsqDLvFwOnU/Ga5HXBFOfxfRReT+USmUHRCu4TQgqR0wUy205tD6El
+azc+qHXJk2oma6zmiHNAtNICPyLDpSFH+uhbjZISnV9Vo1JiQPdJHjRlCJrHJWW
iLSaq3DwdXQMm0NrX6NiA1BWsZhrgXTZtTE0eWpkRKk8LGMKgPvdl11QTlHdSOzF
B18juR5cJhrIy80AUbxCV5eDsquZarFQLlXaPTe6imggu99cA/6uqWrqGAdIXL5Y
8estwob/m1hLJcy54nyzPb8EGRljMjdreDg0SVTkbhGnsKvzNpG/453F+KlQbtOC
jpOb7iwqWU9mFzEacMGRIj8c5YumQ1ijIY29aRK8DTl9K98uUPsCfGZJXWjIl9dG
A+SGCnA8Jzosaqq8EsiBcBa6t/pIhSVOWAOdrNQZ3pQt8gL6lCkDziIqebxUOAt4
YWM+qS3NRRG7ydDCFjZf9HDdY01MTSg59gUI8SGzYvOp+P3ZYb/U5F9SijHIUJHH
vhsoBZlJvn5KkCYBtSZmSiy68JGQa8PuZkwps/NEU8Y9Gc9XPptb+GttDUgVDoO8
wIc3FJC5m3vJQn/XW4GWOfk3bGGiM5rM7UdTP3ZeHhbj9UE2BbcrFnGkW/xYSPGa
hpy4KtbncZsRk+PMpJqHlXQW+AuAyjAOvlsYmwXGJW8CUS8snqpVYVd0kRy+yTSj
JVB5+EuvydpbG9IR+rnNXzNSX6Iw4QE7aqxki6cVSIxF/dMvbJdn96rMPh5oQH4M
4Z3xXrtvgun7XVMljh0BhzPo9/tDeMslDH4IjkVC4Rvuw+9pQcxMMizS9AJOL+Rh
AxmeTG8uv8R0DJb4p6wbPOnpeqVJM3bHWV5GjvhfGUi5Fl5+xPOoFRTeEzIWzklf
OGVxo2ZqM+vyTCm3uYwT58TcAV+PUgbuU6gWG799qL6BD9vIa5Ut+NEb5ToFDWrX
IDc22HiUrCoUM0kYkXpb60hC9hJi1yJ4kn1fTFPlPgnkFx7zaAiXELSywwuQrmkr
j0S2MzVkVVQyfFbwqVG7hXfM+LQauHtqFh5jRcOVnhVINYYC2Psp/howE6QzHZap
RFaRpe91AEVl3KM30mVKnWkJ0OggsLva5ajEDlIBMdjub6if2JHkhQ6CgzOfv9VY
YMXXvBttqvh1MANi7jIU9HkwRmeQkv00z63uEmlaRd6UxzGtomwnof1PGLblERn/
JU/gsE0XtT7O0rJJqWrRGBo3p3GVCqCV52B55NVFPu9G/HaCOesB2mprDzLh90NZ
jksxlfUr5bLc/LwlU2yHGz4kByZDM8BV4jQ8UIO503gN/sA4b40Sb7+hJ+I8d0WB
f78wDkxFvyhFJXvtVKHRaY6TpMKXuwzoQCaTQze2PEVLarqJTjIkbPBgd+ys1TKk
uzuWZ0rMWdcBovdOPM0D1fwOHeHLxV6zuzZE3f+0gnRE042eCkLP0bDxJ5ySNTZV
93H7Wmv8cQgzEsGaOi+GYnoNBnfHng1oPgfRixwSss34YWJyDnD2+LEZEyJBEMqg
hyNnwXI/WoLXMVEzebUqqJ1DhH5+EiRv+xANn07GoTwmr0RmXW33/HIsglUCv9ig
KrjJQ1ApTLyJiHs0tOf3VmqHQ3Pz8p4MqeruR6Fx6p+qyM4zjY2bFqvlxRrWfHDK
c3fqqoP7BBQrVYxQVypybd31K5lyAGVIDQOb3Br7DKqwTb2Ij3HDUhaE+uic97hg
QsB+iv7rxb0HKqaMAqYaakOSM5XYXn9hbRAC3dywxa89Rjn0AvqgjlosMfMQ46lA
j3gyrpqzCFvpUyyxzovjaIOjHcqbS7TPyj4fkuGKBYJHw9Bql1HVZcbso/ASk4u1
noWBGtqHZ0Bs5wGAMUTyIH9t49k/5r6Enqyn9cz3TxuY6u3PA8yyxw8Btp1fbohW
JQ9yiqlL4BD1lYywogzcP2VKkU/cU9IYSY+Bi6hF0J6meP9chOdfVLtv1+XrMvJq
IfODzofQ2bxY4fU5MwpoXkmf9LpPFo6tJsefEt7M0uX/j3kkaZAGr0Ocu5Idzksf
YPFDjroC6lUlm67slbvEqGJrQWm+0eEAK44MAv0YU/h8loc3s3Tz/urEMKc1nwzq
joL/mS16BlZ/eA1WHArend3la29eU/oV1noXsjC22SBKqxyj+KEtVcXQ9qxeeUST
+wy4do5VmUSFD05Jm3UhY/outJFtgY2bsEjy8HyJsjTrOfvnb9PvdHS4LxrFp9xo
34fDO8VMwGiaU7MmDfICieWzXgiix4KTbUlKKypNLoETUN5Jzv6Sqw+Q2xidJbEP
4KwhX+/iWzmRhcUvZS617a37KJBt3vFabBvQnvlcaA00MtmnAjV5w8TDMkSQRW4z
vg7KNoZ/zpET+/LqrDY/oCrBhyN3EhqBQyBUbg77nSpkXp0RqWXZCrmItlpCLizx
7C4GbrJ1lC1Cy7D2DE8tM4bFxCecs+2rRV9QuAjq/WFQ2Y6cnUikcs8PNtMDop4v
ek30Xo0ipQYUl5TaXuwWq+7mAHTNoCRmjWjbRYGJ6Sdwa5XHyrfg3pSsmudu3g/g
zHToyaIZ60UDIrdONoD07YCzG/aZZ3PJg1sPp7EhZsdm5lSIFRy4teUae1hEihFX
awj6+pIEn8avdGGujEdK8DcyFa9l/pjy6NZFyZDYMhDuY+p/xCNS17JBSualKLvZ
o2EJHC5xQUNCTPgDmXtcsaUkpXsCsdffKfhm+iGnJA/lOCQObbE2Jec8rnW++2ex
eoKREm/VjF8q0COzgJWPCpGQELxjfhSs+gqBIZPVEpXd2Dos1fLb/zAibXzKFTfT
WxCHbpaZM5EGZA3AUwG7+QuPZMvb5OCVeeRQzXGV3dwwoEXMZSHc42Ls8AQrllma
093zOxThKsNEgdCNfimp4zniaQl/ydGYhnpnGLvTHTQwXDaUBT1HiAsuPw5dTBNn
lXQVPkQOOVqYgZBhKQFt9LPnAUZf9jnEg+CpeR2q00yVphBygOTHus09YxwLhog8
sNUld3mkHL0NGjOUNljPnmuqPc+aRRWJnW9mByICLdg64W9GsyRJas6eRyENwcje
wWw9nIMyslLL3N3didMyMMhLxHbP1mI4iJ0scgIlr6xETwui1WTGt/7B4MKID6Vh
QMupa0F2qcndLMBWTpuW8PIMhYfOhihdp62wmpDHjceLIhwPylCcZfc1erg4B4a3
+NBys1M32cCBuNa7liSz3aVsp0rKF1wxi5hWMxJ4gzziKTutVenGd8BulsXWnX0h
Jqq5AG6dsfolwmWLF8APDqOyEqHixcBCojmd+bQ/T0OqejJD7mIcZJanuWreOLqS
AgMKPzw7Mwm9nvqmFWr4Htf2xBKqjXDx0ZcP7H/QCxo7aUOu5HN8Eah83n1lDcRh
wNwQkYTbGX6gxvWFiBRHJyGAgxAJ3h6cQn+WyaQ7PrCCZ/0BuLifvFagq37fcC3H
77NytBTn5944sENCPT52ziRvuuf5zDCxaAo4nqjOFdpNWGcknDkZiOnITYpKKjm3
YtrEt6HHC0GN8/ZTODfBVF3hHqdRYf+mHfwKb/y+6iZWj5UnIed4VPJ8wv2tEVd4
me0ZSr9PEW9bqQ/2u+xRk5aStxIZdahZgdlcyyimByvaOwNOziwQ1FU5YpL69CfS
zvHe/Dy78MsrgSQU2rGOKfNS+ILJbBZDFXZBewdeiSutV+2KmMzsnSbQTBN9rMr7
10km5wyGMvYs7S5hJaJvb43DONHIU48kEkHctP7xvMCCNsikA0tp8lulCN9ZwEIU
0h9AlTHDEVzP2MOz2m4POlwbzO63MMkitZg9dQubLbFdgpl8178onVvPgFuiZfSm
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
icEZ+KjMmbpudWwNf4e31ktuOd+LP4urPRQ2ZheNMAzkFQtO7QedafvSYBGELlguUXrbwQLnboDb
vjpzxxKW6FZw3NBbJlrAvkeyeEiYUXKFBO+4USpa5+cDk2kBYzYtaJBEcyI8p045sVDiGPYlb821
6V6sxNYHVGnxbHD2kfqUs9Rdf/HJZMt+FkawgCBoQc/2KZENnoKkbeRN7tsdGDw9SSSRWlRHhy7e
56rhc7Rhskkat2iPfJRAFhcZY4OE3F6MZRE6fSfFbBXV9v3lCGz8Jeod/eHpONpZgGT1MNjcFYjB
lk1UbMBeBLdSXPHtDpaNriNc4OMKB6nwCSb8Qg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 6192)
zGHyrRbvLA+0T1A3jKmoCxgVwAqEKB1YJX7B8ecxk+bAVCgXTHHtpgVDKd91cPpoA/lzkov2tQNQ
1q+vJwPzdVh54WUschmL+6UNDudI5lHNAj6YrNLXuSFPF+heYjyGpYWDnRnXXxuY95UwEhzIC2GX
3V3T6ODJ6gNc+V7T9ghe/uNs+zOzUz9CMqRR4ncWGbfJX6MxnrKRAR6eHI/PVJFe3pndQKE4cD+G
foMguyibKTHNCzcGNyEXMHi9/Cz8hJAnfwxxGdidHh/vxBaZdeCRvWLnxLSDHrNoT+Krtmc4dAxi
1nY73vdNj5w9IwNRtqJLwoLpmakgjoB+meq4M38X2R94/w56c+ckMre2IEb7paThV/qtArrzI69N
5ibvXBa201ShfUrZbk5EGKbF73sN0N+7mSPija4SY1RZDS9dhT1P08FL/Vfdj/sSjegBV166fboi
MkEBPS6ticNTtndwu6CevYFtfqtCObcaUAEKt9mvh1wcCmB2eER6QyK0CEEH+H33r6QjPKzblUWT
2lbRxhQd32iqFkski5OmmPjxzOuQZmWco70b2bb74GrJOuvMzOZqa2UUNNzDywqe9xIFW6YrEty+
r/BtECpV+Urpp7dBlD7tQGn9zdgNxjxAwcFlDQGLwyAs5GtBftHyFEQrZAoqU8qb6aH0iUaZDYdJ
JWRuYjxwLT0fFKhwxUcEZrWMWbeiYULwOMT8JF+2AECrE55PLYti91Kr/EXGXkdoTsOs+fL17/sh
fL0KOoRi2+l+p/WLrWSnZn4Izr02+2NiLMdu2zhx4w8/nOGHTXwGzxsI+oJDujkpXRXPzGQX99Ht
rN76R4KF6E/M0vja/BVixRCF2PeqOHWU9OTu0sUlwaViNb1lRxBIIohGp3Sprb0YZtOwE4eRAejA
4U46n/h2GMhUMtzSZe+bq6MAOULecT0V+Q04pm1Zx5LDjhm04KPb0aH0ie1RK++hPB9C7MBgxGZb
C8hb+7F38IeKcwHl3enIArImfDnYEpUQkAXKcH/eiKk2zzTXF0KQFzzav+SFIqoBPebaLQ1TFrEi
S+WJNkBD6eK2lQ2wr+YiN3EJQaS4EeJMj5gT6AjXiezPy3wj2KoJbGWVkLP1R1f2IhOZCicPz4Tu
pjTZU2ajB2xPkCdrF/MxfvUN15XQLpHpO3SCBK7AUhTj8qD4eQy6rMiyV0epaV6GBbyBiYvDle59
A/+dbn/h89Nby5AOOdjhnW7JSTtkSQ15iaC64OkwvZW7p6bUSNWXXV9fu7B9I25XlUc8Psn6IGsB
bMpTeUX7QzrVlhXZjMfVKqledwWGE0IuhPHNe8vO8ahUqUMcymxeVy9eG72KW7+Ot22wZQmeQGbP
PH+ewEgs5fQDM8BTKi3uhDSsUpzCVmh+TsqDBDwGSLUWtviQ644HC4n7hdSds7AvJNwgClYNgNbO
BXm9Or1CDf7MRavhFMvJ/RHVrZL6G7ezYBI+Dzz3CE2Ul9mwfkidC9ONqR+myrRYwDddgqm9e2aX
Tr4Rd7wYWra8PpGu9o0jU0wgcgfQHqEINO20gB0lbhi67Zazn6BtqO+4eTB7Y2Pi9j6+hPThIrX5
fh+WNzSmbqY87Wv3GMB+Xe+y8ABNNZQ2kS4qCZCm4Cec6BXygQRX9NBjP25Y8clgbUBPiy2zFw3v
Iuk4rfs32pBQ945/zVdnVE85mwanCI4fte/jLFfKZoJyAG9jJZ1FM9NE47PJx/eOLQ1eOF0aJrpF
/f3EXnGYMvQhRqM3HUkLEknmpeddoCiA/hSNaBsVFZEbXGzEldSXnIYENHMSqRNboWwISO7lkp7w
wyF90zHlRwtXgogNKxE04u1ZR/aXbA+eOui5M7p5H2+NYVMvEFyBl7Zo/TrKdoi7YSYxO6WW6bKy
wezqmDB6jADEq6tj7aI/77ouDrq1QTc0qfpGAckZ5Sdlulaow+LqFswQAvnf1OVmDDRO0u0cDiec
Zzb3HVF6Bs1T2s5aVYXIdSN2RpFiRDqpWTYyRyQ5ywzpKL50gNAUEI46yACB6Bu9GACzJGJahHKz
WxAxyIRDGXc3C0AhU1w8s2zlyFd+GKmIOcDdbU8FHSEcpB20SC09f2kvA6IlQkv78O0yVNWAL5zg
02jf1GTtjkvwi6PaFMHabNimsdZzg/lPdbaZPgSEwNASWsMTgoQgsAUins3rDESpqhzYJdyCU/c9
kvoZCmiplKvFxNH1BfA7Hs5EOh+5Wqnky/8nl/n64TkZeODOdG5oCvmggHiL34pyWotEYnZb+LK2
Wm5pSx5hPZxf3TnN/vVwdHMaufYbba15fyfpBT9b4jR0jyNruroZGmEHNB6UULHwWvRzlgqfJs2j
uBLaFZQt+loYVIxc2R4EyY7kVKXXmFzAz0dZjy3OSFxckaw9vlt8SEulvc9PrVSIn3dgaqmId+fA
KdMvUPAitd9gkzOcJZMi9PoDOyVcINmZMg3RNnyj95D5GnDU1+pOqq9Ie1SFzeuKZ9GUO0fe0cSq
V4xk9hZhr3hmJJe+uYSyuskaA0Znx0lyY4TJTs6n5iUCOZNwQjAH7Taz/keNSGwhBZGtK1Wyz5Wf
QLu2VJdVwhdFePSjaBBqkJPJUCW45vtB4K2lI904762UZ9jt6Je4lLjq464V0MSokkpolmKi8p9L
URIbwhnRRPdL5bW1EOGnTigLEkGt2/t/l4CekBoODWBOBpanEql3SuEMV589JyUXWDBHMvs3bEOV
TnZYm7N6e87bcHSwtOjWZOAqJQlHXYXmgJ1fwgWpI1O4Dym6+zZPwe5x+OH4u0ROT56ut2gpwcKx
OumltELtP/B+qkMnUpHL8dA6zdQ5CY5YNv6eYbfVaoUUg+f80+SbjtyIAilMqbzaXdBic0Mo5W2t
vTd1GYEfE1tMIdgyNQlsnMyWiqeUQzFIQaR4TBldZOgCZSjCHKe3PI9a5rRXJsqvN1ZVH79iGui7
/DX/ehdosF02L6clxXPK25zIqff+4COWeKCU9AaaQQj3PLuQRLEMeOHcRRMGLrmoPX3vsztQdO79
cpV2QBrVk+uUMufF47IBMZwYCSycYdqsr6nZY2G54yakrwxAVxvM9DLYw49w4qq/gyaVTMLy7zmw
TxmIgnUJbwFsPaRqrqlhesPkWxSmbqiBsUB8GzQEqCzR6P1QBFCrkrobiV4HNLgAy9PYFvt4hSUa
Vs9iyS0G5riU5l/CWi/5jf6kr0K9227LKzTuA+b0NMlCOsJGQxAfCEpCPvT6bUMVHeDHutCxOLNQ
LJfgQNrKRcqfWNoKM9/WxR4ottiVJi4mXc/j8OWbaC9tCeWTTu1nLjXwlTekdtVgn6YdZ7MVKNQ5
YZAFF7O4TuV7LEGbB9SQFKojbqCtrpDLrBJGRe8KCQrsxstXrslt3FKHtA4P2OnP5k6rvW68hXjs
O/qJ4R6qyllhhLARDC+ZbnvpTmi8jpLpyEWrX5AmOA4PDjCM/9ENUivUiPVJRzShLXExj59m00ET
ra0zUOPkWJTgqFNXmqXQVU3A0UOy47VgRTCcDBgwKx4S7tfYaKipXr7Aji2a9AMY/YbX6oPcoWAy
c6sPyo9jR7Uvomyl7kDA90uRlj0t07OrkYwRyxICsvZT1p1IwOVLuzoxu6LalMQ07nOb/jyb7Y8u
c1jHM65qAozmqTWnYS/V4fO51sGjrnRFnC6Wyer7AWn/oJOS3Igh9RKjdVgqsEkOFhi0QkVYZq9i
0YlzQMWQaz1/01bghAGajD/h+KD0/7feKqQ/cnoYnxBn79ZNO7qNLGsnFTkrT2vHwb2BcVxUWYnk
tCN0v6a3BUShnyZmRX/OGXorvIbIoP71sRPASn5x9seGqpTgBvUlKEEGgdkqVy9ZDZdhu/CR8z1s
YGZKBJGsfYvaDiygTk8sUFc5fTxSfmiM9sVAdPk7SrWmfDOCUAU4hT7Rup+qMQ7N1Ocq42ahZJIr
PtTJG0Md1URoL8yXPYpI8mppBNRofOQbe+M5xwwRrZO4UGjbXiSxVaiC8bpgXsqM1QJ52RDV2GTJ
OmUUEuIWICddyk1cdlN8XPJRX5Xa9OGPdDKkXGW7VEZXz34HXquVeN8V08cL9sk92no52QNg1C77
UdPb7NP+j5QO0e5tEpSl5lca4NhzQIrg9GibdwMj40901CR1rT2QANPd3UR8YRDwFt5YGV1VXdG6
dLz9og8qi5u/00aoQM2ny5aLtywASNhsJemXifx8J89hgchaN0pHc+dQXsqJxnTPlRgLMULz5R7U
sDVp5qCFtyrOoht1pNWd8D4Opctm7x2SXNjaq+vvuP3brkv2C9GaCn5gND0aWZlbbF8PS5ZeNHym
Hzcf0WHYRjLv3KDQiADMe7Mkq7IEb30kfwCNZuUIFKs4iM4SMeW2knn4DyTWQs+gjaqGotZ/vJu6
Rs9vQVHNnVx+Nifv1iPNC95JOUl9BU7iEBrA0kNdWK2C0zk/INWrSKQmMOgm3BiB+w+c0yVpCdga
3kl0TzfXitUDU6mjSa+A3tCUwRCFX5dtDbD1YDuSQoZfRE3tvgXf3BX+1ImoR4v+bpOPr5Ur4Y5A
BKPZnDrNLqeUM0PpBHKfscREWANPqxFwVZdT9/BzWcLLB16Bb0mA1M7YAtPCcVh+JoJZ4LnwLPmA
xgspIRnfkRssw9E9yPC1Mi6MXU3VoGR0269cfuZGYtdZKV+IxH88r/TsnLJE6QUv3xft+CLHYZgY
98rQCjPN0C+seJbFfwv5KniIRXHFeVY1z7+VemPtNsmKeltKL/xcF90lWvQCIY9txKHFfKN2Cpgw
7sGRpBdrhpsTS6cwltcAvNt9Dq6JDSaTdC+TeGkcRIrjtzEu/s29uNz/KnCunzZwBuoXxO+umbcT
rsICuIRA3grtZ06on4SlERDUqmeR+mw5Nx1JT73QbsYc43sxZcCZ4+BoscidrJ2eEirB036QbN2u
32wxRpGXZNDdC0rQb01/aghgQzq3kfu33W2b8IP3lfJpnqTIM+wvEhP+2VitYKpzbXfXvlO3Eq6W
54riJzb1PPovNvD8RRNSIyKoSniWr2GHu8k3OVginYvG7sAvSmAGEDaCE+J2yz1rXPL4knSYWE0O
CpLNJ/ArEuYmc+IVAe34FjV5m5w5LDRaTlqw5DrzVvx/0Xn5X1GddiPEFAGuKvcQoUj2ybqfpT+p
3xz8qAT2pBBTHfombEgMsrG2iwrbNxxhHDpX6aXLgAohQrGviS4ECmilMLzL7eq3QdWjpTRXTIS4
eRp50ArCv5OPWE9cl0Z9eaIHjzJbzmBsrUBJH46SYcOEdcCYO5unWFW/8b5EaZ2u/Mtb1o+lURzi
F5mpOq8GNjLYrMfilbC6JI2uslil6eUrZRy3aat0WgBZq6gWxm4vlvSua8jnCH+IO7oi896bGgA+
E+ya6PuLEYZusb/XuQMO2doGqJjHhCNAgEdl1gT0Sg3fCTitxDB5hAlJK+SYeGvrcr/wNBDYXhod
Rkv07SoBXGmyVHtMMTDHvM3zACROUCJ6pBKMPdzL9o3xXnz3F5PC3G1YJctiu3KsfzdaSLPjCOn/
00q4tvymDaus+u1VPq6HnwLkLG6Lb82o3UZkB0wkP+UUP1JPv1HMGvXMDAQ0nGSd0FrmVbl9+9nd
78HUI3U3mVmhLOyDiinK6zaebdYIq/QTG+hM8GJn12rlFY8/JH+v5PCnAwQ+EUNy1ig86AemTowb
rNAmZFlK93fWftlvZZhKMLH9zD22xS5gRgG9G+EGvWxwr3w/iO3JiFX/fx/l69BMCK9Sz6hEms5b
zPA7TXwbZxLlHMBXiDqvimhg3+aoRt53xZRb/w3li5/lW4cbi+07trsila2Wab4lwxCLhlP3T0EL
NePaB7kuQ0vFV3PMQC8fkdCMcCYlczSQjEgbN0GCefKhVXlptR2NJlYnoc53kkKsTUmfoJm97245
ocYQuGD9qqPgJuN8lKHvABmlRw1c1qjsssWwWWbHUePCP++7yMAIbG+Frfthmk0CZYOy0cMYx/PP
O7+xBuuqFlovIuYN3v4nJj9A9csRX4asFTKtsyv6o1ldi0+gUeHIb7YCt7Zoa+r2fhmQUtopDLEa
ZvmC7qzQ3iumHng1/RJQ+m+DDFvMEZzRuLfMwL+9cBe0p1aDX5c7PQxW1gwycwD16wtVmh/jbvZP
ZaPr20IMeqsLxhzhtDrjxANaqZ04crqL4tWPkpHvdyeB5cQ4gnRrFr5Li8Auh6bVJXRJq51z6Gl5
+die7vsMRDIviJBPZTWhu36Ale6xMyvTRWT6cDp2tW19gAG0JbyR/Etx9OWX2fRmopJMA8beizsP
yeZKgk9jjVxUyH1AICn9n++0nKsWz2wPVW6ROnAdjn1mqFH/pGadR5Qn/QqoIqsCslxrWO3Rqa79
CzPmFVffk8NidZ3guL32XiBLkreD71NT9+C8XtjI5B52WogC6wTRyefkUl9Jvq9WVt3nzrzVay+7
e9ndaINqlCmEusnf7j9wW25RDTAcKXDyEpjYt683/tANpfL1ED6r7ELc52h8VuCH7bp7NIUMa8/r
nHadeYQvCx7xjx93Ws15VbqxZSeVpV318tgphazAXlPBg6uQMJme+kMmn/sWAdQWdxR1OzMr1e3w
vJUmbSI872DL+QXXs80TgmD6yVAemf3U9fA2SkFzmkeJDkmxmipBNX6eZ66ancX5B4dAraK6Iji8
2oKZzohQ4crfaVRUiszgJFZraQLSrUh8yNoU7yzp/oYwyBmNBVzRNn5+s2Xs6ySUHd6CWM7sWAK5
+SZdJUTBR8Gyranluo5yfzHzOjVZrBh7qAn+8AmXH906wtLEQTYxiUjcB/3Yl47hQeed/AUvWPZn
qPE5Pfg4Je8b2ChlL81p2Uc6la/hp2KY3MtIwzIaJz3084QeJKd3gb1twHIcUwu7MK9RW0PVtOUy
l+7pcbt6ce7JBpP2gGJKanxWIMHyaX1cKXBtdlt/Jl+V/idTxnqypp1DNQ5RHvTUa8GWVPJcutIi
PdXFvq/FXmi6CRC8jzuO9m6t0W578i2pE3C4pgRLLKo05hiMTkk2crIbNQa3r2kbvRbutdGE5exW
2aF8Llb8Qc2Yg4BBinr5nhNAJwnAwWnSbFg8XqCMfLMj7oVcw9Zj134KRMwkQzGBXXPPwGgDpj84
P4xuj9UxqsNLsz2JEIhllPUML1OwKAP6mjzpMJw61ZE88lEN+2fW3WOEKV9fKR9dPfE55PHQgh2a
7d9OWCo+NTopjW1pPyAsy9n2i/xYEvteVV7z1CXRn26g37Ab6corYzvunLqGCOfsJUKXAhkjiL+Q
T+DCIbhL0aTkiLAt3xsUwodW+Xef8bj9atBrbUqdDJyq60eZOlS/K/UdOXDPAT3bkUSBKJa9jGFq
zmWMIcaxSqUZqwlNjWxXYn8T2OBUhPDcpa6b6XldOGmr8EijIlH+t0FvS9ZrQkMMlT4P94o16ygo
ndpVgZY1JVl1IilXf7VHflRBqrJvvmVPIYHB6jIVuRl1vGaMkgLLnmwB66rIeD3zyYQGudbXpujd
z1OeCeyZDqdO+qrJVqVc/Wn9KVU6rbTuhe0uBHhJsVqQj+PJ8sD+ZNZhLuKdN+Q/43+Kgy6qytP6
/FXLgMViuRxejIxLSButxcuZ/sjftrE8g96wFMn9LXFtnND0IMGh6c7q7B7kKU+Qee44c608h7q5
wVCJwQd2mlphzbYS4zcUQQ/meZ8EThIGv2KHjzHgfCr2y+mRcsKb7padEh4NJOK/RXWQJPPMTRyi
NzSu0CebQzrLF0V1iK9MYeZd4SWcEJDLQY81g3J9SquGylVyPSmdlKB/tLIKaod/O0InnghfrAJ6
tI8cEeq79WqcfVYy73ivInyhKvK36/BATtCLdxmPADVtUp9u233see49VTA4f0cjKJu9GikY461a
w7Vyj6rrhUCXMls0GlRYvo710mRdV+dWNm6nOVWRY93l1UQ0/oLCWroYFKb0kDEw0YzdEU5rbUBF
vDka2MJ8YLjEoaKce+7Vl3ZYbRZi474UuxPaW14ofmrR+Z59NaZSC+jjgviScisF+WCJnDOKO+VT
OliUdl7Q9uLN9QDpzGE45+UgsgxiHb/rgWLvr+l76tCDr2Os1Px4f1+TJhonYzhmUK1KNTFQu19q
EhXutUZkU5PCPFr45WhAGI5VMrqjJRTq8UgyikdRt7vK72VtyWSZvd9pfdvD9lBGpwUWo0qz6rsB
FPfqBNTxb5xz17SaLlY+TUEO3/IrJFkMRHTd+/HDivVd+cS8
`pragma protect end_protected

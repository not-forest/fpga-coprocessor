// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
rvoCTEwkS59VAPSDRuVm0PhB6kZ0sd2798dyfOmd5H3cmTggR1wYiTmEJiprv8GT
V0d7gDbiZO17/k8SFJxQjTFSuzoeTxZfhkLdmLDw2DlKcZx4c5YRtCBeW110zWQ3
NgydpgDkgQjdeeiEFD89r0eEO2D/FUkzi3C5MM6fm7w=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 10864 )
`pragma protect data_block
FyIhaW+ZxNKNU7vjHnV/geoN3gNW6ESIBwq6wgyiAnthFbyjPOf4Z6YiFbOlj+IQ
QtSjNpNcGee9I50Z9wr1GSco5ohoXQG60/OPwCcmWw7/zwqOa18+4sHC0saxfvDG
/k0O9os0uG1X9+BVRUJvdpVERr+Evy+gb15f3ZaPpIoqkH6qaXx9z9UJIsCtQmx9
ZngBPGppWkG9d5HW9FDlm0RtyjeE6cpYP1K/gH1zabRzxjYXlmEysTOddEe8Nh9c
AH0zpErY5wWFDEf2XzLlF0jaKF5UE7Pl2DHsq/temMTtsvIc2M3OQ817QBcWkMmH
+Y+V4dEE2dLK/2BHRLnxQ+vjLEoxLRRs+NGzuv2rWQY69SL8dFe4phfeT57XGKKx
7z6Jz+2qkhLP+pNMdanBRaGFnsGMqgMzjY9PIrDNEijCcvSag7yXxLpkZeBw9EKN
9l8gCO0FNaWyUaaXbN0oawSQUeY96L5hrAq2QVb20d9fdWiLq6n7Lfc1hKyPVNsN
ihL70CNAD6NHTbEyveXDwLKCRuu3T7XkyTNnrjGzNHLNvfOMoQ5M/ZWktOpIyLbM
YNZ88+vNWTxmP2eqRZTs0GyGwt8Oippue2v2qDchS7uRbTMKTuI0KezGKjyytUPK
/iX2GVIobK4UyM/BpqQ8ATOfRRaNVSDUsRmhuiW6jzjLB5494cNtZoQju573gRn7
hlBJQ+8zYzBcGCj9kgK0n2BVTZPWb2baEH/WCn5UElPS/YJsIrisjHxjcRq+L/uV
f8bRrUsDXd6cz1uZG2v/CouC/VOXenTBN9cjjoO6DmIt8ilx2hiae2L6nX1kWpiw
CatR9U96gG6c25X6A/MOqFhKW2Zx7un0aVM2I0SMbfJU09ZLT4eGcGUYPjEXiAr5
QGLCLVwduS6AkL/iMk7DCtQV0jKR93q1Cf+m+BkVdp92msmY1Bi/CwhRZdQSyBCp
CdI7ploaCWVOx8bxVCkwxUljZ1ViyzIuPhwfBg/YoEKUMUa2CdYc4atDRnc76sBb
vnKkLmsV+a431Dp4LnDtYAUai/5eyZ788qw1D5eT/wUwiJH/Y+JZ2vmB0hdA6kB4
or32OYiek6ds71kR4cSVD2dFzICRaf4Hl470rOWM5Z/V0S3UgIFJDzliixO6Awcp
EConQSTuogBt0aOzRRrEO95749iUshq4jEcdYmnlnc/iIZfQv+qUFVS+nXLmb+Ww
C54S3pSAuS64BbMzjDx6IYKcTVOTdumUAfdp7TjOh9Fwdq5HNzCGQReSpShalvKe
JtFtUnNFTX6HcN/t1unCuDOSN7ZbnRb30IH9lihjGuJVuPXmLt/ACgbmxgU56O4L
zbQwPPC9yarE3PQL3Kxt1OixCIa0+I32SQn38r3Dcd9p7Umr15W/lI0Op05SmKhc
A95EtIbm4V2NviB/yFH8IcxGVOB0VlAO9HANa8g3WXkvkZNksmturyLvdxCvNolE
qk5sUwlBRwGEZc0sWpQAZfkY5XW1BXDo/fiMxXi21vnFOeTkiW4KztJn/uPpfRcW
0Zh/7rLs87qdv4ISgvWaQ6EfEan1edUWKrF5AHw8DHd+xgiOgI7FD6pnrk2HE6Vw
qdNhaWwrIGR4Wuy8soPMCxeTSSPPj6hr0AIp1DLA0XtLLEnM53M7EOkBpkH6xvks
7WxyIrYt7KiNq26xbxNx5LjM/CBIKBb/MLfX0D9v0bIpbBU4076zXIAMtwmSzwS8
AkCNlX7ughHsWjhfB5PzQZfzFFUk6ZtIjam+jLDVAELiBdo8dn9RAdZjgfjR8STe
hx/RVdFxJrSF5gCHj7njEXdZtSs7GmK86Dh5Hxm/FK/K3FnaSaRFGHFknX3hqdJR
AmGILzMAK5W0kCo/MgZdOd1daf6RDOzJY9dl5DKJZALfm48vVDfTPZ/yrTL1LHve
MEn0sSDhJRd0X8HprJoFREr5h8voYy70lbnls2i4sIbljOGctIkqIyhQmTjK8PY9
Fk+ZqPhzRq65/4OAACQVxm8++DayoMZdf9RXxeFvESdc1sdygP/eO8A+2b0vmlVd
fODZiICK8rctAhTwhQT8ZsfppOvibW5OCMHb9YkXNkTJkmGvHKtcH/8ioNSVjMSF
qxRZcKs3Magh6jrXjmKub0OFNXMzUXadvlCvvM5Uuibuarp6jpVM9+hSMnF5iUkR
c+bNWZJ7zdM2mCAUbH1bxN2gtcrmB/szGG7yjE6j/z5tHTGwXMMfxhpGQSOaWOjj
Nz8PL725EBfUzyT4+jvGCnAJhlnJMck1qZmH+Iy5BNdsRIwQ+6LzoprYjzDNRkFz
z6YC+qwYon1wYDnRbMvM8AVaANk6bQoKO3ikhE3i6/8uMMzYlK5yYq9qKoDdHLN8
2mwbYXFXufoe7su0Wk9QMgTU5ui/lY0tag5bBmha0heV03gPel3HHFdtCRxK2puy
1i9vmmP1JfLQF1bDWM0X9oM12o19llj4MyL+lBa+3me6tTjE0G7uSO047Fg4T5f+
XSEgOWevNVnigIgGbpl32nWqdn9X7sHJWpa3fXl20KGj3EZy05zdwx9jwAX8ZJ2E
Q94NNsP+XpJ7ivWcVDym7tlrZ/+5lNW1/xMTA4JbqqR+yxqJRP4ABTBG4YblpjDo
IsXXmkJiJrly/WDrDWjC2T/LThh8h3a0wZ/099tfECp5gt39VvDn9Dry3J/yGKUV
Ehk9+4BdDO8YnFV4PKcRvjRjx477tTL7ZDc0Qx0BfOnqgeeAYYQozRLwBAZA4obf
jeTCPSDaz5ErZfmOOy3mSGTetS+QG8t12bP+J7I+J/DcvTP9clskVjD12mAKvlT4
8A5ZiqbAirIvEcoTBWMTquKT2lD1DhfwxW8ySGdl97YG/PFqyZ7KJXbaHoVH+vc1
9Ot4nQhFYbHNv0kCGGGt8bS7vfipB3Gx9nu4KyqFHZLhNPeEuXj32S5UURl0yecO
J8rLno7X12nRdCLCMhtB07g/0/PLEkeS6jn2N2bVYj9HOX9KJj4YdzByE8lA5Kpp
bggLUD47hgBxo7yhhyvKz3Q4vNv+04y/JDUy0eDAoJIH2uVrN/2G/kTIB0pdNUh8
1uLCnLaxvyBCI+ptU/sFXBaO69GQVStx1RvT+j2xa4GriQyOQTdk4LDBLJSZrdaj
jIogQNcnsMEQwKqkCpzCAkf/nfnS4Qc53tfmKk7piX/XnPu0iHbw+HG+CEsB+CZS
YClrjDexBaPWC58II9uTyDZ3irGYdTesEseL44H3ZMF/Qi3q6stUB0u/ugNMZ6+M
xluBbJHPmq8zTF8nfL3AnTW/7zbZbprzV89hyrWqHONaLwsDk4QuSbn0UICt0r1m
7vOXcPRj2KqAmqE3pDUbXxYJKoivK0vLWZJx/FKcJOX1rKQNZewhwzKRnum6cmFk
RR7tSWsTidNEbWIt3y4Ix8pdQcrA5LhUZpYMO0wwUtsBOoOWnMgyZN+VK9RxiRYi
A4Jk0f3swDlNzqKOxbQvglqQbdvpe27zHaKuBXCiDuuFBVDb/YfyNM5/p/MnDdjS
LEwY8ZjECspjmDr8AwgHBqGpNDOCjuPnBjTAatAQtlRgpnGM4O1Yhm4dKyPT9Ege
UsyVcZqcQCEOc1kZAQuB+d2EeklUY0oecB/JxQKMQWuchNOHI7ISFS8kDvDimzUB
Ku71WXoGjB3zuZPcVqmM1o2/JVLvtA1oiSXbXux/HoodKMs93xOPe/CxySCz5DaB
NiYAtlYBEtpLMGilrNtdvDXvXTLqp22SHusA/K5TGXbOlKNSsrr/I1sYGZNbMPS+
rbnHRPMms657mLKsGBxci7wfLxsupr0fYYU1mkS8LXE99l8dDSCDVhlZCZYT1Cei
VgnMUya+uzMC8tKyTRhkiaclsjaQMKSLVhEywl9pZS3qE2VU0iiRRKd23sPPWWcZ
w240iXOKdPxXwRccFxI7I+wVVLuYk/T0UjHTRdGYC52YQRSEek1bxlkDj0kYPIP7
PCj6L3ipP1e4wbLDWYtSAyBuPQ4caeGMcZdPkA4IyX89BIYCoMTfq5OuKWlytEBg
1wIjK/mmSuwLax3NZDT+hbDfjBPaXRaCUs39X48Jz2b5hdBefSRavb413Ht9dfTE
BPCc2TQ9ZVSsSktFVKc6g8Ip9RnlHnwkbou+wk+tYiZBW1ZfRxt4DzYXKgJ81JAJ
GQZOXU0MRWAW6I3X6+lZTBB4Y+11M5zmy95LXUWvpuMlx8+CJkFE/bpqJro7hAp2
FVr/YOvv7ZMqv38lGuusyPYFuWfIeo3FcbeCM2TXLub113qLGBq3O764ec44M/Ju
Op9n33cU8QXa7xCur5oZD0IExqNaxuOIa5xPR6BkLz8nHJIKk0gwi85bUzr8JeG4
IzEcp1w3HDY4KFCc0lbZuTwyIwdiyADWDQOSjEu33htrZ0WODNJrR13Ubfrlo606
KkrQ7h0iXBmB0qaRYf7MSZ+sqiIHuFP31yNY3OlCm+EJ1RkzH2KCw3TjfS0qc2+1
qdfbmpriFLxGGLHFFjtb5hX4QDibrBMdBvzmzvXIc143CR5bxEm5C/gVwj1WbIr3
ziY8x1SeRQe8T34VSJRGkniR+KZ4lGkHjGn0GK8zpoX3HEynt1QlSl2BVNtc970U
uhcNrCNVlkH0r9rMx4Hv33LEJNPGz8g/VLLthhD4luOeq9WKVI3EkUgDA0PTQ+VR
kurBejzn8ZCG+zblqZDcx69hkG6XoSn3goFUFZHsFmkhZierQfDRLAqGlX+s4SF7
vbC00ZqJU9Dhc0e4YgHaFFLcQjhEh72rcgQvR7Dvuzy8eG33UxIuhUMfCNCkMKG0
s9Hx3GrjnfRkhZ6mPfo2b3LlTxwN597HTSC+qq8ULP0lKLeq6XHXuMPN2qA0FPDm
vzYPNXRWVx6Octc18TDT4ImMNskI8Ra+BeBXnfICbaileHjej/UKWtFNeoF7f0uh
QA0+mk/FyKInNnQ2IwWlNehKqM6nkdUZ7P0+F1WZHSNSWZmlp/DptjVRdLS5+9/b
v01Bs7dvEd4X+19VRgWG0uGBZi3x2tG7dX1tHMlqeQf+No7nC9Q4YPUwrjXJMGk9
LSWt6tB5jkvkhdu9rUD1oZhkrINYgZcaZdUi44hEYOKRpdMToDR0qAVG0FhRCdzv
xvbssA5y8Dcz8Z7CLPyn9WKfk7eEzXZCJt0pPHrWQKYKJfXSWNhxCOif1kBYytD1
mk7AhGVis3yfs+Hru6bXxbv7MSMQj5kE44H+jmnMUl52qM6x02XzOtg8SJqokRja
QCH8PEC84QxXEuhJ58N+Cg8YcMxksGYsBUPx2SYHaK7Du5VdVdkrvfh+QYffhRd9
Yb3rhOh3tBTfB9EOtS65rIgVPynMkIaXTy2feG2/CshghropYnqYxaj5Svl9Ym/1
eqIp7eGenrat8Zw8ZbPZoCs5KUxeDk3izcer6E1WvvmM4Ch/6JwTel3ZMbU9AK+4
0i4E+tjr1Oa54GhoNG2EhKKIodsRFl930xj5PC2jnT5/TImKyeIivlLxjMmqVidw
um7RYIeKKks7872+1S+x+k3hGOTz4PkWDC9uTBLUVudgDG6msCdvqcLIYOV8nbLZ
2DUCZv+QbZcFEtfmNzhDAcUMQ50MJR+bnyy9unIJcbq7jJ/HWmtpCw41VKmM4US2
vmGR2OXZaRiIS+uwlglkr8gP09DDjcs//DyU4swo6LedHWu1BXplHFJgefzRBc14
pqIlLNY6hubn/+iw852Aht8oxws3ZaPfbm0NlA0mUt+svJLm5VsCAK5xMwxbQPvW
CT2vuVqAj53tgr3euXmItCjKGy/fVv1LkXPb9AF/YF6LyEntKelZBIJ+MAGva4Ou
EWg3hlA0iT7Tj3iPg4I7BOHHcsBDXwxZmAVEvQwIzEsx+k5wDlmWFuPMCGF9Phgv
DLR0TUKq9QO5IOKyafQB65bmpHxKmyPFX2YWTlCe+V/t9lR+qkGiMpqrD85hNRB0
MYLgfcbVjvR6uX8huuQQeLDUeBpzN6kIfv1V5uW/l7NFjPzjx26FXLFdgk6fHb9E
vWLvRvZaolMR3szC6prBPn9zx+1V9J9vTEmqYPFMeofi/fnMUJ4nnSuOsej/rcsV
D+Ij43ZTRGI6fnIMro9wqHq5XVdATktwx85UA7Hn8uOv22lMZXfnM3gAxeJrD7qf
IlaLpwkEk55NNh8ZWJVFuajdGudvtEE3phUyOfcRwT27kL8akplAkdw+niVqNFOM
yIZ//MSRv/PVAKaIhPEWeQPwUOuoSqHC7y+E2HrOidjvKG/Gep4M+R2IEqR+XjGQ
tLAc6EOSAIIxmKPl1PQ/m62Gg/0IU4UyLu/ElSS4RlshQoD3A28hcCA3C7GvXe2j
IWbiQS+IuBay1TJbZqdFhzl3jmdRloZXyUcp8L5Nl+6IXzI8V+BIXGEaQUoJKy82
WYyM+b+Y1rMTFameDLepc3zt7iqrwRfqEOUTTZZSO95/0n6dvKhaSq3w1EMc06oj
4n5flVFINwCN2QUrOVwqgMse4vG2HSstF3nD2/dctd5FLG9zZenHUxC1LQyXYJc9
zT20d9Cfiv4dP6LOV7mxFvA+aHoLLFUc69T3W2CNbEKwnb3F9Nv0OLw12P/cCzG9
ZAcc1nlwYGmT4xDlFDIdYQ7ud7jAp/3bt+dfSiTJyw3dQGIsjB++WBJafMgfIZgt
rRMZ3T6lwp7n2atA/9LBt4pw9+gbx7qTFmRQlSzgYSDybHs/uRkhbtAlxBsKtJfs
Fk829TQDfFrxy4AlImkHzTGPHXZ1Q0bS006iy1AecRuoAwPy4fre6CAQ/zCq5fur
y8mbSnfVKdibIFdVPcMde4ho1P2VLY/HsRJg/RYZdzh/BkPK6gPck3lZSZc7NRHj
zNPVfoYP9y2ftBf2iaBNiNjG7l45LzLTNNyuPnlKHzGOtpH9+2f0tYzELu9soAKO
K+teOPhaZ0RdcdOB0MLewWTDo6XxGkGG7+hTj95ttpCtX82wsTmvEPwViSohokLt
xHuJXjdQD7vo5X7KhW3Lb2B5yrchV/Bil6lry4w8HupV4EBs0qL7K6TzMG+PiFLm
QHAl2EzYRl3uNt35eFcEiluNybfaahfXL1c9lVcmVh8/oWRzXdmjZVdTNNQvzrsu
m0wd87iMHryIVIAteKoURW3ohw0AFQ6xGJkXga+X6/AZGN1nvpi+rItI7nbtEvwx
wSrSnxCKWuFvL1QGLvGc4bAoT8NQJqUtjabnzlk+ZV/yzjYiEK4TfsrCFopQib3a
Fe1/YdqRuacE/li4EUccSfIHZNfjs287stQzUP+NVDLeZyw3kCG+/eRjIdMmusYh
p3mnFvap/orE6sGhXZkpqv8Tt05FSASV0etQZvRiiZlfgfnM/JrYQ51/dbHr+Y/W
V7rnZNTtcFyMV36QfaW91fBD3lWu/fRC0AwlIlvahrP/GE4j56sIAAvJI8D3cbLo
yUP8stRqEovDPyAt2Yrb8HlzDHA8CqXpggthZGYT08TlGuUTtfocZK9MjrEqEXfm
9WVyxNMgw5jgQPUFiqSU1AschgATV4rAzD4opb21kGj/C7iZz8B3KXNcOlYMEw1n
BXEfDBeIYbZvhnGH/fucf2Nr8APsrXDRt2MJb1ZpGNjMATjUAuNtQLlo4nSuHXJc
RwKbJLf5qOjd0HWCyG2LmLZJ6K6GqIZ4LdnXT1EMZeiysRzzWrmAwE7chZ+L5Ebw
X7UdqtKJWawBBv+BJehcRCxrmLMfIzgWEgBBavgKuXVQY9hO/kwLFutBlYRO08Sg
F00TKfG0L/VqEuXXvDt0EVJ1ivs52zVDhOQ3kc0Ce78NYTgXlyBp2YeTSYsgKu4v
2TVh6sm+dJLmQC7iUd63pEw7enBHv7vcRxfO8Gmfh8tMPTBwEycKmSdsznhBA5JO
AT5UeshbAeqw4zmUnntp79aH8jmiAfack/B+hH7kNX+61oQDZVWhMooh2lS8bfeR
hUjrYiHKYDF52SkRFm3JchkqLxDVGy5u0FtposfUFD/claChI58b5fYy2uxTWT8A
wQljXU32EtM2LGle9qqzH5aOuxORjSunB4dzwotQUys6ks3eXS0BypP5SxVWEddm
YA55L4DszSz/ZU4fB2+45FImy5xd9nAu3bX2Q4MeVAlSh0KfmAoLfHTba/i/lcML
dq21zLVi1RHIHvpzaY/s3zZPQqVXfw1tTQNYp1wtfR7UUTPkD5kdZ2vq6yspIbgr
WyucFExJdf0PxSdfTBzlY4OqT+lo2GWrD/FHhvXwElMjap1/UBG02IZsIvpLGcgs
zs33FD37VQMVxHIA/pjD0jESrwnZghBRogAmM6cpiEfbIeixh1XAAy0PdG17V1YS
V9nfFdBQT0WSgCi7f44RdjCYx3aq3PYkcia6P57j7oupBpneumVQJHY7uAZTISms
GbuJHK+RLsdDwslZNMz2CFjUvgFBT8UJBSd7qoFE/EE87veZL1gyiOeGYJmdA+Nl
EAzjU97ddYAJaDSq0ypTPnmLbRcysj3z25fuSHk+1BTnJNwz0OdSPDnHVpTmd4bR
neUPhLaMJEx1Oo1hDNVb0DevQcf/vOaFTjxuFKVCG8l//xoqDTuIJljUw6NbQu7R
6XZ6+J8HvlXn2s15GCAmHLKksBo4ESis5OFGTtpHOoLeTNtTrqVnNpjagNe/cizn
g0i3nL0rFTNHLAelyLH2jWPzsXmbYmsiHAWtfclcFy4V7skmrHKOsTOwuT0IKvkn
SwRJ0q+S9Ou9nE7pFXRa3hhCsj7DnRR1aRkN060Vi9XZfizu+yFGNvSLnHXqM3wn
wdybXU6E0IsiU2YDaMbx2/GwXwIUkq0+WPVKrb8uO8o6ykAeDsCjv6tmgFaAr2lO
66lOHppKWUmCsZ3SZBwKBB8gKkoORsk+fTkkCBRRU+fja4DD3NUCp+P26S5F/o00
oE9gsYWqzbXmSVzG8Mty1McPE2rWbYdiat6GougO5mYS8AV3vOIbd5Vr9I9x/mtc
Cggq5kfkiobQalN7CKMWtSa8y0m4Z0PCHAwXM5sA6OUp+gk4Chbu/EGFNJUjCNg/
cdX+XU+VhRdQ8KV0B+EsPhZIA0NqC2OGrvbX6Yx5De/X7dj3V/mIzJl813miQcdJ
dwUFEDOjeHH1RhlyP0/AkVrgKwn0LOJpxd8nJG2mrkHKaJkTx49GJCzfceFcBeH3
5Zm1efY4msb93w50Jn8Dy5jNu5i2q1PF6CheahxbDMLNxQ7V1p4yE1HkVSBPukrt
oO1BdqkpiA+qwvxA/3/cf3/kIxkUDf7PsEA1RpG1HQ3CagiOEdc3ZnN5kCKpYMsT
XHh24WOjDG4kOsHDc+lLublMtIfNGg3dgYejh4SbDzND2jxAbBPdNHcKUHjSTQKL
bhXkhahGVSCRKwAgiZLaFx0aVfp/w8mQIhqp6bnoDYycLQKhP2klSjJkBGZIbwWg
APDic9IPX3yOIegs0KBUDgaB02RrgvjZlqzXw8m3lI3hvQJk/LPdOSN8LSJEgzQg
DuaD57hC7s1lOLajrMd+8odNECZlms88rUWCp36/35Wu7A5SVwtALEW30DZGEGiu
Cbuno1KhbI29x4LUFiEQ8C8poMgX5dJ+/Daafa/Yq3fJYDeuuNVaLHoBjnWXYqHK
MI3xkMuDmC2CEoBvQajPUqDts/60eptSB+9W+653lHZdWaJtJTnhn0gZ6cnqqm7N
eL/DLW9+FrSQYslO+3JzaLhXfbqR4gqJ6ac+e3klI36csZQ8fzAs6WmXkZS/5MpU
W+e86/xJil7a6IcAAFTLmAnzIAW8z9eTZvTFBns6TafDIY/JMOpspbqAiZeGRcGo
v4RHDj8mnjWHvNCT7Y6TJqMQJw5PcgRAVzS+H8prZIuNhxdbqHJi65OztExnQWAW
/ITDAASWZgAqnUHkedb9GVFqNQmB10KJ+RF6xXYfElwWgVOdFnGwZAVMsAEz4ePa
R3r3WPWj3evqSPuLJi1phtWLghDa0YThkHDWgIHzNkkrYwYWGIaaxJlDCn8USOxe
3ujP0D2rl/qduUVptI2tbVgJyqAaWFNeGNXZWHORh97ojnoL1864sCzJuO4OCwvz
/4HFhRF6W9KN1B4Hp1iNaN3FhvkqpCFs8SBdqaS7TDaMmtsrQmPNrhgLQScjd83s
acHrRc5WL6Jb8SbFbxCHwTulH7nbHvwj2nHVEUtupc0jrJijDFBLX4txBjmRWSW8
LUggLyeIheEFMOzS98W77b6urL2AfLPZD9eaRFW45JI4XBfT7r+HK1/jBo7RUGLV
n1qMdCR/90qjSJEFeRM0vXKE0cl3glKe2r5I9dSaPWIFppfCr8F6zZs9sPkg/9wA
IutDRcoZ5V+BKlpItMf4s05ZZb79QjpEUdE8/K7GmorkQfZDQ37R5J4wyLkAXK30
LSeS/QnOcIQfEUGEgHGvzUz6/fh1lC/FHZIUVCtyysPuF4eQCVTf6Jhse6Sw/NZl
e36CVUZvpvvOS/FVgW1fPwLVnJx+CwLCNwMiSIShCmIRG5X/rO6R274LNQhG0R4q
2w0wAZxXaf2J9iRBtZBCH9V6C14rdxoTunmxEpnKPaqPf/UXUXgA/UvX03MEMrAi
cocl/dspiBVmYMybi6cbBjPsrK4DubscE/cGY3LE0/XY7WE/+5zm/gplWwj8QHrL
vJzhK/0JTbAjz8ph+EqyBlcZsjG7mVOfS9lD1ln3apiefE/5GhIygwImVevNLdj3
KxiKRofJTg/V7Ho+YlZgFyO+ALxX27i+AHFghZlNI1/criUocEY9rqvhC+5DDfus
YbczZtjWdI75sXHpMpsAnwx3VU77NtWRK1q+kueI4+2j9t34Kuo+jS9oa9hrH5mg
58u3GdC+4F1w0+JMrrC1QtWldQVpjVkpAUzpYqBvz1aFMB1ftWb7Kf/m2ZJSwYNR
qSbr2AnOyCWm9H/XuLIkxgVJDU4tYAJsjKwYxx0h3PZJXsxEjgQjqgghXuQHO7CQ
P80iCMYhREy7RfmMTo22XPP91mr31xWk97uUvVO38uuq8zMsiVQPeGoeEpSfMl50
IJvG9ZhAF9FC/FUlR6ihltbLbRYTCZsn7WVZpBC3bt5Uke5Xxq+yN0UqjAfuZVXI
odymZkYbohatWzV4SDtL/oW1Lyqjr39He7NQNs8Xm6NjtW6v9q37rr4PbhFMK++J
8yCgVkK1ZoKMLfaidZd1bDOODR+27UWl4vWIc7JBeRRaEwoIupIv6tNfqVkiZ3fq
PAgRZompPAG+6reDBYq7c3e6Nbn4N4grgrH+Iw/tf0na3Jv5rQ2dI0O4inhgRLu4
Ct+WEOilvrCJdNxqADoNm0yB5lTrEUnSLpt8H1A0ZTAVEr51qwJf/2sjwq44Cu/X
jof9ShVY6vvjNWJykETmS0ury3XDNyUR9Uk8/erE+Jdlx1imZyFd3A1FAwvBhf5P
f2G4pA4czDyZs9OX9x4ekA/lCtAQcuroeL1q2c4Bzoy3ML4Vmv2graTrVIZmCN24
mAD0YKpnwJaAoXJ6ow+xEwAnJ/U6bNt3Wwwp/PasLB1mNwCdbw3LXaM5cRnPmIGj
VE/QSfohP5zFP5Z6Ps0r7nVK6kdvp93fAfW1fYKPtwPhFZl27qKkq5uy1FaEyoxl
WqocUSy7bzUmSRl/PEsap0p7lOj4CAvH/cvXAvv6BST2AfUoyaJIJIOi0aJ0OkG0
wtLxi4KMxk0CJQtkroUa6J9F7aYHR1QKmCotVgeC5dWRSHqoGLVs8Ka8qRaTfp+B
SQYx1O5g0KsD58yvgBhkhWPBEoFkIFXcnqv2qiOEBopjh8EnG8R/5m8JSAT5T9k0
4iJ2buvJEBmDeiJ9/9vZ2XGIqlVHxGYGbQcs2/btgDQCgp5hvPjQzYCCdgSZ8k2w
hMwcGf5ekEEGrp5Voya8PXts4F6BFWjFVm5akSuh/VbYL4e3fJRllOHvkrSDqtyt
UknAsoidlhKlSVetv3eVjOlIxw1VGf43EOUnvdj9DYGQOOvMZ7WGJFgnvupl6040
C7UJhGYAp7oAadWlDsJiPYlkIX2dMSWYduOd86J42VzfQaXeiAddT2Tegre4IlLH
rXcjol76zsVLgWUf43D+HAxEffERMk2MvKYhReXpefv5CsEi3BTdcdi/y+jV24A5
/MJFmv2C1gThTf6V05PSMGokqu6wJNYRHK0mBnOGpETzC3IY59+NuBlgeSS2IQF/
+V/f5u3xsBJ+r3jkwraK21E4+iVpRV6ZJVVpJlIzCu67kmjOqg4uEhWti9c+IzT+
mtRQWshKA38TuL4NW6yGR4xuWQdsZrbrnyziWp8l8OmHDVbECLsMzaA0bDwcXF+D
We8I1K9+hVtFIkKjYbAR8BH4gW2hWQAGGRwYvTRpqw0V6Z2wwQUYh+rM+qEJ4IWr
xDmFzowgNTgcbWcRUA+od9EX2Gvci+E7ldNtONe08dr/Kyn4ReS95LSj4y03isjT
P0J1GrsTv4KPlcK+HC1K/sEbYfoa2XMKNnOdJ/kGwUlqidZxIQtj/62hyp8PVh+E
Z98EcP9ztLwrO1FiDAmhaEtYcJG4P3rvVAN5+TxBlGfsT/xMi7SiCsrpZYVtHJnQ
InS5xNezZiQWikk4nUBnlU8N9325jneOhhWSukeuS2KrUzqcij1x5LAwMAwvyoOG
9VVzpwVI+WlwcQrYM58/0rlwQTUnHIU5oVBMDyRLCMD9+WIHeWAnJlD34RdssqMl
meHnqLYPjMCJFKHIg/3iGRW2KWnu2WJowKzoyqqrPO7UiuqTYUiiLW2LwatoebN9
MB8FMvnJAA8aFZlbossDX2z1QaEWV3d15rDn5rHI1LCcAKS0268w+80ECiNn+cLX
lzZ0GnTtgeGjItAOLfrm8H45FMu6xTLoUUNjNLsDyEYeKTz9GrjhaT8TPfjvqHDo
W97Oa6kOlH37DAo39v4KIdgVXbcXH2fA8wr82WAhFRUBY///penWe1wUo34cKsiG
aXUIuYhcEGQ10yz4NxER60UB6oqkmQSIEkkNcuhC8TrBdoTZvd0JP02ZyDIQgeqn
uw2E8XYXj/g9rJ7vtm7Arh+Lxgq58gGA8t5WYWUftwK26u7iqkA0d97b8v/A5y5i
28vGWWH59GeDgFg1ESespg5eoFzcpdKC8uR5C8Fos66+FjLVG01foWN5gOdHi+Wj
FyzixbSCuje1DQuTrEkAZ9hKhPQWyihHSc/qNj0OG2bAcDGuU3f77dhN6DbHSA2t
HYvoN1+8+Qkj8WqGJvp9q9CofYv91eQV3CS7O37LQRZqqONpU9djReizAbkV8z8X
r/ytQ0E38v+qdfZEbmdZ0HT8Qr4C56dPGnPlwujzKCORX5mtzQIskGtqZNOENMtB
GYKsywdqIAtRE/BbSg6UwKmc3jFXUxW4FipEPa0ta5nRIFalE5/8sJ871qAfolBO
MxS/4IPUyUU/BESqwgUWx9quxxWgzlA+q5f93yz8/9xFW9gQ9ZIDjz+1uHWY++F6
scEB0lODdc+5EpOSKxlUsAzyUBX/3y9HtWWZTUARidh20WpMbCcSE2obrFL4AhVF
jlIWc8qonNkqsfEcG2cvuKR/pG3AzgkOboyrid8nPH85qfkGmrIUQl8UXmZnKH/v
0LHHUov5SVd4F4UfMPha5f4iKeM/59UQpG9hpPcCFO+LDv2j9LeuT+GlhyVFhc3P
dUOciwmRbeBHhs+QnSVOSKMa5olTB+4bD3h1NUP9wRvCVHQ91Stlxmsj6Lckwt95
uBYMBAmBgpbiRMa0sFM5icrO+uGXlwCK4UsBuaDnp5fiNIJL7Bcy3mgcBLKgjDEq
xAaAyBQl/5v7GNPlYMABP19Z3AOUzm2glbvd6KQGGRwT7QmyU1OYx+QpHQi8j/2p
qr4xFEbSTqFlsH73kUGchLYdyD7PvFA7YI+/yhF3kRbkBlQx5q3V8XzNPdhzu/Hm
ONZYvEsSdv84zsuceTk2ZOsE07gSCSfD+G8i719auREC7o0Qu9AJjqR8voEWS3wD
D+PbIwtD+5KtPF/iyhpgYu0VYKWHmr0sxCx548X3IUzUXvQHz29LwF8qkmnkriKW
gpRfN7kIQJq97zlBi0St9BGtpl4rcBuXnrV0u74giObIS1/dyS32bsiHTzfomnyr
PnVsdwGCo1ZINxfDb5kFJVjbS88Fq92tslliIkdGd+1ygQ1Kve9w2BnjoFZdsm6T
Jsh7pIvnoKDCHcaLDTA8BPP2ryjOQ8CJr9ah87Xz7ibGq2BO8qsX88iLq+9Apge6
NPDe0k4aVjg4Z2w0DNlhuebdjmVzFEygyqjb+ECGW15bUk7z58+p7OZsHqB4W9wg
QdgAo2PY4vVQ1JRsplIOHklXfMbR6DUEDbjoosLhOkQBoZFmRz0HN9dEuv6uZ6+c
hKgf/wXhQ0/FOXJkMqOKmH/Tp5a46QcvjEvWX1k+t10IePYHflRNyU62XfX4p5v9
hFqhrI0fClPK/7En/gd6k15iMSbQsBDpxI9z19Cb5rzkOl/dgYIHRKT045XYeGTw
McSXXjciuXFaoYgekWi46Q==

`pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
qsuTa2yZ0bxpMN1x7INcmFRgTHYB+zMefwLYMqS4RAXAlgSUMx4UusFNfb5UM9ay
OPwrgbEOIj8ei7CtonEVSB0640+vyTWndwiqhXu3u9bQyYXfX0LW9+nThxsK0kTe
SirstEdjaNj6O8h5KZEhpgE8dcvKAAN7GX7ncLEmdxU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6496)
lczRdzj8U7vKZQKIqkDo2PcQffpzdHJVHJeUmmxNg0rRB70FEsCcR0FhEU/98vwZ
6+yd8rnYEuktBbPwwU8dCe3cUGOytJFRRdyIo80IgIz8PAvksn4O0kPYIJtR3Xim
c1UE/GUg9/CBMy6oCt+z1resxiuv06y1HoglYBPgsX04tWbBa2fXzr832rK+rvVz
0Uh1Q4TEqKMS9nkwWdqDeL3Buvu6sUjnhu2WK+T7ULMGGqGl4Nmj+Ug1TPIiKkip
w89y/7KtmtoEGFzaiHZyKJqLvJYp3v+wilS0u5C+1uR/JE5CrIS2pnhakiQ+Wv6a
NGWXzUZ6rVHf+sbxe2jhIec0aYapQKUCuU/ExBBUKgdqJcTbRK4z6FwZbvESyakb
vhZy9bP5PtRgMfywX+ocZhlseJO+pJLyJW2JNMyGPfrXPTFcV93qdluJuZImk8yG
YKmbSMmaLXQCObQQlIW2q3kNc9ZD+c2dnmDvD6R4OTjdTIqjd29/poOEfH0pdmKx
ChktjzyGHOA7l8XHecx4RWx0NLpoaSDHQ/M/LlWgCMEDTjrhehEwdWND29VIBIR2
xg8V4iFJ9JAgmWBbw2SYwPxaDO3OwAxa2xvbEaN+CjpoEE/3U5kroLaAEm/SB6p9
E6QcmnWXD21gMNjvMDDJHqCpvuVG3+XbJD5WV84IF+3h6IaymqdRJAKNYMGVZo1p
MhXUaS4oHzrNIhxPqe9BAzrq88ugFioCISljA1JEhp90OxSlZbpBTbzuoAc8LvEO
noSGb73KtoLqnMZ8SywjRz+lXUNp8C0qNYnyYOmJDXhy3D7aUrCD4K3gdq4H4bsm
DLEOKIErt0X6z+gu1UHG8+mW6anPrTHRBn2FdEK9XyJenrhUeHTAXuJK4TlcXgmG
xb+0ubUIA3OrKqoxVSUCdktEg4w/JJygXffY1I7kBjnmMVpAByU/vFmv9q9S1vkW
yBn+N79CDX2lFCdA99o9Lryzmwu+ycEedqTQ7hmY0PIzlCUK/8XJdAAXxJETkFez
x7CCGntc/aH0uYojb9bhPInMDwvPt4MboeSkm4BT0+EoMhcQka8AwKSn/IG3tusi
weoG3fB7t7mUibHsy59A6IIiYR6fr6lMow8decUCyrBPC4vErIlsT79Vx62/Acdi
tkXWYrrUGUkbrDea6Nd7Ahen6l9epm2tqUJJPdgTwpck1hSigev0VCwvE8EtPUM2
Qn/BIDFmIU+VLuX69CoCIDuYZd2ytNRF9UoZTTP4JZsPuY7F7AW1kWGpjEdJ/fzV
m8Z72qWkdeBgaZuBFiupRoMonBtotNToxdxZeQpP3vNFNFaQzDy6DkD42Vep8Fhs
Du0FeTBTnPoSmSghfHVOG4qkzaeDZmx5EllWj5PB439sQZIMFoTPeeVyeQZsp2P0
d+dxI2Yjk56lR5rCdbVC3/1UcSvhLoR797X2cvCMVN/hWE9gr0z3vBT/FEfh/LZB
n+uVXvbFsQgKQ0OcLw/Vk136Slf0uQtK+ghnRmaI5yAkGnQRiuur4Q+IMa2UFQwK
Hley4kdb8z4qzBYHHPLTg1D0RWOSqAzWiECpzxMAYNnSU/q7DGgzR3sD6p+wh5Pi
gdwQ1l2fWarUIeuvGpCB55WbueaKAxU5LDR5xJhn+B1VkASFXxViuKAj1QhkRlF7
NTFFZfjfIUX/5OR9cm8JWypgqHJqBiwWY3AX1OdPt2keRgXnQB4LlgWVPsG0L0EX
3mDl8mWKB05jcmhIdS/JzC3VR6tjhYChtbDnbA4bTRWoRPg0WtopzukmtNMx1ntI
S441wke88y+gBDO5Hiel4LWJeM8d3WtQoqU4SIn6c/3shBNP8N23VwW6vIA03v1u
T2bfWL/VG/4PTaT2OJpP4SrOiK5xpgTsr8lJTrxAVy479fSpFTEXTRoHEZBGhhvL
XF7KYC0c182b/cvG/nkJVUBOGfL1VGzOI1i6P0D1OiIDz+FlUyxrpM+Wjq13Cb3s
xQI7jfrLSba5yUpihJcEZTkos+Gi4a6cn1Qw3RFnaqevJYAiujp1Mt43A9Xi7Jmx
2GXKfNmgdBKs4uXu8+rE1CE4nHDr54B2qWTfPXwigDUwazDizjYw+S6bE1tv604U
vGcZW8Xfm2H41Lx8gJ7CQkDxt07tzyfQAhrJ+iJ1JIwogCMgXjEyQ5Pb337mE80k
+FTLaR92HXNYI0MTmTg3vIiks0qnrdN3XeKD25H/XYfUOp4rPnxZ/u5fPCeEt1dC
r9Lrn6z7CFDjPRvsIwtme8xoZU+wMZiQe30Czkie7kzLzoG3Eh/H3TxjEAzLBK+k
6+xmYmsBEJ+F2kkIpto4GhYl7m12rdiQEEd4SAJ15JEpuux0i3/BBiBP0t7G0ZaO
VDF0/hY6+EHevyzSkjJ3rK69wThmelunh46oTL2S1cPp50CS7HrNX1Hx8uqWQsBO
G2SKHcavOcvYkWWBiUvS7x985om+Lqh/+FiWHhMv/J6004JE6d8TvnOAY9eEoj0C
lWg/FHhUURltO2iYN2NSpL3e00BnZ3DEMxERcwL3VOiPNyGsNlQo1Ubc+YeDORAz
RRbb2yUYF0np455XkjhoMGnH42Hn1o8Oswp6VVOUN9/mJSBOeiinH5xINViW3wk9
gGpvRl9FDtoaYyXnTIdpepeyzVxzo/5DrB5dIINlZTUtUFpDYPtp07l48QHbeq/Z
Nr0ebe7dQnBug+Wp8QKigkq4ZUmlrepro4vBvldp13rO//v2b0AIwCnmTmDKtKZJ
RKigZXgFuHExK+QXPlqpJhgDw0OVOiqw4GOuBu8JTKIR/fCQM0Xyj8Kpq2vEcl97
n5oEewFLGSHUhpBDD7Rj1Wz26BNOA1OqqQn9tp7uqljMBKmyFXgvvpvW9Kber8Pi
jEc2jkmehgEHYRLjN02IurWwjPCymAE6acbfr9WcIya2bVcIRnltfIOOB9Sz0n1U
RvrmgPkLgH/JVIgv90rRaKw9gDNV+VQiXDuLJAIcIylhRc/I0gZCkTOvydCLhGrO
wHferiAWE7EUbVb5DCORAGstaHwiY0n3tGEC4eybxJsqRW1M7i8nWCxaF5AjOkRx
ar7nUwWLEKlNxL4rZYPFKxBneIWqw3aF8snJ3vmHuxGfuKFuBMDecj8LJEIlIp7C
Q1t3laq7yxBkUs0aqsJctiUU1waHjkMVCntblgrKMJKYjgcShHOMh/xwrC331Nkp
IHTDsZnvo1ErEX21gcEEr5AzvHcmBf/e9fa0h4VnSY4dceuR4YMk0ihhoznBmj9Q
wRmKxjXfr/abIQV2mATFHIw99Ne5QdnZb/DgpyauEg6rLqDVgCWVhheaAiFTIF8W
2wJK1361XMP3DpcSZlCcIwFX9JzFEuKvam8gace+iZ7eiEkNwEn1Yp71eYji6scE
PcY0W6txaWkcxhgoVfr/BbRi/dAHUHvk8e9bQfDNfgzctkf4AkeKeJPJMfylWI8D
tlCXQ4JhbZysszwyb/ulRR0zABBRlk2ad8eURiL1yRA3lQCzh7W2nNhyWhakGB+z
WNfqo3ImQBbsN1yVSbJOiwu0EGof2+KryUujPBZuKQBKgIqTF/0GBG8GHvLmUm0A
dQaE6zL3hEjBakA566/Htr3AZ7BarUJ4gOLYjfrYSdVhN4qsclm6B2wErePLctJb
78YC+oJKEd1AUh+GLp9XGXXXb3xDw94gqbMsSyN/ub/egs0O2VmfhyMBlXIOTDGy
DmeVIKS9xsdygziH4t1ECL7NwYuKegiQlnntzSj7+ap1CzNA2MmqeDNpBZbdLL2Y
GW6kwMVZvDA8zOAGC9VbEMdyj+KMaIpu+9zEZ6PZCFzL+97WUAOUx5noZ0DhNiaN
Vluakr8fTiFZv0JTYUVwaKcSJ2uR9EccNs8DDb75hogvcV3qt/DT2YhdktGQMeNx
2BPJ6l/gIRi+TIwDeyvC8RU3ZvVmut0n9J6G8yfN7lQ7uY9ur0NiGce+QfojGor1
X6tt7UsLEjEIXhPRZdrj8hG3Ew5vL9pbo8cF/S95ppV8iYQXXlEmpw535ODUImMj
ysUdzwRsd7MITKZ3nWQ6581T2RO9uAszYLkIwQZIqmAXP099vB83O524bPEX6sTd
A0k/gARjSXhseUFE1tQO8I8j/XFPR8WhYlzLo7Jg4+H3/DjPC6PtSY6QOQ6Khfyc
AMIRbHZZBTNUN8cpE3WT15D8NDlrDZqc4y1cxo/VfiwpSQprOIMmaRmNFFyhL+ZQ
KGuQPgU8ptbrBXT5Dk/4qTLdyVmC0GBVTyhYWX70lVG7+9XIAI4YE7fToRz1Mwr9
JbPJ6Dp8kOrtF5yhu1jxfvWgp++68Zqj5gNlM7x3A4QH0kksckMhLvgyJ2dpAEp0
Week5cG6Xc1SOUoU3ZM9dro3VhpKD2kaQ2vmf192W9JlkY8ds/ydmhrau5ncrriw
jx/FOB3PZ8y4v9lPrPSMftttVPGRXgGDLEUGZql+E56GUfOQGkS0prsFsLamyzE/
NrGUUqSYZJRXRcKWOkwhwWTArf2ZYF01ddrY3ycQgpgpHP0wBDV+tkRza12iwtj5
etttV3a67kL6cWN6hkc+oRU7x07eHzR+4Xr+miOmT8ghbLYrQWMzsWLrTCTPZxIV
JXnUNmS1HR6uGTtZK7nQ40pnbtduAn9yMQkstMNgpN5PBHPlfgnRArwBvDsg9t9d
8qtV//4CNY3V4CLxBX1//nyXRzA/6MSQp+DCK/t7sTMCcUh3DFnXo2T0m3Q4oCWu
u/t5s5eLUV1AIIRyNQNZwAnPcG/hPDsrA9udixvt0D6rAAemZfNVeyliYQqlquPg
Y1qeQwA5pPdLbh6aTvRbO9T2mlau2+WL3CfD1YYcO5KvZ/EX/Jf5sXDuOJ5JwGWZ
1sMJr9g6D5xOAtev5E+ezLl2PM5CP1W1yG2lBS/PIE/tyPwJ+dVQUdCMIFHqAAfV
Pj5JojsAoaapkn8oFxplBYjP0aGCfaWRRhzMrjH8AzVl2poniM68+C4ptxotAmb7
su/RiHqfpsO85EF1edkFoJC45gMA1uGkKnmY2xvBzMDdSDVb/x9zf33LemwBvKxj
DLqfDo7xla0DP1R0cBCNzCwJro3LIqu/VSV1LkTyDt4IvOIWCDMwU8IPaelGMe0c
X2Y8NiAc3kw2csMjLKgRZmwal6HgEEZl7LdN48v5FrdIzP4kOVAGEpDm+/+wkt8e
jdqX0Vs3wrxN53jgx9Yj1GlauOzX1EuiLTjY62v7/I7SCGBUSUSdv8OkN+hil5Z5
1zLoKooyIRMUJ2A8CWMt8QtEPpNO8LTaAzqSDi+H8lBwOi34zw0rmRyvqneq/U9t
PPQIVHTLBj31+p3LIAJMNR4E5xQUHljrOLseRHhSb8T97sVXJx6U2H8cI5KMutR+
0L6AjWhXhPW8k/6fkDkQsHuaIv5hgI0uu0dlu/3rq0uY7U8N5FkXim8MIiKUm6Za
PcifxOfSGFNQl+OvGGTi7HSmjJbVYLWzGN1An7SjTqxWG80U4caFteu2KhH6NVMC
NfFKOxJRj0/2YW6r7skvyvgaRTEHckjBAXhVzHv9n/rUCgBtsHUEErcIMf57Pocd
UuSAAjRt4mNftOJSFqrsgfiF0b04bn552gF98tqK/D0PK584AHeAHnZIvsrYKpYQ
qz66LXvEOctNZXN5RksQSwPpHAE3VYDPqip4FKQbVjopXgOCSgjNhLNe7ibi/pGv
Ky5ivM3hpG8MNYuOw1R/7bSGD4d4rbQURVR2cvR5UEVei7ht67Xt21fTKkppYxYO
8l01uPTYv3oWpKP+7hyu0toQXzejbwmdtTJ8KMvZ17yqgU/zyUbjIRRgTahsKftp
xtR3g/PYCmMhMqwxuFD3FMTc6lFLUgiofPjNezyjTN4tzdQ3Sl/CA/XHeA1zU4l0
ycwIHL81QbfBTS8b1JiyfgUy5IbZiXFXxAzvqaQm3Xix9Ea2dY6vPrHaHCzj5RUF
Z/lU+YibRSzpjotJ8C3DUJZ+07gzgfiaT6I7SAIK0Zw2r5PWZWcWYtTzJDEqNBjZ
UXEdnse83LIvYBUjmHutkJAngitAesYA6EbwQFubWtXoxr6uq268KCMwcjEfEk63
cLHuONcnJVxHqzXxEAmUw9AIPn7gN6G6HfZrPMzms4TFE3OhcrYyYEF7MenCpNeo
CF8bDf7U/bqM27JTT4fIJC2i7z/BnCgACV6ok6OQ0SAAQHknD7CbFJg4GzP8N/uL
b2UXhE7ni00S0h2nVaqqw931G3WpuWPOEtHJsTPp6usLB9+yUzxjbGhxoNlLKQ/+
4FbFgMIF4m510FTTk0oZUync+pme5ktfEFMw/X0zf/urIFH4CFPX6oRSFkUgw2el
Dl3RvyEdU2FFeA2dGbPevyxNfOV7UAZw7Z5M35JoeqceJyzaMlGRPMU6d8OTVpn9
rSqa/kIt3mXM3Tg2DzqfiLDDm/2S3p269ep0NSk48PAC9fcI4PFgX2OJ4gE3xxOB
VeCbIxnuBL91NDbFzEzYaW8YbbLDgO6wome/9RzGzNMwddVjsfQyWDOCH7wjYKGp
qJlfvK1LysLKnLpQQ54CU29OmQs2yPKDaZCSNBkmfaMSWzpGgFC7Em6ED8vk69aT
DsZ7n06+jES23ypt95THT+8h1uB2cri/Floj/Cme7Hn43wur1gdR21pjKmfWOPNF
D+XCjlRx34TtvFf/KRX5n5kbgKVHCnYwkqujzlpmOnYtZBZALprPBBsDZ3XWM+3T
ArBbJ8ixgPDiKBKMLbhMjM1n2Q6l0nNGpPizqmVPw0RYVE/70ldYvWUwBNso9OVp
sdcsbWuV8s7pLeuTgGYo8jWjkcavQwVJfXFwWB2G+75geIkykehx2QJgNOsOZS8i
wgcGTpoPCZw3S7QDcj7b3oq0HnhxJ5q5WdWxebPG1ZqH3+IzSRAk4if3y8iAxy2I
FCwE2OAXaC9+MrqXwwji6geKlzXRKsQw5KrWPgVx1YQKLxozOgqa2t+RLKlTxgy0
eFDkXCBAf7Fxw67FFEih/tk1+LfsXqfplGjqRRkMMrWvzSM8wX9WKI54UjmorpmW
108u3myvDRQZDpTKWowxm/2fuBD/O5ttXLYzm5JskPHCh3THe33NENu0ML25X9tZ
+HqMDgDsTXVeXLZZfslbp5LTEIxFchmnxX53WsDmfWLq5wahJUiTTSXrijCNMsyU
w+PHaTLSm0qyYqGPYqDxvIc1EVRk1ErmCB8NB3HDNYVB0BWBhsxAke1PxXOtJPCF
9LN5QjlfxWkwuxpuume4eKcDEPVSPa/RMPGuwi+TogKW0YZ4lJlbPh53Cj3ZYOu0
m5H9opX0AOPML1nMM2khJalSeqXrQZtCBERap2y14EkgBTvx7qtMo/ERBSKyqx9y
w+dA3oDc5djPfdj5TL5lH86/fuzj9hyum5HnvlBijisv3FSE3k22kwZLWtV7yew2
EWt20X3T9VnCHv8GZ6Vq82l0te81EQ4GLJSG1JMmBEU8HkMJPmgkZvQj6UkuoS5t
yeWCDSyNiN+3usNo3XUTn+fZ60j/gGM0pk61iJFz8GBlG7/LzyaZfEgPAxqv1M3G
Cx8hneo2Ord/seJTuhaqIPswHavsUq6+6bZxVpRwkZNvYjp0tu31UpEGYJJoejFF
gODcoLLpI/PglOcVCNk3CYgvuhdnqPBjLMGRl1gEd+fKIZE7XmisE/t1UaUIxh/t
4Mk4Oa/g8SswfGtMGHSZ3aS04MAz9xPrTxVWfIY/gsRgQADqGX0hvIWMDySQqDxv
ZqTH/ubLgkEZPz8gdk++Jku+0p+i1dFfwUzoBggXoMEIPO0/wgSV71TqX42nKkO/
VO1Wav+egoulQYmW8mXV4FBG/I90QITBOro5uFISfOoxLBJHOgqznWEwC4hPORvY
V81QRUcrhOM/JFoMXHmM/8S4YjkZTtjaly2Yrb1UDXUulVhLeg1s2/KyZyXZ1eL9
Er6SYMncZUBFoH0pzYs2EKqnNlgeAg21Gwz9pG2cnOegNl9V7AxlQooBxDJV92of
mZbULXIZ5nZtHis7e5h1EWUF5eTgxlbxTJGZWCUmGi3yT41dnww9AQJbBsoELcLS
spZZrQ43joaIWvMOqrXrNjCccRgcwZ+Kd/1ipHO6/N1kuHhQnEcivfMg14FPRvyc
NvIObDCCvnqkVGTCznaHrq79PhZgC5pzKLWcTnJjR4cWCra2D6E7Fe7yKp2MAI5j
yiTsZ86C1NiguWndwfo7zeEG8t1w3yXJtqgxm7RlRhFXg+StDPytlS5sAEToBvbk
YQIN96I3HwZtVvCqGkTJIjQd7lh38aPtjO+Ppnl0rWyjM6ADQmI1XbuIJLdKyId2
b9tFClGYJz0ln7XS4+K7GIsc2c0KACczUZfNJaVQmLeos7mHsKWu032jt6+w8obe
nEVdR9AyKwO2yteUrXCagXT5p5vD70+MjWc/Jrw8lMnpeS6SxRplHNVv3gqX90R5
FK9urwYDqvVy52rCFCOXfQ6CPggfd5QPTT+vgCajkRY04gF/I193FZyKx08be7bq
TiDuPQnV2/Q63sC6/Sf4QYtDlT9Q96xnr/Tu78owC0lJh27JaNMRtvLJzMDvvxt/
3kxmDUPRVpiLIE/3bZ9GQoV8jo7xadAh0NdxWkpSv+P18vVAh722TuevwJMvAv6s
Xv1bNuhqXzFK08UF7pwxvw==
`pragma protect end_protected

��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���X��f;��on�# ���5"0 �T�PL7T�0����Ǿ*�Յ�'x���!�����*��w���0`>���M�I��M���M�At�YY?��w�/��
��D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F���Dx�hH#5�% �_����|	�}*�s#��A���#N�d��x�+D��D�c�����O��k�Ӽ��;t�6���J�Y,��M�Z��<�CR�p�[?X���Ӱ2w+�D�ˑ@kӻA�f�؅/KU��փ(z�(+ω��8}���Ԝ|���Kj8�Q��P20@�5���"�Т�"*uo�(;��V�~����V<u��#)�Ak�A���)���h��`��ȵ�j��B}�����|��i�O��@�2~��0����X9��3M=��w�z��p�c���sge-��O�,�,� �Iy��H;>���t�
�nL���g�O.�f���۪=��X������8L相�ƫI�"�s1�&��?
��Am�`*3��P�,�Tz=�H�"�_����3�3�x�ZF��4��K72V;�$���t�d�'c�� ���{r}Ǘd�͜� ��BS덴�W /�;��w�:���P�L�oY���a�8�I@p@<�x���!���N��+>�?�<F͔�Z�`0~��"C�����>R6#B�U���_�Jj���,��:��/�-���]P� O�h�	!5I����u.t&y�J�H�3V�b�����x<iK�{M\'VJ��&����\!�j��  ��S�k��`�Ä:-w� �&X|�Ńrs���|�ڍ�f�['�BD��51�JG�E��%�s�z��C��y�	�0K���0,�g�<�&d���>!�hF"�U�*Jo-\���;�BG?�N9+���g�}�Q׾�`�hM�� ?�0��$���à `��8v?�W�)$t��L�"Vl����BvF;�TՐp&� 8�*�y��$�w>����?c�5�AQ�J;�r��z�������d"���j�Z�,��p'�r��$J8�6��G�T?��s��D��N|ɏπ��1�#}g��jƴ]&��b@����3���	��?'\Z�z�a�"�_���A��}�k>v���?��S^�[��r\�8zrC��B?Q#jw���[@���,�v>�M�r���b-��
e~1����ّ9;v���\��Jb��{�b�w ,����kf|���,�̷���B%r��Lͫ����1�j��ؠ��^�;����M�{i�ȳ�u�P�U���>�<ItO�פ�2T`Q�t�>a���NE*�b�7���?u�i%f�!�>���_����C�
ߔ��2S�xp���������5>��:f���slJY�2C�A�Es&��Ao��Jx���+{�=ma�-���Z�r��	g��k��H��y�e��b�k��y�_����>)��~Z� ������ʥ�+t�R>���B�(�-n͓��3����]��gxA$�e 7C36]P�*7��v��{]�&�� i��RD���$�4Y��s�&_���nm� Z�U��[	��n~�h�!a�&��-�ͮ�����Ŭ����ua�����\��e�FuD_x2���lٔw��4;��kmf�;��mK�ݛO͈g���f�#"��۶\s�g8��4�7�}e�!�j�������J_�S]�	�,���e��疸�I��9�m����P<����i�X)��d�o~h�P�+����/r�Js�m2��i��׷ma�<�#���EC�\K���A{�<�uq�u�Q) q�������r%��	���k���PȜ"?�l{�F�TL<�m����[��̺��B���Q��'��a@RR0l]nu�S�Mx9G���O��,majv@��(��_|=L}�����������F���%6��}o���U�	*����d[Ņ�!�b�'����`6Ow��U�`�6VC/�@$
��]ƃN:B&�ۤF�(���lN[������0՜��ܹ�XFM/ ��uBA�e�>�y�3}!��ۯn4��[$�@�Q��"��K�˝i�l�E�s����Ⱦ4��{/��C#9Y�G��ɹ�F<q��	�4�����>����^��,&@«XO"�9G��6�6[mu�}��������+&�@��_��黢��09�Jh��X=t&�Q��q�	&�-�>���
q�X���ʷKU����]�7U�8�́iR@�DU�,��3z����N\v����Q��囂O����'Ӡ�iR����"�+0�P���^��:y {Z	�h�B(z�#��B��Da W�4d����Y�{T�[U�FZ= �A4e��]e�j�V��$��d:�h�/W���O	��'q�K&�z�ї>
؁�?�`Ao�(�:(G��p>w�5�Fhr�z��E����\�W]�:?Z"��Zɭ�����a�r�D�2/9wE��!�ꚬ�.u!��#�7n���(p4���L�͠�j
���saU].r�^����O��Q����S��YSU��B�U%��̸w��z�s,ui�F�<M$
�dL�X��1Wð�<s�#�#�'����B=K2�װn�qN��>LS����1�͢�)���8x�	q��;9���Z�KF�|䱟�I��LO�O�ZV�;���������Y���V�F�=`��tX�Pf����æ���=�u��#N٪&JQ��a>`<.ӋrX%��OX�4v�jKcA� ��f��Y��f-3�C�eq|ƾ��|�ֵ�sA�Nf.�l�tW��u�F�w�-�ߠ�j����L���6�e��&s�>�j��=D]�*��U�U���U��>/��;�oD
��EU	�����Cw�6)۝z)��QW��M{Q2�`���9�2�g�%����ᨸdL����!�i�z�i�1ħI|��"z������*�_�F���/��F>������g�1L0�0�m�9V��j\wQ6����#��.]pE�����Ow����y���j3A��|�3h�c�㔸w�6��:���3f,�,B5R+�;N5��6OH�퇟?mA��?�+�8���.!����p�*m0q�VM߫#��+��*�1R�<
q��HЖZ�˱�*���:V*����py��L��IPF��*Y�Q�)!'�2�륊��y�X��eٮ����� Pi,#���S�:3F�$C�o���>�������,�r����e)��(bPb�*���7;ab��}h��Y]���cJ�IɈ�uis�h���\�8�~.L��7L�(\?b��?$�ذ6o�.�{DJ�Ŵ���7�9O���}�(�"��m'Ա;f����V���.R����T�O���Ғ�5��bE�����N<��0���~�mu{����V�K�^�1��%M���d��!t�(�b*�3L{�����ȗ�8�-�%M�S�Zsrw�5�`��zP��;a��P����t�LYB��.�n�|�9�.���"�m����];��98�;�5���x�S�ƣzX�Q�}2�M��)Ra�P�����d���="���+�w���� X!�#��jPO�r�U�bZ�{� ���0�BG�/ENf��%q嵅�:����B��fF}�p [ي���6�M`ᢆ,3��x5m�nW����"i����lzȈ�8�R|�_g}q�.b��2`D�����^�5H��:��kb-����,���ŵ�L�Ī��m�Lo5 ����ַ��Y.Dzl
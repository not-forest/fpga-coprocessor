// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
M9QRo3vKLXjUctzjs4gcaUj6B3ISyGQIhmVOzTo5Mx+bRIDcl8fOn4WNFQhBsdYVhCI3bnSKvijJ
wUgNjFB2rb4hs64nrmp4xJ+IiVzH3+XgycmYvsmbL5pcbmylyxI9qpiC4orL5rnAG8Xy7zfdsVtH
LZy/WVqsrS08KVTPKQLid7rDeSy0tAU03fLkoMi4kDMYEl9Y4d0piU8eC5fYMKB86fwx55rdkpA+
T9Ylg3MkEVuH6gxaRFI5x4hjDHsigKVBM99KmydoB6b34thAnI4JdskF3RkMihyBIj+8Kh8TnELy
oywDLDyRs3dICMlT7KjLF0Fwqy06xIZOeJjW6A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 48640)
ZdElihRxaH7AOqZ4yCP3yBFJqCHVerYyk4Vpj4tOmdTpbdeu0brFL46orKARLwYlv3+rTtFrSaef
DYyThurpCA8R4hhCzYmLkoZqGdsbA2mg8CkttaEEfcw2HHi/875tGKW2kwjZx+41qXytSGWdFvRW
ixg3kxoUFS6U4i9b5OvhcB0BiqxDIju1kdhhE6ZPsq1zAVoiQDPxm9G6LUDGAV1YBb1BgR24P26C
6nkMSnfHUK6nrYDD3cJ9nKX2t8mlybgV3+VupAEae634yK4AFNRT7CzKfhQ9y7El1Zf4JQSndegn
TVffyXxNJ96wSjAtivEnTvrcKo0qJMw9ZOA6yM8GrAfvpRkpywb+QHs+sy/qhGU44c9iK6C2UdDK
ghGe0gnDCB5TTUNGf2cYUavYJ1L7QDz2+9UXc/fVhoBfqbJWslU9DVWQ3qWhmQjwjfeMHCzyveEX
iZay5PUfQNjJd1YjsQRaVTd0Y/VEgZFODtS3m4JkBeSBTgfbeInBye68VWx2TriwSqbwT2xtczt4
h12E1J125YH7ex5EBaLL2P7JwMbop7bJYJ6dgthLTCm7eZBFiujmxs3cH5tk+4iJyqUUZLEoJrlU
um7Iz0Pwn40WVMmTqFBdKNTsMAQfUBo7psp4lj3fsyuQcAPGZJdafIMUCJ/sT2FA4sxrmPvJlLrx
O5Eu0CdYxEWKJaACY7HQFVJIpTk9gXrbGgPswZvJFQ8eRjJxhubjhjYgP2K9sPrXawt6qzBX7xhI
x1wm5L7yvnEKwI0tqf+dI69XNxA0g8UoHEad20ERvu6PXm/YLOH922OAHg9OABqXidTD/uqtlimc
M4DHNJAxXqvlTJvWvcud5w5bNHiAk95wMA8KyFo/xp5GvJxQv1VpizpCQ1NPKJwWf+KMEnqRkYET
kTS+vg9d7zd/HHNfRFD1DRtQEUwbkrXF7A0KcSSoCeUXDhEtkXsdO/dTELwle3177ovQOb3nWUEH
Coi9N7ftfUhkXGP6b6hyzPmWJHewn1zeIF2F0uq8s0fBl74vfn/hGsVIrnYR3irg973olv+87R+l
O0/w7QWe4Jv7OCukyH4Vi0w9K0dH9SsDTlijD1zP//G8JpqqNPUyJQzUAV9ZUIDo7LNLeWfqiIFB
oh3ZWVCGaeFA4uL1UIlXZffnftHVxMRfeTUs9VhuBdUeuM95KQImDE55iLaYY9QNXgUCrInibI9F
4qSDlWSUiYheW5DBwWaT8V4A+lzqap6d8CfLxZwa2iBzABjOhWrPavvKcmUJl6VfSoOwygS4+4xI
/TJTTzsMgaF4b7yUSLmjl00D6tLCwAcX8tCtNti0dxqXh4cfdo3Arx6d7Zy1LlfYsFr6cC9G9Fgr
DBmS8vDJ722kra34mAtIdApYd/5BoEfOXXc75QVK+5ZqMAk9RCpgW/I1mnrdYRlKfXwK2UHrj8fc
0ONUykjNFtVQUOhrEd6BIV8Dnuyp1vMXXgCcquC0TLFlOWMyDxHXZt0nJwE79+Py3DhwqLu/0VAW
ZJoZy+QVcx1EKcRpXceJ+V73kiHJqpbLn5oc9mc6yYvFeTdvwWQp81kKYPoCRIAK4wY82fYw82bT
yI+GQucYHW/12lMVlsdTTdvltr6uYsUqcBsxnTz61iwGSPEvy59RgU43B/hed3O9jvnbxG6AI5FA
14kfExfBRoNzYvaok72ekAlTImkSqHoGO3IopelLATEElPWHjJmUKxczqoMj67St3RF8RhQn5dus
31npiEPjkO9d96b8PqyH+gzgsLdb8PbshEnl5zUFgoTMeK4fuCtzVECdYVSB811DetX6sTz60BFN
Y3PLw+1DxwcmL08J96f9ls0gTJqm9Nfz2GmHQXfXCndNgR5OkkbZy+WPWCzEmCAA0z4IFQq05l/+
4ZoEb540lJqL6qNieaE1I42sW34G5uFcU5lNPACEAcMPr+D6QhAKGntTlAHNqtGZhc1r68pN3hwC
AclPffqSkw3XLLG2JQHKoJ+xE+rbO1new/xpNMHaWrWRh0/mDxC5zc98gcnwmbMurB596z0aOW1+
f0f1/RQe3DQNZTptLjYdnJ52IJvAwaSjmrNRBN4e3M/UdvWsY/koIlHuZSUQZFPtc5IKHowNURyZ
WtDzATlCyDQm0nxvjk5NkjjLFlRSzJMmqWAPYsctExqYGvvPP10n10aOMK9tEJ31zuSgxmB9wEU2
ohDg2hnjzwmDLShSCGn1+YNgz7ruBWAM4nv1/0phttssCPcfmAcs2yBpC7QCODVxGsDhUsLTYZv8
OTs4Gk9MQ98HeJi5A6l86gZR41MOMtuJ+a3EGDiafjb897r6lcY/FQO6IgrQkCoXvl4k9XgZUggp
qq9YOjFdJZEeoziuT+RhIVJA4ASC0tgyu0Z/4vSU0p4YoyHa8Ac2QaxHHCo9JaUZRm9szD76pVj4
/Ft4bYBAZV7mqEXk3QJ3SveHnlfbEHBRvWfvCk2woproiaU9d8sz4Wb3pLEy3OQpvl+N11oc8+fQ
HUsFcuUFnTTOWPHGDb7VN38Fgdtpp/QolkitHteaCprCjW9INrAMmLKrQHeJaNKMtoxjVXYrksJ2
hCuxwv+WpG28F5TA3nN3ZaS763mR1iaUSc8R1uHjGm+fN8k/JejJI3AsN0n2rWh1XJRhHbSYJCG4
P42ZCjvEjZJk7hZ7q1E7nKO/tRw5HhbP49lIVbmxWumhYO4GJxXiaQDOhU/iDOIB8uY2560eG5j6
AIQnmIbn4Tehnf90jPH2mX2obauwSeLgw6aLnBWIGtH5/uO3NZ05hG2YG4em9s7BKmcj1jgKOoya
UMQpDc7L+sNiIslu9ZXMHRWs8XiASGnhfl/PeQKvaaJIqtTWXaYPsyeecyj7nYtbXTDLsiTgQUUw
9YfaSGE5Vmml31AOnvv6MIoYrOBGMy84J5HiXYmavIPz4NO56IXP/OZTH7UU+LqLzC+hstu/UKfL
Qxe1ZVMTifxle+j82ymrM4NtPL1VkKvQNKFVf8esZ/ClzRNF/BFS3jMgzRjIexHYTCHMUJKyPIb6
PlkgH/DrdCtKEXCSjOoHOsdtFP8OT+RITQhazwQRrtxHxI+4iNxRXWEPZ/ykKj70QSEnMcKiZ47G
kmVnphzoJjRxSefdMMbUyZy/MG4lRGJVj7Nlg0kZrtEKKUbkE3Zc9bBFdKMV+THTovgaTMv+pFcF
Xt8SPZh5o8quDLH/I94A0qCpaYzmAvCNMBk6ucYIb1dN9PyoH7me/UE6QxjXJYa0KrX5zn4ecNia
SS0ri8sk6SdMArrpWyzph+3/IdypRliiROwBXOmfCvX3N0Dl2Qcevn/p8tMRVitEPqsa3toIcwuI
hld0GIq6LCTuwkC3f1qGRxf+atZi3Ss6CAggKgyuVPhIakTo5i4w21CsItbLUvDA3DvFWDFqYI3R
Kbk2bE9Mclb9ocjxEh83R4XPZW2niCvuWiquAmaWYINl4WUOH1INAXLLj+CjKjBBP3tOaBFrwY+r
FLH1QRbzl8vOA37AxX1lKU8vFJ41z1xyC06+GLQEeq1m+2wgMVeR1WTNbBWO/yTR3NIIrVMesqQ0
KkrYi70YDKkYgmosq5AMvLfukxNRTupQb2MGNkMCIgQLaRV7oTwY+Wou9HaOt8qgI6uNP5W4fJle
5fLbYgHRv+4S8/fmLFHVXAY3W6jW0CrXokklK0AbjDn6xZEq73NwtMrdZAjB4S1twNXTuc7aJtcE
futR88ZFpFce3dQr510t+d1Oswv7srPwLDUzipYTIDkBtajm458zpNd/Aq1xI2rKZ3NhVjtOt87v
3JqQW7DS7nreMh+rQlSUOYMtPkFYfUnuhINOT9iNEJimTFHEXKaU13uRR7daYx9gPwkP1HggM6bf
rwzyAHkIFn76Xv6QG0zUDQimmgYofZxYw7swbLU3u4s4tL1JNIzRpZDyo7UrxpZE/bbXsbhDI/7e
wfOTCoH4CUJDSidJYfGXK4h+tC0jH7S7/MXWvG3dFhmsvTYDwlcedu147wKRwo3YZZ5kM24oBJFS
BxfZUcTt+q6CK86pCZPmkMEiFQl6q5mnKClk5EwvZx3C/oRY5VSgIlu1oK5SEQn9iQ5hStWW8+Eo
b9A67c2B1wT9hlXQETqcxLbqJoX8KxpqJg+qJj/m6ZiGiVNaUA/XdVgp73P+Kt5I+W0g+Q7xPamF
UMbK4KC2329wW1AXkAiegcPjVXMLnrg2Jb3ZgHM0LU9Mu/CAMBb5UDWMjZBSnGdCD8UtAZ3GdNnX
Wwf0n1ZcMzcxu16OMkx6KigjlRu8ZHKl0EsRBEUJ/o1l874HlY9n6VabID6xdzhstF9slABdWse9
TDhTJ7AJSc6I8Y3OLKyTaSvw2nMDclP6zYh9X2orXb8LmmOcPD2pkxN9xxAM6XkRx2at5KOV1yhV
2ISwa5ULMN+PqQcrzoaE0BY7W237EbWySCy+90bbzn65/0qFcObe21c0gb6gozLwsMbAbCBPo+fv
IegW4nfZFmpWKxYKw9ozWXRO+1MJ8EnQ+zATkMilQdoz2irgZ/8Pp3g2Eh9BhLqZ5FUHKuG7z75w
7rYlERa3/xoy9pazto4Jnp0TzE8Uqy1Huz4TDlQWzCqGTZAaGMfi5HuruQrras8iRttjqRgkQ4pl
rSR4hESytlijOLynxzkZ32SMkH1vXfEAURW9VBp2P0dw9FtufR43dKt/JbQSjyR4Qug7nenWWsvb
nfy6Dyh/lXC1PH2lOI8EMLtR4ohXVUAwedHu1XRppaFyKH0bkJh0Xh93bT2sGmLjllUdKD/e7edT
02bl1rEPd6Th9kaKIwG9shWqmTUXxyrtiRdV6xETfeijdlsoFvDrTmUPHAA18snFSpS8WKhYI1Jq
g5RcdfsFVYPBkge3BAXr1t5ldyn9S7xB6s9oPhsqs40tReOpck60kJc7pgLiOQTlknXSuO+eXRIM
vU6d4jA87nPUQNZQ0JMnqkEJ9x+R1PCHme6xilsK67vCDnR7xMr48vMOZXwMh3FFAcgPxwUBLViC
E0iMNkajpugeM54co0SJP16REeitXD7Xgn4siFTQMNXAvGEbrVPPWnI9/QbcjMpduMkU8vKhClfm
j1WkhKceiKoQCB683rqVXVQEI7m9Pp8Kyh/OIpH/Rf7KmI7bw5TIuXB9B8EHBAta1pGkNALAaRYH
S7mQ9Pt0vC5qR3ekR4Lq4R1EqRZ30jRAS05nrcX+RCuo2JVmVL1eWCOu8CQkCS7eHLYuGPvYg97V
6doLA8JqVhHt5jXbiYFhM7q9N4gvF34XzqUO61PHQF+HYlxaCq4BXwCZftPvfyTta2mLuGt1ugNG
HZuwwz0AozO3txltEaDsYOR0ZuXTBwYXMafqJXD9yVWnCx1z8DsPiZGeRcQGr/vd8s0NB1h5SuO8
9CmWa8VemP3p+gb2pxu+IChswYE/ZrOZ5Ovcg2VJPzcCDbQzzO5nEC9dKfh6nqLZTr6KuCWvrNQZ
J+9dme+tVjjlNKqsPxN+UvXndR/j0oU6HDtXR02RMYxLGg9pIST4wmmemLkKiBpJOrY/Cb7aja5N
4qqxos5dJHACGa7UuXFyMaz1/SnciQZsGccEvKOlxSO5g3bB015tV6X445wI4b8X97iETyEsHEaS
h47udoiyHxDKDqGjsO62wpCXO+pRO1ZT+4YCpmsLaxFJ/8vK8L6/zj941zlDDD6uqZUl++Cp51gb
NgHehzvSCacqDb6zFlw5E++jwC00mGqUPtk2C2Z8NuopMb7yHImpOR2TyRliJz5LeyQ7aOZTZsoP
O/BCYxJB6zDn9kn2BY+nePJSDqA969RWWu8Fr1Ht11Z57wEHibd3rWblXWQvfYnftSP9Vs6fX2q4
ENLARrZ7oZ79qLRMS4ROI+QOCBZunJ0nPUN1ZzZZxarTqOJsTUOb6g7Lmr3aqNSAOJox74T7itDK
kn90+jUeC3YJAphqumroIrGoTGCGcS95nHV8z2Qh1iADW+KyNlblfLkpUc/FDJCBYx2ONiH9n8i8
qrKSxRLeTgkaxw5jGVRY/CXTS+W0xbM0gdruwUdH8AXxbQktXa4egqIQAkjZtfOvSLz7+L7AHvYc
BnohEvuvBmffFUH2WkfnsbX0a4DsYDL+9v+DC4h/QfB4gWi+xntlu/nXaytuzquoaQSpjGNkHYbd
1yRwda4nJzfiZBJabcLUSEFLDIeXSyNW4ExljCHxggr9WVBlBuvR+t5XcWHzzzUKFnJtlr2pMq6p
utGEMkZbhv8EtWCpyUwRQJrR6Jz+xWXGstI94kuGM7FOPJyqDBjonUVbkGOFy0mxrgNwGNC09oO7
wPMCbAkvNPp8NEC3eKeJ5aa+U/w+HojsA1D4jpBTR+JFQaDMcJBAomNliIjmBx06Kbc7MV17Hqwt
Sz/lMWzjbTHTnfR2Lol0/SuptmO8jKx5Gnjb+WnW0Mw02+Ggs48dp6Hg2GP3BlgF6d0+BsBPV4Ve
FZ8xJxkHMGYy5kjrekMW6ic0K3bE5W2hN8KqmtQVDbKuxDKmXmEn3A8W9L00mQgYy7dv4f3axhsb
2s1ahhCEcLlOmkMgmFT7ZkfHe79Frd5lFO4xWQqUyprvkx47M6oypYfbFnSoK8z8snvw94hdk4Bu
//AwARYLYwtokN2BoyV8ancA5AL0iFjb4uwuICxcSZJfYjANZUG5v69GiD/deOtuew91WibBt1O3
Dl+UL33hcwuyrpTiQBfQOTXcmSrJrUHoSSi/bJJzmAdMKOiVIGIAnjKFQIPCYRqKa1lxk1xYY1BP
2Mv5VrrM3JK2WX2SV2f4Pxtm+4YXsIcbh/WYYDWpIHWBFsS9hPYsS4zzdOT7JhXOsL97+W7z8P0C
lK7S0kRqF+01Fgwh9F4t6is4Ny/f0K7k7uKvhMUwGiUeQ4YYhM7RWXOkzEAuLks2wVW08nVKjwrm
DpQ4QQYIPLGjkbVUvIQeDxeDTFCsz0NgUZeEQqOpIDeEqPhGN3sjcSyBe/EqCL2sHEGwz5hea7EE
DKcfawhMLroVyhs/dcxe0/pEjN9BYHu9eVuH+Nl17oliY0ZH0XlVLSV27w9GhzaDZIiaeWU4bIyf
lE+XBkC+3xF/G5+/gEIRN1g6hgcAxQk1qr4Cdplq+p3mUFMaKsTkLywEaqppVsEnFIgHmswM1xwz
fkgsaoX4x4qMZ3N44IGHpHZTICbef4I6lvk3ruC1k6WFBQTvtYbmlD18twQ+zQgqXdpT3d4qukiQ
7ZNEnUtg7uDqPifIvTdtFbO/LxYKrChX2FSUVoSymfJ6C2uK+VMr//oNHveiyadfp1+qLUAPtUIV
jPKLSIHveGPxyJdfCXDi+iX5uK++1I7vjvjUCckZUuaJ9RT6yJpQsIi8fsEJBWr79mbPhQeT6Evp
DpWfSqTE0Zz/rq+dEDEq9GQFP+FlLzxKs9q1vV3qxRU1X6xdSgmliEepcGCkL8xqHykLuJ1GAmcj
ns+GKeJHSwzd6vtDGr7LOxCZ5Sn+al8jZ5fqFjTpd9jonu3RZIZJ3aopzVk4jgV26vXFGsuwLCDK
iWiYsXgcEC7T0oCNjnupgUpnRyRucFfh1mqr9Nbbpy5JxLhr/l0TA1DMlcvvCRHTgZn41z8VsHxB
2O5JKhkytHrQCY1L4wXkZ9P+KXVWKjAwJxvlkQNlQkCe7HwY9gUwcZhRL+sinYB97oVsDhS5bM7O
do6OlaXVgMAPgCiy7+gMNG4esQfM77fy0CoEAe0L4tBetqi9OLqUI1GEUdNJT0GuZaOewOm7vSzc
d0WEy/f+6+MNnuj+ENAThWjXsOiortIELndgo/Zii1ocVTAZZA6glw0G5ej4qWqBnDVn6Cgau+pH
tBOBc4bWejJtHcrZFszkUzsIgJDMZmNED+SJUZyUEe6ycwmPrY0qAhmk3Uow6eV5g5XA0KXZ/+Te
yNHVgcqQtDbgKLHN29qjsyRD2syPJbTSvltvj8kR/34CYDLqyMgh/1zzXno98mH1a34W0QyfszDz
dUPF+QtwpdomPI6xse9M/Xn+9s8Jioj8YPLjsRSfJuFUXJHP1k2ZXTdww5MRrGTcw4Owae9IyoXf
Y7PfNYfClnZiK1w0gzwwoNK9o9JM+H3bq1Q1LuS34C5yCI0PzZ4FSHV+1u4Eqc/Siu2EDoJ+syYW
O2mxdI0hE/SD/4Z2PyhAiKA2d53cZFn5X3ePh/rdYvdfq336wUIj1EA2Krt7JECZtjawqj518tmp
PJ2VDqogMwY+LMAw7K9bJ4Ut4a7BNUjiGILrpJlJA/221cRiSgclB2poZHrasVmzfEs6TxH39nGm
cIDYJy9K3EPIxt53rNs4gBV0NqBXYuq35iGMiafNSbkmu8GTFWzZ1XVjE80ICjMsSVV7SbwpRrt8
bbvoPqZKQM8+wLbWa5uKSWMc3szgrQLSYhrK+klDfTnm5ywhX3ZjxBWuYMtnwm4w1Lyr9XndLQze
tKbROnxC6ALRZT1OraTg9SjpKxtOtC0UE8s6j3Gk9xeqw2AmsF7q8042Gsjatnuc9kVN3lmV/yst
GUesUksCVDFE14g5Qh+DJisEloaQ9JX3cntll6J6ar1QdPoRrC175f6cLKKmreiT3ZOBMD0r1F1N
jjaGNmzj/hJy8VlmAfq7sEtjPzyWfWM6VqT22Iz3G/o81xCnjIfvUqRHV1P1k7U7Q7Gg5OaIP9km
LyJSCR7uhoj020EZ+PLDObStWoBuQgqRkQJ6zMrTxVM/GdaeAAHYziNAOmvNjjbbfvY57I1Dd80b
wup1uollhxqG8AGkxYzHAMX4HirzUhNTHcYh8aJ94mhnQmsDSqvV+48ChJr3XAoX9OgmnBnXlgP1
xGYnbJoUS2DutvXOxfVjTMYNcsHDCNPO53xWw7F6S8/qD2E3mIiZyR8X3T9ibIypO6fvXIs3z5aY
hlnPcfAL5CISpbZyUoWfY1Q7eP1csa42p0EvT44kPXCABxQCyq1/R1Q8qisgACRiNP9vegGUahLT
D9upZbcfiVlmyl7pq8JbCzLC9pzVOocdEGbanh0nYzhPPwykm9bw0bhTPwbzcDTn1u0jHH9ShwEI
SbhE9tiz9PcYJX+ikLXxRkIZpu0CQZ/a7dAY4DmMhpDRlop1WETyp5VAc9xQgUIlvOMdawJG27Pb
VVC43qufZ6LI1/NbnT1hhbiKkYBTL0uEiTr4iYrSR8o021/ueJxIrETMBj4JymBjR+dZKfN/xcjf
CFaXqqG327MpoeLgMUvHfwsarDVQgxW67bWZSe9tM/9ReLkYl4PYiVevaSwKfR3SM4tSPF1pl9U3
6l9a+2XOhHdurWxZRA6JqQoh1oOooMVJvj8n+GQS4E/E6sTpkYt4NZO+S+xgnxxqxftP0Js+8Kuo
HlmuCYRJcnPI4R0mOEfnIkiNfcZEI9mtSWgm/bP1AQP67LFuh81X2LOXrTri/UsJ5s7dAi8L88dU
vzyvKI9OgfWNgKru6eu3RSiKygdQjpUboH9hi5ogXcukokZiqA3sS3Gq87wgsXoPdkTO+wKfkxXQ
+JTkZqMfGQvUMOjK4jOKqCPOLgUlH50l1kYAqSvU63ADJ0tDPnlvQWRE6wy5xTNfpLinrRa3Xyfv
6UeNPLMeeHdGrqdrPLp2HWwV9IpUnIIDTmwsASCIlAA3V2dyqaJ6M5QRvgvmdcxdik+07jXhxOom
1NmYNWS/DYruyEycPJU+A5JGMniczDwx2Vl1QaIcI4nzo03wUejKzRCcjRn4BMpK6pOef4WX0XSK
+ohi3NNApggEu9tuzCqdAsgDg+W7mfWqU19lBRkJzaoomiuBSkcp1MOt0Ew/ZaEjVIKJNtx2Kges
rSHu2N8BxAZNeJXa423XI96+RuzFv98u2ZSw4rZWEEPe1adE5yeyFiBM9iL97n07rz5PJ4tcMsvj
BoVXH5D/wqYGU+/huL0Ekw5AvSRQyTyDy6L841Gq61VBUL8xc+mkHHNARPH8oYgdNEPHW1hIwkij
wtvZSLZvtLBAzCD8U16PUXSTFFXWyRUM3n/k/rFKQurLka1TTXYNSJ3+rpFaf2TBeCw5eXTzQjwS
FJ3dekBqWHxBpD3a8y99a2wsjLYGZm4QIqxpjbhXVf7rUTzQOho9fwyoEdpEkFF9DjK+lrjz1ZIa
EExJpI80hm5ZlLcVMuF4yCG1HZooJbwTjdoRBX1XA27WqnIX/gMdJYVeCjyJln/PJNZV/8M0rEYK
/nsrQXOxR+nmaHxQ5LTV9ujYqkm0AApV1cFVa7sEfrQGNhOSND4jh8dJSJZAMIACFDl50/SzgZM3
q5xi0F1CzbcFaiudRm/XIk29oT8Th01Hkf2Y/KBxOM+Kn3WS3Yk1jM/HcBss6CPlZvUgUcHeMsr5
bBGzaDxReZcJU8ZDtBUYiM7hF7h5UkkDLyuVnAlRVa0G3Km9twrqh2hE8iweTAM4Axm2y7mcwrap
Bcju2cV2z8zc+Dgb9AAVDzll+8KzWQLoF0I3DCHn6WPOvKLrz1tlWnK23OEj1FDr/jrDvgXxw7R/
AboRbhRFCubCt5ulRZAgwIuETsEYTllnY2+VW4VJthglqYgAHtsKD+J9Gf7R5l+kxXG7dYji4w4E
Lu5tGilQ9sS6UfYdH5HkVQPUepIbRPtqjw0lENNa9dNoy7uhKOpJdBBXK86gfDyVZAj1vm3r/Z/d
iPiWNAq8K6mlXtn9fiT8OBiiOAg2eDBMjx+AGrybPETQaSaNAW1IYG8YNguvCV1WjiC8TrfyhzUI
+wB2JzgURKiZNPtg81i0D31FHyH2+BOmwtpIRahJlvbe/zmphA+uShW7rIa10UI6Mt180L3vspvi
VTxyGXAJeGvFhY76aODLpIoPdNouD/r7VABlBn7aySps+uVDucHwSVcCiqHNDKIoAl+VJHOlmYTv
Ds1vQm1feXWmY4yjRYDgFrIMgEwZ5EgfNAHrXI4K6R1RBas3yrjfoploHcZswg4AExIUwKQvxRih
h+odYcJ+cF+5+jvU1QcLH0uupem4U6h1dKLxpY1kIj4XK//WX2FkxJr3xItY8ohP838BaGT9iUse
a9CH/hFAEB+KSlW9aTBYAdLIkehim+/xVi8H0SfWuuhx5MBYCG+xwdQwWFjHBy9UN0je1LB0x1Fe
iwDfTrG9kkpR4p69wEFY1SrUymEbhaS9JLbHi6TgpKR6hq9AR6MEESKkbsszfwb5GqkC5V3uzuFo
S1+ySO8mwIM6Xf6h/gvpw6uAxd8Cizn8OCdyMIEBuA5MP5fZlmMb1Y5mXGy8m5IaBt4otfrz+5Zs
uHMQFjcTmo07E0JL+ogjg5aYLz/5//cm02StEzfD3uVLpWdRU2McVb47ZFtlhb1M70CsK7TMbZT4
f9bG0/U1RJyfhWmZq6A/Sf3iFJwc2jlGX60dtHEWMqWb9pbXYlmLlsSIYPkSofeSt5sIH9o4O5YU
BBWhrYXW3OEo6RCiZKJerhyYjz0o1P+Bz2ZlxrkAChpHWS5tBNsTaDM1YWJTLnoEzWJ5t7QaZIsR
TE0LIyLahcZXbI7Owa6PyzBqTAhJTNZsJzEVIplRIZaxWghY4nASQH8p6ovj5nKRiY/De/zI0EuZ
n4/u/zzSzYZpsbheUKbqWNi0AHm08RoNBC0uHTRUImFGYxDd464/EbObWe/t/Zgx8MmhM9hVQd/b
y5C78NBiyKHtfAO//pbdcB8nEIwars3W1XnKSqSMcTi6orZM+KBrLYrrP4GtzVBXYSfiYxF2L2e9
KJOPOsTnbiHbHn5e6eOOfaviJnsSs8biqciz7765YBZUc5CmHkgyoKKKtlsNOlllBF6SKOkdFOJG
drqFshGM2xrEfJEqoV1LsvQCpS9on/WOSh1E0UnfY90dK9MIzpZX4eN4Pj3d6JMs/GFpon7y0t1E
v5vRH0BobefjMgvGse6Yn2z1NYWMTO2uSKXYMzLFn12nR8rle6nfHWUN/ccN13kQUKCoSKsKTJtD
v+JqfA8Nl85CYrW/7NLfeQImaY5RX0J5xjg5zUWAnvTIvwaRK9Pt582jV01I7HX5l39G4VnSLWAD
OKjyuDsF0d3CdyddqYM916xhBih1RrR5FioM0+MMBKGV9WAUMzv65ltZ6iOM11Wn47wMP+tn9NLk
l1GpAAQTDW5/eVAwKVQv9BhNEDD/nqR/95K64g57CtL4JQJ/DbRnVhhIW5fbsYjNOwP7AVaIIwwP
KZv02BsOmCd6OG89bQMTk1M5f0slSn/s2bnrRGFGL4yes4cOxukEyDLP4aZlH4/bBMbtSmCwNcOn
vGEcH2TZuuE3V03gB7w++J8I6i0IE2pOEeBVutgGBcuWwSqnuNVVhuD8dv0alKEWYtB5m3QDLzqo
+yOyDjOHNOYCCOsSSeFauClO4afBNcl1aVDtbi6jHFDDuKc83DgNPezJSKScbesAI2eaFCIgCEba
MY8+SUbrk/xLDJzgia7nCMLyIxCgpVlkHpRRjoYpRKC0Bff9+2DesgBHd/u9vOQE6ILdJO6+nKtv
Jjc5SI3wDymMfqkrXQ0Fm86iA8bA+7kqvOi0mUTSX3fhHMrpeXO0IVjamHPLWocYK0lV/+1fms+f
TzaJCjpnq/wQGC605jHk5vvZycM5LxQxjMJFiVorP4wz/gOVCL/pYnoWDOJpA80jViyWN5HLoZan
VApmUIl21LjrGTJbhvovBxHCBFu/WrubidQyT1+AvJ6kRCswjnzjie3rjVQQN+SHGGPdUwwhVLVx
bhXGZUL2Xqq+8ioYw709mr3dxVQiywUOOgFmybUs+i536cZDLDwaKubDVE+gC4U7h+zlUcplHZph
H8AvZC+CiZdl8zh42IffVrBSqvaTWDJqJXttMaIgHJPyL8hLTjVodxoGrHS8KlvkXvSGUSndcTAC
RGsySOrti1zi9YBxih+Z21CC5o6jlGcj8PC1u3DdCeVdt7EFC9eIiMwYgodBbgE6CA8SC3K9vsYC
Iu+18hseZtZA7cTHv1HJcm4rnazf6veNBJ4mb0ENYDeUewPuRX68OOPdmiRlzvMeeiHxbGxFCxey
z4o6FZVedXmFhSTDkVlLJ3dJOP7Ixq9mlR0em+Us4QDGc2ahQLzEp7xU07g1dc4bK7R2W5DVO/TG
GKBOaggbyX9IcKw5Mg3u78n5oLBQMgZNCyKVQTtlXEdpnfesRbFZkqbFtYNq10Zrj3+jeCd0ApUJ
10fKjc2jk9vZ+uoE60uYdcbpdD3/9za36W++cSsrEZj1tlHDybCeJ2SoMhjV3njqmsShWjyVFTcF
yoFlMMyoFcTUxpAYxhlAx/HzeuWBplSGS6ODCvN93/8PR6rDcaxMX9TAE5tcGcToM9tYb09NkUdF
f7JNrocAnZl1ORp0ODFaLHgKh6gZjGGPU6zFogtbHb36CUTtLB0V8eULfh9qHDITmXn9H1pFYm32
67FEPDZJrX+qY5/EvP/B3WFC9qmgvhoqR1Fng2gqNLJYVq4E9t0lMucx5HELzLVrjPOWMMCxqR/l
BQOiEqg3XtACneV8H+2kIWt/XM+VzkRaO4xJhagiRHcwBh310AW9OcyF49D1suuxqRCxr17fycVr
43evSE779nbPZoeSO9lwCzGCztJKFi9SJiEaJTaX8xMdz5XMdDfESsNM5d9Jm7DqeFDEfPIMkD84
Efka3f1E2zLMm1CUlcUsUqzLFpEEgvDBkS7bCz81ngsnfcyKhTWx6t4KCD5JFwEVY8W1D9ZZXgwY
mYRRSJLsza1qmB/moVyADxAYBlP49fT4P6mM8qxuuFayO97MoOmBavdBElpXXYzXV4RNANZReFXn
u6YRuDy8+xP42GbAjB+oC9U2I5Or5p+u2vnm45dGttgr+5aGz3NiChHqGHme5tcWvT/2NioKNt3i
h91LciCkQrin8mOJDmQOc8YIPkjWpfWbNi1fZoQDXaHUWfunIDSZ24fNp4CXTw9Hf7MvzrgnbSdx
flE3aWiMlaFkRpuqpOs5IF935i3pkub+kTVAk7+vV/GR3s7eki7wWFrqH1VwGOpbuuMg3aBAbFTp
M1jJE0xzBbt2knWNlyeJxgN3OyEivu+6ahy2xbh94CBKM0tUOtase2JFoRnFjezXWy8xLhvzQ8cK
hYyHkOBVoVDFQkKxj36vJxShr/DCnekzqbTgzEU9BaRva9ckqRVSk8p4ugChniz4khv+4y4V0BwS
Z6kfE4p+wAV6zRpMsURPESv29Ch6UUxC+Zd6xhEABjtT51CnrMe8x3enqQRuRf9md4uaXXNv84KN
elZSmzQpapSdrj1x1+AYm7Q1+BW1yDiHPgVHjQ8zCPxdRU8MBNlpGoySTIGC5aeKs5YjblmuUKfB
fDVR5igfXcsC/2gS7LZjzt16eciBAzXdjiA+ys8rnMYl1lk1deKTOcTKzMdMMfrh5L5JgWFcCTPL
zbVQiJbGe3hYiSaAUHBEGaY0wf0KfT5FJo3SW2/Ew0WApn095qqJ/yGmQzePuYfphWL5BfS8fWQQ
ltb7wXPwGUd0cRDYkj3rOZS984Ezcd+15g+tGRuNU3W5BkTTXS9LE9j/fOhujljTkvauYpQIg7Mu
WE+ZKQExjEVbzlvJbrXY6rIAcYxa3Ekpj4dTtN/ckZQ8+oVB5MIJcdZJofVG3rb0lW1Kn87hqPJa
WTk4P3gdqNie8SWi9+lGrI4KJDhAyfr0UdUOFr8FbOZ4U9XihH7YqiUayyopWgPmraKPOeo5HFfM
EKvp+jwEX6AcyQZqL55NZ3DWlXVgdPLLWCtCR+7mjkucigC9oZSk+Z4Pl1GlXxmNkRdzrF5M4glA
uYK56Jh7k15MRt82XRK1zXwLlkUgtVf2JaRB+5S1BQtAkD+3JHkZjcKBS8162aGk0ygj7qp4hrtW
xRF6lZBxHL11Jb6J0I85xCKwIvzSlwCaSnCLrXzcftlcBmizZfc7aBWWPvfJy5iUnucQ+/0cVxB9
Cc2z35XIaM5FTanL023ffm/iFVjnt/u4+xJ058pv4JH02CT/5aVNjjjY62Jg6pQb0nmZQiJkzjnG
NgCcdQzFjc3dUlAZSqwH2rl4j21uvDCrmrDHW7Jn2vFLhMD9qZVWZbBN8XepeT8418RhDMpfrfBq
bex6STBceC0Bw/dzZybBqvopDZ8bPfFkUmOXQxf7bwocyOwLAxNrDFF9TcZPG8tTc73+fGI+roet
Xn27dvEe4fFfmPsPBl9VCLZP8enPniTx1ntPLMdQXM9NLAg03PSH6qRrQ1EIsC5A3wqbemZGqrBh
1/l6kDIU3Z0C0I2ax5SlhAH1OWC4RESsZjOM+93drikCy9xj/2o9YAoNIfBDWn/wVR8agl0tEtX1
+1hGi0aM+gxF8OV5MNezL6k6GAFm+aHUllVjRiuyppvWW+z+r65YauGcoPiVr+thsiR4ljobL10y
x2IX6s89v5QwoaCB4171fqS6vVIChmuPiolKV6Naa/x5WFw4ex/cdwh/14eDxH+K2vc8XEpvWMKa
nAFuxWcsKoCM8+UHlF4Sxzqzl18bSigrA7UYmsaCb8You9DetoAQVaJ3XAKe1D8shdlgtRvD5Xkc
0/Nan0LGHTVkL3QXoN5u9FVypOIgd5V4EzcwfV7WrquyWcujtP14vI3r7BrpISsrHGWstTJHKOjL
6LMx7Vmvdv7hPnVjUwPEebdpky6x5assKoO//QSy/OtNOINgH8Uo2HMF5J/s2wHxFMv5RrnU6CIx
1TQu9U9+X3AcShzZZTIGkkYrpqxiJ7/l/uFiF4HGln8Z7x2ipCVf9m4CpwpcPiOY61slFVZBql4a
CvltYfjDxoID7JIwpvb+C6hcPIWlumQrS+3EXHqVC7XK3QazdiwIb7EF3ffaYcK9BPgpYhE3hyqD
o87BTytzJqXDhXRrW0h2rvE62FHSRVYEuGQRvLAEbEFGdEu9QTz57Pw4kVq/lZHPGu0Vat7wLdAX
H9Etaf9WdU6oR8w03Tl+JcHhDLK5B47HAxPwpVqzquBVDZiHgdmSXKxRFAMNW7KQXEq5NS32Q1b+
ypoKHWkL59Cd6YLiVIr4X8xPcpdO5UXSXt5DirDpELqJudWjnrpVYJ3AihfPa4dQUCsZjdpa5uOK
nKTdKoKqyjzRDu1ka1IOjDVqJlnXnFwTEkY2SKrCIn346JXxTyseLYy59L6uKtUWTOuNRtFyf1Dr
MsQMtDEBGl3WKJRnteHYCuAmmlC3jyKldqs0gge1pdMKm3Y+iLj/7sTsynUYHqFS3xvn8iZOT0xu
JCXjqVznRfHX9Z3FgpxL3+UP8Vpcwvf53UPkU7ReawebLO4MBvLdBAvVGY+yqkyukcXgn8LvWAj5
a9EcBBn1zAHSDE5v/o7DHoYVSdTqb0vuDsEO8KC1DErfPetZBn1dEXRydBSZXArocKZCsWWPeoXA
t4bxyZNas9XrqWxhrIuRzVNQ0J1oPbHROwoYboa3k/m/pBoKdIv+crCsD7V62M83Bcdr8dtsQHN0
DFKnXPIMidXC15rtwqyBS6lhOg5e0iyQInp0rIfF3AQYMPQzgMCUi8i8Lfns0VLb5KCuoRfwr2oU
xhGqUVEswVM134vLwiOu8lZ6OP1qKUGBngbRZ8amaU59BGpxbsGPDJNq2xEnBWA1kBm3QkQwGewH
jT7YEmoRC5jpPgmX8DmWPiBqpnANm+qRUWP11GRaDRDqATwOu/knnKbbGQlLG0f1q2UHcKQgoqZ+
S7RU0lu3xXj89MulIPVvsixu72f8SpHpDK8U0E47ulraMA/CtU+ixtGPPzK32NGBWwpFTax4Clbb
j08RliyRtCZ/o854kRhduypwityAcEU3EHOT47746zayIJxQzmbwQnHazvyx3hE+6TDZE1O34KSD
IfcJqaaoB3JxvWM63CJHp4oAoTP3sDQf2u+f1z02abuvtaliC4io4D6JkDr5I30J2bs5iX6aI6tL
uoD3Rd7QJgoG8NJSF6lSH+nWwg4Z6gIkqsctEe9vXhRelJcoJWiTo4+L9/ipY8R6baICNm8xC3Bd
X4O5mQPAafXM/QcgQQ793MCWMqHfqNEqjGXe2l4DE6kWN2U3nIjM4e5uYhTIRvMuY+SsIa12X87o
9/W8zbIX+DAEIXLi+KwOm617bTE3+PtbzJTlxdjDLOxCUE12UHzPaxDEnPhIHI/z0TasGAc4hkQB
Scbk/PGzdYiLY6sdAykn4cDMpveePyx6cOG14Y5zQSm2EO/puxNzZzaPki8WTm7K3qQYD4EKsjhz
3P1tC31Z6ByWE8/spJgGeP03IKrWdNhIBWX/IOKKPcV6Lr/d1tOiSeLvb+/3hQW3avjK1fWz75hT
DlLKLfGgHovAZe5q53Ji0JUMReQK2hu0zwo/+qNJi+22MPMitZXH2ZD6SXIIg+yKuBNAP9y2eo+s
zDPiD7u9sY4nXC7yF1sTbFhqElfnLG/s8ftLE2Hl1mvm7DqMSp/4eD4WWtGTmVOQmtIlJHfcH2QM
G8m5fdQ43bnkb6Y8OthbsKye0RD4tkP5xL5uM4pZTyxvFQJMKzPwQWlLMyGmpLRsCXBEIen8B0vf
wMgzGuCUq1v4BJaDCnXST9PQ+AKwNy1S4AVRHLwR0wQcXOncAF/OltClDHIRP4E737DyGY0Nj7eb
MygzmyCTZO0AXRTj52JTl6kUSHQpe4PZnlslnsqu/kfcl7sK4X7uvcYKSJ7bOCyH0NLRprhLhrxj
wGdpAWE/Gx01bMVgGasUuGl91rskOWxrDa99RkKP1T80jSaLoArkZNeqjRbEo5iQrsJWGsZGkETl
ZIo3jTSsVaKe+rNlDgDsdwR/6EwUJsrLkB93w8uhJZI0Yc6B/hBK/7P4Q9HDUkTiYAbelJpU2KhM
Se5Wur3OEkTPewKJ3MoNgCWHqfMbxON+/CHT2oPmBbHEbe8OWScQOLPVd5zSOuNzetUeuxmI/tvF
OdaPaY7BmLvs854p+ayiWWx4yBrpNcpIGobgr7VDvPUAzJIEFDR6O+9aQ5KSzTtMCSlKt9/ksXwI
C1oukYPvpeAud+Zdt/IppJv3MeAbFOxxvVSzrj/kBvS1qfxKkOLftDTa5AWxDAES4RZkO6GCVdqc
7E/OGptlJivF6mWESB3XIRhMQsxysFPe616sd+uHNrJgkZ+S1rXSWoKd0VXnTshMv+ebgZ1px64i
41W3sZzfVn3J6atw/Vf6oetzTFaFmBVgjKapzGmnKznnHxxrXM8KKdWv5/tMSxaHnQPp8lFMjuJX
W6/Gldw0pmbkKwdadiMv/q3w3XHGiR/hcEOVSeoEkUeqe90Rpf7HwyQqNY/R/eqnh4hgr+gBlYpm
thcpm7MZFWNcJqFzieqfWKsweHuRgbNVexZaO3oOcHEinTDGcO07dK8SzBTdvXoxW/Wkpg1vzZz+
gRxg2/uzrzEJpnzayP4ryDa/D7MHKE/FZHTAhHV+QaeywksblZsxFHjwg1d1KwDIOEooNI1vQsci
+GkPaKnhY6GNvGsEKeOPqfLU3khLIK7EMVOQX0qoOR0QlLKiMignXqJwV1LElh6wnorWaILoI1ZU
e+XkaBPa/YGKoUD089uyltA70nG7nsBfElRKXuKVbYkHVA+D2ojRXcOQu1LfjDhc8Dpalj4ngbQ+
c/rZCv3JORubY7koWgbFHBTBY/RMjW4KjqgevYsHbyrqRs7O/Lo2CTQfloXNQ52DIZ5qrRFdHgv4
ipyvMDyh2uH5H1LXKeScXEp1gHQCNCDab1hOsHwGUVuyXjAKUmopkyVPmfo0c0+mjG8OdS8RmDPq
q87lFuDTBt+2Z7eQLeAqO4p6qLFb4N7+01P4BWzfcAZD099/8ZoPpofbJMq70q3LHLpL3MgXuw+0
SYV4PHj7AgmO0Q9ODjK1CXnSSxBUN2RVHA22TA6XwFoyhRtVkuCl+JZuVQo41bLuLqmaPvmqqvxw
Jibqo7UUwO50yt0Je3JDpYk3mp5FsFPY0j2zL0Qf9pFU4pAHMGjyYLJxf3FZrQErvom6LQYbdZuB
BG9laVsuoicCUgQUInj2qk00m0IVJA9eEMaajMU/oezgc1SPHCp4Fsx6jdEXdKfedWIzb917ukj0
UUjY0vdsFtPvBl9hik08YnkAT/GQ2L6E8lVPsBFS9r9zyRMb76lFh8yIdSqpctp9VR13yIjNLNDK
BZroMA/m+HEeyL4SkRHPkQbbWkKkR8wX48cwsNqgcCA1oSAhFB/O7Xyf8eaRu27OG0x5jtEBd54m
HgT+2lUPI/28+M2mXXxFbkjTw5x1LNJz9E2hO4jGg9BE8GtvPXSORxs6T80EzNbLBZXgTavlygxF
DQOdY9HEJZtEodjpScDm3aLIHD/fLIU0xlmKL8fcq3q2KMSYlvmu36zNuaXp+byy74QIXy2iKCvp
kqP+7fZ1KHficWus3bLfcutucVXZoJf3aOQSQfFDrQXJQQVj6iR7Ue7pPeJW6d65apEnorHHoqQ/
KIOT7vdd60+WTulHXZeKmSb8vsT3WGm0NmKSLD1OszyQQDgvY4hbvyG43U2XhFyVgH0CakNG1001
/BozZIljBW9vxoYbpoNpeMLK+/choJmirK0NfoDXc4TT5dnhaFKsoXkyo1me67vQM+JtPKY4sI2v
hz2eWj0no6vX6C66fVTAsMGIc/1PWCfmUsfd1OLJR9MVGoDDsvrftdSGzgJNDc7K9igGsDXALnUZ
Qn+5gnJkE004udTpO6sFidijO7n+6RWSU7HaBI6vHWiJxJGBT5HyCFxDi2tU4JhN0GpHJmRO0F5/
MpB3wag4SKpvq4SMgBGxXRLwtVCJR1lOiffMh3zbWggp680pYJFySvOIIi6BY63aHEq8QJD5q/7w
+tMG5saOafxAnAtsWZZ9NmdH5wrUtxbmCTszrg3aNLZkNcL1mYIBaXo5I7TUi9SXMw248ZjorEpI
cKHYOiD+gPVQm9CWscjS5tsw+X/XfM22abEUP5oJhS8iwR4mcAgF/yi2/4u1hH3kbJSRKQG3ZFa1
MPR6CaYtZvw/YWtKvB9ApmnyUvy66JbmlcfzWVGU5lMLRqhrZjmUL1sUdIBeHL8Y58A2YjAT9jmj
jIcHorbytdy/614oS5PwRYOvqDJXaYVQiykQxNlPPu5F8EsW67WawYuf56/nFUbkCqYMiKFYvqyi
VIrTK3WHCQjbbJvDxnq2td9rFECYxaM3b87Y1JNwXyVkQIWR1SNslT14a3R4szAsiIIKOEgpfXia
tUHydDAPEnAQjpBp75JtplvfQ2dcG2nc7UYXbW3ZI159avjoygLJK5lJIVedwa5OaczWkUOq1DIa
yKHme546y/LjfQ8aGHotnTEmfBPmfC7BY2RdsypX8+TJvyQBVhOV4ceBz5l5OGl6JJstBwDhid30
pfdgvksZkO0OPPMjOMg6viBPM3I0G5ipTCzidCHG26oWTZ/WPD+PGlQlwCu2j5ksf4zvpSHkR466
v/3HVyudm9W+DgPleE+alSM3u9ZBovJ11y/NvkhHzkf9K21cmAj12rSvebh21QVWkxLELS1eNK5s
tLXi/MWY5ZicrZcXtskyRYQcj9BbOlxbRyUGxUmi/FWtyR3AMx5pUHWBrPSKe1vgEY+wiOPpIs96
bOuo0dZ+NysuvNKucm2vOJgxPIcEwz5y9TH2+5buEdYG1x5JWXF/xvhTiGOUYlWaD2/tr//NM2lm
UWj7a4WoWpUZ62b3KZniVG9R8h+CTf1aPueVbs4Em0e7qYmZVH796fRiOSRCeIvi9EWL+xvjtrZl
cn7gErrOrvYcdowbkaIr2Hlv+BXQavEhmUefCnLUtFqU51HT2Kpqlv5i5tIycThAGguEGHte+K0L
nV8YRgVDkzZfSzPxUFM8g1Q5eyyCVJRSeB+Zrv5llmiyNdz8EfJC0XwATGDXfGH6vnFEzvABabF8
XQqRlTsXZ2LfFRXNpo19zUV0fHY6ib9UsJvkjKMLTi1Wa7ZbU2HqeC+9iDCBFDwmjFxDsJi4cv9e
0qsluFyiDqhDSjPRzkGXSRUW6GgoMiskIN1VMdafXvcqhqjgs2ImO8rLw4Su5DQSJ+kmsbODdGUc
fDR/SehExOe+an6oT0E0sVXqQtchqooLx4c4PlPaCgJoHodX3NqJxsKt4yR4ZD6He9MzJ8v7SlbL
gzSRZi98M9NTOoUL9PPDE4MpzneJiJe0o2zNjoMahtmem44ZER2Y9gCY182FuPueq5VdCEXjTttY
GlAGPeTfqyQUE4WZRMN5Ldvivj/YwgaHabULGF8jdrBXjsBceFcoxhOKsScqFPfc+gE0QKSz8sA7
cjsZIan/tc7Sa/zuBAy4rg2vuXFJ4ycFD876fUC2m5kyRnIQTChyfY2b9Ddxa2M3VoFaSm+DaQnG
LwOdZJkrqQfqaNRDLST5yLwsUGxNQcgfHbRHhLzpIvkui28GGel18YDxpCGDmWcyILouklWnrg/W
4WFGU081zxSxEauHbC48z6bnNFl9+ZbFOqiBkELRzEmPevDtgl+4m4sjO+nEwKQNK8aLWG7zNObL
PsoTlUXmzRcbTzE5N80CKFjQrkRtHE0MuEnY+qgwfwgX+P5NdSl+ygUde9Xcniy5QeAZ5sOVli2f
uwqVzrOoserZhEDOro5G2U39WUEnqtC6QDwPiGueeNgL2g25oxYWh/Prn4P+pISEesO9k9+3rsby
A9aj2DtBqREx+soz+1boGfLOqopysAAlMwNKgLzbWRygeO2bQbGwh8o3EjOQz9Be8brvGg6Dq11u
Nzn1mIrCveAiW7UDFS/BDBLOJzmOqrLUOx20vDHIxU0otGi31seI1Vdi3wWWpwARzm5BHCKnIEEu
QgSwQ8AfcNootr/JygJbYjh8h0OelIoeRuQxmSn1FF7GGNVO95prDcmKZPztJxedS0k9mXRrY6RP
HfAwVaAQcH2waVix6odyNIsw+G4YTN/VLKqYd06JASbEck/z6Q/xnr2jXlIbCq0U/mBQ4aF6BauW
6cilqZuTyQwc7b1woyVhMP0loCB1/XeiKtVEqa31TczSA1FdWKgluhL34RtuoJ/acgg6c4CoHsON
TkZ4iQTZqWsOEsVN57Pekd000cnTI1hEMHSbtR4K6aLAAh3JmTZGwmll80fJdiOzq9KUPaHV51Ms
8pCnJOjDBe/7IHcCh+ZiQm/8fEDLRlBrHpsIki5UjiMWkOlJqaah9Ivi520UFqecfpg1FZzYo3nK
HcFF4IDd5WzztTI4gp4+GHF+AbBCQfHbeptBEH+m5Yo9QENI30p0tcmY7wUHqbkvZibAwNYoCF4n
5CwTQW0uEFNDL22n7fIJgOFHT7xC6tKXMxisEeBozlWAUrMb4roE5TQrVUQGagsb22BoTlWaWsHY
u9RzXVaK94NuV1R7e357OvHq355q9RwvBnCLsHsZdUxjQL/tB0W/MB/XogET2CXD8TJ9NcOXGb/F
OWC/f4WYMj/679sYZQe8mKMjB0UzDn1iqQTWaHwhLK1uP/cp+DKVJqhitvjjVDiCFdTk7+TUBRIy
CYrTxfeZKBi3SNAn3ThVlvbpZv81DXjF+WeNpUdzXSXYCy6b6vR+JLW1XnL7JOtIuZwQ8SQpFVWG
ffWQET7cCAOGJUc32dF/JIevweEOe6CU+yI6ykkDvhnJUICAN4Ug8y7fZdWqw4FG9YvEQVD2XKn6
LHkH0XYpKzrbM1gbwGRPG401Kggcv5AlSe/4UTlnCsTDM8zfw4KsuQbP1A1Wbxc90SIxZyzI5RBp
ICFq0+Y9qWigL1EFWkfvRCaaLbSEf6VvXtPvxVG2XM790l8Olb6jYCaK4Pm4BCc4ESM3Fr97DO0v
GGPHJG18Ut4XynIangfZmjATJG3hRdxtQGPM1vQ2sYdKPXGW2li4aqOYmr93DAX9nMQGdccR12oZ
jTplUzSb16Rt6HK/ktavX+2/B1cf0Qhrn88OT/b+BSoJ1iuQr70qBDr/20Fw+XZ6PhkSyifX3vw7
Ysj+YP5SkSVfAt2XvfHbd4YyshkwBqFfOcx+ejxlk5CoiL2rCVQbX+58igZEHn04MZpNQ4XjV+bL
RCLVd+X8XXKNfMGtQAb7V0/lnjI3dzPAC+ek7vZ8egcnAwdg0Z5Fn4Ow1OE1MGyqFT3labTIcMGm
+QfuveONi6NEjA/94nSx/C+jzJyA4vr6iX+m3JciIjukw8TjW+DYFQnYoYreMd2FvGDtci4OcDQg
fNrGmwYT+l5dX6iaikgV3HBlPcHu9CRvpGsRMKy3Px0XzxVyN5ukCrLJlsdxRelh9w6dFBAqpM/M
ZXNWpTgzprpMw4zc67ZXfhnxj+PGt7uCvCXp46GCpjDKWfm8/PBwdAuFbQ7jHZXjKFcK0QQxbvxh
dSOGs5amELWcY1FyxtH+2EH6c4Yug0HUUk63L73RNRJ5O/yxY1FeFMLO2AX7I+FLYJIlIEV2Jg7k
nPA9t9Yv7wtt3iJY0dp5I7TWbM4CU2MJdajISmCCk8RY0+sEEKLFlfQgtXlzMK/8hxjpUEzbldMU
l/YBqShEDeWEppVzbf9KIOtLaR4ApeB7PaURvcOEUNMl13bnw+BOUNxbKcOS2b94m2uwzA18Ge0U
HavXMNznybovO1hF7d9cECQQXKRdjPSomjL+HwU8QTKtcEzojCP80687zf3SA2FOY6PPJjvxd9eh
cCf8rtRH2hzWeYM+KwltmWJHVU+AOK8kxzuRBbhTfpZ4wlgU1oKOFSBvGSlfbuHNyH4xSnLJuHSt
JnUOTnnPKsV4yezQd2IFc7r05+NQE/rDMA7PYSqhO46vwIZYUWJHsGKTnonMwqKGldk8mk7FUCdm
lMLb+k8wbIVfaU2BR/RzXQWb8QS3SBdR8/6EVmA+I3c32wuJjax5JBNg3OroT80DZz9P4MzZW9gD
NC2Ga1MwbPsaxuzDkFFyRyiJp56wZcDrTxxkaQx84u+9Yan3OKX9z9FklHsaBm0NZI5M/MSWEzOA
wKecLx9TmxBXiYw0NDr5I4yWYO202kAaBH+udmeXntMlDBBpt+3MgQByWsvmeBQhgAHxRv+l3WuD
YeoNo19GrRtCCPAv7K5qXKfXPrxSWb4OZ9oNgAsKxJYgBqrgSbkq3L/7pkQCWA+JkXSBiafwg7O5
WNvIPiNogFQijJ7GcF2rFjF5lnXFC5b/jUgAm1oyIxXZkuenpYRjMMMZMABIXu3qoi4urK7bSXeS
nLEnvCTN4I4BUTTkxfUfQvw7YwXpbAta6ENsl9m2cEyqQ7Uc4rDLCV2ZHrCfUL6ZQ1mHHFs0KEw3
sl8Du9fe8e/hsIVquDcEGdXk90azARu9NB/YLRa+45cwfI0ttwSvlPz79dTwg6MlEmDM4QapXWs6
m+v3X0FhunKCk74MlChn8hPz5PiIGuDrgtUf9AmI5zFq2sOXHcYWbwDMNaHAkHABXc8QazwCbZmv
7Ip4LphSRx6vKi1C7aG1HRMUWTlPifiMwsIN3efOnSn+W+tT0ljWWw/xQDtwl1lUQgsqNDB6Ln6x
fwoBPOxsJ787Rs2y9SLGxUwbBLe4KvMVBsotNEUC7X8Eobl4qTUVaMGliCazWgRunHYvmqOwxaD+
aoH4r9xHK6HPM2IFWrecB+nu8HCOUgjWjkRTUfIWfcZJ7f39ydTyVE8Ct3+NGzKviUi21sJqO2gz
WlWix1Ei7MqkZtD08nqkupKLNDb/joZ4v1h473+6yMlVIz5TCRp5pb8dW5ODUCoY2ciKbW6/bldA
vQWZgoctM9/GlzxeIf8nzdyYD+gnbJzO7MhYfKtWAPQZBSf4TDgcX5o1icFjW/HDj4SbuSePFntR
joMMBW5TLt/rTREyUl44/ubKKIX1sI7Bx25A59tgwJPN4p1Od3O+0WnoHN6sX0WCrcmmPUPIhHrV
F2l8m331AVdIGf5YMexHY2WgoXqjuOjqLVdV8NP7+hibCxWq05Yvpsd9yQ8vGQc0ntauhzxzEx6B
CzPi/o4I194GXThJEDBvBVd1QKaRoODx0OoQgwkr7VOfadr8YOHt1TAuc3DAH9f3MqE2xc0NH2PY
/1ygIZM8gUie435kl5A/iY809vdC1Tx2wSZQTAlogAar2mxphYM8WSa0A4eM5elSpM3rO3kQUuZT
BIp4nKrNZl1WER0A5lGJPs6E0pICgXAAe/Nlb4FfWWN5szCnlkwsuKtFs0uIfaRyv9GxvnQzfYMb
G2qROsrZDAG/PzOPwRK5UzZ8HwNyHbASBAh0uVefchrews22g2peUThYC/BC62ukGyhUetuO+3A3
WPCNMrIJRTzpWO/RIUAsQRZuWRLJpW/LoStYpcJi8nYfly6NCvKfpLZYfZAscCtbWFLoZGqdH4kf
GIQZXsI2N9XmY3zl4N45qifyFoBiec5qJy24/VAuB3Inlfif9v+49N5/PkM/QLASW9PSfmWAxXsb
8XH9PMUE7dBdUkhre3OJfpH8BlcOUAqqYo0cnlRI33DtIzt1nT5ZBCCoJ5s56n0OrXO1y0CHOvcN
RcPihvc+BQgoPoPGEu+YUW80VmidQb8JyMkTAxoU/jP8PWyeiHzffIaeSdaiYp0AKdx6WmiFw8nw
lcg4yo3SqZ6uFv9YpBPdQW1j85DO/yaDjjghWD91HmZCAMFAkH9wsQ9fTKk6otpoYV4Qv00rerAq
yq6b23Vno7+j8AIUnZI7sa1h0recbIJCX4Kr6hhusXemZIXfepiSrL12NKMSi6yI5ur6VLdoZqXw
ADgxoTRJ+aSGpumVPj6S8hMUW/GnMIHYza3t5zm1wVHnXchm/hH/9a6sjQM5rBmh+szmdrA+q32R
yj6m/odjpYvjfto0p0FRIx6rCLbTtMT5P0Q6shqQU8dOOEd/BogQqOKFdn/800mAPGWl0PeX0PCC
SpC1X5/Q2eTD05YXhWmOyctQqx3liX7QSJzESo1z/hXVGBkWcYZjwGEozZf1kNfKxPh3SeZ30ZrO
m3rnUJDZm66lxhEI72vOzD0J9bRPV6YHOI162ARzRH+A1Ksd8HItTK1ojALQd1XBWLO/Ij3nRf52
HdBJzroNW2HdyBhsEe47vVFKiLv5MYPt9E5I3YUWDXHYfhlHt11iOyg1S1l0c3Fox5eCcaRsFTfE
ugthiCd1jE8hkhUHIwZqKZ0/8F+Np1tnwExIJpbGO8MNdvfTcUA3PCYt1j5esviBgLcMCXYPn4Eb
tLawE/ALiqtCZK/AAmPg/FMMI7GSu612Q5iOS6uloAFdgy8AKkprwnB4T968I2GaUkw66tW/kTCE
sQh0Qu0XM0P66iR2isfS865Uu6xJnXSeB5yfOu63VrNHc+iBoMaCcALzXRUbovWthso6GYa/ZP72
zl8fstSf87GDc4SB/Jtsusc1yw9CnjXHYAIAmHmQC8sigQ8+OmOrT3+6sjgBZdtMCOWs6z+hhEvN
P6yLkqWqr11n6mFDF04jAfyByavk1/QHKAyHTTsFiXw9lvFNmL8z2BR0F0VlzsNXjQJ7P5hF4XG1
J6zqpmJ9dHkpk0kEApckWhZPsUz5TP9wEIrN+n0dzWTS3G9XzNjJUsXkQ18Jl1xTvrrrIDHky901
e+5ziO3fZxMOnizF8K8zPWA4Ac/9McUJd9hqKsLxPrZ3Cb3Y+I9lXDwAEOJg6mk7MCQm5de6WtF0
IPAG6CK4jfOBQY3tt1Z/b1aVLAUvq7pq7Uwe73b1jmKwBb74wgSc+iSyhX5TxLUO5sJ16SbvqZLC
CwI262XC/CmkISakoU/XDXVhUvOaqx7rgtay49U/HROInH+J5YBBwgo3dqXWYMlwYK43szpxBFgh
ZWLxqFsMQqTuKD34v95mlNj8WeNHEAvz/5piPcUr8sGImi8w0jGtTo8dNCvlatJHlppmde7p1MMq
/7he2riJkwL7xqSppe1ZpdUMCDD0yk5CuUgKhypLxAe4QVpY72LaVpwoccYdUipmqKh+qPIYiGxe
wXWmtJWlQ4Qnmb7jc54ePUi/iU8qD89/6C79J6Jw4Tg7LPwK16R/ACynplOKc0DFxKigXSmuGv9H
VyixE9KVdtlPC7iyG5g/lWUZ81gy/RLiPtzVaoGeol2nnc2EG6MXYXySxMQA2koNNoj+HKip2L+B
JUiUeJnBXZfJxbTHRKW7Jm9q6T05i/IafTlpYq/re3iPZYNfUfklFZSWAs0AVAro7QhxneR1fQDM
Re9F5AV1rIWyJP1daJS5LhK92IhhRYyMOSHkZkBz+D4riHP3vsy7QAjXcmQnI1j2CWsUG46ZC5Kh
tl3NQh5gTfUsW387QbC/WbOD61BR3KVBpDl2ArgoyQaWoMfgmqMYiWJOaUdKzQbWhuLUwfBtXdgc
i8bsoPtSbDRl77BxhGjXRsylg2hmnzIXW1FLiTrXOPvHAkO7Kfc1E49Q84H6cIFFTaewuZnZIpIt
wcuPXVpebjWYDktZi+Kysfh5MfRRqa4oIOKCbJpYhhq4EjhvWr2yiU4WdTeb1gRX6rnG7R/5msYk
hGitVXEXLdGAf7lBuoN6uNxxWNU61NWhOSnAoUZ1g20Q+sxtqv/MYDTpMww7YqfBb6hZ53Rm4YEo
7A0DLgoS6H3OTxbCP9RPGXRNwfGEgF2shg13KWNuECKUsByyZJTiFnb2jbMzXzdiYa3ui5imP+I7
yX/02l8qM/vYt/2lsyGgokA3KtizaX8n2PmCuPRxqq9bHHl8j4jlcdOjSiLqtST38fbPPvN1uOfW
5w26hjCyBASZk8C3zMnBWp16b9qvgUeD75DynlCXfHl9B9/IefG1C/8n4Ra/uFWBVzZbVQzId/9x
pXZ5z7BvkWfWJ39zvIm+cdKr3Jmaq368hl3jpIcMxGlObJ3lAjXCkOkWoXuo50fWz7Wc/k/Haehp
K3kpXF4Le1cDuSykKHVergcLM0qXHxS/zQaS/jA1600LW1tCLcGtLwHzRdLq+bJhikCvwj592T7g
qtjp1nGLlKtNGQrzS8G49HJxWoVhjOWAgkHvcmpsptuPxkICH9XOAOM9/XX4eWuY+QW00ksSQZbd
Ex8qsd7TdW7PNd/YyK2q/XVQqii4BFROO9lo4vyd9VxW1A9tBfQfjMCTrTnb2E/A6crG1YhylgPK
M3PS1O/XWlj0dsX5M4AmbkVLsX+v1V0zmVaz4a5T7VsMrFtrz/DRipTDuZhyCsNeFtxl2gED3oep
yEB4MfbdVSGnmKl4aoQWlFZ6r7XFENfgOfv5Mxe7GQYt/wulWVS6Nb/Bg9ksb6OR/WZmtwbaT0Na
c+dhOntxwjEeS7kc9oK/oJO9n1cyp/yOKGzx8sU2MJ9kz+s4Kl4LSSNNOd3ESzRCl4zPb7MCBITZ
s1iv5uMo65u+VSPVdRe/f1cLVjaCEAvbf/7K5gropCwkvLSxFI0htu4bI7Y4LmeylwAXVV+Dz81f
hj/vL0T1VMKc/ZwZbA3ccNLBPonpWcH8RosaJqm0ZzO+TQUaU3WSe2d9cVaLenPdQqZK4xKtxUxD
cyb9g06SfVrVFU2M/4fVFq+TOXkD6rPHxdeToIjSaAE3Ny/+Ye8M6aOOZ5L87elHSCiI8Kvi+J0L
wiODveqFdvy4yJ8EnzU/ZHYxC1LHUPeDfq7LuU3RRKZv9eViwPlr7PCioTgZEYIovQ9k6Ah3bif0
ZYU6dhJfTGTPhYN4vWLKP5NjcavDH0t/i3wg4BT7AZwDw9RKfkPryowpaXzJ3X4mcfheTsOhQuys
/r9az4RxK2s1/b3R4lvV0lpfm/2EvmlwMRajsL1zkTNnVLgOl4ki4w3TIBR0acglxULZrYwX5gkm
o0RCvALPq/jIxH53LiceelyTcEItaudKw1Lo7MhSTjjuTuNdEQ7HEbzfrOFhbHJvOn1UcYprk4FA
oN499F2wd8I4pqlJbHsRJoyFPW2I3H0JJzSx0eUwmHon396ogMfbRGtZqp74LiOhpcDLAN57Pg/z
4GRgM0hLHt1nsez/a7FFWa1CBQP19eKW6BJOYTg7SBcoRcvjVWnB1QD2+4NiFUdLl5aukWu4G9eb
4Zp7OflZD2Ww/4/QpUcEnDQ8V1EsbQ8v9jyc6nWGlgtLitaEHwsW9Wbi0QVBpHRjTRHHhfCuoDEc
RBdvlOCoe8EoOsLNKY+UV4CTzC1HEXaTDenOWgPxq68VuwJjWFsk5c2FYQaRP3X7zqcazmgNEALi
gufPn+0NX02y6BzlbCl1kRMFXhOxvPa23kbuvKvFH+kuejtqgIEZD9ISYqDdE0bKCNe6aFzSXGql
aS+5ajnZU9ir4gF/YanGh7e6n50OuLbFC/Ty0tWaHJw+RiNjTv2qGwO9FF9XcgRZoClJkVhrMiCs
zQTR9wYeIGSgB6ITbCRKPjUMsaq9ELNnvo3VhmoMPn3lr0HciHIZhZNGhhSP4jgJowwpzyIsVXs3
q/LKXx8RHj2M/M2UV+V3f31hAtbkC7YaI5OQ+ho0d2fhksjTG9K78afrn0MnIS4xzYtT53UEvI7e
rPYAcC6zhzFAwMdgJYbQReHIbl6MMfpFLCPXy7e+yGBiMzPyMw29Wc8E4ROi1de6lYu1qwvcUdK0
HE+HfDjDflVDifL5FoPipITz6n84cJmXpP16A/gB47NC1H4emDBMYRiyzlG1Hum1XNgXFFWUHeHG
OGWuEyxFNEtnckbbnDrrrpGEEgvaPCS/uvRbo0sF9kVBYA6lDTdmtvxoDuLIBFzs2BTDTFcaurBh
xzlqpQ3b+mTuEV0Kk4pkzKl0/OpKPF7vRGqNsnI/99HPRxyQKVBsuk5qnoykT1v4Y2o556jNLH00
CKBGIWD4uL6XqLPUo0Xsnot7Vfk/2rvNTFPeaJfOZ9kdm0tfBGKBD8tpaILrwMfMooC0UAms3Zte
23wS1mwCPlVmjnUxQYqOCWhxKLLkmn8Lsfbp2w54SZrpHl4M9LC5O26T4Emv5fo19wLS1SQlPAsU
M9dzKfPSiR674Cp8gVcDvGXFrAB8as9oSz6r7xIN+sAvV5Lw5TITVS3laEo5ahrVEvXGahZuKRMO
ZjtewMZu0WXqHcE1jLqp+C6jsmSV8T+EOBgarjG6qm+F0meoIeTOmJaoZMfQ4H8/OzxaY1L3nSkJ
opd/r2kH1rA2F8aohFVqU1aoy8jQLzLHau8WkBv54jwP1kZcNPDHKLYWwCKP3e1+jamhkVoQiDd5
spl+4inp152DA5zCnfx1m4WnEkwE7xkLqCq1HDiFVA6aEFuBp4sie/QJMrwInxdlxHh/Lk9cKu4n
nwoB9KpoirP7nKWQhBp3dmpwVB7aFRqXwr4rfM79GBPrbCg9bOjbE5nH4QHtdIflTq5zXNiYK9i4
coCoh8u71NMn1x6/fhI46R6MoCbLOh0RnIZD4O8bkx5Lkd0Ho2cVbLFUSZQ/Qj53Jab4UiaOyR5A
NG7uw05zRWaeEcnfPJ3pWi5FhbBpq+F8cJO0DAgWZnaDNpJWNwVLrX1ENYUJBH/z6KKWzQBAEceq
wL59hi2jtC4WRzCO/p8ASyqeHEhzcchtLUQ3DvWi+e/MGHhw4+cT+uqSDNX+0F6mxhAYoTMAXk3/
Xv1cY3BRCT/+aPnTgBvegq83aqXNgIEyT5jxof/LjsI1bopeJ3ygbFNbJjJ+S0+krCoBpUA7y3T9
1N6IeV/NLz4Z7+c57FzJVOl9O3H5axf38UIW32/bhmHPTcjOI/r1HLBICul5keod+WKtSwLgaAjz
zS1JlxcokxyYKunt76XLrnxFwJD3zlDkowXWyTX7y+2Z2Rumd4w4F5RQYJZNC/JL4gtB4x1f2O0p
k1zM8GsRIUe0eGmIgsbS6E7sMdVJoozBsHU+EqUYz/DSrJPkPzckNT8cng4clBFbITAYD6XlCuh/
0cI2NSP5uk0kjUCUeUrhk+cW+AUwOS3oH7xE4qdwmyyRNbuvj5yxI0uPemLjrCEXiNUNen93Ahyo
fjirqwiaLxIu4HfIQgnDejpee9eko7OEgJlcp+Mu3g2xGgsLIr8sYHa36Xt7cXnblJ5wlDFdZO4e
QL0ZqVUJafkVm12+e6PBexgnv6/nCpgzi8QLCnZbEf4us7c8jrLzj6kdaxLHckgn8f4CsUnA/5jg
7UcO3MiFOvIE/uf1AXVosV4UPBXsZ74fAP4UfLN05evHPNhZGaFYDk7tlReEcfhAE+sD4WtHY5g5
eG7FQmPIMr3xxRvI8bw4fzNv5iHHisRAJMZVRZCudkI8q5V6mrmZyamsJB2FRQvX1R1qk0uY4NPU
6eBwYiZ0bcsyFPfAqJY2MdXWk5YcrjE0yGO/Dfd03MprI38Z0lIjCW8ymwTt88eLbt1XwVvsBNDB
w79qglOjS6Lj4cuRSMBuW3BOjtyeOniGZdYDjxImBhGd5Oty67XcjtnUIN2hnmNN19Bef12F/pgi
fwOj98PElhqwaON+LH1/N+IF7mVWeKIl1BRazFs++OLxjUMoEGgyQMuE92PM3k5n6y/J3e1u2M2Y
hyi+Na/oZU8fE1Ka6VZf205t0A+YatWyPZfzLCiXwhxa1lgQgyWA0CntBqkH98gjfZxQ7f+LjY8M
XWd9pjDRYKrKnz2TdmU7SQrrcKOYkqkzheRpijhWJsruKyqviemQUN8LGOmyzvVH8XwNLg6XrIhS
T4j2VIVZR0D9Jpn4AIuZmOWjkzE87Nh2vEbz2DacDyx69lIKXSDGSOxLiyDHayp0JabgV2iNcJF1
6LgYWtBV+e70JfABaEX/+vAToLs0uLrhE7WmYx+0A5hrsjGmphZO9V5jwDgXCCn+M+XtFq4wBAux
yfFHsKGOxkXJDOh183lt3coweiIOFnG64ENBjyHTC5Dq2dH2eu5VOdgIWcVTxtJkvb7vTYDILkj7
l+CLjjPjrHN2Blu7ysaIaAtiHtCQs5z+0/Ow3/rKHm8WkjZSYoYvHppzA+p1PZdLwY3sS8VLQJaA
Vd8VwFqwmmz5MuYG/g1aDGFbreY451RGLujWMSX/RgNrm7uPr03/ImLl0804g8NL3g9Nn6RrJ93M
5pJbeSQi90NZ3PtiNEhmrkevkxHGlWdm2swiRlIOTFQAAarvuf7Sy2Q3RpQXHo5uj91e6E7WsSr4
QTFF+3knkfkVTSQda/6JqoMW2hE6K0ZHsgyFhwCD3i0l0NMmE6O3k5jmkorbRXtQX9P0usdw9Zl4
1IFgBT/CbtFRjJwZySJrLysTVRKh/gdK9vcwJo0it8nAofjbQ79KgfHuz5xnWpI+QILoJTfo2o2x
BaisEgUP042/4+byah+j0u+tk/7zymAqvNb/4G4BX3nEnOo//K09l3+s6uSpN6zBT8Cs+HHbJqNq
G5R0FgZcHP0eUZLNyq0w9fF4IZxnbFsZcGt4x5hcrY2Fpl5zg5oWJ4UtweD6Sm2h3kq2kZzlxGh/
XLnaOsBay25tpZh6Wrb/QZ4YfS0J82eQhpdSOLeDQOMghWsb49sRSnV0Q1XUL5JAr1a4tU3E/sPd
NKtIWOAczjv5Hv4MQoMApRl0uRB2dD+QK/0CNi0A5SHYkiRJ8HnQGbxG+Vt7aih6+P3Uybnca+Id
1OEBtVURrlJUBCaZFH7cEhbVFkFp7yCq8VnBgxzylI9BC3grLcKx+3zZ9fH8RBhq0Of5xOYFSzIQ
LGr3TbdedwqlK6SIJkAGDFqe498ixvVlT8to3GHbW0P4RDNi4zG8b8c+ad29j6oa41ZgQB0IJrit
StbDSAzJFZo8L9bf8JhciezWx0wnXw9vqMyimRK8ihHPIFI5yZnFvqUz1pk6RtJgCJqm952D22oN
mjheDEjXMPblb2NYMkMeBXwOaK5Sp37ZXj768LgE/O381s8BZSAbt8m/WVoIviVtf7JIEdR7rpvY
KxpM10yzqNu9mCpOP13d31MMUYeBr3n+hUI3zg6+Epehw1kPIGM4VuOHVUoNf6q21hsNJQNT1uMl
4h/Wk3mR4bdcC2aqZ/GuA/HVp+6bwzaEnRm2b8Lq9YuPFVShoG3DqW0rgnDinOfq8cSQgMpL7mfd
C8Vt0pS/1nIvBxI6F95hztC6jJ2RDPT04qL0C9xt/usC3NrADRIMmmY4lMb8YE0z2O3deJJxnucz
8zrP2QX7Bg6pHj+5kvi/1SILxo5PXHgtyMXyPIkGTFpcT5fU3GKTJRZnq1SaR39n8tWyjb3r7vC/
hNVdd4bo/tkujHbFyr8RlG16cxh0aVTm0TGGOEPVIAeEq69uQ+UEVZktzxDmFNyjPj6P9Dd8QJeG
Bgpybhy9kQsI1hMgSlw3XVikhEQHLwaSGHcxL2mhfc60y7GdK5F5vcNDI6m2+WzxlBssCxUWkVuP
d4BVn51AXsl7ZZoBp5S0BkjybNOLNzOWKKXI32krse51RwAmWy1azJME6xaeTQhfLxohfXlV2KCi
B5FEmocvoUaDWwJX+DFFm50shKfOx6PmP75X9KszqDhzHpEo/9DKoZ4BwyOzDRZXFZAMN4LRI+Wn
PafKzGaJlf7oQ9rEdXOC0fptyxmWygk1co+itirLHunin7VaK2lnWNMOWDjoc57CzEM2/2vM0/+C
jbT1Qs+2wVqjn+RL27MLlmKjYalpONq5Gkb0QNC6/zhVa+6ZvLkrq0hgK4/rVXeY3cIyIK+vfweC
pgzBSQBPAD8W4dplHfmJ6CkED63PEJjjAkE7twbmRs3vFY+Jy1cMf1Whr7sumYMVyyHxl4dpGGv+
Iovzzpk7sxkBA7e+JCaX/78eZYICtdvlFRpeX2I5tTkfByGFyCtPuoZl9EO01C3RL3PEDEi+KKvN
LC7FRK7EiEkI+SRfqoZuKou07cL1MlaMgfL+2m4/U3DIwFXzjwW+G24su5AHGulTdNDa28FVO0yF
542gUIOqY2oeUCUX7/OmG9+XG1ajOl7PaA9qw3Ga2aGNoenaeJjiTxkwQP6ZozyPbaY9oQN825PI
yYZuflmN45bvfd108oRm9d00r79UEL86YSpJiFa17YbAaq4thCNVy6lYEUnL8T/SOZagibtHZHiG
/47/bUluSbh3JiU20vN1Pd8liwlJ7tnFv2i36Sl2WbfAqH4dozBntZAWkjnzUIp88XIA6nOAIlkJ
vq8m6X0MG0qZPn1FThhzlPvGr/MfHZSR0ULyiRd0a4aB2oIfswuxwi+kvt9k/AiVOWhmWGHJmjX5
pRLubt2svx8nBfosqaO01iG1ZnFFRL9pknHQyX5PVj+HGs+RC2HPj94quOJOiSu3AIB/f1abPShm
v5e+BOmAQO0Ji06t8bllwInpN+IZdpLATfkLaE04uXe+QSXVVfnkSyS1m0BDcUre5HIqd3ppa8J2
omCmyYXl79Zlo1OhHLPJYu88bIs3ekLCzlSofFzsuP3CXQtDGdntux41aFRYLaxsRQIZaOW0AA3A
mjqPHS5glpiXXo8VxHPOOh1ZCwDoICPkK1CpRKLCfDLFwUcDbLuiedANcxfAdDJ7NH+Z72o2IJ7K
s2UNR4dexdFNB4BUBrtwKJtfwe8hhdO4AP/nExqc6wJwf0GmB4fYn9YNU9kAIsvYfPc0bJI9R7Tr
f43vTo2TUCgZLDy0grDmiKfNc81JMsXzAJaGBVQRFXIJumB49wmXErCdNVzxY3iI7IJ2Qam95J6l
FqJyNtqFCnZNFWRABxrnCAw3U0I8nSeQQivG1Wf2YMxmITTDyMwcX7kDb7UXeXmAqaD0zJhWLJyd
5PbY2uNCcEACJcY9IdiaatOzA8BjuIfdQKuvbgRXc6DqCaLhtusTio1kDPLMLI70RISgtGxLXQM1
X3b06y+CoI6cfFGPuKP8VNNCGoyHsshcFAVxkQjyCdoxM3gvcitQtCA5xt71NLcYsft7GBjZzgxp
dw4G5p/7VJIjJVjiL+Z8pIanHYgzAKwTOMm5YE/XOEP7ITdYRahDUm1PLzCdU4EfgtDFj1gUvqog
TX/Pe2nAXPlU9xBvREqo1hjR4sgmLq9ziaII+0KF2BwhNUCfz1BQm/2dg82hJPq6kZL6EEXNvD12
JR3LJDGX6cwv6lvg5SODomOFpFMvueqbIb8dyvxla1opkhVtHadq5EVScVd/T+rjhDWtU3Mbla1d
SPQc0YRCSGXBSiJ/E4TocG8ZiqkIyA4GRQrZnBz4CYliiZ33DEAS79tou+iMxADDaQS+p/iJvTv3
zbcd8YwLqyKGWoxIt0CqWVWqR8WbuMo9fpYfdm4WbF90XmoYejvfLC7CXHLMuw+AZ0UbfnJTYPy5
FTlQPw0cT85W5+u5nmMYyQqpaLjAU9tHAcwcvN2PTjoivtm+mPamHo22RHPJBAJvBwRVrJn75oIZ
mbq53dhMvbbe147E3aFQy8xjTJV5h9LM48C9olA6t6Oy5+wozolM/5KNi6GHjvezJteSma9VroWV
8NhdVWRwIaPugwDAJ3Wzeisne5TD6jwSJT/yinB9aUnxU5GOxO0zjfWVcMOXl5kpE/YLM5hW65/3
VusfYo7invY+y3asPRew5LmNfQJ9YZmESek2+eyPj3rcnhyeoIHx9r2UHDbWW+etVP+7ngPpP1Tl
QLJ+O9Irc48PHE321whvlCZwqnzuTNNHWN4XRgjhcyvwLG+FCMDRUx2ae9V5szZNag8rf01laVMj
51yUm/4YE/luRPyd/mpq4BWplnW5bcyg0rdvnt1oZbnozQ0+ZIm3Bnhp3wn9qJgRMDgKVFeQ/7a8
BVgKoGgc8fLBaZnrqJVyHGf3HHc3bYN2t25GPCwBD1RQs26RS/pkwHn7Ntd4TRw0uNo1msozGDrv
U83wAN0zIiv0oCxexlx01OiyO4hA3u4ci/+pJWFh3NFY96stQOhyePv5CXqm8sOEL6Z/wh3FlQYL
4qN3HmTVZnwgTBSeY8oJXEe9PgIiOwJJNGHGMtO8Aw5Oih7VX1cSrfdhXlKI5BMuV+AaKbhQkfwn
k+7VkhBISV86yNVMMC7VqaGQgqI/eR9FH2U9TrISsCXCyfp8+9E0i6oASxbVgtQXm/0tJNVlr8aq
CYrQg+q4sOoJYMxMjnJyGelNXdIidJuDyaNh76o+OeZCeqXg6FBJr8YhpS+JSCtIfCCO/6UfmwlX
6LHWO3GFT1EYEwkweyrs6oFLcNOo7pEwpJCWKi+tV3Be+sta+ch2VzU5689KUXSUrIHLLbhgJPGn
H9RMx7rjrzj6THuTLoPLpObv+MusVduE5G+FVTUTjAJ5Bz4Wz8pOTu0i0dXpgGrVy2h2Q4DnE4UE
ZqNTo6mHUAUhpDLC9DkwIEwXUTwe8NfilVRavAttCLQkuftknJv5kU3M7yxzAAitQv4PFaf3GgFg
/g0L64WL6zJMJPeg6FK61lV/H64JBi3KIv/jEtMDbgBz/h3G7sh+qCEQ4hkQaoMNpjU7/6pORqIH
CPBr3tMig8DEk0jknZVJ03IW3FnbF9G2IxgnCqesH2ta+vh4xXjvWZ6RltcEpe88rXQDLvbGu+ss
Un4CVIGAqGndtGah7BUkSKti8T6wbZwoHu3omUW6s4akva+1IVQRxiq0Iv1w4yFfUi4SH13u/AK0
9PwBYhLATFlevlAlqpJeoHsETJIsJwJKwtGBvgzfn0wMykC/g+W6U96hYRW2OZ3eI5AG1DMgH9Rg
OYloImLWCk5Kwc5cXJT88nNq/0UnV2In8e7ZXx/OwqUlUawaeLLTCvI8HYOmQD3nVg58F14dzfgv
9n26i5W1gc3e2YIEp4CU/S1p/Fl8Mj7CcEyMfO3Q4lZH/pgqlbUsMWfjXHhqlsYR87OlBoNjEVQF
6jOMhMYiu8UHiZonx1PHjhFExixU56pu3m/gKV5RmzIOUtSZZ/zfHz+3XKAyC+dtsOMk+xxPTo3P
wcq5cEdowMI61q3tKl0kkwzgxGcVMRFjvGPIz/Dikz8hPpV5h/gv/aKMS31nxOlStJVMJf/FNtbG
frHyI+BHPVuM7Yr+lbGcYZCuGGwKXmDUl96UVy9SXDp93r2zGGa77a9Qd7z1gXyi8F2QWq04jTUy
G5s9HOZpIjhK5oxVNmm4Dyqb6PnCT7KM/493D3A8CYLTSvhB4lGrZylR0oiJqJ+uzPn0dgpP5pgm
QeopXAJbSPUZ8UPV1lTX2ck6VbHq7+RxSrF5CGP+1l/19fY/qLESFAH3my915cKJsi/2ZwGjkf/a
MpUGeQdOfbuny6pIw5/PfgvozIEwFFnOklPibnqGCvjG6EW0cr4QSK5EszUrfwFVtwgwYMcR4KES
d6jz2ZZqsMHi1WTN2reYFisi5Q6sN54bwVKOjeqvAi+OUvugD6C23PVqCSiF1/sWrsmf4EEtNZFm
RdXVsYKu1goBWEin+OZFGrZMVmMqMUDdsqyzGVS/zX3GUs1eGci3wCoK1f225Q3lIp6kvoioimbW
V0C9KUTZp0C74ykVCD8qRxqBRz0IDD2akUFWPAh+ImDspCR+ETg08gP+lN2tH7Zf+mXQu6AcIguq
IDUAekvchmdGG8srtUeFeeI0slXtXO2gMIqx6svJ1p8qAOU3JCzAiXd0RxTQlq8hiOHtxOFuw2A9
K6brczZXv1CFUXUSkrlh2w0etaqIcrMaum53GmrirNziOEU7XVn6wiE6pXiaysGQsjUIZgKmIUjA
3oZE6nc5NvFy/CO5yZ8iS5SUIrIRPuPFhqhwmZmi0mLODEnsh1trzi9PwwoGEQs5at7HPpQJT4Xw
w0m6ml5++WgRBBWownPGaEiNsCMtwWyS2+y8W1ugE5KhjIO/5+Y/ESA5rnJwIyLAeTrvLHt583en
bTNvfkjZ3zaniFiDitFGdXipYvQAzK6IGatnfC7YVmw2Vu6pprVceQWmJw3fH5GRKor0ORsb+8nm
Ns9D7iSTrZAdaf2GC6ot9iN4b0JgCiLAaXqkeq9RyYylgE6JnPvrVs9SyxQVWcI9efGSwxWc8u0j
XX8OtUU62ygMDrEzYnXe20uYRvRZymdXouI+K6zDhhjPrGPZ8IWifVELNHIFdjuNWUvRSDlKmiHe
CUz0RwBRdBWE+VQ/aiG9HEflQLGCJ3kfux3fDd/fVYsEBM2vEXZ6Zcu2zx7vLJVynDiY3QUKUtb7
MZCqgLF0+M87mmTROhYGcXhPldRCLs/4rNCh6+8SRmaKyrv3vosPS8FODFhPLgTyyGlSsW1GQDop
Fv2iIbBHrV7FXn8OC/7rDNnAhcTCaCMumMvVH2C+yIiVpxhokksneW/1yuaTlPo74eBAaZlFnE+n
MoGgvIyGO6dHPsPljSKI0rn23fPSBg1IiRafaSQi4Ll2HtyWOP8hqHIQSP3qnyyB2Qh7XItjyEYB
Q8+CrKp/LnYkG/mcIxeksUYtOSrW95FYJ5Zi/PyEepROAqlZNhTqckdUEczGYYlfCPydsMfXN1BL
h0Vlt2Q4GzAO3SVJywE6Ul1TssJgxGKUDn5l1iSBcAT4S/b50XsdskxoCmp+XsJrZlSc+V6XQ7Fd
twEhgozam/Qnmv6bFdzfkc5OqCGY3OJhllc1LO6F4Cmw8BrYaXuVl6GRLCpfxyy/Y+jKP4rW1Iea
op0bQEW7d5ubXt+5CjC/ArWhZQONULIXyEaNincKI91sgc9Roced7LdCjFEeCiYrEtcV8MvcqwVs
mzvoedAsK7X69dstiyMk9bK6jZifBJ15Ws2u2eiiPNRZa+w2e6BxjV36CyQRLdhrtV4dYpn6WXbh
UokGANa7I6upMsvG+JFdUmHQVeZ1zNItJOkT4FAiY3NSgZlZeDBh+YhDDFJNBrqyEt3nMySpUQJy
juADNbAl9oqamKqM6+C+F7e1h64gdOly+a3Od2+NIT6c/6dnRnsjux4I1kIfyX5nKdeWHlNXr+h3
1gWeiQIFO+3JCzrgGDI1U1wXOc3qZGr44npwDNJp1uZnUCKY8OQmmn+IaWG9kyCUdv4YymBebfMr
iVh9foEFdWZJbF0LXk4TWPq0+CTZnHPaYAkywJFjk6a3PotEfnpGtF28GHAhcShqzsGbCeJT1vlA
mRZ9iNDSXENBCJ9pPREfoFKszTBSiABa4Oc3Q3J/BmATTFhK3G80HlsTHhtOQGbmRlgsg9DoMAtB
YD/893aTTUuU5bHrcPMSYLkAYTZixw7OGP9Xqa+y/KDc7YKZeXCRVvVr6MLlfnEU6xVNrfE1z0ky
BQdTyfEnwnJo8a5zr1tWk52XVDeKdOkAx675WuIwt24La2TIi7kRGaotZeidQJE7/mFIA+0qEZGu
PJQ+ZLbAesQyY63LpDmrgGNr9lTALcUcb30cy894UIfL0w7+y51JIEABGgTW1y17GUXAet42GE4i
wq0bpdz55IeC74mMu+9jTeguADDK5TYYjOM9nTTjC9/NiW8erU5JzQjsUCPFaKefyo034xjOMmPa
Bi0GsXhpSRLuv7IOyagtJtqwmhvurb+9SEPMPgp2dpGoRVEp78bLVwVieEY0a1YP6LrrS+av3dIC
dyMhFRe1QkiSACf7b/LUTHmgTlVoJFibGsB+YaViYyMnm3lmNo/sV3tgbXOxDU3qUHxY6+AnCFGI
xqq7BwxPj9dvHgotOdSNidNjHQGF7Z+z7cKtZgmtW+AabT8/cLPBEY4Dw+EEK0wwHHIxCjl1DjhN
gEQaq7Fz45iPl1LKRyctPFBNyuNHMcrtdLczC3dQbe72aG9jmO8LibWWe/NCKDdx/udTiVG8yh0n
YgM2M7x3+MvZSfKC5+Oa0VsR3I8u7Kf1LmIJekfb2DXi5ZtZQEZiomv9JqWAZxXv2vfKePB4+0aj
fcZqvLXZenEvlXWRcMcLo1KEiG86uPTWjsbSNATqaG4X0fQGmbyVec31LF7TVvHP4D9qBRJ2xpp+
4UXpMcXuexLF/C8YTOcpofJMFS/Qwk3CqhACvDPITElVukCrdtbuhzwxTjngyxNUGt1KDQC4iwry
HOwDXjyqy5tp9LXjAj/3RueInrAu6LVwX6vx8397ykPMs+Flznv1NemsrRfUHUvVCiRvePJCtkJf
z1cJ+OfO2EI1NdhHvJyk8dd7/HKWDM2NqqZvUQ6xSOXdRPnsZNMmdw0pT79nO/8vOLD1G35+PJsE
GzGLsi+L8I0oK+nZeUAkPkzDT4nZtu65/QtyEBjSNcoHXTkfkpYOioU92LEKHqOagvzEHvnL+XVO
SU5y2hrifCo63oS4DSFFiUHB5jASuz+Xc9sOLEbTjTZzKtk6hZqLCWYF6nESP9gSIR6W7a/ioqJK
lGk2oZreMlyFsARtE51eAZwpGkZPV3w+IKoBbez21J9SisT1AEdrpz9D/x8q2SMCF3Q4w88MPQhb
RO1fSF31WOxoK6U531vZ/Vp2kUylEPQQgbHXVerdwUyuU7irSFvr6Do40skitd0hE+dtiUKHaw5o
71hfG+f3ePfBEgbfi2sEDFCzJhbFFKVNuq8w013CcybeeHXh6kWLbCNLtsJorjBYNupSMeL1UvyP
ato3EJNiXqmFAvisQN7OwJpOydPUwg7yZmd6gjwFEo8H+9oZ3OSTQ0aK0YbFfsx3mouQGfopowt5
P4d1GAhE86SsX9wVVnMFqJ5ZdfZa/R1B0427a5FJN9wjrtufCrbEtBipv2StjAaY5V+CcWjSLxYX
3mY3kbVli1ocNBcwCYyndeAEVyALaX91Jzw2Wk/7ln811Vp7hBKaUrp5mRZfMQf97n0PrdRoucVE
BP7BPXH+VVNCzb8QZ7pk+1idVNqoEx3eP/eHggAEKqwGHjsd6MjeayjULTsuSyEFb++R/MIua7WE
gUQf6MQKGE9294aLba3Ydl8FIYmGQA8x+4zM4CUjI+N8XD+sX3r9BUVX7Jcb5+3sFXBvmbdec/wJ
hppwosCzG7Dk52zjF2C1Swb4nP/L6KOTU/K6V6wVDMyttjMLSWaGAYMy+n5nWct9HgHud5VIqAXI
W8pRf+MZpZO2z/x1xaKzYMPXepTO31Ah3F3l+MqE/WkiIfJ5vSkIoWzSXR4Qr3uAUec+pS056ZNc
2BeyvBHOLp+2SuxDAA1tbP24dWI0rLuLJ4lRlx8WyDnXPtx02QRcArI7biYxBhdgmJ/SvVCSsWT6
zbDVT0Pv36h/Klgf6WWA8OQbXUBfo4x+CPLRHWqkeIgZDXv9s0g3AKuNQkNENu+h9NKi3xIEnTA8
nf9EXRo0/jUD5XvMP4tNW4/0Rr3u7/x4WknTdmYm4Vls8hWbX1EWqoGtUucZ+c+uKylAseRiEO8E
N93WY7Ks0W32xok2Md3KON3Wmxtim3OqEsjsc7LJFv+KzeE6b7EfaoFg+dt2K5sOUoAtLlNOetS3
IkHH6cQFeaUut8H5QjsCW7sL9TJ1TRRz+cH5lcqMaM0fPNRFUj/BRJ5JuMUZhLr9o3ddDu5imc5r
jqVVS+jIlsJ/ckb+1k5GxU1/dba9ArmVkdd/aDBhVx7TwuxRbQy9Z9pc9vFBPXx8kIFECYqzQ3jH
BXfTbJuNqajryOSjDefa0BdFEHtVhwfLksdEHgNQGu702oshUp+anBSMr4Q3lDMZFkRfMfHCDldC
Mhkrbv2J9U4hejln0tdoQ0EVBjVTOek0a7okSw2zEja2Ew6ZGueiDCW2UqqcXOrc3SIJczfkZWei
BwADTJZkllarMJInmBtUEssSSP3xaqrRDgCnwe6Mvh9lR3mAiSroexvcVW+qtwei0tOru5DHr/D0
mRNgQpin+JqnnHazE3+3MjWWuIMT743brzhRYhYMC1wz1sZynrBe+MwKOm4mKguc19GOeyw3vZfi
vzvPvzo3x5RZgGjJSqZO4O0naBkQXYby64u05r3/aHSOQ5Sy8usqcvZ3goesTZZSIIog+H0nBEgO
nZk16DPEBLRkNIe13HlsjsnRrT4jGZ7mh3DSOQKHvFhWgeAJcpmEZhmUcJVXwd5FSxYr6iQueADd
Yj99PVIpX/u8RKzK9fEIl91x17NBnqfoWFaXVDo2A6E629hIHyD3VF/MCV/HBtTxUPaDx0RT/Uu4
IaGRWJc9Au2ULRQ2vClWrtswg+f0Ld9yM61ul6GtjFJIEqT5nokllT8IFQSUoFHqEZ/r+T1d4CWo
CvoD+leB7Gk/xp9+326SOriuu4FPi1lOBBkTq2sGuG6ITO+29Yy0AyyvaaRB+RB8wSprd9tN4JES
BscPbWdatYgrC6z6XgFwIYyYuTuAme7HK55HozRFjK5hSlHbwXecaatC/2PCmjYbRgL2LCp1M23a
ngk9xJtaGJIfAQ2bA2N6hcygYCTVJho/EmvsH1e5xFCz4tvfESodExOQJN4go2qkGM1tiSO1Ctar
AMIDZ9XCX4ojsweLT4ee/mLMsEJ6X9FzILQ9EWrbCM44FUZofsS+3zJYRmmN9DGuWe2hibh5N6fU
8YCfOOCX7RBmidm9P4xfutn1li8KZ9pQARykbwdh5vWrgkgu3SDzwLbz7xLV0lrjAjO+tmkdb7n4
GFfcR3S5srmOBLUjr2MTe2oQ5lc9gLSFoKUXmqgGoNYXLczrVrIL6fsjPreZcnY+YBBxIiOMe1bo
FkXsD5t/KwM0EEtHGGKaNfc33yEjT/uDM1s2EJ/+A6D8QS37ytGyq4MpRSENof23BwWwg4WS+DrV
xr9Qg3pFm7pzlcha8uxjHlRqrrsSOBQqxLYVevoXcZjtUwZd0KMgt4X6XCE2xSoAli9SHVN41tGG
xc+QkN7VfwgF+CeKcH4YcCqeCpnaYXr6r5LYMZhLiUe4AmYAYnEtis0GdPvsbte904owGf0R0k/I
WqKFG1FTYxp5qBuYNqpHJc41gqdu5+ESNwiwDudDCzFX48PKufWHASSO2CceAnPE6v59ogrpKQZd
r2x13k1qBOQ8SLdRgcB0MJr1hV2fi9hUSLVtr+oo0Vc9xa+eUaWpdkR2CfVApM0z2kgkpOcjEQb6
IMLxeApQUtVD99umvaLWvAYti0wv9VydCEWS6vRRfXx1+RGeV9v5fc8sXQnAlhyLvMY5m8Epz3UG
r9sz+ha+ls+f3bFcLU7/O+Cq+ZOEqFeHGHWB5nMb+Zqj4HXVZRCyjr/h/Bn2x68h0i2hRPIZSLoh
x6XrZ2RMIBOzbjJlqRhqFKaxDtNrj/4GNA9q7RUUotmnwkyU0JoImsDiyLJMFSww9GF/0sbFaNIu
Z3+FBV+IvGCyo3fTw9/+ot6ba3QMlwfM2ON6vnp2LuEPrzmoGb2ROA7Rj//46BCkKTfZ7/wGpxMH
teUTOIkV/qkcam0deg84Yw4XF7jnw+INqend1sJvzewfcP3J4625tWmdyUtmYgyUzJTBWiY9k5LI
HmR8V51od/9/2FalB/iSO18foUPaU7oTBgkGLeo39JuSyIN8EymUXD52/5FDUZiLaqtv3KSY4FFI
+um4GcQzQdjYTd7ZgLAfFURrGHbfOQTTRAvtcKM9bS47F71gibQzy7/YSeq7bArtDhMELr10N3HI
Z9rs2YnmJDiAf6nVZ4XO5KzC0YAbtPM3dHmrkG8LQOKf5WlB1xsUy3YPvWuq0KIL+Zj2zkiMeEKu
IEG4L1BBRVmHlmxCw6yd1w/sywdZGRMg5WCG6mHNXu6vTRwMzcolfsdIUVXQHo2y2InqseiKtXtT
Qm2+h2GK7aHA5daGHKzZryTOCCI0O34hvSYzOQdZfYfQ+1MPZyCGK7zmb2ODUYN2+5wm0UsV/jys
MevzankLKepgGD1JqQFcreHkt/t91m3LbRaZxMPM+ao3kYTD08ti2exgKwCQN0W8ARFD/m6O5tEQ
iQDc9YiIVdMGTzs2FlEKkgjAMKsTFSefOiu6fxYyljfuNIRVIEmhdOW2gcRwu0TR/05qMGTMlQGN
hlTdqa0zr9eIPdu46KOqihRRIu2cE6LAZBLTALwnggsG+BnVpfkDBZdOqe0xYhwIyvPKN658q1VK
jyyh0ST+1R+WaHp66FTRxzWFJOdQUDYHtFb6T84OGLLwIWSYFEJnjRm3n2lZPom3G2OKokIfNc6m
b/SfbOhsLOLuQAOccNGfZ2eWv91rvRzFvBysn27N0jAAoC7IL4PwIsbDGEteRfsK5t7YoyMIwqLN
MHto0NTWeA/Lt1ABlYe/gY+PJTdeFeAMBC404JQKlL9Pedf8vU3ac2MrFX5Czf3xrXkMpVKDqk1B
eWAU8koWQjJmQw53BaqmDdiRm+CTIr3lVxi0lVbNyO0QoaBInucUrlsp54JRFpRAHRwTd/fjfcim
7zijn9LgYhfd0nj9t0Qkp4Z5uRMpk9AHQlmzifcmy2CFIwnr52NfcNZHVALbTb9uSVrZbiYweC+V
2nmbbPUwopO7PA43VPz/AO93v1GtKIYX6aCRIJcO2alVtE77Gcti9fFDZKMMIViFCCzMG1coZsSA
zWJ0vA2DQy5rx6rkXvmbc0YsrUYXUiEf7M1zXHPlHD4qp2QOT43dcFDBprwr2Mp2CVKICHePWAwW
Nn98o0LGl4nx0Y34/HVXBvpYOKD8jlGyXy/IbM38299OKXLeF2+dhiI8SPj6w1B48uMUMMIWPPsG
GtTbhlG1ANg0pB8wjUQ/c/ze7itINDz+MFkWovj1RNS9TfQjjmb5XQ92xiGANks+4fDKw/ddunig
RfOqZ/61GgDcgrMdmmCp5GQQ7REhtqR+ro7RZ8Irz5jlV/3zoDcOy/IGY8F55jfNw4JhPRxuqvPB
EEDVGXHn2HYxjjBlAVyqZokFMSthkVS3ledk8ydQhDZ3LLGNoOH4tbWN4ekZ23uWqd1WJDOkuPxK
oc14t6LYEH6s6GPUyzGRag3DtTEIJL+HF1OIOt9ee7ye2dwyThZ2mXO106KsH4VYWYLSGzpI1Dwi
dOJ7r3tiJXuD7RdmRLO7ANMmwN24qGT2l8LB5Xa7N+V315CfVmnA1Q4sEnbngmPEDv35cROlb030
lI47rSlEb7+Zf264n7SVwTrv+IHwJa1u0Gs+S4MUVeUQ4d0R2p2aoZApi80OTp/zI6EfxvR+Z50Z
e9EPGVknW4+dvfwRh2Sv/nX2K5el8+lPZgOvJtJWpYvrG1es1q14Be36nEjUkz+f6kiojsm7GfDu
2CBpmDXqunWR1hYL7IStlV1DUuPOhy3I2PNVd+dImeUMdNRRqbg12ZuJj4vY3AL/lRYEpTSywffp
bJyfYSmyquOdrka0fSTxCFs/C3IkIWj1LeLnP0HOrhfkBmqZc4x1EeVNcInEPtlJkvJoFMTCTbok
JyTduFyp6muHD1Y/MNbDyBwlK5I1DW+5mcPJEVOjUnWsFtEq3tN4BHaYX8iAZL+U+GP4HH2fKEia
xs4YxuGvTe7wc+L+C8a7HJx4MFKFxgpAMHcprijuDU4IzM2yapsIJSEvfEgUaSVYpyrUsg9+d2A8
eY5zjcT6wJ9yplbVzKKPEc+WD4tREwm/IjcOwaEqXbrMLPeeGhqdpsYg710+Pq+5XzZC17ZPh499
Vd2vevB1ui1j5qjVHOKRQVT1yb4N7iMy18ZHr3z+U8oqESDqw+/PAz5PuYV3jdwrQ6pfOjw7bEi2
ZbO5m0KDJiyNIM+h/br/wb3E6dWjVJzbp/L3JDdFa8IIJ1B/BRA1TfQMMB0fNYX4f+wC05m7gtvA
ZIQJ2Hbo0l/IWCqjjR8BwmAKOOddfLCYqlvgamKC6VL+QcFywF1b4iXlMg6M+VfFdlcPyPwCnk6t
krVzpOpVO7ELwdHf5EAFO5PkMOoLDHaes2LmqLtXyD9ym+KZVAY8s4IjKwuch0Xl9j31IDBKORcb
AulfSMeDbs5kO4MG8nfAVJGXRpSmuHGSdfDUfH58e33ORiWoQkXSHxxmf1tPdO+K81XXEOY8C7U1
bDby0bUOVaLoJM5zsiqxQBLtlGMGIt5ZY78ZNa2TiWGxT5COqhfBM7ikHNQYHhXfR71e0WVKuKYA
UK2dvStFfoquF8WYPI4cToQewgt97cNkCIO08O/oXs50YGWPWLinZp7pqxY6ohzmoL/e60Cl/1qD
ag1qL6ip1yVx9+3WgWHw0ualgjhDR2W+7UPbxZcOOnHALgS5RmzYfma+juD4/2lnFf59cTpKuAcS
nLiodWJdv8lsYTXdpfIiJfTvj8sB7byyyuhlBq14QfpbcfG9Ex3y4GPlZfmR9OfNNfLTzw9lDqxZ
evbZ4MRnxIPljwYR197gP1HnhlhgFn6fbX+DaeDtMEQ2VRbxwSMf9mdtj7CxMRIehmlgZyX901Zw
0Bms0EMmrjY6xsT6ZBDs2tpEEjD82rtvCOazyQHEk74Re/vZbhqWFn5xJrxGZy6LgzZ6lkxeb69x
ASsk20CBRIc1vo1VmkZ1sSfcEln5g+cDpaWQDG5mAuQemRHCqkQanM+lcB/1Tv0NLQV9AviHb9Ct
HIKBUxh56mzkR4AylcxJqso/mOgNInWGm0hGR1aaVNi0HldFZypiMPLH8xDM7ElPDbhJVPxJfjP+
lMhRgLqPyOPslfeZ7rH7tH6mrx6muAQ2wIxktMMU+2hKU8msVbmDlp9XihZ5yWUh7eToLdH0160i
hxm2xYSy3P5BkcFEgR9URTox/JMP6ywXw1uwPdDDPslDoWLNO7peHuUosqnlhaI2zO8dIg8SX1or
KD4GuFBMu1cIoYTNw1hIubOSPOTqYB83JGrcDXVqCV2qAYpymzhmv32zUzBorWnSixKsv4OHzXWT
LDmKUXrU5eiQ3qSzyjPznWkfQyIMfl7MFFGjE9JojyHR/RHQ0ER9lc2cMsD4irCKt1+mCLPE23T4
gU5fLC1N7Qd9w7LL/I1oTV93ZRggC3IzjDsutGeJe8Cyou2zbZUDF4P2m/KYNwGYep5Hc25cLtmC
gxoq5n0bQZf6t3mJqyjDXQHrl3Kcj1qpHhCsaGLhQ/z45wEyIpdVS5GhcGDiPFdZ/r8zN23tEDhq
cCUmA2ei7GXV05jIjkTFkXFKgM4JAaIzkOCpUfQwGX8Ll13Y6a+yFOfpWLA3/3g9xJiXmsVdBSTM
TM7VTc4/9psIGXYrCZtk/k0PGrcpjgtzkPnXFOkL7NVUUyHx2DGlW9bKzkRJtdKHjSquoWTJg7Pl
VMD7IfkFHS26DtMTvJh1MqzPjRIQG7BvtYJrtkRKOzZnYdJXHs9WtXFafUojhXdWrAK9LiLGYUcJ
BGAf0MnDpHeemC86jKoEIWuVbN8JRjiTo0atzLP84xwoCFleaqEneHYeHmdikHdLOjeqGUfawiO0
DeFEqDZsVyJuVh/61SkrI8Ei/cTrBAOLoO9L37EykGe+PsY0ADqi74b5Ay78MmfOYkGbCoX7e1AN
7TGRCq90ElFrG8GU+lmpAysWXOd1YS6FgPCp/w9LGlv3CZQWJYMfyViugC83ZndL21VS8M7lIo/m
r2e1WYR3b3vxoJmjp5fIBBmXq6IXNYbj1wSuzH2Cpc5k1/7hpgab+cSmI13M/stjcOfH/m5L61R3
2Qprtvn4L+r+e8Mlg3S/lsE04GRYg5hhxOPy43DUypMZ44UCZuHKmpheC+CPB/IWmuZD43HSgzDk
j/bnKfUhDEd8LsGLFkzBCBC1I8T4nDPBXPt08ZgBn6EhMgizqDT1oKVTCGJcWFUTVJwVpd0ahUms
LdQHcfvhh5AHnNot8ASpsKYPang2BEyoTyhiaNXxeiTxxSM97/DPzro569WwIJPG6bTIyPHkBKqV
0ssFiMqAdajs+34RDHm8XDAFH+m5N7H1cHZvorwG6WMhF5pdM+pDaBHdVDISWQQ9NHTJUBkyn7gu
xXLLrEWa7ct0YqVpwriqGKsoaFkUdzB6pvpShbDBD+0GJQu/w20cHB7p8F93H6OO5IqNZWIm0I7A
/efIivmgbOysRWYx7/DK5nOuWOHFqmNIgZaxTVoL7jTv+66eAjRGLW4SPTR5eot7XuaJP9w8EFQG
5prLVUTfqnnDbSDlJaPeRPl1+TjECoOxmTCaBbJXP2SUIkGC/Ougqdo+EYfPHtuwy8y81hdKd7f+
vLezgHtu5sKSs0KHDOK81Kvws77m88cDV5nvGDw157Iy1IXyJh7FJb320VjeP664mZXkRQHoiQRj
S+JjSdDs/T1tpIKvAwVEgPwiKdfrtoGx7BKClEKQdt0K5JHjjFSRXZ8PV8Ts3YUhIasxl6HsT9mT
oI06znLJ/2nvLAPi70mrj9PiDxCChkxDalPuvxTSw6eSU+DyABs1FzW6b3N2dC7WDgO6GmZenEka
dw5XY7yP0TKVEkzCx0FYRyc2cBQK1tJ5zn6EayQyWWl+HJv1kRe4ZcRVyH42qfEtTamQLKvwGX7l
yae3G87cGz+nKGco2vWFoZ/Ihr5NlFu9MExaQxs/7unaDiAbVUOIhML8M0A81IKRdDNg5ftcJV5g
DmzGY29BZtorKFb/s/oXnQ89T3ChRKC5XfmDuBLIaa/KOUr7m+GMv8xf5mBK33tXo/fmOUw+WROm
sdoPu5RlZRrf4QCu9P9AjldwEYUGRt6vrCVl5kvGsNsDut4WR9Ojq3aBPv45Ur58l3TY5iXHVwb7
07bSXBzV3l/6XucA7Pvxx/c9n5KS4l+tDbcyBdY1AnTQx/xZ+p/imeDoIPVMzPnrUadiOp9Zq89s
eaUPT2qf78zsObAp6FE1gGUv9KtSpXd3RcPLDuRzAvFOL494C48jycgkSS+2Ec+uSKw3cUr0rlWZ
/u/HvopDmFuMkJ49cdGXOhfsFcQU7n7iBt8tezwAM+YydUxwqkXH4fRLysKYpw4vIDGCDFqlKzfL
b2cGVxYE5wxqHXUZ6cUbvGNAIlyQyMyAzEhuP55tgSFd7tXyOEPFdgohWvCrw+qE4RVnE0EsuBTb
nZPKNGhLGTrY9tqLGqjT9lw1J8SsG7A2jPNkhHpeWCJ8OZzSGqWQ+T+swRsp1IszorZf2JS2670L
FinunQX/WEuyI7PWvKKPsTnq8LWb4oXSvIvocbTew+a+RRVpgVhREE0CkF8VtyRNpygs1thXL4iv
8gtSVvkZHkKSvOdJY5pA1RY/VK7CY8KuQmS1eHZoF2rgSpNEyFDApgwisspox0Mpp2Utbn8z1M34
3wPYO4paS1VHq4mnslzneh51gD6vSHxgikK/tr9/pKlZYpa6m4Bk0dIkdhoan5SbFg9Ojphuzp4C
QxGGuUW5rIJypPqWwWAyJ1B0XQkRl3JtHPGsrxkPmqDTe0j6Z/GYPeyAEVrfkBcNeDLGVbZ/6Y5y
wGnuOhA3kvS55ZaWOAElsIsWqGWmfv4x9N8Xr/57dKq1ryGNj+APre3penGBclG6h82mOxaC/fyz
BxKhNgjyyBM05qwiyY1HzQdE6a7bP3fmi3xb0TosWWAbDuTNSiN+aM9MowKwPSNAhp58LmO6n8G/
H13ZvzbSsp8vdBsYDMyEyGH+C/NAFH0I7bo8fDiJzxsVM4oM+xK+hKnUlvPY/pHl+L77UfKvDH7G
Kr0s4pcEAAy3Ky38AOeZOvY3DwIBEjIO/F526fG316zcyt9gPhf/l7x1vFhR5jTIYC/uTVJAks81
8sX+u58uGFJ4/pINVol6WMRqe+tMjcXdqxw0uqUTOPGqT+nJxRSiuSAX+U+q/uI6zLbWTSlbIePV
g1m/wBd1ywNcqDm8wCBYrZSnXa2uoMU74txfWViiGuLKQo1uFFb5CjOCMnLB6W/NnybVLrgINE1J
D4XU0OFrdRyX30U1PvzweQX+I1mhdlGt1WhBVB9W5f8Z7PMGTre2lFvlKPnf39DSAC5rWeTlSH9P
95PoYuYCSR7du/FGamhdLBkIimMU7f4qReMHWovbxxex0rMqC/v0lYtO2uU8nH3dA40QYsTpMjVz
rqLegjTsEdhc/YiY9vKesa/2GTzasBdsrmmdVm1zpVthTbYq4/UGTgki3w6xRE30mIkZllg9S5TN
oYth4xf0Ova2Siz432LZidHvd679AGbF/eqKQ9zMiIUx2OL/qAAbGCuDj9nl/JAKGc02k5XVX5ef
Pz7DCAkOai7cTKL35a67bGo9CSbjmUy2th66ADBAK5XRQDeMzKJLRbltV1K6pf039d+nZhG3CSA1
vXVQTY4MgyRZuItV1TBnassbcCpVfMW+xGrQclfHWPqouFVZPRZrNitbxy1OCZ8YE+kuZdAzNPlf
ONaTlD4PVU8vLWfDhgeoVkZd7C8G6+loRZ1GxvuLKHljZhZvlQLu/SGEc9GdJYbHve64OE9s/9os
hV+kJ/iuyyR1qktdmbTZp/sDTKRN0ixg/BaIWq604Vfj+oF56GH0dqmfxeRumjdPqKhV9Dq2eU7u
F0Xx+N8h0rxxeHCW3Eb1Gox10sK5ENup3XPWJX+nI60DC25Yt1fe+gRzPlabpP4kEpo/yxy0ypam
4R63BJoENx5c7xQu2z8B5kcYRz+iY8PARm8oFMpjYihFh8FU4ji+e9IFX4TSpH06LPh5Y/JvdZqo
9cH6Yg4ZCkL4Xi1FKiKBQOZbilDns7GFAfDuSSS1zxrH67qK028n9wuhpXe2WDqkeqLlnEaGdvSR
4Pii1VfXPiRBAQawgbxtPFQOOKDY0Gpr+EiwkkSRc22E+JzCQ8GDQ+9rE+x/mp9TH1SFC3cmZHL6
9lfpCFEjrtMwE+3Mkn+YatwgW+N/LBJsU005nJ9pvc7E0yQfNrX6afQFiAC2eHotqXPjqmqvdzSr
4NfbR9Ct3ltYJwzCIVZEyvj4BB97vrhQbme2Yd+aPI4zdAdhCRntyYb4S/kW7nNN+VjEIOrve3s7
2zLW2zeTemJjq/C+M2yJ2B+xa7nPCbk1cmfOd/ia0khLm6Qlq4ox9cCVLb1dhGi3Nie+LkoaLaYW
lVHVr5AkF6nvEN1tyRPWacjhAM07zCxx0z96RzcipH6ZUZOt9bYJraqGt7EsraurburGwBsMy8tj
RfKobODgn2DI8PWujChxuR84vBwZ4YCwHWi5CNUXQ8TR9qKqwMJblXtqVmMEfyyWcwBu8IImoV0G
TptaJxmJROqSbNq6SiRHyKEct97Z9h8K2/Pboc5LpG6pg2xgu4FeGcQzbP3ej+yiZuqdiNeNwJwa
6TD8sTAw+IODRzHi4r+Pn2C+lTnJKquLWnfZga1I+Glm4g4csDCymhjb+dkeSjWx3mMsJfK5UEY6
fjFXdJ2LeeUULoAP8/UpQaRAzfHv3ulMJeIki8j2QwroFWBwV1sBKCT6a7/FyELRoNyT4Ng6QsLd
9SgVQTWf9Fo+KBHkwDWR2SY0Du4zIAxOsbNdpvvCc898olnwuquqAr3YyYrR0SoQOcDFv/5jv7yT
9ut6uMpjRo5lNekaHWU3kg95FqHWgh1NsMrOtrTfwmOKinkK8Mc4OdJRDUK7+1vCua5/Wqkkwb7k
LVf3xtQdMYfOTZrImea9L67mOctXz8hvcUHVb78Mt9EnwZjyxzOzIomXfW935TyO9pYX/Iy5yq9T
AvXEz8bBvJVwBliJa1/4KaP0Qv1RTLPt6cwvf/2ZHzZfR6b/CVMWUtLBWHQ1LTmPygEdRXzWkLOr
V94GGAykD1e0UP+OyQBa+UoTXjpzbETP+IW7E6CjCSA/x6zS6Lkv+0yoDRMdVgHb3riaod8iryMY
Xij7m27zaZcOyP3cZuh+RIbXrByzZmElZuVUUNdTdwx5YynWqRaHg+njoOubmdw2eGLCyTTAAjYW
gF3ola6pyF3gjxojZ//KJwL3176jAmF5JPDU2VRp03Eb/jknex60MRRlx1pLQv6IMKPD7OcxKSd7
Lo8K/ZnQR+4bLPPd7iF3WcdDShVTJw/6KnPV56GxqiHGfdnIfyH/u+Vts5bTftXDHfrZ/QaFxW+y
Lx21uy8Ur67yA9xy00OGD6W7O9oejaKL1aTemjLwKw6WcwIRXdYpElJ4kSjNm66aXCzUeMCkCLiM
fQ3LqpkjuhQOjBrCmokgc89On7QtghBU/YeaV7Lwh44QqAdygiYFTA+teU6JweQM2UlIxt5AamYh
kmS7yJRsJWiCDlOoZgLxjQXwb1aRmxCIZKMhKqksCz58RIdmBRzWDyF2xZF+woaSZgtVlY6jB5vf
5OVwJ/S7nj+stRlPrQLaQA61hQXNxI1G4y59dMP1Z3wO+ucGAxsNLG5TSmnnJ4SqXjBKIsdS8WyK
/lnewh7VK2Rgjguu4zftstc+9dyurvgOa/sN40yaeQ5TsKPbkd8Ms6yM9GTHtyJUcBQdUHAJeI3q
iIlTz7kw6KalLsiKMsV5XyoOz09V7yBldEOgTZ/+PHGC1fWLnJlQttmO85kg09BpV3nHXLwVjsft
QD3uIaMBW2KO6NJXNIBW0FxcckHLkGjVZrBtMpVOAJvznHlLKf8ezZFAy/O04t5CWLzC24UM6+ef
rKGIbMgt2bUn/u+tTrS52MEq2ur6eyqYPJGckPFxqKM4xR+sgaq5+4VPLzoL398KRINphYOEqL5G
S565rkYtLNIz+cweCRZpD/zgEWvGLObtSdGjxZgQD3bENhYnJQPBdp2LAM01Qk02jJX8PGkgN0rG
60F8fMQekFo19WHz8X7VQBRryd3OAaLGtDym6eNiKdk/FU0FJcE//64AZmSe6uJG1W85F3SPbQXH
UzTtkVinDBZVCGQV4NchaLD5i4mHRCcNvsLCWz5UGjlZ41IDE1L1b3Zx7RxBlC07nKJ1sv2/CPuh
E5HoFYFUl7beO7RM8Eqp6zHQaWYGsgsjFTdWTi9J1pFovYh3RZ4IQn/8dnBwHj5yRCFOcQJPjAK/
8XTwZc0wYyv75EkSRiwmUd/YsQptuHXfCQczg1WwGPSLlpY0io+/zLflTE/TD7Ednbo6QzGulL8v
ZhFkENLRqzQQnyRGe2aM/AiLtjL32Sc6IivNOip4Tfeva6Hp/Vt+6EhINfJqogBv2Xsjoi1MZdFZ
/3PIbeDHzxw/+gg9wmpFA7xjZQFU/l3UPFjvGIbgxOj+EmTwPQI8G/BB1O5xtKXogiynrYmVqrBr
MyvkoXkHFx1IEXMO9KNN56VQTw8ylMc7zIYO8/MnhnK4StublmkADRT04ZFu77DcOpOrjJN7+GMM
rTtOfza19v2VrtvcsuDyUC4IhKMXy/F36cJVcs1NVN63X7wMEtid7mrWfyadwlKuPVGsBvgEd2d/
LQDgacGKYIUyTlY56cjwYj8M8vDbzGP/kK85iRrp9L3+cxC/PFOqWnCWFcZrsLGIKMiMjFpAPbRk
5ItRGBSqaqrDlWpjgRL4bSUfVwf6yQ08xK6Hxy7Sd9NGEKA8zOytsg1f5n/anIe20VQKeHHbqclq
1hVesuRMjOJ4mrgXleSyFFgfV8q6yyHwtpLS/fNqdsSn4vkCVp0DPur+W1scf3kyjk2ERN+1IGK/
W1dnD+R/Xt0eNcb6sgfNdF+9yJAtXlO99f8v45XiT7bZX3W7JL4pypmgDIegjcbLEiln7JbQLrCx
YWwWCzDQhzjg+jraMixTaakYqfQaAo2AJY3bZ6H6V1VvUXJDxuy7v+W8+L5SIfvsNzXVew4MWQks
N0hq5IAZzwflqCT/nUoLB4cp4ZanBNkehzmhIvMtfNYxC/UZ5+JfyNF6fZJO1O1huF2mdbX01rlJ
shwI9SZ6qpC9QYlZmPEfNErenO8fkR7HhkfkGoQTY1nHM91SsH2J8h6foZOkxoVfMatQQOI7c0Ez
zFAGe79s8Nj9VU8gXtyBBMaDTTAnG77I1Pm3rh7XkSHii/DdAZzjraQkUdyPczgl0rKecsR1juul
m1n5h+dErLbWeuWMxDm/oGRpErHtJEwSPP2LMOAuat6qV0qQpj455UH0I8txnc8rdvNyDHBHuwrP
0czMuxzZFpGQcdFPrcBMkkXfIRgYF5ohCuoCgsd2HDx6I/BOGJ0FbBVkIRThuOojWhiFdKhVpiXQ
1X0IYst/Ku5B5w6wzQKAB/Jh8HNiEujv/Q/xHVOB89cv0AcGCuH3pGB7+13ggkL104FXnDr3boLY
cOAnAHENg/urj5LUsG2rKsF7YvqLTb2U1NCFhbtBf+yEZGFm3UJcV48E/AJqmgopwCprIjCIN+9G
wiy1QDaxr6gMup26QCdZ5jFTck0ds5LoEo8DKU6YThescR3GAW8XmDZf6RN5+DtLg+8+MknZciuD
emLnkbwmjOm2BrORuxOAjTk7HRO9yI1tfg16OxA6KZjH1F2QeltJvje7J1Z5Q3P9+vrx9lwiEprH
BSVDG90n5Dgn4E4lTa83zZTowQmQ+Kl4DhN1ZMtswn+EbMmHo4mWBCTJXRknJpLujfDpKGjGcAZ+
17MKAu+dQSYHjr/zDzUMr78uzii1ijjShR7Phkexbt1QwbhURdHaDENr/ztZ6KmVvUocx3nD/no+
u1ztqt/cICPo0zkH97xF1bclPuJMIM1kLxh50re37lZ5JTKMg/+p/momzLjqc4nO1mIyQ4Rn7fi0
gnCiKW2A3qTFGzZOtDwCzdw1JUggJdUdu8KDmiR8jRKxGGmt11omhqe/O0fYHpYDWTVDPSDHI6Av
/1EuzgukvqoPRD2Gt6YUUGyBSnUwlyZFl91EYvhWmBITWDajSP5KLHnVD6lbTQnJewSjatObIV91
4HWSa4rxCV1d31bJs4VL3uhEeL9QTf+f+mm8PP7lTPItXSEItzpHE/vplUDg3D3Ckt4STReUwtkj
gkbLk1U+vRD72dSaKSGEYIIBQuDdm62srRUsC2LaaAUsCrVJP8DT0Y2Q7LWaK7sCMBHRYBfcBfDz
11qsLH3ZgucuIISfCTcwNTycAQOwZ1GSWtGownHc4AC9VKa8lBJsetLG22UxIFJfkvE4aUkYNOCR
yiBEkiz6VQYHmH1fMl0y6+K3iaElVuW2y/IFlsvBGRuIElzV1tgQ8NkC2+qkGgfc6Ta3zPquNujw
ZLU0BKT+C3MY3SGDktEkf3BNuvXwk7JMCfy1E8Rnhpa9BYUbIQvUbmf7SOupLXDzUyj5/G2GryPT
jmXazIVIr4fZorMWLof3WpFpqv+oe2jYpA8SRAlhuqNoOsJytiHcxgCN9CqlFJJxHQZh/in5JmAS
YJifZC8hiW1gksBAMw6BvD7EsMY17S6gOEiRplRFOl1+hUIp+XJQ4y1+vbgVyntlUph3IgmqLXt/
5F9irqvJ+6Jdc/3o05UmFywm/vANLrEZ/4k95fe53oDtu1kRbjv9U/NoTKhbZpeErOPWtOzK7Ucl
xPvW1mMUk+/2xZZ80PLmdXoTp1BCkdwP1Tz/G5gj7ODlT5r1x8PsZwf8DVfA3rYzzvu1X5dtqDFZ
sPirXKxdDpnG5PYDRGYQYtMBP8lViEiTgMSqgUVPirgXGYIetPCd2gkQUl8vlQObXXXOuPL1Xp2M
23fw2o65K4Lx8pG+I0GxETPGqFVyX2/XM4+SO90UhpqFf8n/6UWpqvInqiDSep88QD8l3g895+sk
hA7XBB0HITqX/87FI94w+AnOYeJ61MTHo2UfVG1NJcEvJakZDeTV9fm5PCccGCo7M0DFxRA31TWJ
xk1MNIdZbIs1drkXhmrwStvelK1y9xWoAVtUH84mu9H9GLIuqEcP49Punr0rD5qQHkT//HQNLGVb
Gf0OYw7RXM4Qx0V1y0uXsaNm64c4niyiqjQ+txmk+FwUDHu0AnIvqEM+bcjBDyl/uZwIfL86jYNH
89uI1Z0KNhMl856ENhW4P7ocihGAJ5IpRSu6FY5CNJFxAZOX3kcdXd/ag5ii8gI3VKByUg+c1lXD
d1lA5febWKW+YjlgZ9t6l5v/LIi/F5/lYyCsj0+0RCQ+3pxHZ6/YMTTMazJ9orX8R0nTHLDPcSKH
2m8/NHw/6uJujOeyoFeKhKr5EKW5S3TmwecQBKiQVUeGFYesX9bY4TwDGeeaKevjtftfbO8inDoC
L9QApoX+hktwmQE96TgIHL/2olnVjhoJDBr6iTjTXyUXgiFemINsCdewFdLKM1QwKZdo2qqrwgZU
ALkAnISHBBFQYl+IpJEJaotZQPjyGi4X2/XSM1CFKbDqbqgsDEf4HKsGFYaA/IZc1S9D4XJTMS+9
IAMVa2PPyTLc9o8xX6ZS58inSz02lR1OlxsFHV9MDOlal1qMlXgrCHoxzE2NnOLeqGj1CLPJ1e8m
hb9XJZ+RJlbBM/P3aD1TbxO2T/t14ZdsNFJklrCgf7Jnrh9XbcCKlwYu29ZGgXsYFju9RQATtJi1
NsoMlzROOgp0yiiEkwMiIS/OwznVdU6w4cR34kpol38TFj608NHnTEB/NUl4kLsUl2mb6MxDgCMp
nPcmVYw4AuY9XkM9JmCvfo9396Bupr/lNicY/VbJt48e2JibIoAo/FVL5Uty+nX8KUUrUxpO0kVL
HY16g7q5dsKVSM6/ja09lERQpii7j1Qf7XFVFzaB/j3x61yuEaXogiqUFwCYoYr4q0M2bRcOG4vJ
AUOSjqZS+l8AhMCtWqm+2BA1j+t80bFREySoYKAboIU/TtNm7DxQ59RGe3ohINvx187T+ZAwcXPB
nkSBFv9thRgfjHx3NPtT/mZSDX2S9lybHz+QXC+TTke4qn0Viqf0UyILVEWuUQabECjQ3mJoyaHv
5gJfofnVWKhZTeTEMhQWNVK53UaWLxTUNgnO+zzx2zOSkKCwo4nta6EhEXujWVFFVyszVP962Fo6
kjJgXOgQSy8kLzjcCkBPrK2O+fpeWjC4NNrjQo0n1tx0sCuiW9G/YulbNS0hBZTjQkKvJRg6z1jm
GtMPIplcoF5un8d8+jG4oXXJ9u793aL5zrKnK0k0SsKowW1vL/MGNnLGq78/ONtRReD2lBA9HRBt
mLUKSqTWY4EruKrzFx+y8KtpQ0/UfVY1nmT36Inmvu9wX4YVH33aZW3I/BtHihyIRWXp2gDgZ11P
tnFTjhh1dDi9oU8grnBpELsvRrjEi6ajM8omR9BoUXrjtlB4VdHRZbqTFj8bq7J3hE+OPGMxmUfa
eMAtR7hap+AcYsirXqBe1FSx81lw6dM0FC29a3nTy6WM5aK8ByJaazrO62gqONo0UIq0Uh0I+T9a
254x3koV3Xrp4oCfhsB4VU/jrhjvibw1RigNjwXNaEUroMLAyeGjQCltqdLGbOSmDgdvam0BEkO6
K9d7wIPBBPDsperAyIJAvdbghN19iTHIV9z3+UYAt/l6+D3PR25dM6tn4jKrvU0Q8ubDOWsxc1NE
WdE8+pMKFKMAu972A4zwoE5b3xbL9WucRNnHtBciIblRt5CMdMUmd0wKvR9iaTfhkQOyoA1NoE1o
HKDi3XVa7hHfaKhI/nxGb44LP6cjSCZmm6kY85y0KSDC8VF9vZxI+AknN1ud1tAnoG1hE6RNkWSb
mniNDBp3T2Tcf9KXL4oyyUYoUwDiuSu8FELSJPDQvi+lCjcSnEGVwbZP9vU11y0K6wOeJ9DLkL6c
cdivWQvJu2tw/P1RB55X+turMIBPyE43uc/HnVWnIOjy1r/MqhfAaAZGF4Fe+Euma9wMFLzj3pGC
hY+BeYdVsg52RJvG0MIafbEVoSt+WsxKrWZQc6gSXZkvaqsiqm8WbwgCdlAUI1wJvtngO94Aa7WA
/yaN2XwmDr4dvBLgjLmQLxVBox5Rs4PIpx+4mvv7og4kFHFoT46x9yLBQCNOsEQ4X9aIM/1ts7Rd
bgkAuASvUMV7YjykujWoVbRpFAwN5pxhhet9oyfA9CDrXqZrp6X2B8ZTQkNDgv0ew6A9tGlFjpQc
Eu1EAG1X4J4K+cejgPfgG6cX2f89gLp7A435Re2zCu9TWz/M7QVSKrwwne3yc81LkU2i6xbUriCs
m+ZuljWSfU2eN3M/+nvkjdtaeFGP433OexZapw6QcuzFaij+gpVQT7qs6pVBf5YRBC/sLyaMl19f
ye5JP8ia7zH9g1dBrYqWQ1OLWZDfRHV5gHbMOT0YFpGAr7gu7QOj6Vq+s7eKIzfN/+mgIiU5QIXB
Odr99GFd/1rhdXwvu7CdL1THMOvVg9TUTdBY8uLhr29En0L0/gvYnCfQ4YJUMuTNVavb6oktsqeB
XrXFFj2Zk0TkuBAYI8WuHILItBpYTzQEmDidO47XDBtR4kJsbum/DECJ0Sx4zYJIx3KFvfqC53oY
va1fwWT58nqxMOtWYLtd2vMBFIfPWoyOXBbISfUJF6Et+aSruxOWUbSsMksMdI/BsSvZi6nR4eY1
kyCHnNFvO/cQ1AM2Mm6Pb5x2ma8mD/IsawW6nY7DDh8gIbA7wwxMGHRJwVZ0OMtIT96bqqgdbT0C
Lpqq7GkWIjpeQsbJQGCeif1Tf0eNvSxZXCvGAfQdGujv7RSgh4AY9Mq+R3iYlS+i69j+ZvCM7Z98
eZ1P3CzNAJ4nG6tzhId+PwI8kRvkDflaHyOCMqPhs5/V8hABWXmSeGkELOXn1rEguywzDLkycjgX
h8g+ZbGZpV2gl4gqhVWw4t4m74wm3RrqVIzWuQB1K+KmdkPPsVRDTIVxQqeXmfNTC8KW1unvuTRU
QU2OMAtdNlCavZSuIkEsSGLhajwCf29dgjpgG9ciGi3VdwLCCq0PsXTtlLSj49+n6iSw7hRVCLfn
imC9IVrusAThBtmUtOPSJD+gOFzEYYBjGFf/8RaOuReRVz/0d1ucHvOL5YBi4AHQpQ/GEUBECFwy
9MMbEtiiBrvXqhfiE4D2G3ofynkRoMB1XYOePh5DQZUHwDo5S/tm9QrYW18JlSBlYPruHmXq1XLE
gA/tXf7as02QOP3jGvewkK1kovnxp0guUVFLFRRI3QakMryLRc9ikfT3DVJB1NFWDzeuqeQ5SPSP
AZNVbMIALSG3WKEeOd7GfZmUGi5ex0HPJChg70wP+TMP4weYfG/HVcmvVugGCm/eXk6fzA0bBWwi
HINFIQzbHi9o8vxpu7mUONlRxVsaCP9oB+WqZ7lAWGEOxfwXnWKIfeKNdTRLDZ7zoCuoWGkgp62a
VzoZf+jQW7OrcVVGzvomIxgCPMWmeODLstiN+nTrD9V1PAtVgDWENLxsDuJ9PD/uCJBnYFQ7JpP7
ivz4yz+78q2L/kMU98jABLFW2xnjSOC+I5FdYc9zuhRNYeRMSt+xUxDnhZxko/7tTXpdawWPGKV6
wAeKXj/p6jZeFP7f+U4eqzFmgZuPrXL9toNUCgsAfTbd1OCsvJ2ZroSGQKWFOJ6+IcMNJOcvQD1V
br8HXEMucT/2GwzzrqW89DWyAAlxJcHr58QpCdb+9g3/ui7bKGPdn5IeVZUzfqoOt5f05SbsSum1
e1LFw8rEMinx1zjSWiDbGcMjDTqd3wrdEChwRnwmXEu8lf25t4T/TZwTchPUIFCxO5amdXpIodPJ
q2MI6+aWladbqwl+9GxcmPVvjmmlJSmWC6bTpU1gPVZk+IggxpjuNAUyiw4KbpIMooFLYhg2r5FC
MVlILVg1OboUaIc/0/x6+BDSDa+aJerfyU8RHhHUUVgOooYn9PJUiPW2s9IuiZPFWIC8Yu61OKcD
89FCxTAZIsOWFlUXsdg3OV7G1LpBl/wa2adqpRhTlT08TgtlJcdgUI//94VekSe+bXs1hjUiA8r9
dw0qGJ6WBFULnnyPAfRXy+GLC0bBGNR1qnhw8JoPoLvy4Ad+jo2OLDoZzyszdjg7NSBZm6XRSIfT
13tCRmN4c/nZo0Pe30QvwqTdIldiGX3fGooYpqdCR/BRFSP7sAhRrwNZwATIoHpwa5uKBhr/ztS0
yPTWJKeJMh/8/y+uuPQ4CZpkhx8t1tmdjQ7IBtbnoPgB0D+GIuIUG1Msj8kGPtr/78iE0WK0WQDl
FEnlrDqSEN8bs5+lMRjvaNsS5Hucsmz+srljGAvVVPAQRA9Ec0Fg23dPvY86NraLfYBi8vXStXeU
8H1TMSmIr/m1z8RfvxfZzL7WFkxWGrHVHRlAxfuINdG0ARpnyoD2IwKhzcgluVEoVAUoClsWrqt4
iWpVj5YI72bXu4J7MRhk8SlJHu2SE5EXFhgOb2rAmEqdDw+ohyjuc/aesGWdqusCK33E05rgMrEG
SwLFAlpTdujDGmW6t/s63qVzcFXMom86do64+GlCQujI6HOC1sUOGUh5yYfxZCAQuSKrxDf1NeEA
jYQOdbUPsHrPqcYZTa8RmeTqfMwLTyHUHK7OaT02o1NhBrVBAZvjTyeFGMzvyB1ddvsbrTQZouG/
81jb3osZ1CDMbYvsOoXYVjlvERPYtzS/1EOuFnXnAhgCbpRCsjIaga9XEvHXdNlImjhFl0btU9Ns
ytFaEDj1RX5/La3R+UwChFdo11mc+bdggXKNanNqGn2kqvZRYd2iTx9RRkfKki/REd7UAB6qh0Gw
FP9DKwRBCcOPZ9TRravwdmL/+jTUQ+w2oQdt1+hgPPzkdLHkq+08tsP37MiGh/HQ7FcgOz8duiMx
FfXfQJLwaeCiOKjU7NXV/RxTsUKatwEj8TqS3FL4ujkhBh7jZQ/KWktg+GIm43uLSjT5PXAsrUVT
L92ID82tJkgZP2uJXAdAgGhMrCabURXwwPEqhukuvNs7sDmn4EYzzKdDNRJ+4aWf68xx/RyrkRJC
LLwwxN/QHePKOUMX13GaNDHi/m7tDsm5Ud2SyN9uKCZQYvt14q4WDQFHzvFJ88O1FgVC2j2V4gUd
KQgKj9JVZTZTtblrlPHbe4i+ndACuJS+rRmqX5mGKFyLCOSHomPrttkZ8agSSi4UCzIDDwzuHMM3
IUz6d8MNpFOsgjaWPyb6w+BvhpvORB/FSzLmsh2rP8eIuf6M//LR2H23rnYSST1rEU7Vzyof7dzs
0NjFD8UMIb0+S6bJtJn7eDpjmpU1xmBSFGEZberS5vqB0F35B8/hrBpsZhPyUnYlO2iPlpOPXF1f
YxIq8Hj+vgt1ELFxk3879teVyI0X+qoONe74lOi3EgeR+ZvOxzyoPnqQdVSK2m9AvXAHgt+pqwF7
tOyvIxQw79lLRA4Fy6hE5lzm1kfQcw8zJUMhnOI+pqswbsJGUTXBAN0du0ral3QeybnVrBQOOYO2
Zy05uXVG2gS5R6Fu4PtAqDJMKrIptWza1KYUWhnBqUyk4GF/Z6jH8eMBIajCUAdromIfuNrC+5Sv
EO4fe29iNGFl5OsnHKXho+HceaMrtVNAhpduQwsVY1AGWFdPM97QXQLLLeMoFToR1TBrFTRgwcIQ
DGMQwMT36RGj+qAL9QduyWpnk/Y05KsbwoZlJI5VQVW2j/q1raiS7WpPzrJ18ww+CxdfU8ltBm4E
nlk+n+7ogVm9m8zOFC1VRRQwLtEGKEkVbbI5T2h/ew8aVpnQHu1UOHVfQtLtNMAgUyMFOBpFUz3+
//5XLRypavj0s+gG+mbyKLl5vDNZ7loTCqKhe6pGuE1lzLu6oy8TJuUSCd5/3YLoLwhhohr1G8Az
0VGJi1tzP1LUHwW3UBUhJ0bNlDDHeh7LsJDx7ojGV3/z5XVG7yuOUk38C/thKDWY1YzxOyt65+kU
0nD/RMoA1DvGYhLy2YlMfudh2HLZRMgmL4/7J8IFvTsdvf92Kmxixz0XmFeHYGjk1T5mTK1niwrq
gyIMsOQsCvPdMLajEKwSMR6NkhBjmkHIm+KrFSZIkc8QB0Jf2G6vrNwqcNLcu2cq1gaCKq7hV1kh
b44yjqlE2nlV1Wtz6WfTVhumuS/On99D6jpMZBQyk1qRYjjXdUriG+jO3JFemuOnAl69XGHDpovo
arcc601didVU0jFLyBisVJRs+VRYaHghB4daG3WNiM1Ct69PHFoBkI7qIV4E33iPO2M/NyVSbyZD
ZqRhpdeaXLTkMpCfCNZaAHZ4zNgr0c+Q3AmXjpI5Mwd7tHJfvbYpiRHMEgAluq1d4hdc424Hadak
yqcBxTjXQZccCbl2KcidB2nhBxpxdA5laUghccDHPppjJdJdpa6Nx2WIKzSSaPYuNATtsQUhjoL0
qUiNTER8HdpbmWlgAPK4Eo4wjjBU3pOw/djPWqIrxpk0xUaAinqIombhjMmTHpWqLdBZ1tebbAz1
+dcy0Wc9WjwzuIvRZds6ETLxSWlLVY+N7A319PWSAUQY+EmEGqtOwNDQzTpMV3c6bGxB2n2b8clX
AjIgDjJHtx/h+XAq+h9Hi1qQB7KyvTfNMR59KFnfgXCbj9ZWarlKUiUaF/UI0eS+ZC4upaNWbLKP
mXl/JVpSy/NRCspZPETs/WhBvGpJZcM1CRRmezHotke2Ou88ymzqiGsPxrTy9l3wyybsQ5Q0yMml
yhMCjJvfLO3etbY0Xz7FM51A0mywkg5K7Jy+z82kG7u71RMZmH/0G6yFBYMTm+C+rDH0IH350ZH8
uzXD+whxKYpcuGwJ4GudPV247Rrk9iwJYVtEyShNTmF66sGXMn3l4iE5xu4NnZzRReAfhYS9OBL/
Fxpx6dcCUFIE9veymhwPuZGABBDgut7Welsoz8f9nGw1Of2C9ywO+ueRdvTOgcJCBgez+w690CvV
/kq7lBHbTPgSTjpSO1/2hksmMO4wmw0N9E2IuapSMCdG1C6wuq0whFrkDOeno0Ui93jkuqQ6FpYo
TXf9OJW/OBnPn2KFG/sAjrI0YR5P1PUCEq+WojHN2+pMJfe9Pxnw/tfu2a6SjKHqTu2Ha3jsYPCK
KQGRyWfStA75NjCDFmoxqtCMtujMUvHa/nH+0LEqWH/98cRnPEfDCGHTjIQKruKg2aISbF0SJmZL
kcnoWMTrzHQXOXCZ4tMsYSsPiSuCqnlP1geinEX6Mg51BZlHOxQKNeleRYMT0m1uCdwxdbNywugk
bg0uqxIj6cueTloc67Q9JaeETWEclTPxIbhcvwYwQieaVAzMWvv1yPT3lHP4/NU87vOzhLHao24S
tsJNkKjufz+q/0HpYqCR1K66E/bGpZEV+oPcMPZOY4Q1TTIE5S4ttorFIDd3KzDi+VFFRwo/ApNl
fqtjzjPiERzLY7xYr+y9i6Lv+i+C6S9H4D8Qh2/enIdjLKs3FtBJsedM0njP5vW4e7s7733DCYzt
HpTYbxmaFuLaj2fDQsWrHQd5Kok9ra9tddxtiFmrJznF2l2O9ELA2jUbzNYADQO69i2lzoonK7wZ
G3YFQHxOCslCTaqDVsPl5p9SEs4Juc4iU3LiwJRzOJRigJtqgNDCc9mN8yCdumAaaOUkH8n3Tylv
LD7usaGe3mNSp0qeQZKHHKVxd5vlSpX5tr2hcZlMvrt4ezkgXUvd35ODYSDbqNbKAUzypb5ZT/PV
r6v0GwCwLCCMI977XwRKSvooIDJBmxSDYfV6OEDWPtpEErBYVPOxsGtixhvl0aP3FsNpUdLuJyYA
DPK/m0sXeHbOJ1XFB5a7JN7gVtIxdVjHT4RhdXincBixN6OulqJHmZFbXdYdtvdVV3LAxUkEIVNn
z6opDAcVJxPhL38R3oqho1iMJ5vqANHh7q5AvwePn4qFdcE0kHfiKqLfVCQRcMK02oTqj4P2uoPG
WDgCsKSbpz7Ztc2DR21+L8ZnNtJ3glEF3UdxTWHzNeEkeo/ALm3kNCN4Sct/7lLv5iarpdPOFd/+
x4Eujcc2p4w5jxKZwbmnXdDlqD476FRYv9aosHeXYWIdMdVYTvFytaX5By05SS6xeC8gv2X7psn7
E0O0riiObCyzmbHRQT+oewpEKFKdCzAmLCg7e1E3dNZD8bc/RJxdNN4eobd/g9tdz0TaRoFUpNtl
JhicfqwAeKvFZth4RuXogFthrNc/41SfWn1M+VroJYw5oCWacqqTwSSvILN2dlTQPqjgWbQDxsqU
57SavsXw1x/fQWYpxbdNVY+/KGsrq4o0GIH2661PK07oXtI1BnJTnrBlR04YExcisoQ+wX7QfZnR
xmnbQ7y949DYoh5JuMAv9vxaX2WjRHAHnxafyJCa610qSo4/wndNXRQp4/Z38jeAh40dBrstLejk
JNIaL9aVSCXt5cOEKDoyX9ZsBFRKDlk3mGcP0yRxN0jclHBp0a4dWJyVa9dKMcKg94lkDcqNxj54
8nevqdR9+uBuHv85PpNL3bTYliDu8Znk5sZs3fX0WZBmh8OZ0YNNnGG9xHIB5OFmc7++/fxBlNgb
1rF56Jgg7uzDE/XwPC/C7mFte2MJC37RWSqWJQwgsXh0mHtpfPD37xiwVmALqk83nVzygRRMCHc+
rjOrvUYD4IAY9cRMgSKUjWcOrUvt+O2wwXQ/59zE3bBgwoip8pcK0JnJQMXzxD/wra52++Fm8pXS
NUbBd4LoXt3V7K3nWhhced5vuUMmgD9O+UIj/UfgL5psPHesAvv9kzsBMM/4JmU+2Y6R0jIaN30c
V4HR1m3r5qT/0CJzvTgB/z3k4lJ59ocD87XrvOrs3vawigJSzJrLmhLdWL1Cdou34Jykki1wueKz
Hx7Y1iwr0DaWgHCeakut3bY2XtxoLXgaOMKJ3mElZcyT6U+puFbRloy54OkQQGEK+wxBGsICpjoJ
XOwVEzpvolGjlRJczr2FoDFjYHUoMEFip53BmIMnnP0cYf3vho94zsnNpsqM1MbzU5uAed1h0GgX
3V2Wi0BI4kDCQD/k/FUG/USTtEVlnGaiS0Dbf3t/q+dQOjUUWBvS9XHcX6OBdb6IVgLtx39+VjkQ
mx0/Zp/01acB5Zlj5omQaGFvn4JlDfhkDI6JKpwPe4KwNDAuCGXwIj3EHEPZoQcs5Xh6k7P4DFlZ
JkvGqEGMsZFej5oKDjbLEN7/+d+1/Lbt3i6P7MtEroPwWMDWaMv2YV0SkzQIbxF+5s+pJyEgMNQS
JjhIo4r+t3GPFWPalz8kwx/OMJHnrIeSXaITOTq9OKA/Vkn2HUcQ5ST2wxhJTMmHPIOij2tGjcGZ
xZjokoJMi23EgTbFMw3PDc3fuRmuO9MU+cFTSVbGOE3E0mtZNfq0yA3SY1SLt1ykfh4bQIKVlXRh
12m/a+AX0+2L1lZiSBvwwAs0p89UxJSGjvMUO47d3BmwAfLK7rh32Z+xSwtQdMQfE/mLq7LPao3k
Slz7D/stEbYT1+lkSRtv6jXveH0nTykPm0Iy9IFUDbnzJRIHVbGYcs6mI/J8MtaamiBwuSeJ5HYD
QiF+B5ogttGHtcOnG65kFlxjsJm0Yicss/xOmjWP6CBlzw/TYij4wUNd7ZohBupMmG7azZ1YpFTd
Znr2PpaeY+MqMYloPy4H+rMJ2k/u04pWTc2OU7zPwM62ZMfiUxllLSvpdSycjScG0xyf5VUyY1XT
ylOWdFrbZoOY6UESVRRK40w9rZtESsN2n8wxJNcR5j/Yh3xUNleP3cstgJJ0eTKlXjSv7XRR5exp
jTjOSchHgk8swt6yz5v15KsqPw==
`pragma protect end_protected

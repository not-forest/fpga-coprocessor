// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
JVnCaxMldmysQB/7YOJGh/RjUQvUK5iUbKuFAoLLxarIwMbcOq1Q/lBbvCg39Pj2
J2DY7aBPI23nflaoneA9f4bnNuNnpZnTuQpJEoiYQrMm9LRDsSESTHdwfrgKODZg
dybYOtBt/tGp27DFs8LinwHcYad1RHLm3qtf8ehvW33cpull6BbrHyhZFyIysZ5l
Yw2uG/1CeXSrGUI70rUPWyR7ll8ffsZafXMh55hTY3iP3DiuK3Tnfe+TCVxIs9J4
yc28MwBcnjml7awRIGgpcrJbH8ESzkveGdahQBM/blh5c6A0bJNKMnSKVfwP/ECM
xEUqbi9b/1IimbH1PAMFKQ==
//pragma protect end_key_block
//pragma protect digest_block
V70IB5656v8X/mfxlib8IMsM6jQ=
//pragma protect end_digest_block
//pragma protect data_block
PUOZVgrC78CS4kSayEgyfwjv1bL5KGVveY+f8MTMaUnlPfzknoQfNKRlgnkM5/WQ
3X6hBrVrJ/ZpOURGJiSJ/JZZV4SEGak/BPLPx1qh3OV8hEwTM2FrVMEJfvI8itQd
GDG64RTYv/d4sQJZkdJgtEy90Dsj0ln1QllC8Fnq7WQVgCsjO4jYYXB9ROVw7J0i
NHelYS4Qj0dk5/NNsIL4wFo5pGmawmw7oAcd6fW5054Eujw9EmLiSyP/okYXq6iQ
9txQS6zh82x9eIit7u7Hp7XB2o47KV+m8Qbo1RpWaLsaIyyY+xdVc3x8DZE3+rl0
8cKktPwFzBXfgRbnPXyEXfLcWDbX6OgFdR6MnOccJzcmq+zwErZ/xn4o3cbuDeNQ
OkZY3zVEqVTIrZNyM6iVmT0UilG+Pat6jFrdlrc3pKJnNYCvFTL9oR9e97+PaGJB
6hj2oM4RPZOyIoYUN9P85QjB7N96MNZLSrmlthQ2ZpMVwTBUZ1vKFyU/ol9/wOn2
x0uhBNJcZDN7Q2Gz52gWc/6stL3UT1zkENOJqMWkMJdWur/BVKpagzWPu9OMTUGy
4VUgO8pLuTRwRR1jXQrL/SxRuqrkucLkKSYIJIBEiCN9dN2PbJ4YI6nTYzIqMqeY
5oZtqPMMBQamTHuS8mHksAjR71DmFjT0NV4159aXNf4+ipo40j9Z9Dqzzdak0QX7
aQuzPnG5VC/7cbXtbwvTLL9YohZcspsxjkGartgxlldeN1+c5cpyqvRR5B9ybHGA
7bD/h5zTdAEEa5gd7IGLPepMhjATtA0PhNsH2okSahwECC5PsyuUl7pcvt4vt+h5
yDkk7T1P1R652TU4a6azkrDWkxTxigH/10Y+6qVY02Kk9ks0shacE5D/dPKWPVme
Ej2qgIVTsRn8C7HNRjDphdDqoqZAjg33wIautrOw4ncney+4R4nbu+DouAlYC0ZX
XE4ehxG8+ANyxBdqScv1J1omiObsKlxWOejaC1zeSdipJD9PbOuLMETJAFMurzbk
J7V7QvSUYc0OUqpHE8T+0dGfCifLk4RoY5k0y3NTjhz4IPMF+KC1+a6GD60iGFL1
m9p+G1UYe9AqZplniteqb00Z9j3s3Q8VI8ndvdiuLx8YVY/5hlhOEb2rR9VAhDzH
slBbK5sPiahnbpXRJUHanPof6VLCoKDqtoWQb3S8G7dVntLQlduJAeSag7Hases8
vRNzN/9KVUAaD6v8CAM8rl4fXXxFJm0Yp46QVjQrwbfnc7cMRVIOfdP1EPlXQiD1
z/H1F2dj5h9umMGsi8hAO5YEddDtxXi3FIEgyLu/j/XAkDNfFZZLw71/LSfdVPIo
mCjZnkGjfyi105b0BtPL+gFQNJ15yslyzsxJlQ6HKVp3WV/hTgzdG0s/OBGlqZau
3oyEO/Rh0kRBmWYrcfEM5SoUnHrt43HB4QqJdMTKfkHnk/lcPv1b+s8vFQ1IF6B8
lXTXA/W7Iq5XMX6rLHZPA3YbQ0IytKO1qayNx+8HqUpagcHl3Akjc4ApJmkNICE1
liCtlhxUx6LrK9CvJv843jODTo/EkgHKh7bpJGNYDo9EduXqFoBSpYFKQzkb/fUb
yoLBi96nqMLnW/L/ple/KTD6PGNWnwM/IoaHTKUzXKfn7zbU6R1Kl1vK6bH9H9xP
8FNuscqbTTu0jQrRHVbJPscsaYDHJJM3nihsxDiKJUuKW7KApOoaEEwmAz/kpgN/
BgFsJ3K9MLWc+KIw7GHf+UDNgYV89Jyrs+gKcd0Ya9gTZ0LygMfSj0lerN6vkViS
1eY1mg0RxeXYqUbo5vaLoB1OYuumJAampyaW/EkUuomGWJyi3BvdRlj0+sVcaNnv
Zs5edzOFfskXGfQaZPktHRfa6C9b73GxjeMeCUvB4gaWatd8B+b8UMRjVvR1b8tO
Euv8gK6ON1xVaT8OqMsMTAX4EPVxhlPxHFUJ6i8uMi2uWCBtYyy/gul6lRAN8CqG
CoayAZJT7TqjaugSxKO/FnF9YXq2lwuC2J6Mm3wpR6G5ch7IUaWZjJBNT1HzmH15
UhFmDQOqhGXNTynOdnfh/bb+m7fzE3MhzYjKNpHp+wCMYpFn6P3b/H402w7jNBTx
DnbjOrZexHY+8fJD4I+xq7io1BFQsQSa968jLPFUPgVz4CjViwn65Ejy9Z2BYI22
ImeybZH6qkT3nngIHJ7GZeLTGfuP8j2Rl6Q2Ek3LJPHXipigjFCxPqthms1LSJvD
zGA0tsEPJ2ouUAOgGolZMjcXA497KcyUPzf6fa9smBQB3veCOiMOLhOybXYP7y0K
F7A1KGedQ7DRlrx9iKD1r4ifXFUDBRCNTqJutVYfZV/ZslX5cnW0/t1EzDScJoAw
MPP9kxYSuyA3z1prMRAhk1xX4VTyL0ldVfIjxDgMYaUI/4r4q5i68ukKQsNC79/X
w2IQNFoCC0FG8cp7qHH422S+a9Kv/NNbxOKyuhSYCKKerx8/tX+iYgPdk7V5+EOg
XJjkCCfZwt8Nrw6jrgKg9Oh3aEoUeAFeU+mjwv9FgX6SUESv3DrnmVQcsdbq8kOx
iUFJ0pLo0R24nbj+WH4PLcpkWjtqB3haHxNB+dW6zKY6Mnx2tXJiIpRe2zel4jcc
UfHVv/XBbxHiqLFbaWh3ZtVUYEMbSVILmDBVZ9DHLjnEQPd7/k29qp38vpIjxRrl
9ZdLNQPcecmx/PRFVU7fGdxLgq0OJLzpB+ylExLpZUyEp6znZFtCQo7LnQ+cuUXW
8yzZzrV44EDofkl53mbS1Rn9ctPB8AoK8K8L6aMb7AgprUvHPH8irDyikUSs71GP
wtT/rco9bT0x0lalLr/0suTq+RUuIuwLIySwlAn2ubFJL9B/xyTwiwFFQfI52OWm
mXrL9llmKASpd5fFsUI2c1Hb4/Rzv9EPjP6owZfEw4Wi8Lc6S780IXEjf9EZIhg/
GPqFeJBVQ3T1ZBoJWG3PQXkjE7kO5tTXk+Q2Kqwvx8NXUNaEE+m92toLl2ugRxPu
lGf+a6eQiSgmHnOdXA1lpygphRFBEqcnKsZOYsAzQUTlUHS9lMEFEHrwBipLIPOh
+E2FJUHq8oV8Nxm3JaCnfhxWPvJU6ObMnGaxSTAOLj6hw9az3Hn+qsHZF1X7Yv1s
XCp/IBL5WJHRS1zduxP0fuZO0EPx9NJ5nN/DM/EGcJMjhWoXh8YPow9p1/GbSicV
Ech0ITwYLd6Ogg3iJ7wiVvIB80NzdFlE2120ib5UMG21RvqC89LwGm5pslyE2eaS
r+TcYvNGGKkG1DhjbrLz35Wm7sB4bSdxLhb2gpuDihWkWTG0JJwtpZFSrWIYvySm
Uw9jcJZIb2SOnNd62I0pAiLvv5fIKelpvPRh48maSqBDpsva+LT0/MROZgNO6JhU
8cjcoq3pnEgCEvbzfydohHkpoFZc3Gry7VPa3WU63F6xo1MrPA0UNQXzmm4e/TKk
gLkYUz6Z5foZWsUPrFymnK1h61RSjiTGrC/qH8WZnWz6crbJe05HRYLa/O7Vlr2Z
8ZcFYdW96XCj+74WiQ03alNIPsyEjjxzie+qYvhuZX85ba4ja0jrdtD7O097Lpsy
AhegJ6DTGpBLqHex5QaFAek2ucARxNuD2eP44DsSYn0il+09eiE+BFnHpgwVcmhK
9rW3WmqPAcWQt3jmhGW43j1YjmC/4EQrLhDuF93GOjBnUCgYRukvwPa8iBXLF+Z1
wOrj71QOwlc4CvfGUP3FpL/y0Duz95ggvxAs1veOnEF2OyyGc8JHjx1Imb6xqaaR
41RAs0shuD+FDUjJrC73nkRNubUfE3plCYgFeHeirFIP7GQRaph4RANg2noeK+H7
+OP8MhvaaeNGJPodvy2QR2ZLOMtgN+G+TpVcrrWy3Ntww/9o31g+jfCJgJmgBQdo
Vbx0YUXA7EdiDu+bpbRU+W9fgk2aVCoHAyPwsuGug8kv1/eXX+Hp9/nIn+MnYRt/
VvK88E5UBomGOdhhd8QLpf8kq0gK56QCRtuhwjp+NtocRkqH2VCHKIkCPcjdN2p+
sLawJlHkvYbdvR+u4fAio4Xu61/XpeQV+QWk3J6TWo0T5YoxVS03sF9g9E9l0NOM
2KdgAnXZgX8NO+AUGFx5H6NY9dukP+wgatOJH4ufSFETPv5JGZdHI2Vn9TbEosmV
Uy4z/qoRhFqyxOvuyNmZuZLAO/CC+vy17KGpZPogVsF3DvHKSRR8A0YjJSvDcwgL
TL+E7ZjUQ1iBQoYy03Tab9g4bZTdixBOWXyN4wqRDTEIZty7AgAYfxokE8K8ON4/
v164l+UePjeLdLLCkBhASc8mAXu0UEmmQ2cCMQjaE7kg1Kimfa5cocmQ7QK31BLr
+oIAA7M3sTBmsdVxv6LkRdO6H/LmFQPLNGQEjq6rll5MZBRy8Ba60yQnlGF1sJlo
N3+GA9KrSroWtor8bpfPKEmZNMsPJDsSG+YwGFLFfnEByNB/E4WtYWuGBZMKx3rX
QHToFD8XH0DCA+UI2vmfEeIqgQGPuHYS+lggPSzR1kxiEo8X5qiJ4GSNbB7zF6Et
MkMoRVTLPjWjNVrfmIgJRQIxGvf7vcSIk5904wI+CvMwES8+xtJK54IsJZ2J6g33
EgF3jQv4WzufzbGKmsMziTxLExaZPdGBovJ6JLgHRbfd7YfAOe66rjhTKyaLfvDA
FvTI3zQcZ9HaXfRkByvTq3HlmLybBq1u/j2KynW/FDA1sY8uZIEN7dHDDynnGfAl
+0nmg4BXvEiMeiihuaYXwYlFE5REeqFH1mW7jSg29DGkCdP2AzS112hmnKe78Wi+
3nt5xSe9lDHcUohVmuyLs/TLt2HZy6Pmrf6hoIxMm7ux2jtU1r3In/c79LINq4Sn
OsFugaGLAeWTfzaxCRA0/azWT0b1am7PCr0VAsKGqunlXWz7kLYlWjfCQa0hVURN
7hIPKF9MasCKVHEQ2FJAEZmgYlmbiOAMg5+kfMqcD5xYH1GMuWlDZaLfCjRS9cM7
g4x+Lbb9ihSJGTHuEipkxTAByBz1PcBRjLMOsQ8h+QvePPReKIEOWEl+oGE0tokk
KV2+jCbgFQvPI0UHp1PtNTv+eqjDTltkcIbm0Z1fbE3htY0OblTqnZEBzqL7eQP2
mD1Ng4YnqIc302FsBxHzZ9bqpkOSeWyI+rCJcSyPQzuMiow3txMVRrytDeqvStOl
relJxfvbIvsap1tu3AKeiIC/A/zk1in7DEuiv8z4T6E6RgJIUVGBtDLPo6zd4FaP
htR1xXElVfkDKgimJTS375yiwvGLVz3lFX+1kqMWEKmprfzEcGbXwJLfmpWHlfCl
py2f1Bg3imy5fReMNhp1mvuOKOtqq+X1LfijiNeZxg66m0dsfryOkUDGXwZJuJfV
jrVD/7KcFOuazH9qSR3Fc4qMG/JBHCjCWvTx4GDqv0A997FJuXgQwTdbuaMM7wAg
7D+zKxVflqsH/OM7hFHLmZpUiKec3eEE85GXeVQd8QrLqrOlHRG61IEX9xW3gOMi
eyGdaW0wedd5EPbHRadVMi9W9fpiE+d/UCQBSeOSt8ykayH/+SA2uJMh6An55yVf
uQ/2C5bTxhh7a1Bdt4STtfQpG/4uHualyluz53r76NIZh9+DhHc4QpyUWiCGKEKn
gXjTyfaqqYX60J5b66Vjlkt0HiGHOhOCxIVS2viRrN+l46Fpp8vy+Q8ZE4Newf8g
vZv44GVZ9Armg6oOltb3GywsT8zQMp2jBT4f1P/K5lpcCuIOebQ20UmQkXK3MTd4
9Uvqr+9RVr/2jSWraFuejWH1hbv4JVf5jQvMm8NKbEPo87dWLfX+qHi9zPiEGrne
fUxH5T2ok3rRJK2gXvT10VljlZO7L4Bt+iuVYG+I8Ep/u3LEhKGEOtH/FgB+BpsF
LnSPlnpFz8T2tSUJcgkd0lIZBFjgxbW2Wtb/FkCIO/hYKllBNm/nzg6NojDaBqK/
Z3+rigvwXXHL0yCN3nV8q+FHvaj4rxbzFn0Om5w5yuSV7O+Bz0P/qCoz83NNIpy8
yIU5YMIZ4ApuUVQYPR2dlPMS/qG06hNbHbGd5zv4hiVKgfiNJozin77DJtavQf12
2zFzv5Rb2QZnMWQz56NLEDokRDvBkAXs5GbcpIqUzMz3P5We2Ly07UeG+++rXeuH
kmgcVVG2BPW5ZTkwmrInHuMQ1A14jYdv+2BORtoVh3Nqkwy2LU5kawJ5CO+TSEWQ
95vV+MSxZ6bs0XH9IkxjCGj+1iWDY1xpPFx2o1qT6uEFhy7DGUIO/AFClm1QYkyr
u/iPflVBVwvAqGFwO98Zpeg+xe3v6smCCvXfa+d6UgGOubcEwWab2HieuE7l6wvd
kxRKS0+lrjw7JKQUzFRD0HlfP5Q+DsF9UehENy4AKXHwGugxbgHRtwTuYXJsPBK7
wNusUrf7UCD/bKlKJcA2DvQoh5Cp4rujtFPnbMp1YBNjfRWajoDyvH9o+ZFM4l3H
TM/rwuTtkNmF66Mzd6bttqJG7IDdJWKXVhGkvKuNaUBh4ldTouFPiejV8mFrykQI
PuSbWJr6VEnsjjZ7k2j8kF1mGGq3Gv9RrdXu0RnkQSuslKeyAd5HyWqS7EO7fd9r
AWHkPBm3jXND3tRprr0cmJso84mXKCFKNcJIjbFOFzE/JYS32t3YJIgZvft4IfOJ
39nrNLgX4hgkStIyHB93Mkt7glpn4jF0KmkoiB+C8i5Mj4T+pWrY6xjU77mtWs3Q
yZygAjOR8Evf7H3jitM7H6SzOFO70EJvsTmyRb/jSfsTArrq5uLWNmDtSD/RDvyq
zgADi8p3Rk5FKSoCvGZfeACTZY7B+0nFsb9jOWTFklO3STZzb9/JL28jnbbPKBZE
Lv3T9KhIqHi8nEySWkUY+wgCvazXhq3O6OrNFIH8FKdidWqUAPt09HCKSPSnzDGW
PbWGccyl2SE7ZM2960evgVScHHzKFZwKP3s7w6HZQoFYSPJ0zPSa3xyRl/lOWaeX
I22oPPjxifgy4m1JYhvZxb1iEkHOXirm4bBJDvI066h7RjLACNbNJNmpcaKx5J4m
cgPO/FNEO6aUfSlz6tBggoEPiq5Oflpe6nGRKuLaPHxutr9qPf8/NQxf0b7jGPeQ
STpUlmRIgyKnYgq2KP5A7KBRBdT9EKDtQYJcPZaNNfdFrKHod2E4sanLI7Lz0zCt
V1m/0TwMhgqcNkn+g/ef+JIWO7HE0n7AhbbPQuh0flwlN/HRSPWLsLi5g2KjGW3T
Ai0h4fnQxQ1FhRJRkFf8Y9Tzo8Ofu5C4iF0ofwtviU8mRxoJJzT03sXafnAqi6TZ
39aSkcxUBev3M0V6xgBqprqgVk7oKl5NCM+jsTkVrIT+vekZOVRQmMbfsbpzeFWF
yxTPBtysggr7jYTrEjGXNCd2lcLrM7bfUUpntFkwNgzKiTb4cS01mIys3BjNEVwC
9/8/kBD03jKKgbBwW0WD9B/ThEGywye5jKLvLp98bE/sax0q/gkFSeKMuyMxuXJS
m8J9Hibcj+3iWfvJoGD0g2gK0mSvPOEFEHk/M8OgT3KvQdvaBq7F/tFsUNNtNJNG
c7iuICpP7ICiuXuL612bUNR7LVXWKYDIMjuYxJl/uJWr7QGM0xz4bWqAV0Q5kCvE
lMmH8mUYPTyap0ULzE+HjKGtoIpYg+LNFtER/26eLblKWKeCU/nZQsi7Uj5Cne1P
N2J+M968Alx3RnCefftiweNV1a1YMUtP2st1k2Xvfd4mZZHdx0J0PfRkvZmSeOHo
EqfOCUWcQFOVBY8JW6VcIlWlaPPRmDprjrfRisI/Mqq+vY4/QFq+7+5/6VBOsSPc
cJ7aiEGpgV6/MJYuLxzHca7H1tpeYOCWV6zHx5RvsDcQkIjd3AlRxq5s0AtX/NNb
IsTCwWlNNddlcDvoivNHuFS2ow/fNopL/oLoJkqcuFFl2H3g0DOzk+FcOxU9K+s0
PcuMkPypz9qgfH5FNN+zN+U/3LB2FEg0psajAtG8SJ0nehhjfca5MCfu9xvLQ8Gi
LjS3cMDuBKuiQO0gFrYcXyWMVtp31Y3r7orfFWiG/Cs/bFPTLq0FMCErrqvdGaxi
UgOU2Vi2pvmUSL1R1GcS6Xb8lUremaQ8YYDHtmeW699RsdULpDmVlQawBY++mjqQ
RRM/nqz6XgBX6d9YJ9am6JpxWFRCh/G5dcnga9TIId5R/PvoWondng9Ju5cExrw3
lyVhRftLgMguC+eILibUvFRvU7FGBiD5B015Z2Nej28bVPkKycoWFc89SrqRKHbt
UsbJgwm1ChX4RXooifMIP5oJON8GPxRN7IHl+rVFT172Z8BGEM0QQ4pPz+1yemCD
aeV6lhg7p6XW2IK+3k6J0QPxJQRIvbgFc785l6bF4SDYISlI0BPui4W07Mj8NR8w
Dgcc36x3dlHa5zyCikM/d1tlJGy3uLA91H+Bu6U/uHIcJkd0bX4jaZwXPagL6Au3
kJK+yR3xxJ0+YxuQLCrZbU8K8TeYUJwFst2gG8Rxv2H36xS3+a76hpgioCYOaeTU
nitJP/skIz4TW6JQHmY3F0kf1YEV833FHN7hSZ6wJYtbEvU61S+c4tpRT+6dpVbi
UByJ5OSzL/P/WFvNd+a8w+PLE1yZoxzZdvyx7E5FNblqIxf+xqM3dj0+YXCba6jt
2zXNXLJzwb7Uk+kf1nZ8mEdapxPLm9SVJG7AFUU3lJhgjEzyv4m4rRJ+LMaWIOeK
/Cj7F6dJiL4ULDOl6pL/BqFDbQ1NRkxRxb6KMYPW/uur4M2No5Hyw8JJoU/NwUfd
TS+z1kgmIwJmbWAL10UoBTKObCOELZCyEeeUUwRYGGbB4IKvjS1MJvS9lsYI1FL3
mRE+34OVbNQ1oPdnApCiIGq3TiKd9VURJoup/hbBvUJcRVOKbuwDm/ESZYxb1/4R
o1Wqs7fVA6F2Jg/l3XbOClMHxSToqKwwj0AJTIcsmizdmvAh3U52UwD/T+DIii8P
Vx+W5lbbB2mIk3fbl5Oj9eDk52f7X+FSB/RtwCGbD2Ha7uGGWYocJxYPGSLWxECK
rwPKi1bJpQ/wu8He4VhtNctem7Jq/pHiOXzYakx2aAgBNzSEbKAWGaUQtHmS1eo7
UH+HDgJX/B/gfKNn2zy1FEo/PpBYrJfNVaLeplc8ULW+lvT7/KiQ1ISP1JJv6KJC
oiLiLH206jtUdtih4XLXD9qRujsvYqUEaA7003Z7IGqUF5E/HJy/vwkcK9i4ZqZK
TPho38u/ehVkDpTYoLkVqMM3eiCZrDdJkQKLJ7bNghvKcWhY1ygBRIbeux64Q3Kf
Pn2pLHLB8NquP+K6xz1lyw==
//pragma protect end_data_block
//pragma protect digest_block
RBt0tnTixQWrlgk7hRhbt8ug60A=
//pragma protect end_digest_block
//pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
WcGoUOO7TWiwsxlnn9yNFgHaWLuGVN/oDLH5cDryREGeYscMqB4GDMdw2/H7NqR1
4fL3eR+q+n4f2CCO6+4wYpFyL8mFiBLBPQ/KawuZcFYZqChG7W8Sc+uSDHUlLQN7
IVoXB37l7mtFBEhbY9nRyYeuAF5/l7gumBuwDr2dkro=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8816)
46wS2wZtSeNLgt6gvfbMn8pMdIMgoQMy3vXLUQ1rqCxYg7gxuR42qOhTbksYMxuh
sAfPNBnukHBsnVh1YGF6twcWX87n6/mLyQAp2K96Z0CZyQ8bh/0PXgggxqKi/wA0
pAhiaJXP7QzNIN7RXl7mYJwA40ftH72Qkjjh3+azuIb/CKLO4ZShN8D/Qog822p7
L0d2KZA5FpDcLivQIcAnA2eglKls64XrNku+E3Dh0PVZDcu02lQEHSkN5nrZ+PXH
pxD1D4R2KWkvHDADSbidxcYgZVuFzyKmhj43xYFr41P1Bo/figW2O7LhZKSHYInz
RVem48YcOwNyA09QX5aa1noXAAHAZvuBFiWjBT+UxSLMG5LORdZOC88anF7z+gk4
RVVt61HkHXmDyDw/B9tGNk+rSsyPCiw+RuXRfzxN/czkPmv5Zz+arVchmIkMiGf8
CqoA2bIdSMNtL16J1pD5LStQTeM13rJJKj9tErDPqSiJFbe84NemWTQAoOT+GOPJ
1EHbpg/OixfcxceW04BOn1KCU3P3nQITfQEBTC4JYn+wc2RjeUNICp5HXroWDBDD
Vlj0DmGjbxXcMpa/Dd3MZsiGWtnzOAfiDp1r75B7TCgM6WVNmcJO2BeUi/xTtr0y
bEkB/B70KZEjW9Teu/E/iGxJDSnQIl5pzAuk4YsMNQuf2gPANMRG84y7Mq0mYyBA
8LI7Nr16FrYUsmEdOpZt4erQt80Mtkkb1KEICPs/Ro3+g4KkH8WwTkMJmpIKsc2e
ph6YW0aGRdxIaYnRM2Ju1AuuwfC8ad71QsQT3GHpeXVmZ5DBTZ0g9dqtYhRXbUAq
MLoDngYoj8l8z2T4JI07uyHcNVMZa68814KgEx8Of77lEZdtaRwJY35eG3XrMnB5
66L+CAYmi5jFGM1Hae4hnzNX/HUdyoBxIFQZxDif+FiJB/DbTSInZFWpE9liStTG
aDqcDMg2oTKOeHXNdSiXlkIwYrjZbl8Wd0BaeJLgjjTwQYFK60W2eJz8FZCvC7Fq
JMRfxk75paF8e1LQN2ViWsDrsUaMQtyNjaOdOL1HW1Q7j2nTAYZlbKeARBG6fG4E
PSWzBcApBg4lHwC4SjGbIUY0+awiv9fKq8iUkro6rey8gOEvZWO4vP4YiglwVn2t
+YOs2kxKIfJmRkYiu2Ab/PRrr3cRt/utvQZDkarqjPhL7biHGBRorENlleNn/lbH
7Cvgy4+eoiEK+y1v+vxB/4PTcs10YJcpK2o0enbMg6WEDxNPUxv7KpJ8Pa2v4Vvi
mGYHDb3AeZnjlVwwW4vITzSAYuxvOXPO8xr6s75VV/mKV08/2H0bemqlFyeiYRkQ
Lg2icS8Qc6vI/sgSLVOHBFG19r3vDlGVD9SyONRXQtHs3sBrO0TOYP8X52MnFwqo
C224K3BLJkyiEc2E9p+dQgAK38gocbr/hqvZfpY7VWQRWDduCK0v4U1QjvCDOhCt
Ru3Fkzmp2dNo5tDPcMPMayJ+EGdKD4cWfyTyCDuS+01wPQuyK0seWodF2ih0o2Yk
6ptm4IhHRIZZc3ntdgGFAaP6B99ZuLPJwPTiOA7ubyU7o9PjeUbdFJrDu5RpDglE
GLYh82YeddWinpHRpLstKOMjo6v26Mw2S/kGE0Npsxqw8oxkONdRhWq60+YDR/UM
/nn6J4Bpugl6xTgHMWMScPyDGF+CSjYQeWxTq78IL7C5s7O46T4beR87xrcOjVDR
AoZsEwJ7WwKd5theQOjxMB0inqCHD+4kU1Y5fCNXQfOpJgJNzcLimbJuYFIyJuvB
rJfPw1Ak51HcngLbDqj/xoWYWw+62tOfJPhWEU53Mk2d45GK2hNAwrajmUjw3BBM
Ieb4cLRkJ29qI71gfxrMV+WI/bsvNwqrxFV7t7Co9UGzOdSpqQnNCzbzvhYCli1l
YFF0hGAlu4v+iEyRimjGt1Z/AYjlgPWDi8jWEtwcHbfVQTLNGZfSNuLICrOUGB+I
eoFTH12ky+aXApH/J+fup3fhNFpX+2O3Akmz4CTGhzLsW8zbXrAI4ckXAwckelu+
Nz9Bc+XEmTNU9fSWDtrG46vTHdwdrFoFeIAhmxQ1qGQXQQE2CfPneh5EY3eP+58O
PupotQOAaX2YMRWBcszNyJMp7gW1a2OmHvCcMfpFFAZrnH3ZlK6g749oSgWdlBFx
NhFSWHapXQELTYHreuMJNgeWiEUHAXpgv43KLLwFBOOE3LbpVPK5aTLEXKjMVwXs
OSUzV/Zhw2x1w1lhDKz6WY5tHI5CmBUMOJnP5/DrbTSs1osv6qtme23/+QxjCbre
SWwtClyFV8WNRXhTSbicIqhooaOpfNMmE9oElBJlsVV/4aioKQu9iyYiXx/NwMmx
r3AurL3fyuWTqUCE3vlCh0HJHdrMIqa2+Aokq2sNtixEP7MRLyleqZV04AbYWH2o
RJ6gQWWCcQVBLfucLQduv+Y/yNnDoi2CUys4X3jE9GfFVYqWxVA2bC6Tz3ZXEW9C
CHZm7NgGQcQ4b//6JjvEHkg7vtpblrBmG5SHgowuMex61CgvfamruE+66IZ5nR4F
l0npGHlxyBT/Orhjn8oEVJIP00vgQJeXoYdaN7oJ5sQZ45fnVWw6c2apZDoCrNt7
glzBu7jKQzgpm3wbnm/oCjxBVOg7ZPELSSXqRIAeosEWPEMWv4kcjmKnzfZ01LBE
XrfsryU/GNg25Dd0NLjQ+So3HKzThQvUlJe0IglgQfoq9oCtjkJ300+3KCGiHJhK
AkpDCdV9CjWdoU6isY2PnzVhc8mrtZAsUDGaYUYiOeNmDSA7LAWEzXKzITlzKFyF
+Jw7HNQMWm0Sq05NkOtYo9LPdjJJlw0/1qmoC2G6j5XfviW1P2vnAr0xms5c0rbU
U6yvzopthkLzjVmWXx3R5LqTpeJ7dqsa4Xq/fRWNMHPZK1M3pykV/OlzDISrPWDo
SLyW9yVmkwOVEMf7tieWvaynwSsP+p8a8u5wZBJ4h39pe5PVCDS2N/GyRynfcIyu
jblIZgQyvjscj1SaPylVX0kOl+/ey3d/GMiCykDUfe9Jfqoztp1bwmYlNAoD9AAC
+mLtR77o0Nqs21n03c5wiK6p3rHdW4rLCxjoXLF7niIw5A/AGm4coGCPtl5iDr1l
+Q68VAIhyKygkTkmT5w22YB2nYCJ8PCOyyrGviX3JUNRPkyMxNW/otIB+Rdsj73i
d1KTDa+II3u8AYcQZsp17IWSRH9sE+jumiKhjZ6Zy14rIil7kTRHNAPn8LVYVjY+
CT94VebQ656rvfxK8pBUhOFHvnQsyURliCISECQFyz2UoJFxJzRZKlTc7Vp+XQBr
qmczqYkBBfjDqh7+hIqsHp4X/vcmnuV/eXnxuCz8A2GMeQo4ZggnbE20SvckIOXU
DVOeQbvYV6yBJHRmbfpZOQ2UI3+N/kO/62cntteXXPhvjRlR8mZ95pJxZTsO5mF2
2Yelp72UG+WQtV1AMdP1OXOK1vRo+GjJeU5Qa80BpeoeXV9XMh9vLpHX59s6oLpt
vol6aSF1dAysRSqrvh70zr0jw+O00FPplXO1u9viEpqjkRIxg9DSBOaxIWm/yBq4
Gbk2BXQoe+dkKdSpazarEN+K0qQU2rv40Z6LE6k+2ntMqO7WPmUR0kDv0b6jXJpZ
dBKsqPhnDG0P6uvv/LoDmThb0VoanpFFJN5Bm/pj9BB9dQHgfb0nEhRnRIFX9kRP
i2Fkj4GWfI75VS7YAas7Qe+Jf4Y9cfbJYhJyJScPQLuqDzf4wTTybT9xx3C3TJ/K
FzHCdXSF0rWFZ3WX1iAVorFBaIsKY6D5LSyr2aqfvc1L7H3tj6Pgp3ZrstfYuN1k
gp4UuP59his94EKi4D5IeK7an35KHl6WGgQ2ZOqjTeGo2+C80UJr02sf4clipnLn
ogzhGgw0iG98CZCZiaqBMdg9cE5GMoSPjbJ3/yX6R1Fx60JQzVQ1/BJBkMJhMezP
OKcizbk9cTrbVOMJz1kvJSqBXQqIQVtNtbUUv0zrenS9gHu/oCU+a/VxzXyKfpNn
2r6ur7214alrhcHUT+4Han3cpPpe06EBczEzEuDZt8sIgfT8ZdrBJWeax6OdNeas
H08fbGHGelulKA/eyiq8l36N7vLuIPQob3ZNe252jNX/R6szlzfnNvawP5FA70I+
46/pz2X8L6vQdA+OL/LtSjqkTKtBKXryLvMYkbuoeADTNIaHvoaPReS9OByNzGey
cb7sInV5JfKouyDSXTzwwq1LY40giTl7zmjU5QNEfnCqazzl3wEcKcBbLOzpdq9g
329mkMf3VckBOcMteDoqf3FV7dk8zQopRUpeDDRBfAyurdWxHqxXbE03D1yhL8og
5t8/hkPxnE9efeon+d/aR6tAAUt6HjWhUeChJQcCimVa0z71N94pfftz62ThCoPO
Cab+8nxmnXSu+7tTERf5Ji6mvgEf9VjVNCPKaqlWzMyONc64fX2e+xtJIOS1p0hF
E9F8BGfnNGUJ8fR4HcV74n2SXLsaNR0kE+s4G9oHczkpdCEFncxFb/7IiPlvJmh1
eM6OmP/0Sxid7DHpQBzwtGLAu3tteA13dqb4pzjbvEPT0UtbxigeOSsMRe84i9cb
QbRuZBE3yMf3qhKJ3mbjoiu2aiFtkTeQMCsCRzwnXEo9SllKr7u53PscIzAOIQld
ktif1tzdUR38r0Wcop3hBPk00KNwrmtl2bknYnV66zqa8+BhRqVZU1b7LRKGLmAL
maeOw4Wf8yheBMP2uSkMkDr4va6tX+C95hTZyk7L3kySjL9cQV2RzCe9TVLX6wyB
PvaJM8o4EQE0Hs8huLLaN5Axa1pu135XmfRTWhUDJThfHH3OY7wjD0C1JA6Z+HT+
4wWcGurSanqUpYIJwkXrCd/bY8pe3NVCvgXn2F2jsPfuDY5Otqd2kFDo+1+cB2FE
yvMvi0k88CSxU0QPUUOMhDYRTEpKnYdwWKtC8UMrbsPS8K9+gNnIy83HJxatY445
iXqkYvQuKupYkpW/c4IKqgSaTJ+kesDrynWNFhiPHYw9QkjSSG0JCqgoC4eRzBxc
UOVrYpaw17B83fXdftIfN0d2dzjBFupTPXXTp+oZkrdTSwV1rk0ITS/wMopxDArY
+ie1dxtqUVpaseaUwuDvxEBoKnDRHmdb+X4wPmMUL1masTDaNEQ+YaznBjTnvLEy
OjSDizHW6LxQi8YSpKoz110akjInw6KhR+ocOfOYrr7P1SuO3AO+H1QI4VSif2JQ
+N/nEF2QdFDv+VVo8SzLFROLcK9QeSj/JXojn4D3bl/3O8FZy4y31XLgoKu0xu5F
y8tkjpcqJtN9WIha/++quNnyLSYV5DQQ6R0IBmB4j4z03x14XNz/9wBfk7+PMmbT
WaTuhkoE4BxIPJIGUkXO1KkQD40OwObknUTVdHBx32W7Rf34Ubi/XdbcmCxow3wB
mFl9NsI240/sspfdA9gBRPmA9YZCgPHaPBAChW7LmUY7SXZZE5kb9eqJBLQ+PyP5
04J7c37ErDKayyTLpsN4oz4v982rnrHatC3RcfrU8T0/i6siYmLpKy+ZMUXh1GVE
ZugUTQ1UWPS3fiKYaxIuixDJweXdD6E6xRh4J+UBGrTXHC9fm7+LGUACBG4CqV1n
oixYtCSk7idPUWINiZpRArXUPOaEqB9LsXzxjIDAMilsK2MPQdvOY4eh1wFCB5JL
/66Va8l+sMJQkpBusEEdurOwAohwnJYHdLf/23bv5JRBJchti2xPGDOuhaw4t4Yg
LgaT9GIYXTlMcDkSOLt+NXsmO4+tXUBte/L4nHOhMp9QnPzV8fglsFFYY4WJkJ03
yfRv99g3IGkaGKBa5JbqZG8F7sHgpiqI8RQjD8hdpB0ychTxd9Mn6QuSCUpMYbV1
odqmHFzmgxWdXVqFtA7PwDu0QgspKp69KNTGDVkaU0G5Y3y/kYEfq7oR5HymB+jC
0480dPufxfhSL6xcCkmMbjjHoAw3hkLvV0NZIzBbTuKfG5MFuGqWDqmozTFhXfpA
tnDjmBB8yB5mzxnjeQx/ey7P8Mfw2O+jTqtCmlczi/62c16c26mUJw6kHqVReSQM
96lfvEV4MscVZ3jHSGi2cFESqOz8x827dqCr/sCUTuLdeFQ3ZXmoWBKimkhVu1LX
VrHkcMQb4ohX8SsVQPmq01Vs8H6nDDdC76rFup7eMYztYkWDlHjYykD9KTq2sMs3
zFilBFfRNcRij9skNHdaDywZ+AsTmTFyg2nOvYb1cpXVPOkkJK3x19GmlzCKJM9s
Mf4ksLb3+vKeAd8Tbnch9YykVWOH6AiFpRX+Icy4K8IsSZ2602U0IBtFUg7HbI16
JsohDdNOdGwTT/KZ20fJBzvLTwKnlASMGWdz4NKTsK5SHr74dpn2Z5u6CQsRuqzY
JKbhPNSdw6rR71ce7QYWkR9tXo9a3NVCsm/ldgGZeTNvSX6SVSPlJyf2QeRJY2u2
azFDSnN97ZKefu5HqplaDp6zZ5rP/lIAuYOupbP3T1y5TUKxydaYOGcKFn2Bjy7F
s23ps3dEa07j5BRbuvjfo2FtVRRLL2IbPorqC9RpQ98Ns9fSI8vH3vLx/3r6/5dF
p+zsxLwCE7kD1LSabysIOvq+NNvVDtz+YmZehTyx3JZzyKYHnNn1H8ZV8Ekq3wsp
bj/Yoz1mVwb7TdotENshTthkeyERzX4navsnrdatFaNWueedHg2tItuMAHiCfUou
B/DayM18FyFCrooDTa4xYybELJ6xUWHAdhzzQu0RmKfaxTPaK6aqzpGXvicJp775
O+GnuschfgtndXZJY8wgfstkMLCHSGpNnZVQiLvDfrXtj0RVa/V9sro1vGu94Yci
1MIzBea91bmra5esqYhfLWsDJVlyp8vV4q6V0yiiNqX0rx7oVb230D8CJDW1Y85L
Qrfo77oqahkksrH2fUwLsyeRwgu/b8OGm1t2DpaTVd20Vm+GKgQJuXZNVna2s0h9
wD//79DaMCBmzOP+7KwjBLEep/KNN+70AX8vnlQoegiNS/KpdabPbNB0ECS6oWFS
dYKCK1mtiCEnsXFJnxxcPfxYuNYllYc9w0Hg4WnhxHg28/AZOLAIiwAt8MTfnGm5
aMxIj/R5j50klx/nuc/pXFDIBaDMUsn8ETB6TpUsxnqvb6QNRwfxX6JF417y9/M5
TBSU8tk5UC1Zd0EvB2bUqQCtMOUz8AbAdb3OxduBLwFQ163T3QK6WCS8D5Rq50bd
dytU1jurK9JBSZf+SiPNLQCJUOhKsqtt+wWM/6GMvbYFCsUwl4GYo+F8EvfEZT3e
aZXxD/m+oRpORVmwHqK2MaEA+Y3AGgsy+ge0MgMEULsNbtSAAkBgPg1wNRioURkN
WVgtxKJ3u6tLhHVKspUyALeMD5p00ePDX8J+PnyZsluu0pwe2loIZQl20uYqur4m
f4Mj2jMuR1fttAO1zi35HToevRHPxJ4kB6xthvSb/TZByrX8TirKtrjJzd9SHBd5
2m5IoKJpQRzO9vyZbbRTHrzl4KPP4t6k6PQCcB9+rWOcTbEzWasPakgziaRXcNrq
2rbWv3gMixlU01CIIvZcRdkdhHQIy+uCGmt9lpT+mbYFfb+Km6MDzTTKfLsOmC+j
OgiJEdcjFNm+pdTrAp246tSetWffAgCx5kTufz+3BcPs8O3oiW0sbCzDGQN61eTP
ejl233IjHs74J011X4oj/XcJaAKYDSHEVxUYroyAWLVFAf4wHseGVE7Z4xMwOKOK
8aUcXMZw8ME0Ii2tUtPQGALg8XP+miu76ByFUBTPQY3dPCRpdn/e/dKgYDskl7Kf
T33RjeMigLfwDTBT59YOx7CtLV+ee/QJB8xqVUGooj5gmVOPAs8USZa/xqkgAOxa
YXh7Z9fzdMGXQNy0xsKtF7zHgx/RLFRtr1ddFvfiKs5CEoUP5ufAH8zrgJ6GXCbX
UasvKCvn4F3JGrYjYwgMULeJ0ROb87obLNR9+VLudjH/dFEZJZAj9SYAeUUEueZc
o8HkJ1oZStJArBuZxPZCfzt2Laq8xv17jjEzv0odmeCqJ2rET5aJw2Nrx/ne5AYo
+InDIUc0HH47kbmmAGggHQj1oWbDxcxKLyEMGT6HQLF0iweadURwX0GqtNd8l0Eo
6EMBsBZEybsknA21GUFhT17PK/+2Mtlkg6mkgdJUlJb8Pu0Pjs8ycf3kl/3EpYh6
xliDGG/CGnpGXP/nwID9k8l6NjqRoaLeYpjeykweIyWbcAMsaxL8Fku7ALk/dmjW
yXCnyy3qZKbt31CMg+bONDrVrIO3Q4jUdDBXvbhiCPL7LUfJAi+Ne8w+qZK3RALr
lnQS3ZBNxIYh+/e39qQoA700SGxRrEoiC+Azk/BdwDYViW7cw6hyRhF7PZZUAJvu
P3cszy4spWN3A9VJx/9KIpn5bFMXL5ZDujYt+Ik37XwAQrUNFWKdrvSyz1lOGTi2
5hRtnUCZJZM+Wokj6d5NabHJZlYz86eCHuVsyErIwZiNZiHpr6OHsfyi/TVW1BRy
cuON99ml/DBo2y6FYllRcB2OuGTsB7VQCUv7ln1jS6sgKOa/DK7RF4wU2QOsiQV0
g+4jdtNgXIEYPKOSPnyOPfnsv35QcxRBL6RHrW37M9xAYv4eRh6+LIH+6pxtsKuM
GBEYSpj+Qg59UVxpkts8oGbd4dQPDGSWpwq/KZ0MM90iNjU5Fv/d+2o/tFSSWtC/
S3A2615tfMSK2PFUOcct0sxkZwATOEqztPZLxlj+wnCePzKB/9bp++oL2FH0uwUl
LI7ebY8urDu5rRotgK1crSMSDWBnLXg2m+Z3DLIUsD9ge/TtFBZWy6bC4uWpx8a+
BO/XDwCEBL+s1jbRIcmrjeprkxQrY9YYIARZ8uhHDkS5OqhpThPbQCUQfUUvpHxb
LnOtzG+3WvIFKE2N5TUdxUopnEio8HSvoBMLPjhdc0wdm0e3LC2Cy/uZYU/T8Dce
greAmWF+u36srsE0qvVvn7PcUsWgqe//0apMe0fsWGqY8d/MS+REt4Sc3WkKL2Un
mngvnI6gi8b+aFmixk0uO3kwYilPmyjopSa3OwGz9co/ygZfVV1EaJ/8baLn+0f5
5HkiSKH++nTJW4S9XBZPnQycsN1f8PDIWjn5AxboDH1FPU/Zmoa2BajcpUtz2F15
tW35Jp2fHg+jf93UvdyqiKnaTbK+wzOvRcrSreCCa9afniUBFIxQr42It8zqcgeb
DVMkJw8DD7j3gNNlubD7Kz+kyvSm37rMVK0rO8jcEjmR9wbhx05+sGS2m+nxwTai
hddne42rYUgZ/dYXuL3eiiu1ls99U7Uf6hvH7xxXJwI/WHlXS3bg6jr1bMa5gx87
oPeMeRgjxi1NrvgriN7puTZ+EKnDVT/6sLjuVB3tjXWM1Skg44M36NvKKg+x6WYt
HmrWQ8vgfmtXuTwSNTYqX5VXtxkl76Fg66TWFD8+1lzPk+IQyAHiGqGhmGTfvXR2
b3jVdv1LCsRtCX0FIDEwXJRpRLB5iSfQAKGRXq0ISwL3YtYU6AHixR8UCt04savk
L9Qi94vHEbONg0gxgZjsxhE/17IVJsHV9cNuOk1Ul+gSPBNeEP+qwONDWn5hoU/A
WBmripyJCTmxmVe/MprLtPOQp1LLvZpgKQRO81UMjCHLs5JQVShFcDexTIRg1n0A
6WSgFhVgWxy5nBy4VCFUm3MUgeMnz4v5rmXip0IduVMcyKth1T4tjvULUNg9qBKO
ZOAsDyGI0jtVlcBiIpr/LLCCUjGoe1wtE50AnX8SqY89Eb9RMX6NNcPFzPdLVRPN
gr+ZEiMHdh68lHmH3dX1trBw0iKWZ/g8VI5kQEJlDb8FumCxaao9GsNIZITt9kaI
51fbjCKpWZYIIpIhPUNeS3ua20FUePWMEoOHfCazWOwhqSvKoGLefaSKvyhzKlVs
PD1VluOsqEIxjQ6Za448oYJHyMEFmaJg2yyj9+rPy97smQ+6Ef4eY8kkxGDpbUqb
ACsM71QObTe+INzlxEzky7UZtaQs6Wqq69HSWLmGX6ZJT/NBsFznryg0bvR+BYep
sK0Xc0Q18ou8SoGBrAsYaIXavWGGG89PKLX4IuU3CFwBToiH6pnSk15EgmrWyGa1
gaQ+JUD4V3VZpw2UDNhZ+EKuOnAGZgmhiBuwbe+ep+fCM6on5wNfj+xtG789U/KN
LMP2utV5/FzoLstYOwGgYJQmynLyA0wqT+C4g8loF/bCEr9vNGXikVRNhNKHfZoa
q1oRzqftWZQ9WUk9fntEh3iF/lrZUmc4biYHf7JnIh6bgxxY40K2XH1yrhT7lXwY
9kuPB0PETFTkpkGH+0MLzkPhF/EY+crD+mCk6z0xiiff0E61l2X8/2ATBaL52S13
soXTpOcL0oxha84KGJuJeIBqUlOd00IrJhB2dAYN9kyV91f5Kc6B72zablYkKYgy
LN9q5eTSzS1RX273QhvsJJ8p+5g8vRhwkDv9ceO2WLp+1ea0uAFXbAOuvy0LAt54
retJfCieKcQrvEBCXBiVyeel7ShMlDIn7/0Z5Aat8qh7RAuqlDVAzKKgSdAX5q1H
rTlZC6/KmgMRjtjIMPjkf44Xv3LDSxVe6m11MzNOrv9m2uLGehCbpK7qE5XZMwZX
NIrycP5QPP3zCetCHlRreKEtqZmjDw3ypvPD/nHvguydPdZEd0kb3vIptZ10Z/dI
vTeNRyMnunUw1uKe7XcuxgGuQ4OyZ+2eRixaNtJVBpeO3wQrMUEgDXnO5u+rUNId
5gCzFrjfHjKOMlF6K4GFseY+VLsRVKUtrvNXyUnlKpmGzK9yBd0nfa7xDQaQaxFA
9TuTvh031DMZWFTH0MFTTRJDJaSR5GDgVNay5JnRwkB8LkMQTg9NsuNyXrqrg3V3
hQOjFPy7/qBt7GivIjrLFUa28LESlTYKCIbVozx9JeYvydD9XB2Lp5W4jiqmlqDs
8znPakkMBc+djHaQAnRDT8A8F8LOy3mW4ntjI0yKk5KL4J4FNG0AxfPM4w5+cwkI
lnZ6YRKWUC1R+4cKyKd6Ji60SknXzKaG7KXExqdJGsRP1ArrBPCen5GTdm7r+0lY
zSYs3JVzvOa6KEF4xkqusAlLMMH+U/KfYSHtvgfGhuWKvSfK1NjVMjJ2YTp5f3u6
/s1Idhx+pgynShTc9FeUv0rD3UGIL7oqmDJ95EYHQoDpuugVUlsRNUKR1aAfM4Jq
n9buqRvvyhJnxz9AGd9zid2mlm4sdTzsGnraappT0Ajv4bbNLUFkNmjNAP2dR5x2
yjz6BwSqDIS9xqFw562vzH+IbscGH0plAM/2rjSPPiARJ+yx+mwDcsEaIFdIz58f
dFx2C00CdrlQvnmHn608IYrX2uBxrTntovTlNGwWnXD7TT0fB1sSGFiH3seqcXNO
rf7DBaJa8ZiqhqXX2WyAGrdR6VLGF5nSqCv1NWwXRe6bi/2rANojqywrFRLQZxf5
jXy727X6WgxoO/PODEsBj3C0hU7eqscyLX+4y63mFZd/uzy8iDiJ/ug7t6d4qXVr
dWF5glAbE8Jm+t/m1qaG0fcgJz4tPCgu7logMuTNnEJxIE6QtrtuD7MwYC1v1adj
fSU+DrO9ralKcG4kjvFKiTo46HUbBY9cCsID8nN4mJYQP9vyrnw203gKuq5XGuMn
QNWCzi1kjyN2ybSWWlCbuSDf5FUFsYE9Xxttzymrd0vkJ4RFRcGqxa3kJkt4mqdE
/UaID11CPkpKjLSiLEkE0og6JW1Oy5+GNkQxgAnaXLc=
`pragma protect end_protected

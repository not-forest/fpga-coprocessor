// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
1zHro41wgD7fdjhMSdsF73OTvl2SNPP4fV1XmNnpQO1w6d6D5FlmzwT6f9FBDfaQ
NsFqSg6kV5PJzyAYSw0CfgVqdwQhV92h9NILrMGy6F7Zzz78Vsj6zGJacT/2KMit
/rLTMDGbUMebaMYtpyqVimjn7PZ7ZGQ45R9bIpLQTPA=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 15168 )
`pragma protect data_block
2LmB0DffhLityhf94a9RLw76qn/HUF7EpdVedBsM1jhEEUv/yT4tnhR8x3qJUMdv
ybJjzL1QXUqBwxi0Cb62/2I1Fez7YrL0B+LB2ognLRWHaUGL8deJ9/go2ZzpdwlO
sh7e83FC34TDcqZ1ppu9JFtNjY8ue5VF+DBWkzbBrNS5HNxKk6ZpXPU9csgN/cd8
owP6zhogBEs5JWidsvasRW8LiAsfAnFDzL8l8qa6nbgpQkN9qyRu2jAIFMu3XQhp
pNJMjIjZuzuyntOexVAkqVlEhnxPPmlSDneGABEi/mBBf1dAsaGkgnk+X1NU0UEn
mskE4jw5/DqcNQOv53Fy6dWy5rQ0h9L8W+1fw9gPrGiH43xIbMgiET/fEmXw6PIN
GAVBrsuVO5wW1zaQz3nXtk8K1dzC25KBlPg0U7E9m5zzNRJBhWokLGqb0jym5Bzj
BVtYuSGnd4oiliZCLOte5SN0TS8a13GruKoyS+KtuWJ7vGNaYS2inkCNhMTCHwcS
JHhnWhgVvLrh7nwmUE6WD9wJPdTo6dr/SA+C9WnZWLJuVyyhb4N2CEkBzPI0BzkU
ctMZFfsy3z8aKX6Es5CBTf0vdLkJPfRYw4LM496wKVN/b9qaaLuLvrMnQfTygsyb
aGmAzt8r+bFHvTPRrrLVV76EViZ1sRDPpcujs8idabDS8xu4Dwj0nAzvVcoqKPZj
Yj8p+CSpigiXvoR0HM2flTBww+jsJQttFjBMUbM+qhzkNt/ZIoIbMZZfCZ0cKK+2
7spoKxD8V0rh+6eOWVLKu/Wzv2VdiHxUdh3uF7PBHVBwXebrp7ZJkgLz35JJSVWQ
cMrIQH3kUcDvtpfYevf3/+uZnRfzarfVBLVXKaPlf1GaoF3s1hQt6YkfziiPWJ7H
Bfyg9TFnof2zbdw1DhUd6mOWnRq2Ivj49/+1OeodQjQHVnL6iuXjFUvgoegwrvUT
4bU49ZT9VX1hGY+bGme4PxqbbBicQk5shLx3m3eAJuYKks+pvXjEvhB0l81ljb6d
UUVsDwLrYaJe74hof2C7NzaFUhgiBQB3i1soMY2aeEOGgT/wBb5Szv2AkBxKiqmg
DAjNXDZsmsD1wA6SX5KvAtUTL9OnLbidOd012pj8KVlBJq0+Qx42IjeFWd1/F5Fb
0Mwvb6rpNNYCqUoK1eLCKnQtt1NmrTaMxHlSBXhZyrHv4x8DYYT5qynNnQncXKIp
qEH05tMhY3/LXBSiTnspuC55KC/nf1VUk+Y2aJ+Td6lHwXRtsxffpV0y7dKlselU
sNs6V+dlL5bF/WCvOg+x4PYfmsvwHBomilT99dTteAFGV8iJRP1UThlvQF/Wj7Ap
mffDDFmPL90EeKKVwHeondbpBPo4XNatG5jtfUv7VOSt9zzGKJkCkSFfkkuhmXkO
5HEKivhn0ulBxpNWknkyvUBpHiuJeAjmleULIcgXIpLQjhXWPYkWW0G7jszKg0YX
In1QKsnhOprIUNZxRNWhCpngS9KOWy8u01Xig95Yn45eC4xE3h5JwzfOmOV+RQ8S
UT8TJUZlftQqsR+jI3bPz0h24Kk66PGTJ48nLId7zpV+iCYzKba57OTLPyIFOOeJ
bfOsQxiarSvYZRs5p9VHQVjYMYgiHRuyv3KeHHERaKblsh8C9wT3KUzQjpQW2l0e
YnfmuMbCr1/jKNHqfbGcp0vfNAYMQpXH4SZnoWdX+1ONAueijfwFivjR6nK/34LA
r5g8+hX+W1RjMB9wjB7DxdbcdFZt4Yo6GEt0w7872DA3OmwmQsxhFqNzyC4HY+dS
pcz+8549a8rmzpbyD1rcosCFHsJIzIANVS6DVK1mvSobdirfKdFTGHpJ81lN4i9L
fqRrVHRyFuOd1jqh8Uj5qjT8UPzGpTtWUXVLAj4q7ttIYh0o7s43xLO5JRCHeWwr
hZiO1BR95lAybC1T5DJ0skZobHUP7suQEFGI5MVtR3+54pXw96IBczwjCA16Rdrc
oUgo6effQvnuMBlVeKIWX1wKrV6xBBgg2ReQyI3f9A1ETjd8x0nA2k0EEtOa2S9Y
LvMLoP+/9DBOI2Ph8jMPwc2ZIuLIL2VTgf3/F3fVYADj6Nq4fj/u1+m83FqbXF23
s444AppINRBzYTlk5M8bERDyCxcOa7lhf6JxOHyjqjisAteFNOkLCA/85DNI7T1U
F++svVAXfdf1zJsc3F/gDflfRpkUOHoeCrDtnPgMdcR+LdToRTfUAUTNyYFEqxyZ
mKY9QpRo1mD+tOHmNK2NxXf4Bknvou3Ogh+zRC1AgtBRjotAz/CktuW1Af031/b+
GXkDOzHZMSskz+A5p82khcaRODxGwbctnbApAKil2vFfShsIyKRKOBoEE45uudKq
bzCbkVmSnk6w+1Yss3LpaQnnZwuIGMjajwErUaK8zjGZNGGZ9PwzpNmIn94pMbf2
o9xgJUHw7qbg+DFc+/TIu7zZIU9Ba6kcSqjYd7/YOw+APSvklq9xkz+x2WJfkEZ/
T+5bmTjzUwUp6w8gf/IhloTEVnJ0Z9p3HXsoyhZG/GWSwM6Br0EY/aKYyZXrJyNE
rCQWIAtcaOLhld5e3A7kE/z2Jsw4CtI/C1A+SL7AYM73JW/WxWqTQv9jAyeqhQMk
vdOhC3u7/xIbqZT4VL66VXJJGhzSsKZLfFcR75nKz91wpJJ0Zfbc1n/BLstdhuls
ShY6FwU0IEk3Xr/w1XF86cQEbfij5MsFQayEavKEcJqF90kU0ppFo5BMMkYKt+ik
zZX5kqmJi92t1E1dVHwM91o0rJMuDrRmgcqQw7Pd9zDBLQS6VWEjQv5yNiaQViGR
Gi5bewMrOnbwFaOr4zvqsbiZ3QnOZpGpHTQVCAU+bI9MigF8ih4634mAoYTu2xLd
LEVrGYp6YdKD0MJGgLXm3KDMlvXMy0z3QXQeg3bmhvlq495F8OkgIgXmsjOYZl67
CmBH+OILAPCCwVhL4Wka6i1tr1ArnA+hUYWFKY1z4VuKZrPGgOc8wCvOm4uEAtwA
baSlREZ2MGs5WS4VgBm1Ful7m6efGsjjxLVn0dMQ4fJS+pBHR/SW4tGHGEpTX32M
F18S4EF1ixX4I4tc87s3U2jnH7m0ewNiIWJYe8FkFmUyWu/x/IAjQuMlkV8Vsv4K
hMsAm0+rXenwM/QowOxOFVeB1Z9LawHgav6JcelMt9vM+OqBC6RG44taL6t3a+lH
tk7NCXWPG2kinDJJB2kvCtqoKjFzPpKknj9CcykZZ8QopDAoyyhnQXkiTaFH2rRx
uGqJqI2V73b2KCbRce7tkvvveUMp3XguF0EAaXOyU/72CNvWZg3mkAtwoT6chcuZ
LIyf1R/tia7TDC0th6ho0V1IOX0rZANRjsKRkR4/xwib+EOSOMPx3ClKWat3Ucqs
ruxnJpYWdly5P4LMZ37YK2KcYojQRuqNCmC75gbArzK5jNbHq1heAOe3GAItBKDe
wA0Xr/FEX0fPXSj7DDYYniZB8zojB1bBl2NcJsTrRIYr2VVAgVbrDApDM+XUfNPd
lZBiZO1vxCc9jHfzUeh4nTi9ASnhDVvmZyS0QIJpT504ZLba5MeqfdRu+psuYyPo
kqj/Wn8AqX6/UfIIkZ6Iiv7f5P8Oiv1QFqRQ+/Z18niu+zCxNHhgsNvzrP7rqrvz
UDx91WEHTFYdGFKOuor0E4wauy44dRaKvAuaWfwejCkPHqGTJJALdHg5EjFcVALI
hg+Lqc8K70qz98SojcvJxWk+wALKF2/Tr9K4DsAZc3pC/ji9iiesritUtDEFQfuB
GpIuYawbiqAhE+6foL30iX0sMEUh1iGP7UQPMrZitVaiGxcFNLnziBpLeAFK9F3V
PV8HPsmcGWWxu6+y7kP1ceASExJ495IqIXCxEvqDN1DDj42pgv5yExa3+LlibURS
DkBj0SlqiDxlIioWcwYr9woSBwKTw+K+lNdmazLG2cGYlcvwixBkeOCoBjT8Rx0z
+A5/UsF38b4DV3J9jbKUg5DbpiOK6YAZWr6AMy04fCP5ttiu/1QVkXmCT0j8WZsy
AVW74HOzeChPwcCPxTRr/0DYayb4TFYxSd//XnvdPMV7c6CVCI+WAYsWoABcTRS0
HdfQjjP3r3O+kSMKG6LuzCIp1u8Jgk9GVCuF6Yi43u2IVDXYiTeMeGrMoGxFmqTF
T5rLe+2jzVMMMySe6nNecHkk6We3TReiGiMTs2nBMTU6Mx19WcUTlsu5AYZTlrbR
72uIGt0ze39aIeawyWf+7L/xR9dWCW0yc9n3pEquvekGedZLAkC81+WmQ8SDKrU7
I/NHIq0PR9LLFKw/PRCRbVivIlxnF6M/qk9h3sRQeylcmHl4qzH50BZEynnBNoVo
01EMNqQAFjfwrjSJct7i2IpX5yp/qjV11Hzs3XHuqchRTcpm4C5OyW36NSO0qoWl
UTDXw9NWdz5dDjYDhN31xxONlUAqbxvgtTbh4gi1rIjORdxD/UvlqRylu8u00G9E
AhXIvzLx/daH4LX286CCpgr90f4GxdBwCjbFK7dRSuw4UddaOJt+WzQvNMU6Fvmv
O2tVHwEjpv5wsfgVcqCkngO+W9HNcy72xlA8GfNyL1N5x+7zdXgYJgrklC7sDvx5
9i6B1/8THRbs0Pco4FvdeSv144DrBzklneE0Lsokiwpo/qvsuLSM2kV5g7hyi5kF
lu2lPfkqLqfvHpTjIWNkuF7GJxBU7/gSqxpLm5OoHG+TUaNjglXpJDPSrfaPkh98
aNRb5+bjWmv9o977ibPBaH/VGSOaJNADwpdDV1i1Bg4ml6fvOl9oQz86wua3dMJ7
ER6dAL3B54+jKHWH6Au9pu1+eJwicv3n9glXnuJvzepdATy0Wk+efqe6IeIdPaeE
82isbU7ATzIcP1myMER0kRG8OvwfhwNbiazxhYoEZK1aKIbcuHeuw45k+rmDbQ1T
QCdb2tUKzwH/MGQ5nih/WO8eGyz3duXBslzjJlnI/c7fJUAJD2qebH0umbZcwysi
TSw9e7t/T3xTbjWJut04wVvpK0S5QTpKEgQgPe5yq9ZqsBTT95g9uVmfsHFuAVZG
ky4uPUeNhAnMdj1hj1n3kD+V0Hzb3v06ghlUVHkoTaRTXaWuAYexIDQhUJEmCIZM
zdirBIV90HTrJfjF2KAG9HuOcAaVSDM8sR+K2kVObCnnqN0WFkN76lD5grvIj0zR
8J5LbduFXdqE+rVwgTC4S0mziarcqAl4xpyjjb8KuIMb/Vf5eglNF8heJpQ4JzKy
ooKS8EOGvLb4vw4YXGrupz2ebHsEPcWi6cwRV6vqitw/8t+RA3Z5YWjGLX6UQ8lA
wBQRBArXUqbAWnljlnLNfEwphe8zbjbdIsAXkhiofqbo5lO2DxoNxXgPOzOOHcHc
6dyveY+KvK1YEHcHkj+jcTP2amJMEudBNf/ze0qIfl5haY4A0pK4htnp78vICfCl
kR+X4KxFu7PH4RWRdg6nj7KiOMU+4YWUzG2dgc7/FIBAxyqtq7pE7NhdB4ZSHa7t
0kkZ/HO6IEnNcixq2yp/T42ZtHzgXxACBiEBs4yGOJxSgGYYVWdVIM/qB+bbl1PG
2Uwxl0soKjhwMSdMlvs8DdizP74jQZ6bj99m8raHwl8S8IWY3g2NGdr+7Y6+X3cB
/ueatQz4wHtn03DaVh898SLgk4RNJ5baSQ2W5DtY7YJMn9MFzUAfJwnOPQP27y9/
Pq0HBHl2fN/IF60JEdPrbV6SYfbXUakVWXwhUazyQTRK2CWB9j3+anx7cEN3lUIt
1Nqxjj8Jo6rfLJixSvva2iwcko7HdsLXFJNAoKthgVktWu5nH0bTnqsrFoSE9QLW
7Ur2j5f1OG/nmk4dNS2B8eZDNQdevuP0RmeMwx0Ho6OCbfslcDYFFsErMS7Agq6M
eFJvTMGoayedYaZsesKv3h59Pk6XcnJYF1R668gpzMKBOvcuLGjgS0oq5wOI7pbb
vmsamKDbHnV3LE9GL71AuBzY+YmGfwPxExzEdf3WHhxLdrg7w9QG5tkJzT5SITd9
0paiivTKP+Y17y12cd0C6MSBPf5pVzsRTWu/ZouHQrvCNPU+raBvUWWWwNBwYDMJ
3Zn3div1ihaV9jLnJluQSqPGcfduDcLkEJAZhSzSv99+Nwdcwjrods9MZ+fpzHz4
gTi1qgIZ4gWe4qTCZ+6rzr8oBB+YH6bushGfcvDwb+heyQxWkTRh5wiLHM4cKc0r
9Zn0/TsHi5xe+SkNC1Iju9VMxXKjXKqXli1LSDLrBBKxxbVoRDvBVQqUfFU/tPbQ
tmhjQHOq9ZfcdFCm30R1YzKjntDPXYGkA6pZOFtDyGWlqUUUNGTt6sHDp3vyVkr4
SYwElBaxJjjOjeT6CQk+iCVCF8JHfiZqw/WzPEOV5YKv5OQtxVWmc3rDYNZvbIrN
pNRvhu6RwjBRjEnTAh5J/4JdCZIU2yrNLa1yzYlq49I/EdOC0kG9rrpONlJ9MP7D
+fAzJMSVPLfr04ZCeJndgEGpzpmg99pzHpKcsbkV1B+JkouxDRlbW7+W5Of5moSG
tr1KSurcHp6tb6EI4bbUG2I073DitaqY8LNS477lhadHg5C1w7ocqSU7H+pKoGYa
5lj46NSblRC9KrSZAd2/mlKdVU0ExSwE+b+jtnkVJQVIaeWfSWCSB/O30TwT3NTy
aZZll5eFTXs8pDhvRa1VekXyrwZ2uCa5OLpVOmLbOQucMWB+VhTkmhw/SUEY4yZp
p3YAur/8VuvvbTjRySG1KY0gIMYs+sLb5LePTe8D21YZiGidmEYkF9DkBYEfq+RO
O5VqPvI6DTfEGpUS1OSqq+LWIhBgM9VqNHGMIhMpvOxQKwPhfPGS5gECn4gH3NUM
Wyv8tJMc281SpySM1EjWAcRuVCDkhtKu33Vb7dLAoWfpDY4qrdyNZTh6qRHnVm4K
F6gpXag1vWoe38ASzrajiZvW1RJyZTbdC91oKI3Spxm0lk4PyaMey5SPIumPjAMb
ycEtIkfRgt187ZDnc0kWkCV38FsP0xi/FEzK6QqBWU5775X5+N8ZQ6AsLfToKQ0m
hrCwiiUTHyYVdGfXtCioPyqMFRJJuu3p8yWrLboCu04wmV7Qguw741eXoDjJZM6+
a375+dhXoROybNsrQaAB7FfU/aoAGi+u9HpkLNBT41Kx8zd97qal+VqE244nUm7O
egsmEeQguzeBtBPDp73WQzkFL1hezV6D9Er5+ZjAh2pW+3aWHczMzlL8vRmA9I3o
I1DC0/kGAw66yV5UqNqcEzI1K0KcdYGcW5yLCunB4uO5bK3Acynh+ax1/4hmmIzI
ucYwhBZwuBq8oWdNEviSvY+JeNV+IcToWtl25spuX5hhyXGagM1eYstD909+CxWa
3lfwWDkn/fxNT9u8vNMryAt9AY52WOK3o0oPVSKkL8x1DNaM00w8wMQQSaaS24Og
wL8faLX4rPRwPl8tvSd0+K/pGHufB5c3AgfAkopPefYGSLVqQmYJJ1U13pm1mhqd
LXLX9zMb5vJo52ygekEXr3IOiWbODqv6G12qikDEQNRjKkV2+ptG2KqmOKsnPtnR
aXXky46+Z/xwzrbeXORy7SyIhvJqXB3RS5vWlrgXOhGtH9MgYK9nMKooXJOPKAzq
FnbanKRIZPh+CzuXZm8z0oVARwnOCgWUcn5kdbzfQO7VIAIPaMc8bZBpALaq0Pqc
PIm4OCEvBxvJCnZI7FPaTqPJbB3jynWka/rCvEBZOdlvbZUS4Wtrc1/2VQq8pLAK
aeJRUWqH+9SfzgqkONaaP3PNhQT56xZ+vEdsLFLfDU5hF7H4nXwpGqwhlsL6FvtD
WLB1FgDcHq3nn6l5z7dQsOmOaZTYHYDi/fmiVOf/Ob5vvfMFmgs7JFtjzy4uoarz
NdUJC/YdNbrTSIXHQgeIxqSRilIf/O89iIPnVKpN9wrOjlpobf4bZLun1yXY+ypY
U1WPNwmBnZ5yQWAA6oEocv5TKKKNJ9i4dST2kU9TSQZv12I3C5sTxPIHhtftEICg
XHYvurXk3ee79bLJ+7IJIoQk4tM8C/yPR9myHdMjBSahGIQQXhqsCIhP4iqQqJBP
euaccht371NZ+ser3w3oe45T7evtZ0ZpsDXkHFw6gRCOcceDW2Q3pExNhUKMAwL0
LCX3hyBPpLphQ1n3YAyx4tmBedQ66qF/PdoXUUBwdjbS4lhOW4HO+dY1b33ofcTv
ok7lpnEoQaVOOuPlVeL9gt8HrHNm9+Eo1WWjtz047r5S20doHJJzk7ZHDat9+2vD
rzPJcmS1ru3SrcBnR63/9cXJ4M8t5SDGilRM5VBScdetZ4gIeYgex2JaV551QMHK
vtX0WP7qM/2EOHQA8pxh833FWMo47IoOAEFBn+29BETOLhw8vPfDcUjGBdOFcNCl
779JN6uz2CNome0rV/SL7G0Zg00I5cnBq4a5bJJfbtyUmjtoOzlZttEvTAMLmXtS
HiEU1QIdFNRdIuLj2zG35EX2fP5gQv5PkJzbtP+9f30j8wNEX/pR7ntb7dcttBj6
L6T+niTSyw9LKgbCfpP+ZvUlm21yuJ1TA1+40AqErlrULbzw+Zak+8soUyKc6uDq
nnFVC5+3PGlUgj2UOICYAEd7Ahuw+53kQRWmKa5nID+YtjTl3g/cfgDlNSL71+rr
DlteNF1eb/6qTcvrwYQ1eBAOQEycvjZUgeXIs75soB3uWFgjabxNrODCWER//KAg
3ofvETSF2+iKD03y307/Ru94cV0Lrojrq0lsY3dkIEOlLmbcDKD7IPiMA0OjvwHJ
2EhzSiLIH0UuxOi1kNF44EzcMoYbn3p+wAnwJgCh2iJ93WajLz+z+PEqUwMeS4sI
7TQbAV5StidTnVpERp1T5GF3iWIjb0tRHrYfKulrTLZAkSShf4TxyTQoJVlqEzun
Tui/twKyMHnvX1/MVIBWQuD31Ejmzkcbu12Y8R1S2Y1Da5kBmATRXEF4e0EvnkMd
1rN3UqkXJDUalErNYriq/HWPv/dAUT4/Q5VYqcniLlkp/2FPQI1DtUymSPFbxWmK
UOr0r61MGxmK4MsgbvbgVZdY96UxykPfO3X+V714w0LFMIu8+kNtJJLfZr0+F9Wo
L0nUUVWCQVPD/DQ78M7qGvBdfNbQODQQ3XNMeUFu9B4ko7By4wA3sQqcr7y3IdV3
ZP2lAJ8fM3DxuP0heZ5Bz64yjjRmVz+47pzv7QUCEjkGxO0QupodL1RD4sy7exAo
SeNB0AZRF/BmBC5II7p0gJWgcmd2OR5ry/OIDmnhJIRdbeHVOJOG1BcIsGuihwwd
uwBDrHiO/f5DyThzT/T4wTAh0KPTjgjOKi/cl85lqlk8b4WoI7Sdm5DOkX0mNLLl
wOvMtJMrDAKTABHK5uOzfVrkN19bzTthbX6Dcu/aNHbGdFDBkc9PFVn3eAqhBmYv
A+72PWhdC9pa/cMMTMRbaClBsRs4dcsYm2NtQxlTlKcY4PaQtZ8/mPBIrhOUYCkN
cMfu2dqHr/TLBsHRo2jyAgTbz/QpkMe18+nMHEaFfLzU1woErJ+sXMjTqFQN85tY
RHxM+1tzv/Of6TEjKObRwViBkuev61ljtOjYAb/pdwFqg3o2fIks+eMT55iol5Jt
CIAFP5yc/aKap+uDTH9YhjTEIJ7IY9ocdmXdDcFcoaHwjXBZcmLHvMFEWNeHh3/i
IUsjB/5L8YKqLr+hCWc+/Rm4hp1LfJbNlx45j02aUkSYsWrI8CrmegSNBWDL8cdA
WAjuY0LcpT6GiWqc5mltwpjZxR64XK0AR9weE5H9oQEuNw7E68QpXj0nYhd530Tk
G/KUgY+dYY1f6TKYQQbyh54gZOQpwOBtboMlQ2Ik5PNa/VyIJl9cQdGccDaTcMkN
yHZfXn4sPPqAQ4vG5uVeOlOk70TAMfCbc3qcVYOQpCbTArPjRHrkOwJoTjzq5Woc
rmxAzAhQ8xDGfZMUgL8xWZBVRtJJe+QemB8+AVjgw39Eb2RHKrCbS2jzGedgOwI2
mUwedqJamF32Z5DqHpcDtz/vgidqHk55/2nYL9FaDsO3xZ00flQq9SnZeVry7BnH
zwvIqhberQu31XM33fWbCI3uLvLqbrEiYZIyIGir/jfYMEppjV/rDNEyMM50wBMQ
P3xcS27HfZkgf+TVM6PCXIHZMJaXTmckS9FpeyP7ntB05qCTrucQvP2THnpkf5ik
TruBJs2pE2a4q5qXW3tn4axn96OuUsOZ9SIJk0WZR7GeHn6T9BcHH33CTsZHpRVy
reWID9FU9aWGFIYe8hMEU1XWgwBy0Rs5lXOKcU1CHvj2fdk40EyFhYE3KdlDw8xs
7jQju+XRYqtSYSsjk1bH98pnCcAnDPvancsAu2qkVvTdc9UbfBQ2U3sSOIqun9C5
7jPFIZFlIi2iB3TKEo6b3Nxi/B6RU38XcgBNUlvHDzAShWi3nIZkJGIn1na5DXRs
s5YsZUz6Ti2+IP8yyqA/z14/3upLQFZCpXhJUaeO30J6rf9z1jXCxsWnv3oXlhtl
Y2Kplnkq5WxQtOemd3+EA2q8LzBdo7NVzxQM59prcFJAAqoj9jhdVne6F/b16VWR
n4odb9wV9wdSI0mfxqQn+B8MYGnvgfk/tGf0/KxI63KDm1hsQJbNRFEiDZvOrHN9
AjsNnTFKgEW2dHFTDPbAqOL02tsZP00E63NlkAETLDJTV/ol4GmD2sYPnVCFDMoL
jsNuL6VgQtRJ1W2NeehMtMd61GOvrfqJ3P1+7mhRiUwy9So7wnyOSy2Q0faGyV06
6Wi8TG425eD7Us66qQL6VSBmWNdaXo5jO0P4i+3lGtCXxEksAcZhQskkqviWMqNI
U2RGjqgqJxj9EpyKnSHP4wJkn/IlPw32C7jZXSKnDmnR8AbwVddexNMlIUkarTMN
WSIRRLygR5F+11kSndkppxt4baK7Gz9od5r4pSmUCILhkZIg/H2kSDZRHMpqqNNr
U3kR5t7ThK1CDBbM3c+yND2VmyMUpk5vGT/iTowuvmQt5Gt21FGaPu+d1Ojg73ov
1uYMiWfNTRyMRLF76YNn4xURk+nKJPMz1agnx28Kv1m+QvpUxlXKIVVi4Fd0xgG+
R0uYkQG5ZeUz0cAfSYGpP64rAE/IfgMav85wb/7W1iiIMQHWu8R66wJRzpsuVqZR
/Pc0fj1HUJ55M9wPBSkew+rt1nJb9V+W9+YtZTj/ryssR25OLCI/YRLpit7JORsx
8jOxvd5MH+wIlNvbE4kQFGVIHn4GN0SClGSCCCs56fUD9SBYvvtAPjCPkz+j6Bt7
c1V2jfUwNrH24vwrOFwrh4YzhET52siVNPlJDDGxwKOKZs8DcF8yUDDfMdP2IL01
6L6/WEPybjwTzQKpCtG+tQlCGTF5QcYnp4lktOfxaIpOkl5cJ1lE5u2KgkMaQ+wz
oV4Nu9LFlag+IXtZSHciBv1ksB4LgylBs88H3VivhBZ9HI7tJ4jBxgFQ866QyBq5
mvZiY3EWxLRVq5rYC7QDaGkCX6xNTRq6/VHW0I6k5KvaDkYeYgfrUdQZ9iKnpyTZ
wl/CVgFvkgZi+Hil9r1cL3UfsQ/8DBhfTT+ixqayEF8X3UQFPd20u2Xi+J3iPKhL
tUR8wweYF1dB8fP9W9rBwoAFZcO0e7rFHEpyqgPl8Qb7GT1IIy32NIbo8+yqfjQD
ardGiyYzamjWPeTTY0s5LqJDydbR0gXbXbnbn2sXe0azuSQxwECGzJ3ExFpRsVvo
cpcG/DvUqRoI1qvHEb61JyrNAnmW0iBmg2St01iM9SNFCkGpUROoGmYeL6S3fBgY
CcLaD+Aqz1evXASZbq515iynZNxApqGrGIeQXwcrv4XvSmC5FZ9lnD8MUUPvSrdy
o3dSTCsDfttorUfQVSgikBBbIiWElKSji69IT8UZlvFhS5wAT65tk9ppCGTFXm4z
lbaJ4AhC+/+Fm64oxIG0W8dEHDQmEklnBr8iFZPSEDDM1YPV/f7H5aWwyvyTiHQ7
GjwLhzB/9elPPNd0pX++gMRBgWN+D3BDKercn5ULQHW9wu/WeYwnZo6tdN2l91Zr
7VYJmR8Hzds7zLB8oDfK5s7dRDli9JPBApTrxbRurIV9SGa5QXzN4dz4FK4kOUas
WGIo2E2asUAwDDPOmt9ZLCkax7dRNZGUjdCsrndwimfemTHk0q+GcpEe6vZ/05/h
9Y8JDsdC/xE6sY0h/EGjdTc22NorqN0NJaW91WpeGzGwHOfXb2oWC58C2mVhRIUg
gruAlfhjUk89Yr9vvMCUB0ZQsnijdyQs8qVb+jtNDNhYk8GPukVBbbAHzTkLTQ95
IXvYWQRxE/T5XJy8m4OsRb2hr3lq2C+0SIyfs7pobrS2XZ3C+MbZwCGVsLuxnNMG
VcFkDkrqgpbRjOBrA2nThKzyo0e5DXw9CzzykT7/7PvFpe1kTEt6Uxi0HE4ZdJkz
blpeLgq5E1+d4gaOgOA97GhHic0UPM64ZLiQKVFJDs91kHdL9B2HKg0oODW2Rp50
vLvY0EnfRnA36trmzl/nV8yGQT8BmpcFljNwY2ELFBXMnDKP4v6ja92Vl+d5JOiI
f+feGiTmivvBD1B4WHqbPiN1wWx7PtFLrxEq+w1w39f+Muipvl23aASs204kNpbn
RAtfYA1XZDMDdmxCCIMuvbhFiET/vRQ3pBa8iJ8/ECi2NaQDdUTZaJKRY3bnxl2h
5zzL67GSby74MaW96MPLjbOzYCdH8c/8jBVInQbU3h2X4hr6JK8nLADR/enWrtDp
FTJWaJSjJRe8ESlL2OgwuVIoHhu9egiXMKF1exkDR0SZK7o5RaTIYEmQRZcU+P35
SyApbtp1LlrVFMkn5aYYBPMlnKYzZkOVaThrXlh6twbDYAh71/bELUaAnySxu+bc
Z6Mb5D0WZd3T/qgkRvQwzA6TNjmiC0kGBIVj+78rKU2VZfQDWluSAlcGGEn9HMjy
T08vkuNUfNQzgdPHGTJgSfLgOU3l+LiE0yr4QOP4NX3m/T7QKE9NAKkHmIuaCZqn
QEmbU6mQ3x51Nu6+YOn2BZHgPw9p9rNQPLQ8kql6MNhCRVr2mL0NfdVpxgg2zyK3
5Zf5A/k5AfYlsZgygB4I2mJYB+ehRAdfFJ5e1pMLoViQZ7wKLfXto3Gzt7hzzXIL
aAZj4psdg8cSn7aSvCAiQlqDgUR/gocjuhTJxvt3CnRfmJ9FBHNWyqRvM6DTpEMn
KR5fSyKtddbjAnnDudWayeSdmPvwTLaMsN7eGdEFmE7StsqGBmreSfGVawidDLVE
eTz0E92SdaqawSEbTPRrGDBtdYq8w6RcQBSMcUIB8Ih6FIDPYGFlYK2Gk7X0QtRN
Cdp5cc2PO32JXQWHgcwjOVgAux6nXqopnxJmSuzxy5yVoDLGoCMkYZNY3whptm2v
pFu9LjdDmZmsww/vPNn+CzLak3hoY84TtzA1xCnFcMjxLYwnMS01GlprZRtC2bUK
pRuNhEHf6z4p9ZxWav0CxMcseOlBFrG9p8JIKRuQJNY717SXs+lV1YP9Ztf5Jlcg
IOw+VmacGZw/x1OUPO5ZVlwoK7ovii2XB5z+6zLLVTNMlYqC3JQCGAKIQ5g4Jetn
yte6DH8eZPMxyZlY8jcX57TU9FdKKW4gHSlnHhC3UDxTahvG7fzsUH7s7qnCSYvo
6bOoQ6uK8kGV3cYoiU1Hb4rAZxz3zMagdCKul2J91Ow1ULa9geOuQdKOkPdqL6KM
GXgFWUGLZ+f0BStssSNeKphjwhdg7zru3IfOrWbeM2pgQCmGWfWOQLeQr42jFqF7
m3azZ1tXSlENPVZ9U2g1If2uiTPM4xXyQyCBYBDip7MslP4FX9LhoORM+iiDg2aQ
PCwDnteJpeca5a+I+wp+bDf/KBKy94UYU/3CMYn5H82TKm8pbT4W6eQrhwfFemZn
KNkcv51uMmM2bXxZKgPkw7WvHZQz7F6zzts+z7OoR3WcLRrTJdFdAOFJixwOtCfV
ntkU+trsWecx2XZPn46cWFkOZAUm/KeoxuqKfQOGi7JqUac75Y06OzKlxcAaHbp9
9oLQ10nkcg2tYrrfylHqBRnnCG8G9AneO1hJ7vhRdr1DiiptKiGck703nVO6Hi+o
teehYO04LIeyl1tr22IUV2WmxaKBDqU0f4Zk5cqylndSAaaZHGDuFWUHJMv6LErt
EELnI57245W99y8a21SAHclZvG6vimsnPRds7PlegLc/YafJHT0vEFaeTVz71xbw
I65I8BVFegTLocDQ7pqYvNRcALdL8wRFm4V9Xsg0QZUP0g84dUHoxsLhan1/I6Hp
hucDtrRd8ruyg8eMOwX1POXNKQRcYR+Nifg50dc292PIaXiuTp0Pkml2AmPBR6Cb
LcxN8pWT7c3IPe+LVgFLCa9AuR3fUn8x9lrZkgfIFx/azc4oRGnUZTIYrivoHM+y
d/V1aujOtGKgRIb1d8M0Es9egGvmat9ZH3g8BXtaecw4BDyY5ZfpD5igplMvNa/p
GOPt5uP/eJkqnskizFF2f5cm/eptEw90nvjYdALW1qXsQ2EdGAg5kov+Nx8uLKZH
sSi9r79TzKBeFc7lfSGh8tTy1sR+sCO1CDoXRoSskbu8T3lcVHYCJzeDfMwP6xb3
kD6blqRwbjiVCPeLHthrOrREcjlUQGkSomd91849sHKoZdGVu6ktVJyou5IoLU+G
StMwR7RnhLw9MJQvI+SAkXrL+t2wI8R2HoeY6UISHTR7wD6oFJD5M444PZVnE7wY
0wuB+rHUD2uLwTSoCZmMd2QvWmc+e6FXkB533DT++eNyiC/OddfsDsngL2PWhOlF
5+3CRKCXPJjGcMWh69BZ97ijIivuCMEcRoH/ZLeAJDMcul+llhTjgg2yXgHWrQ+k
JHM3/swAtxv4sDQS9/hJkpXpOxpTUicMsqC4YIpajb9TLFWoG1wjX8ZH4T1s1EYr
rl1hjFSoXreTE5xcsJ+6AoyanBUsURMXYNPn2BRMgWqySLh8pYUrceXbAkNCKjH/
KnCzGvDhmb5/AZKxIFv0p4rX+Kwce/uICTDdsdBgLjHx+HDhf6d/xVEq2hcDHJsL
L8SlzRIXoeTLbqpAooCNuPjW0+fpuLQn9fIU67+bELx06Uzg9xa6km2b/qNy7vPk
miIF3U1T8pY6xFSnC2FJEjTapmnTCBoDh6bYljiGw4almz6iFo+ieR6arhDbzKMW
cFN3reR/xLHPFDUrQyHJls6mUGEgUR3NOb57Lz3WYPmf//KIhUNR1ZW/IDfyiA1J
K/mgcT/zda9cYj9RzWYom+aaU7NhYgiqqT0QiIbX32qFHqdbJQ/oJOrqI7LZ6ZBe
gsSes+5ItXCs4jUVYIB6v4CSfYAxUAXxlPTDYOptrCPWdxPxL8P+JGz9QvBzGZfB
+7kF2wirvqJD75QmgEmt6CiSuyrdLO/f/9eXolxSNNI5+PL72FZRw3Qoy7Gfya7J
FdYSegq9XtJT55UkgYC8kWIOaB8/k5E4Ca5gFg26x57fk69Yh/GoApCAdb2PoYsK
vODFCwb0Nm2pI1GonnSjUfsFhuLbuBYWXVcERpvQ3P3QgdeQC54dx/qW6y6TzGsN
ga3z/21QmeYCATMv9KRar3Txl7tpNK4kLl8vnZA+wV39p4QdXgfAiynF9+hMGGfv
eT3XSqpL3yMDW/MWcYPin2nJL9JX70SXMjbkySYBScsXKNUaVKID//PglkJqLG5Q
3bBEB6U+mox3pCOMPUPBsL8EILFuPA72o+y1M5qDf0LkqXX/cta7YLawfqREHduV
VmTNLSUKpgz7DNdmSX7Axu0HZvAYvciASEsvJGyknm9PwvwFMGd1O3jtXRKRpths
wOt/6ihpKRSWpzav2rKF5iVaMiOu/zAAdSAkLAWXza/R4eeSGdt5v59AYigtsqYP
jOSVE7ufmOJKeDi8lex+KNJRJB9DnVwvBMLxS52ZBv757YwqK7nVtjQw2sDX94aS
wfDTT0Al9lQ2+Fsy88Vqcb272JVfjfnZZCyjLZXru05mGFU4Nkj0iEHZO6g8LpJN
u3u9ZVV4rq2bQnrLZbFkQ0TOHjFYAYFyvt6qiVON7vA40i6vsgmP19ifJG1m2py+
XPJwBuP+vrOLNMPPdRA73Kueco7sRO4bjbl/CZEC5cs568yNBUFSFMTYvzgce5JY
Knd1SrSQWO/DIqZWC/qNQgNfiJ/px11FS7FJVsdIHF2mjCOanRlMiir2nMUEwcAc
wF3W36lTuFsn0rs+zMRaO5YflMhYdGwztFD1N+Tf2iFYj/lMvxNINvf/NiilOYUp
/sZnQgxlWmJbaOsxsadtqR3WIRqHkKKlszZQxsxYWLb7s4JDlAdzNKXbt4szyei5
pRxM8yQnk2X5ztXViQGscv2y1duMMjXOldDJwYe1FUAxxT8HWFOq4WiOAZOeLRZO
F1R9qZNAc8rtc+qEfqii3TyBa3HkFlrNHIaw5Vx5t5aTIXDDJslpbhBocenvE7I4
O48lRCrSYOXPNPnTHmQcbb/voQy2pdkSW6Tu2XHQigPr6hmIxttGlrqigKHXvaaH
mf9/BHFFAcA3N5ubdRDF2j9XJfd5FTKUgdiE8622ebNVFLZM9HqsqpROeLVUhePb
V80kc/6cHI4Pby4+0ciXeWGCNtjWOnFZBn3yeKTxOj4fGZHZIUm1zLXDhSZv6awu
TenscA9vvTKLrPNqouPBNWEgCEqaQnhiV5QqH3KZ+CdjjSj41YoyKR6cKavPfA7r
eGF5TfLJxzVf1Or2kWB7ciJYAP2azgfEDNeSuoSVpU7DTlcQ4+RI5kWdkXK7Gi/F
QXtZt7gC/vCSchGhzah1yxWWJy0DaaotgqTIFf8ucQ7seSzF9m3leb4mo+W3RFAj
i/S7etXpKcn2hlgYPfsG3nEMwAhSYPf5Frv9FnneTNNTF3y9+5QODtF81MV51EOn
EIoEhq50WxNw3duPErru458EviQmBFHjXJ4M2wnmM3tAEUPKvQuizTBGz9j8EFc4
T6ijupI5+VYKwvi0sD1+pFbFdRQiz7g81a0vWy6PwxVXFmJidlm0rAIcTi3lAz7f
zGAeuNicufOR1yA7b3CmkAkkRkmyzMOMTB17WtcNIOojMnTVtJOWBP6bTu1AfyBO
c0LcpJuP/YcAg15G8LGyRWzGumyVzGW5rzuhViW9k+1yV/WsAohp801b7nVHf11W
XHHDg6nkkh7qDVf50LzE1dAemoQhGqRvftWx75znIo6iH3bYbkJtmCbFLiLrzqAu
6Qr8GCdQUK94YypqRY6nAnhc2/iqDdPnit1zd7B8JsFoP+xOyPI77Ies/HRraZBQ
qXM9rGgG+VrM95CSHVa7XNgSd5tSM059vThgVht+Z88XkuXqHt+LrP3AluhqkggB
Tn3AIwc8+3MhgcPJbdTKpykcaAqvfbRpS09b8M29un9JgyA6KwEGqWTgV7Q6SLpv
TsLmGvT8oQRxlpwZGWOutxgMBC3AMj7dvH1GS0zFAf+Z4KGY34WNObUMyCIVBjEz
IAASjflBqd9NTj2gmfeo58o1n0vJ0ZjSeq9qMDxe802UXYasAYmG6N9G9y60QBq9
ZpBzmOb1J4KHm4/T9idXC8ST9mHOY2WTnbB/5ZOzetOkSLy0VG3fh1sXlFw0Dyi5
c2qitAJ6kVyvPwpQyo3r77B8dO4yS8vEeIa5BHoPlPVigQ5iX92QiYoVnh0B5C1g
DQTFscpceYWe/Dcyp1JBLmn2wRctYPyrGC/WBvFyLfU/2PzrqoSJID/AAfaK9aws
CI1d/c4j7LSU31t1GzINuIqR9KS8AFym/i3WjehtwEoqfu0J1KHADtQeyVGpUfbv
oGBONHxe73Pmq7jno/2aWuzgu4XrqsQUaQOYOQGEpUXKs7i4G14mjZiOJq5OobJs
tsxQHjE9pbkpTbVodeIa2EszEf3jyS0vblzYAiFUmvqv/NGY8R6w3F6h5TshZWrq
GuCi64BZM0P9eh/E7ZiOaBDCvPmrJk27PPitcoUxCI0e0ixERiRq7quYeGZCJWlS
p49DZzu1SrfTHROl8v06+UT1/nyua21gMNT+b6FzlLeIwecjKcZmbJwC9oENB4sC
DWZTGr2mSb+7kZrvJ7zOec8x2vJAz38et00LlfIcL+zueJnCIswW1RWyaZzO9wDr
cF0w/blruUZDLzEan7YpyHrU5oeI48vX3TTSxlgjZgsmlwJ4DPCtqWc2LlNKEIR/
3gGcVqQ1R4isqZYDxVOvvEtziAKfM4DVm1vSIj+QfGBh22hOI9/bXNMrMc/IygCb
yx8JWkRQcUS9mIzqZZBItclQgRfH8n0Rnu/kwGKfflvq4EIFazRiXxYVBOvyY6jR
sKr/mKJJqdvHd/UzgdLDpDfM2peRhwRKwY0tvS5jJ+72DchSwnezEMAsH7UPzvV+
BrFj2Vmj8d5NuQ7PtP5MONtPDt43ORha0jDWaeaivDkau8uHT/M3WurFtnRfoYSR
kvTZKSHZtKx7U+nNzlKieK8U2esT2hOBTioPRra8WoeFHMmR/rhZrf8jDp90d1qT
Fp6OiTZe4g3JQxiGwLs2KjboSYh6lkv0og9V+CReWa8aZcxkjcZaR9ZlFKNdcMEL
MGdgQVrpMdsR2aVo69kmY46kj0PTO9QiZqoP5BA5hMj21CsawOcddD7RhifLo+FB
jxEkZZUMTjHdcx6rJgi8Cg/A77kQclE02uGaimsfbrLzT+nHIT7StJbG55pYeMd9
W+62ihRvu3wrfgQrLoo387e40GqsJ/BjLbcsPnuSag1dW07EOCc8sXAkIP82MpWd
d2aAlKPlWDoOdZyT3JDNCe9nVjZaM8/+dd/4uYN7cvHyT6fSaixZu96B4m9hpzAh
drbgLRDtZ5/8sDSUZQcgP7YOFogIs/TbwKfH0pUb7eZ40Ut33UZ4aIH/bne2A/kP
ftO8CoadWtE8N5UaChumBHjxSt0aaweVEKZQRlRq69tyfFhvmqmKh01ajpeCiZpV
gLyzMgxhD2N3IDM9KDqaNxiNQsvFyFkqmdaToMLxFnrNpWB4nX61kQ+4/4CR2itI
f5w7+qMVtW7+7WNj/5d3JY0pkjkyEh0i9tH2t6CnYhj2obmgoSJVMB9K6cuOfV3u
uxyWaNJLOBak0Q82Fj7QrSMeKUNwliQpQ8fpTTgiMBPwqmdxJbhV4o1AeczAfuPy
hT8BHVChbtRE42Azs1ZJ8/WuL514Jutc5Z8u87A79FF8EDVs1mo8ZZEICSjQbV19
JeTX2TJqfZCxqc48wdoSPa8dn5sU+ZWfYrRgC7oT+n79OjOlnX69ZYLVJ2V3XKvO
GD/m58m04frWXF5skym6D3pqsg/kRNfDnJjhrvmoq02C1RBM3LOYH89d+k5oTpkA
Su8IXNDEwzIk4qThZ/OzJpIrpAueilJH+CAZnbAGeJ49sT4m1P6cdqqdrZrImqRL
vpEdqRRg+FdfOc0oAAuZCe/6DxUNRwed9UDcw0/1PUtgRji2UiHPOKLFkwBRuBL8
O9x7MINPvU/ivNU8VEwVXx9PIt9bTJvOoJUDeU8KLcfWIVTUzaz6JvXJeVnn2nAu
4x0UkWp3ZpJipPnDwnEXlydKZD+xKw+uF4LkK/31StZADj3pggDi4EkkSrRbzxv8
4WfUUV0EEyREHZ42KIUEEkat5tYAxSPD61p3VTviropHzTCg1woe0B5LqXYtmFB1
5Oosr3g42t2sR2/NRnYf1dRNC9c2E+0jIcPy1Zs7ESwvfJLnfh/RngEgOLgIy+Vc
5r8Z+sRi7hJwujbcFzFwz3sC36H2+dSNUeJ0fF2jN9+/zZtmMC7CzcbG8ZyCjr4n
hAYfvAmYxyoXE6cG8G/yQhTfEfW7JIyWLg9AwT7JpnBhp5JYId53qkYNtQLxqqWI
8Y/UrJJHO1CU7RkMBz7uv0YAxJkKDYJrmRMfviTd/oTxc2mchYUFBbJsSwIxjzop
nXgevorfLodWlRyu6SfusMwvvbUr8ykoMGz6qgzvZh/m0Fr1x60EeMc8QMQ3nfr9
K+nO9adnxl4KufPLQ1F4mEJhotSthjxVvg2qUXTkpGhFF1YGt68ZN1ksNCzz7ECc
5LQn3kv1RxTx5p/jP57/vl39sDeqQyL6+eW9VrhYnmylc7p7f5eurECfDAcN2gFL
hNf7sinB16S8+O3sfZrDX/cak2E73r/6NbyOVgyRkVY4Xzquv4unZ+iMQewWzxxC
CvJu0Es9+PxcaozVPCiqp9fnJ7GUqQBuxnRF6ca3yZcr0+A+JOPBWajZH6uocADc

`pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JECcOMqxw4E2v2fZg7KKkTs+nGERufULZS5wW9d4APHOqrvTY5bndo18ngunBZZo
u1Mu5UmEkVvP1jnNjsdorc0/O7kXfru5DLaOmy25bC97VjD9Wo/SYnytvfbzV4xP
NfA2LVmjpGmR/GaoWUQ4ZreWhLHiBvXO3X3gyXSlj28=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7120)
H4KfTx2nf110PaDQzPTeuMy6OcBBJtdWOggzxorTVy+RGn5+LYhSF6+qoq2iYlSb
OdsySN0J21fQg2OCORb1Mr7CAUB+MOT/QOwF1sTNFBody+wDFbaIIb/Sadlb2edT
EbMQC6lTm+mMN8jsv8Ky7VgruyZxtdwLfhL1tzS87ObxVbsaqYXnoFPhmbtoG/IY
U24CKD+DBCNivatv2p9CceKhrp5+ydpMBDrJNOZhuQ70/iJKhTXt2mFr748sXEEY
ZRtJF2uw7kzkBY2HCZ4iPlHzZJqPKxSxvKZprWuEckKDhXHaarRBYa6HnU6vaYhJ
+ygB1SF4OMwqscYivLA+XU+Dp8/l1rFB40oCbTEcpuDK9QStdsKAmmx26H443g+V
Da8ERTLutoUJVIFqdAdpHKGk4JfcN3ODfOsx4SR0ENTq0jqVrLWMqWbKWqqwd3iX
4hvFVRckWhG2LOz6KMnrFGDESzAGK8DuyU/9EzZ1ySzgWVVilKlaH1PIrZu1LAfW
9n6CeJ8SGZo7xVsnEkoryg02vrv8+Xq177Jx5c6hfGsEIwDEvmOmd9s5xxuxHKm9
tSXTS59BMxtGlLLPWLza5zDQClJHm0HjOkAxsU1GXgYASlo/X4uQgMQMwjes7Ohk
V88CoNwWC9Q0GsqZQjmeCpHWFVAKu1eLX+JBLod42PKLtps4M470cNUDiLaIktdP
UrC8RTIvhY3gfyMH0ysQsGaQu8XEsQU0M2/pv734tx4d8MggD13xdlXoWqJUub8s
eGrSd2JD9nosjaKR/Z5rvtI4q5cBt+m9ePhvJMBIgFrOCJKiL61L7FeDwo5zw7Dt
msZ1L1rPwvqtKoGksDpvZIwXKMCZkFJrvahYxE9nwMsRr6gLs1u91JRvgCIuIdbG
rehrFLNp5yZevOkzxbB1EEoCpW8bXDHZK7N9pqZcONrfIl57VJho02t/TCZND+st
MdxEuQGVnhIzuqGAQ8RGeHjJBqPG6ZBEYo34HWHJGLqTuS3EZdtip5VYPzleMeNv
eXwDbk5e/yxtTrT3OXQHAF/mNU/7fCdFf19MnwMID5WspM2IwSUDKx18T5vJY2L5
9Kj/Q+91cQW7TcVwKhM9adjGH0xaKJNfWPpg9Ro7804UCFHCVv5mMtS/zaoYokFb
1+z/C/xwud124EQMii6nGhGv7/OcrsS3CoZFXoTls+i//ZwHrnM/hn0i5pR1bAuk
cv171CEeZEZPGHH7ts6pZrmaTCuWeRhTpoROMqm/OrVE7VtBBWs51Vunkem+/M1p
RBtKHpwUt+FkV5dhHFwgDPr8TsN/DJgf1PIQxSIYu8xTRXI8yP3LekgC295+zUbH
RMwAEZ1uxsr6OKb0PEwcjwtxus7ClMSUOdEqU1fPwuc7u92VcR5OaAALyzidOofh
wR8IMQN3ex5xO1fnGr5WWz9a4CrgdsEsXR8aB9MBsD4SwRfpAoysPLEvhjQRyUjI
ocSgzTXYdb+egHHUn00i9XNlIUVcv8B8D4lkxUALLnUDGiN4cPdRkjNMWlvYzDUV
89+I8Hwz74qxnYN5rALtiqzsY0gcSF5Ep7P1ebwVf66BBq6tIQOP9iHEEo04Ln13
txQrrdv3GxThyI8ifEZyk49PfxfuWDo0/Yccb9p5zxur8CUXiFS6UUp2WvKNdxtq
7ScMat/nRbyXV3giLl9Htiifni7IHNequkr7GSygPOWDuWSVizzb/z51Nsrd0Bbz
fAXApxB0E0GNa8ZCkGg4dT/iz/ht0URvNdCA7qVY7B+kFZVxKPjqLv1195masSrz
CZDzacWx4WZFiKZa8jS/iNWWE5XNGzMJ50C2NkJCZ26qnhY4TahHW72RH/IijYBT
TviBpgOFUL4J7cu3FdtkbdpXRkHl4lH+35b0Ao4x/1n6Ok0mWVDALyrdl14mZmLV
rr3vP747bQVEIj3935kDXEHsd3A7027Ya3nqOXIXANrhXyptp/YvnSC93flUVHsW
EqskhfdGQhAeESSfLOyPHaf9X3v6tjLH0f2uhuE4SVpUMG83UUxYKU4exdzQu9lN
foc9fsq8tZp/PQ+0zWnB0FCRi2HOLKd17ATQmjfhkUGb0R8l854NoUD2SoSfgvMq
WwPT3tShH5KqePdcAqAVhOC8pWK1T/R/gybPSJ907zB6iOY3jli5NoevMhyDroja
Mm+hMlXCebCwFKwlcGGKiP0OaEWOTtg2CQeZ2G/M0rHHT9sLwaS+Uc5yhjMrkyI5
8KwyJPCZiOqhuqWD1ADUGAPTA6y1rBr2JI0QSE+a+qXNIsvSqpYY84rT0vm+RYuJ
VAn+nbVNY7YxFxVDa2GKC/70GZ81QweWrSbQ93Mk1ZpXeq8vqUy6yJHxEXcz/Ajb
DciqsXndEeE3/g4J7kPNABrBtJbBNuRw0l694N96mcc94Jr5wos6j0/E1Cuz8oE7
ulVRZSWPVMmn9vfO8sANvbspjQQG6IGLwD8GRme+3R5qbYfRG24EiXzxqDv0y3k9
miT56gUaDESYKIK32A5jCA/C6v7LtAiqr0wCziUM669Xod8FXpOnDYwTCMG1pg5u
ErNLGf56ey10Mty5piVm0oGRPRjPQTpduRJ/r8Mh8k1ROtfmntBe9eGVx37L4o7G
BLp2a6zGRHEDw1Fx1+5FZ45AMYBvE5FsOaf5UER9ONNyiWToIhChdxKdWGB8zKYB
6W1hQ6YDYE4c6cU2W6y3ls6r9hlqAfaE57bG+Er+fT3ZT1itP/Du+HrYhAw/hzJM
fRsZB1SFgJx5ZbEkaTX0SWqqm9DXAAjiPgBS6LLRMDtPu+kxQaS67HE97LVDP4YN
78f+WQqrO3Ag0+9+VOkpk4zpXnVN4JY9bhQxZX8zjxxl5n2fhGNjfZgzPXpNg+j/
3n10JIPFm725+ZKr0RmSGlp9EpSLpfChSGR1Jxr4X3nbGCYWQzuvGrx5jGTNj6iq
TZUzuiTK7beQDJT+4qsinZH6Nuj/FbwN8kLetpEPmoq3ZD8uAbxV/Unk33F2YMM7
qZ60s048lQeq9kDXpn/D9DGeaEq6t19nphMp2biAYAQicOeV1WgCOzuU+pQGotaM
+gf7WVRdCLHOlBfMLcNbsD/NL9kbyFpOaGHf7kGlyP4ySzhNMgBXhfjD9arNxw92
9AJeLbRbDwcyaA5fgzNK3WrlZ23oIHkollSR2q6yTKwe9AZ88D0lQ9Tyz8cCdVvj
vTT1hwawVrL49CfFNkW4GNriBfeAAhxrRSdloRceSj7Cx8C24yZcPVmANm9Ttl7R
C9xJGLDmPm14KRBw3MOeOY+oVQjv1wXd1MTYXthu0EJfFCntL5srHIhd5mZMvnC9
R+c5W6XIQyIRatec/91K7pnXYi3CwZia0aP27oWxRrmAJU1CDeXMqyPHQYJ+1Cys
P8M2MkYTPjYGwnTw+ea6+59er1P+HK3ScggkGWt6YwwkLj+yqYRiJBW5aCdxd1QM
XZlK/m3AmueXUQP5govqzM5T2FXGR2TOQKsQu3BBb6deqcMfIAAaVLexUAtDGZ5H
/inIyzWQpIrCMOjPRmGbmCEbtSl9UdxJTH3VZ/vtv6TLbCFL97mkLPOyCvieigZd
6m6tOfxeEjIJWF6FfrYzFW7nEAe607dbzk9P1EpHSM0Izn3dobogmxCP2x6AXSx+
ItNSseldx8U60hXUW+q7NH6qW5lfn0OsrzYzpr7mC4GhBcTxj0ktgqxdx7N/wrHq
sfRmfr+l2DA23+BGVW5bK/Y/PAA70VvVY14aWB6hrev70++HC7kVKDEATbE23cfL
dVIWEzHzYAehC+Wq27hj0KsURhTQscf+NC5ZSM2W0WfRbRVgJRCm0Llktt5MPUUq
vnGmRqgi9Sqzvlw1f2HeUb08ezhplK5KEvrDw//nTBO6MaD5yepcq3/yZrZ6El7f
+MEc9ylbCCjdhCcyq1cICqm5TP//Ct15XUGcflaeBAfQXGPVtFCwpT2kAetf5HyP
r/wlJbWGFm4JFPaefVfgRVZk5OZJDciKXX25oNsDu1mZre4atFPn4sir8ciotRpN
YGLpHFk1VUkrdfY8AJHCcRXYQIQk/L+jxydOVpggI0uLz21Djs5XeFTPiIto2Fqx
fFJG1XjwE8yzpl24Vu2sKsF7OfbHoITSTu7qMwqnTelk+J/PKlioRC68h0KaMzc1
kuxSVwUcMHBk1xZQOIpxwOlFv6dqutJcyMb8M2oZp5eMnvW07DvSP8HK86eSJqRl
ReOg0ajhuc6w3P2WtUwhcIajiOm4Ra3132Qm3QLR5LpfcLjKD0UYUU6ogsOlsjwu
2Q1WgZx8trZNfUUo3+Y+TJ7z+ffeZubc8B7CcynIkBhqKxL7cbVI0fSAItvR8yXm
CKpJDNgiv1UtQTYkB98U1cixe1xH2pyN8xf0LXR+SMXbpo/spykA7z0WIBj0s4rQ
cONPMQwnN12Xy969MBanAiXRyFgzNcJQi16HXxnDAWBKDcCVHNH/z/PxQCVEijt3
d8tifYDme1qvH/qwNjD6rJEp++7erZE5GH1uMyEFlqW7u1pOIQ2BqK3EUa6cLt/c
TRY8QKp6ianw/ei6xTXvnhI7QmLB3C4XLJDeujcE/lAXm+qE0HH9qr705BW5a6A9
y+49WXujlgPLfhvp+r54IQWulo/1WHrwD6RG0RtQxpxT+XHPNGPrH6s5X6JCRQ56
WWf6COpy6rMGecEkteRx9i/thd+PzGA+0Dx2GVATIdEOov9sBaSqKuXwGEtZz8L0
mNK7au4cy7Lsdac0VdHxMzeLHpTgYWHLqnGlED3nFjkzQjxBu2YbGi1M2bAUeKFq
ws8JnsjYEVG+ehyf+s6hPnZV7cmMfEIHu1zCbnDxCvNQvqlCi1zqyMI+DfiAS8bi
1L2//MfEYmtDtJSlCEFwDDXVhC282RjBuPFsSBHOo4sgTZqcvlcwTkECRGs9WEGE
RhlMcJT9AMVmhZbLa2go8rHAHx9kHb8JarjJ3aSRYGSk8NVy9by+v0eS5eiwv7cY
PvDvwIOTLZmhb8PIeDJiG772wGAH6kFwTfGwibJDO+MOTgAwCAOIxjreJknxWuWv
8VQJizPhjUQdnScwzP+cu3R/vOpvMWvu28OGH67FIpjEnUqlFTwD3UV94JR5Cr06
++A5Cbwm6donldq1eWYeaICJaeigLvoH44yYNfNIWg2oIwY/xxv8chQaurYzu71X
OATurgk7/CBL5LfTk1BoWM745HtiRYnjwA4YLfEc67cFcrrq75N2US3Fbfq6Ng5w
/sZUQy/+yXNXq6YjAyRPzBnb0wNWf+epatPbBtuEcJKDrqZZEgX2Mi9geJ41MG+C
CUKlUjugO/S6snCJErIetSKC/UCvGeCTEZU7Q8/of6ZVjXQjUAFkk8dVvA/3zAMW
HFR58FTutkk439Bk58os8rs/qwu9DfBpXUuIXbX9VygGsfttirlUGkide0B1MpVR
+vfC/xxLv3vNwIGyRFn/J8puvtJSfl1MXPMA9DiYZ7on3NZhuc/qKR4wpyCut3Ke
kFzurG0CVb5PH/Fv0uLauDvCOrpAwIvQIfn2q9OwSDMqT7m7OmIJmqxT3vLZ2B3N
UJTkwv5E9f75FXwSNaXKwarzO0TFAEGwBf6QI5yigXcqY8FC/zbDeisdFhQv8/BX
dDHbbAq38rbbIhFci0nSv8L8xIRZgmA76AF91zBvk8gFUA3Wvylbgr5aJDkDhlqE
tpJQ5rZF1fqp270JCE2uU1/hTB4GlUE22PD6KmK9bE6Ag3RXdYvLxj/HgfD7bGks
0YsJ6Jndra1I9Y5Frev4qaVF7EI5Ewau9EamOYO6DrJVSg7mPHPv3NgFIXmKKQwx
FbYZ0T6YhrsIfFUgF9KJSAdiztFbkE5aJTcP7AROogjTRGF3x/BfmtT2psiF6GHx
5PqTXwjvna2/6XeHDlH337LwJTH3ANFB767/OUM1twErSZ8d72VxBzVhfIxwcnE1
jICUZYKS9ZmcoKkAwGOLSUUA32H1w4fi/0D/YtjHNYiMzInkO8O9AzXOdhD37RDO
5tsaiGxAqRnVwyUh2Vj5tVpDg/E+lT3ywmrOVt6oto88VqTADZYbq3uRIXX+8ORH
gjhtiH48inXpHDbO0t0YoSs1/F9fqdS6V+aT7N3NG9ZsqNB0UpZNk7WKtlq5llLK
c/vl43f2EzBJ1m4HSgo/TDBLKhj7uYx8oQsK2h8hdHxuU/9S+TeC3ItmT9HgqtIH
KjhAs38aqXbGWP1yTsvyZ4FXPdCGo4Y6F2X9iYAOJZiQZJW9d7A5WQ4BCXsO3yjU
YJm9sXFi3qoB4SXOBOUy+Rse53T5nqIbXQWF8GHBVdGMefME1rxx2qWyEBhCgeoj
Ef9V2HvaKueb9He5luF8Q/o57o7idV14WqfMWZaeGFlhN+yoDN799h/TnhhVB2LI
vyIHW0t6Xp+RN4kg/n0X8B3G4s5sHj/vVt+e2AC/yKnpzsIibTsKZJUZRTVRn3QS
RgZ0KVQCa/T1uNIGtAeyihmH8ZNqcYCoqW1+CMXabcBYVpNm/yfexDiP1aJcCU/O
NyOaJmagnVIWAEEd2NbQN6qwCGEVE0EvEX/4w9yuQdPiRK2VNiIMeuxy48SIW1j/
So5UvTVsrQ6bbngR9mnPpY+VRLIG5xWmO4Ww0IQU6oYNCtYP++MYqgOyh+WJyh4W
EENeUyl/d/7OK1bBD9eh/a87Mr1N28OEsXauRbXElI3oNOCMCdx870W0zYng93iZ
J/fSUeaKyD9zz28Xi0gd4ziY7HwbZ19d7du8DBJpY6tYK74ilC+yj6Opko1lW0uV
/1kLeKsgPK3SzOJYLa0yWPSdvyIOQ9+RkPR/ZE0HvZCVA5eBEnjz6PMLDvXO/49E
XYKupTGz1TlVdu5lNGQOKKUvPx6XFLtD2T9PzEwcynb9jyvkyeMo4/NIbD/2QLiP
LfyGrLEJJ7ouh5H0TdpJua5ixYdCMjSO+7WsDAureB4SLDY8pIfuiNw94hVCbWoF
u2Bc1B7j9adlL54VLG1ZvlygnPP4o16Gu0UP5GJ+Sxi1jlxSgcF47p4kgk21uLjD
W03mA5lU6j88smkep9547hYmiGZwxwq7PiWp9EUtMR0LLxeq31dcCAgZywZKioep
fMIH7OstLGDZ16qO9WhbJSN/vCyMBVfOhkj/ZfLR7BPjLaPhhVSEoYSz4/+3QzoY
+tGw4p77bghR+fEjos0UAnS9UWCLPfIoMZc4+Dn8rzjshzPiRk9RXSblU9LusRPv
UfglIfnABss0bMhFOvGfbsb92UPLEYZVR3ctST6he7G9i/lGEIa+B9DvqfsPN6fu
nJCIEs7J/dmctGuoA6bwQWq6SC0CoNDMXjBp4KLEK3sGRLH/NTq6JY8BbNHIveSn
N5Jg6oC7Rp+oET2w46nRmYxb9lNA8ernIyNWwPQxmkyA82Q+doa7tigp4RyP93eT
rEPI7NjyMKwWhOiZYNnUzeCYZVy4UsYREXGsKbnrmBHZFBimygaSaGX29QBD3fbB
6IRlBo0c6pg6wevMLPkKTu8H4RU3pCT5544ZimilYmp5thzZp/dzmguoubW+JZ50
JnVGC78/xolesQaND+E5jiQljaSX06zItmcIeYRDG67GrpIFX16KYwkJ7OyI44xY
AbDYWdbKMICUeaMoLzaQQBliNOYysmF+C0xO9uib60i846dx8v8neZsqmyS81Nz0
Rr2HQFUyZbKaICrJxfj6JCjPnRR8/b6ig6q0s/PMLspXTKplqttgXCGKV8YuIMc4
DqE5K+xV2hM9ggGkk972oWtWWH+nx509T2zUWybQpl+2XBFVaA4v6bQfJGo9dBY+
5cM9l2kyxn2ubhU65h1ypKaeNnSzTevn7ftQQxTBJNOprusQf9KFah2WbTneBoTI
DP20v+5aGJLvwb5U9kabPbO0dTVjh7jEhveWAHKAliaMxzrIHvviR9qTdgbvkepa
VcUCZD4ANMkIQRc0ZoVX0LXp/3wXYJCNyQ5Wgy0W0VyBxA253maTq1lrOvu8GQDY
Qu7PMR0P7BfMNSymd2YCJoShmheRyMUnqWvBD53/en7jENXWXkCO7u7OcOgdmzO1
IKNCPr31/7NBLBTkRHGXA1tr1Rfl4g1DZ870d2NNgVsKghayg7vhNdtBh4N6rgbJ
uLGE1Ldulv5Zhbn+BiRIEv0TLOqzxxD8fWi6EOeGQd9qs5WEZ9H7YxYVwNBe30gY
vG97xhG9XQJ01TbnBNfyS9FBWsMDUDg1OySR2sOl1J+MTTGAmEMBztzCigeGq36/
39VXX+iUI9QNnG5EoGx2hiqjZmvGbBZeNuovfWwHmqiP0IiWvwcFtJMuIQxix7TB
iSG9o50ar4s14VBpHKaZ2HfnTRrftBR49/YitdmxTjmFw8v/ofWfYJY3qXXiekh8
vLuBucRCvnMpnY7+/Vedas5EkHnatzZZM2PLbCfgxfiejr94/Eawt65Ml0eZ/aBx
iTD6Srt7P0tirG0AXXu4UbHNrVxA3DYU4vAajnJb0Vp9dPnX7HglBKeVaN9aEx4/
eXRC3DqvVMj/fxi4CBGdmiQVa5F/utzVs/4fMSCb3TGlHF0R4vmmPlwmJiIXlXUj
0ZBYaAuQRRGP0XLfw2qydhPy91vl+5L4FY5xo0Eo+HX06XzJ2vywhDBZvDxyGQ6D
HgxvCRuGe2aLhJ0nrLDwvBD/iQmYiyN/JuXAjcfC5Z2Svk/2OjK5n2vxTVaN59Av
f/NKmB2uZg2V6ezTk01NsThK/ZBH4StXMLA7HmN0FUYMC59bQ+xoaATRw07NfMlw
5lpmGaqdbd0SQ0yISBkRORkfZtfz9xNYYvOb+3EKldCgFSMfp4ki0sxIa3OeOUwX
hj/fHIpdpgaOyBZgwz3NTz3RD+HJb6QmL3fYg2cVhCSDU8lYqRzPeBBXTERMFgIp
pJS8L62Kjfpr/EHTR5WybuBJT8lcRbuMClm0TXYf/wIOYf1CTdTm3936QCMXr0hp
Z6vxKPrzRA2KyrwiUD1AF+Aw5ksWgVcPtV4/YTVr/rWKDGXhW4AhqrXfhBIKaIA5
7n+GT5UN8H8YQHqIeXGexFBZ13KtfvU//bmTnCn7Kb8WEzltRbNZF/yNaELLQKSn
b0xgrqA+LETGqDdVOa/OsDUY3EOM46H7kr7u7yoFZkeXHM4EHO+//EN6q3v8CA3F
bz91RROKekaPgCAIJUKalG/7lYCCBE2WY3vs0dNgtddfhyj2Y0OY2FWhTvzi36qq
bY8x94H7DG144mSLc6cVfZOavNiADGNeBIEkap1ga9gRcGAUqPBWqf1VSOlitWSX
+0vR3gY5dpc3nRsLboumZjjyq7WHCOFl4Vy5UNbdpSc8+YU4hK8K42vpliESWD9Y
xPZJEzmsCgK13gOc8y5Syf+aQ40wLLf8SvmGWckhJGXA34kejjLXvu1Y/oWVJVMA
qP+jZZfhJBKsPr7Z5KMaiIPWH5jYQveDH39xTEy1fvm9ushvlmH8+9kSovmb00iG
ZgNuOONCTsF180PJRr6W0g==
`pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OhTB2rNZCDkaur6U+SVq8ash5xDkezJpLqJHlgmp0HZmc0t3u/kLABxDxBMEWjYZ
4RAgGR7pCux2mMhO8adfwcZ5tXOsJmhWpgshy/F3H+x9phCiSYk9TE9R2wIzC12y
HpWGJHBV/NskYYv1CGJ/nrV1y1V7rNSfGY9LqqyWuo8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3712)
JQ7xM3XlWgE5GjqCHsi1KNZPaBmoCCkiRtO/uQG/SDhgHSPdHuZa883fnc/ID3bs
OQuDfok1ripfbPpBVTdCWtXFNamsxJRpxNFJgdcWUMpLtxTjgEdrYbEhgHQotiP9
f4vwjTzMYLLAuUjZdMP/fOsRGc8wc3sbOfpyFXWL3cosVdG+6UZyrrwVs1jTjisI
JTgDNeCJKj/v2mXmjy/61pc1HCXXvcWTqF6Oj3VE2rsgJRbTCo44B3bp39mnU/Sp
xr+abLTaXQ1z5RAQEXJH1GoA4WRf8riOlvsX0ynKXnTVHtJgEKzbZSDKNqDjZ3IB
E1hGXZMPma/yDqy/A9jVn3f3jOF6MgCfw2MX9pjfo5wVMJHrvzVv26SbJxXqZOn2
VuYQegAjsmOcTJ9uarMIB/ph50ciQ4C2wswbGjrVXnI4RYZvYdTYuAWvkQsYu0Pl
KHVRzBOqEhshfEk8T1veeexRgUKQng+yYoToV+pjfqxixqze7LFfh3Nlb4hPgr8B
ICM9o0453T9xeSg9ZCYSPkx8fjStIqcflYQorCyAS9zABIQlP/GfSQ4m4KXKmVAd
uoIbgrBeURkoq5O/QO3tHv51DSJRFV01Fy8gKtcabAYYIdTQxDjyFX2OWdoH5AeF
I/qsELpQl/qMgCYk3TTv9qShAoP3IiZlXITl6gzXbXvNBbmU/mgJ9OVJjPU9eXL+
tKFVMJfE32R/iFYhi0jTyCSWAAB3E+1gyz0brCpoyNB4lYeV03y+bmdaUekGY940
7CPlXqST7YXQ4zfegvTI6nRS0VlBWYxEJqvP+yfAZJ37Zr6MeJbtrXVbcSLb6k0O
v7TBdO2+b6P8A6xkbx5zDakoLoqSKNw2oXDNGgR7+sEfGncftBewpyP68e2rB7YW
ApdWw5Wfd94lNERn8UKYdqNx3RUYynbWj4UeQjcbFIUTxLrYDEe4af6D7QHX2Nvm
zTJk24JyBnb9WddSTMW9QjPlnovvG6v6kr1900SkRM+nzOchqewiUYvrJ/SoVa1w
BK94C5TRJyYr255QJlue55Da8/7dtuN3S1pWIUsADdO9fH8Z19xzKAVaGQ9m7xao
/R6AlepNACC3jxVL5N5cP1vA960Lu1NpHzB6ZwDX3wdzwyf328uTZrXV+7lIBZRT
0cIMcOvhm/iE95A5wbaXrEJetaRF7pjzxuKhY+1FB4yDeVI98oLpwaDcFF7LRkWc
90qCN0eorM3SedzHlU5LP2ry0XZAKOkqJYsACCgSaUGyAYgZRQNU5k9QCoz9obP2
V5j2lxkEUv7/3daxjnTHQ1fZ33Wyn2SAH4eyecfoPcgnDPhoPYiaoaVc6ZfQ//5a
KpNlrHr/9VjjBCS/tHsqb9GMXuBsMbnT60fd5GLd6mRVNbCR3kDopcvfi3hyyLvp
bYVbCSzsbbjbB9qp4ezKOA33F/4r+A48SRfT4NMqu4lcCB1ZMVNN2VlVGC1zTz6F
/fe7xw2KpgsJR1khBdR857lMroEvBALHFNjM8zgdmyfNxqw7XODa8b0HEWQ18uK1
OxyQ3LxfPOtki3359OAET6AOuOXXf868Lyo4nQpuS19kzHfHIa3H4QNYuCP4tySN
wULk2Ai4LSzBcIPxm4sjlU5qKjO+Yb8EkzpzxDG/sxV+4N85EY7kgsAby9cWg4oj
8O3lS+P/0ymjSTu21pY+4JY8pILf+d9y4bhhIcWYXC9KkuYC7fOQcp3dyZimlfT2
2io+k2ZLOgaE08btG0RDd+QJEfXybeDNPZOv2E5O65O3AMalXy4287zA3XfypBeL
fDw630YpD7UuTHXpH6hGT5oCpFEvs94Vi2Ou1MpkAaJ8lW1r3+WbRv5AtnwVBcWo
96+tCAlNySFg6PQf+s9pEYk/fdLujYynvMO53ZVSxVYmu+KecFzNChATTFuPLqGk
ETcJy0fVq7auDWBtw7sGy+xu+YtJL1PXA0aFDAYXYCmQmyGiL0Hlcy18d46FEDkh
tG4bPD6NsYkgL6WNqPxGb1INZqrGc5iJ+EM2W03D6kJeqIc/SLwkPXX8ovCVe1Ns
UDCxv6bgwGJ172Ijc55XB2hz5pa5Yni6sc3ahTnEREnbN+iY8UMSvRYnQaCj1W1r
FKQS4xiN1PSpxfx7sz9RmHRDYdAx3PXtDvgKW70oKIdOBu2uiZBWswdBCQ7Anzi9
U7K6bQf8aLq8oBqtsFRSsXvI9IUztfSSFZQzesYsbXtRvnRFjrZQkC23S+peg7QT
gBTWQGmAjfxIndqX3oZHy0D4gBO/LBrbREfyS67Ca5wcl/WtS4SaZuTfm3RoSKic
TAoXcKFrnWkLR75WEPwN/nNOdbqa2t6zvGpvUxh7S/blFV+Yae26eSfekuiKdweI
UlFIBiuwTV0l+4V1O4ZrZSw3oS3aOeISq0/VnBe7wc7H7dpEu0aMHlLgg9E77dgE
RPiRG7Rz6nHKwMtk78e1xNmwXN7HZsZyyNjtqySYcz4CdyJfmXcE9vRxBIdoGOjM
BJDM4yBPHG0LeLyHmUXq86W8po4sHGTCLJnvLomUVeeXEpeIOuV9XwwXrpr4q34j
in6N/jOTKWSXE+H3fNha+MfDWjBXUmF8o8DDocKtzxc72hiXVNONxOtI0Z79jWsN
a4bnv75N3Of+Vsj2J+2HRmL3oafuDR5YJM4RXzL3dJ3m/ZEmhloY9p+VkV+YV5vh
sLH1NlEngVelXvabb85ddt8KxzBhLO3N424pa2nTnsqNoHkjXGVf8klt4URFv8fv
Xq9ZmHvFfYqfBi4O0PjYxcSYWErP6sxgaqOzPqeSu7mvvvCi+ohFz0zYJMxG9sqW
XCv0oCnAPQQC5cEyVWnfpyFyuUd4S8JcWaYPVIh48hCYT8ErH/PS3yUjLJHDYUR/
VI4kyLbjZt1NAZcRj50iBAKmdHQMM8eBCaiGxoJOQR8ToCgHtz/TwKFbNF+WjmT/
2qysSFz3NB8ezmG+0S5H2uUpyqGqanSu8Nh/Wstoq1IL4w9Z1RpRdO9VkvpK8TGd
lIxw7OLHfk2olXUnv84BImydcO3QXepek16JwUF5bO1h5CrOwYc/OzpsCh+sgYE4
Jun5ALO/cgsoFd8JZ0qlBMOh5gNFiOworN9xPLqh/+Xs/d711ALUS7Cc24KjEe4U
WGk/qSSfgi5tAG2Zlrc/wM5cHOyfmPmJ/O9mZcEFemI+A07AR4aeusKxiWg95guL
CXJkUXhUPblm/flsGVfwA4Bp9v6Uh4GOFWwgGihmHpvvD4145mLqMwycgYHPCt/p
OeLuGrOmdcbq2U9Qj0ltPpQEz/sX6TUlMWCyMXb/B41KfQ13DMlIg2USIyBgOkEH
m+3nvgAykBtFEcOy0UqS1zY7xeIuEA7g+7S0DUfcZlhrGrrMUGXzFX5jUw5UsLIi
wHxZSi7uHVJ5JpOR8H/T+0dnspmmtmXJiWyh3flTiAQMSvN+tvhS9Pno5rXMJlDU
4xftpdIi3E8z49ZGf9/pG0mN4bubTju56nW3hEqLSxR0TJgdlVXPuRLd3yjxe/dm
6XCkwBIM10P/Hio6EUVdodCoj11867hxCBHTpY6lL9fhBD56mAMDctrdrdKJsl2Q
T6zyaUCeM5AQ27g88HqFcFWSX3pP2GR9XsjXsFqqRZKbGobGHi2k3pcoLvimsHrT
ej2J8g0/iHmIKlM++0FpU+cbakDrkLDmCU19lRc1WJj2APogrmNKqhcTI3rq7Zza
vO9WwBZqYXgrJM6oeL9qhDvtmgsRJRr1DYjX3TEKHIYGMPYPqvjC886hv1laP7j6
ZYoWcOQCOJMawl3ZRhf9WN+8GUQh23DucQtnruI4C7gDVA54M/9m/sedJJ8S7cOe
3coB1D7Jwx+8buPk1F2jMkqSyXZlvD3vLu0eQqzR4onr5Fs4Hro5+2m+EeXCVnY8
ebJXcBAmLe4yUGxJosR1Nce9wUKV/Bru0u5kMDAt38KVoAmbin+CS8SE7amqRusQ
Ap72HEQAPARz/G50ieAEt4XFw8ip0IeyUf0U7N3QKPPVznrN101yoW8rScVwvO6P
S19rGpBm1rfoecr5AxzWtbk5HsdiZ+pvmOaqWNN8MwNexUS8R2lwTip16Qh1hf1r
r19KMH7wwI4DA45SbPvsw1+SZS3CUY6t8zDt3nHqtju6eKOLTtg/EcPVd2VDfcm4
nvr1k9Fr9UNnjc4JNOOUlhXuTJoiZcUVuEwD09/joGzyOLs3wNmHVENx41a1R2Ug
B6FNx1OqilqDm5BwkbEBxZIT3YMWWAqYD9sJIwQeRk63vow8NPD2Qg/lVTJjCYVH
ZfbBA19I1Ey6lxz+6Rc6CvjZ9a5zrw8jesbLlkUZN6mTWkB6M+a+DApyn3m7CZqw
AU0zsluV9vmfA7s2LjMId94LRrTbeAgyZSnhJ+JkHPSdoRyL6EYtZQUBnKfTbbnC
vbkPWGInJxLAIvibI2H7zelBH48ISvtmqbRb3VgQKfs2d/OfYCv6JjzmFuJY0CDU
UNdkyVBMBH02HXjFm1OAv5AhYdO3GGpUqMqveFQbDI2mZS1Aa7dPTpawJQSUfVea
e9p+Hrhc+pY95lQzZ8/ArHP0pk6San98H9YcCJwrLFoyeb1rj+EpN+BRze8Cedk6
j4oizTI0hfLRSgAGRxBpElKl9Hu6McQu8XkE23kql2aZFHgfbxtdwMbLRZumwBnl
9KUKASQtCql+kFOtGtLQ4EFhHxXytP33LGqcVIAsVzCGVjoaPJf48UKV3jXBYAKv
H0Yo+PBnpkShvnW20l1dvMiJJv+Qjm9MeRoFsjeJfWZVq07lDYASd6LMzSWSOX+I
ABSuEj/NRzQJQ92We27eeGnHiyqtu+eDI0WghhBqSKfLkmEKs3zJJicGVw6VG+87
tnkHDkYJLj7D7nbU7JOrmmwjlpCw3hHWcsztwg+xX2G5CY7XijDYzl3cnhncck7z
OPHtjxyuG+hThnoHEY2n7w==
`pragma protect end_protected

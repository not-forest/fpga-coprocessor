`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
hQ1uOo/C+02Q1AQPIf3tPQvmymh7M8c/1DDDS7fzozE0YVAVBR990rUW6LENtCC1
RXfTG1xg1XJhSuMG02GFxiMtoki7OIzC6W/UkLHYkiLZ4AG3ciPOQtivOL5r0ro3
nyknAWVyMCZNWyRJzwASUPpQBtgCG+yb5pihbXlLevk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 67648)
t1GV8H0wVHSzGJlDxIj2rM2E2vYWeRZT96+J/nCiHz48T8AgNHUIJawZqZWSUVj7
buwX2JUbhsqqdGSuni0PAjBx9iFzQaH1yxKq+YvathAh7etq6yMY0X43ksc78JLB
bqaSY6QgAGIafaGH1oSdmXUmk6qxRJM5vB7dqVOndllb8xHh6ZotVCTbIZTrinWg
smanxLYV0Y0jE2TVv8jGyjwKklMi98oIoEeQZs+veyVaydhkTN6C2sCmhByBVt7j
KTa6uzDzfRgh/NYoj/sLynmgMtG9rSqt1Nf27Levypji4uhsQ5q2wq/hgnF39tE1
NXCGEpEik1HlLBhgZaBTdhWfX2moVBNy1ULdq6Hotpu2c1E6X1InjmkSuCOS4XhL
I3SuSV/1W9XxggvgDqNbmiQiJJSx+NCso0o+a1XBRR7hUO938yPPgDsROiU4f29j
nQroy+sQxXjMY6kKQXqKm2DcaZ61h3c9SiSxv3Mnk5CltiwHDbnNA+qo15v4oW5d
pKgyI7V4+ARp6xOTH7WHa7wtHtU+bhbPl4qJXtlJmYCc8onqYxhLGP0codhCfN+f
5sn+ZePpZ/CPfkDgDJj3XE+JsUVPmNyMDUAFVf65aO0fgtTDQ+HCvDMCAaB2om+c
5h2ccQnLhS++EMHveRXINQv9yYiOGquJcLCkK8Te5yzb00fK2hb4+Bi8WURRSB4V
wowMmm9bacrv5aCh6F4hF0P3m8aYMkZNE7fY9H+GAUki5JOI65gLxPt5qM2Duy0b
RQDEi0UvnwQB6M5SrH0hYdDnqYRayA+W1upwXGebTdljf7QqKaWC8hTYtmQBjHeE
dJ4E6ecERr5RJlHhE3kEZxXLbqdmEdd9nhcxO+WXR3K3igdlH6lI48gf5mMqjJha
yvUf6pG+51UeAfOd3XAZo2RR5jTmBTC5waDLncNI61MMDNVstIp6RNtNM7i0xdut
8wZL9QwdC2ZstH60flSZhZtBvJyNtBxcweQACJex0bq8bkEih1gaTGubR201MMGR
pgVq/Bef9CILWEaF3LoU65mo1XpY5IEzQIlCcKFG67/u8nLyIOr4rbdbVCX0STuw
V1VLww3Knj/fx/4IbvvHj4wBp4B1ALKh0sYzNGwpKBxZ+gJd+JwXFM8gFIbRH2iw
2jA9VuRc3FjmVQDJgbnlVOD6WMsyrnNjleqmXRNOsDe7cNmEmg8dzNi9ZBZCsvjR
SPA8j15eWOa0+umteH84+Bpz7E4pOLT6Qzzegwcw03mLMTjBL6mUdfYyv3NxLRwS
sNu29yEETuWPLTx8zzS3aONh/iupiq5gFofKv4ysO6MZWP4zmUi2OEGuVEyMLkIc
MWjXyCLwgF2z9E2pKpcKUavzAoi8Fl+CCTVwgIG9OBJF63HMMkHHT4k3T1xs+NFX
l95L+2KiesvqfWXXKAA0MuE9zq9DFsyzdF1ek3z3zkP2Wu3RBgKzVJb5oOzLZMY+
/rF5TVwI8sdUo5N6C1shqpvaj6RDeQB7WowqPZffRkJIenNVP0HFmkCmjqk3Ew41
YRSnij7HT7958o3EN05pvDFmZYAXA2ee7koK31gmh7+ZfUlSSpQC5TvuHHwKBu8n
WdZYAd+jglzC5YOCfghoo0z1WK7qeKrk58NmP9YSOOnECmbP4+d5Ln3r+W9sM0OO
rlpITqxzOXpl1NC36VWqnSCyzf11UssqEdV86dG0aozBrU+FEmGfi2NAcXCed5lA
4otaDpfYQ4nwEn5mZN1SiieGD8e9w6ETnL9+xzLLABa1xc3XkjhorjInFJxZM7aK
i7MBb3zyE37IO6OgzrVhoC+DzVaKGz+saaL0lRbwciBxdn3/iNj3MR+3azFNIW/U
r/oazhGt6EPGoETj7LOxe5pz3kdDh9vexxDLFkS0drbUGlDx3uKj6HcYB7Gztk1B
pz8t09qqlSzjzWvJzJoXT6q8jiqO2wPBD7skd1v9QST/rtTD5rVF1A35ebVQPQww
HdIral/BzwxkIy7kA8kWPoh7N5RMNi8YGgwfv3UeLvcQTRMyP8suzdshs5LND47H
ay0MT5Agt905+L/ro0rEHN2+MreztxZm5BsESIwcMB8KlWLHqXUEnybhC0884q6a
4WQqTelE8KdMzjDK9QFDXZ/JUdjJ104X6Buqych0vt1K/ydCcH7mQLrk8+4vr9Jl
lomN/J3pMdN0hbduSonhsE4933xAYDIvHCTx3emJsbJM51UhhQEUBXpJ3nZKtg5f
wYUz842tRcZ8kR5lpuaisygrIZKLsFgI3u1YlqqNvDx/vIijKayoSshlgw3Sg9lj
nX1IREuniBBxk4zeMQkOC0Hshcm3lOeRhWT9I6PAGAkKyM1Au3sGLhzDFGs5pc1k
5qIdCz8QwSwz4J/4k8Ux+ICIujOnwSAc5eGPxyYGhMakCCzG2s5/0UclOI9Ld+Rk
yM2soomR+Y84ZzOeZrm3j/zbr9cqzMWhZwHnuV9rGIhKpIN4uT3QF6XhLqBTIOVH
lBy7EEB8GPc+sRVr5JW90Q2t1FJNujrZzsgevAqDuG5S0BuMM8eW/Mc7jqL8TrZ3
T8Kgp+bJ+2gZTsdzM+t7pwh2odsjNIV3aH9nNKK5CLvO8H0+XwNqCISrbcBkGPV0
DaTxlIt6PZWs/iCngkET05YgudU75NZ7Twt//zCr31J/tLuCRhgLpSgxC31El3zg
me4P3+0NlRQ+fOmDd5sGudBL9HH16CMkcmO0aSyyrsHPsPaMf7ecurZqUrp2IvXx
/fPeX0337Mt92f8lVBXn01+7Aztmtmhifjph2TKF/EV/KtQG9fhaR8eCOD1T4V+p
tdjFW3Xa5zDtbdyWWGoPgPq/X10B7NTI7QtdhWCuBRKZLMsxKBieyrZo5y8Gl3aF
2vCPN25pfUs2uMyw3lGPrQhBuIadsHzNxJ2rUrqALyVaUh/Hgij++kLW2bt25uIj
DkR8oexNFC8A/iChePgc2zPOoDDWQAwjL2hF3MCIn37w3z3SGu4eitShi98QCPTk
gvKj70bIZ54RiRRmg83RUaaJ8ndc+TbqPt9pvInjWCQZQANnVox5Y71v5jujzwOS
ZrkubbGYGcB+bR5Pfoh3zZwgdmFuGOhBT8bqfrYWett6xAbaIlNWin0nAwIiGk5k
eDtO/Zx1qjY56QIJrZZD/qo1aZMzXRVOkitwUldbGuAA63SalPic3c73pNTHhdLB
bx5zg5NkX5IAtfVvocXjGr/qgu/TtTdmAMdLkpZbLTf/uPnCY7IwtL82rS2xIjpM
1pFPzkpu5fBCv38OYbXPucfCZQl8WrDjKDmcI67kk6sCd+aUQLlvzyDcJ1nSTbi6
d8bM8OWEzB60L0RKSTD2wHKsTJbkaLt/ul/pTAu+c9c6aQJbTqv+6HqBRDXJLbLm
/3lep9Kor66yKvkZU93ptJhB1Wsgv4SyV8Oo2VluEqfKJBTMq8zf2XXT7cmzCwEQ
3wJuAsGbKzB2j8B73kOmN2bhomqUe6CxFVc24rZAg+7/rLlpcGJ4LWa2q/gGZyL9
12ls+AoBlAALP05f1YWKIlThZ8247drwUFA+JGqMgQUu7UYMcwjCti/PldRqxtyB
K2tcczo1UR8f2LP8Yomb1WLmWQf1qQFjjCOOJfvVKYak21PViTFYhPstnc0Sdvx3
28MstXKPQsRITBuQuIl0oHzw8xAFhb72M+aeY46llkBRndUPB71VIwKvOqDiIsc3
K4i91wmNIYehx3fJ/YQ5t5DPh4a687l/q97BGBG7mnDnR5bIPyvLqSDKHgiLCJsG
cciATAU24Rvw4x7bhilnZSaOM+RWBFk2E+Tf5DYJ3AXcH4xD/MBhLa2KeLGzUPmj
RDamPZ+6LEIuyMg0KDORScsyXD2dDFlaZnd6Db0Y+sXu7RvwEh4aASjlMjaCfkIs
rmMFAhbCjESpCxq8wGbHQ4gXwOxTrFZkzKN4jqQBp5tJRKkfO7NM3RKNJcqkiYmL
FZ4o/jzYbHNTPd0I8wLRUwCiuGGcL796d0vL2SCoP+ZlIWaHL/ixxQSczRTAZPKw
0mlkPFSrdfb3LxqPH5b0SHz7AVEm222jEw0RP4XKij23a4G1CtB9EClAi39JFhmc
IHs6zqKUUn4mrz5Ne9YdyJzvWFEokQQxt0hxPQN0zrfB6N3rhH4EE+KhPVBDOpj4
U+EHpbpDQC08F4V+VcqSuUyMuFs17DcGpUAnWYb5WWuIvVTxAXD62UK3k1Ug7VuI
bRaHCmoBiwcG393DYNoojPdOCkEgfxn1AhO74blCfGQkUItNB/6cOL9cQ67Xa2HX
4fjtwKu0ywYeawPni7zsewt99Uh3OJdJ7/k334Z3pZHKCX6sdJhWaI6BaH2tkwJM
T6uDq1gHnM9vOLl5CAwbWIjRhtFnM1F6m593LyUPe0bxiy5BM7cYROeSeQUyEyRh
6O9CwlLEYjM0+cZaH3ja2RrTWiSvIQcjI0+TMeLsiZszE6abOusdGexxGp4IdpSr
566b2mea9BP3YQv12ZJA852wvUbtBveDIj9oFtNY61v4B3rh9B9NKp8vYDf+Bs3P
hm2PfYneK/R97H8/40h2R/ZoQSzr6w3of+shFX8hlVEeL9+kOnjxrQs8CWJhaPy2
bCxolY/a685G8HJaOIpQxwu3eGpIQfgE4rIS99vFl/q3p1J2HQBvT6V5O/ElPVCl
p+4aZ728uKWND58nygffSYHKYf6HoyhntaL+w2ZXR+UEW5CCzWYI+ALTJcfNNZIo
h77a+Hr5XsGmgAhuokj5e9APj2gpfnsOEgA760ELEiCtYy4B2AnHvVmjNkRV5bud
w4XZYTJ/fzfZgD+kqYMaaKGlO4hk8UpJvvMxCvM1gKivxs3U7dBM5APezvl4I+sg
M1gGJ21l5FF3rk6N4UfjL+3c1FSBc/w9TMCjs73MVEu92qz5RbD05G00gMsLfFed
rgLQ6aGLYXqgqRZaUveA6dE2olQa/ctrH+LwBMQXkSHkN/j1eA6L/0z+xsKMk0SR
owKubX4dIra5IC5qwfbHRMtwtYJtSPkaKcnLGm8YmOJjhsu1qUTw8RyEsvwNVYao
1aMC0NqIMpp7D5ATgIz/D2ig49bfg767YkvxA/2HarwqFYx+OktWogMSy3sfkcLC
95IS3gRnf6jhNIzOwIRB7oQRRpyGP2Tb7e9pWAh514Ww5v6nS3+QrlCC/PHy1US0
oRZjqaqrpY8qn2syTvyEIauEsOw8vN3xjNaCtTiNkmjulHmD2Gjz0pzhGQdpi/8F
uFW2mj1vJWoynCU4mTR2EHvKIpwMoAChiCpR9WWlllBx43q0mQe8ABxCcU5Ph2ju
AN3k2X1IQhySKmEofq+CYmDjMk+9ghozNBUY18sYUCsqH07RHhzJlnITnAOby4qm
nAd8Aicr9Ca0/o1s+HaRGd2JbaiMhnPAm4+lRSGbjPNl55wOm/YoEU96WBmIuMf+
IWMlGk3KK9HvUYSuTFn//NGJoZ3wunSeaemrt+5ldGFIAu5dJRnAsTy84Bdi15SZ
urh0hJTlpGn4nxAKo/HZ8V4ywNMTOK/ooMClMtIzeftKNb1XW89UTqNQKNeDGL/X
kC1Dlvi6C0YjxUsZS2Ssc2gj8ru+W00stZRNrNTNexuKZoh/HEH/Rvv2EBKSg+tO
fQhU7Cw+x4YiXujcQwZduxtxFhlOZFCTWEw7aAig+jiXORs5Hj9peYmuBPIdjRgi
xADKZuTEnoIRXEwOc4zU4ZIKT3gbpC3WveAqPFqb/NE5gbn/Q+La9znxBpQJ420N
QBJ0x9oy2R/Y++Zpw6UuFMzHn28DNVdDjl9iqn4JSbOW+11UCN8kmqf5jUmw2nyv
QDZJq1yuitTdBN+TKwmtlcOE6pKJVbc9JZhsJclkdGFcWWLY7kFXkvHF8xCgeB/t
P3p9b1zky1Luyhv2aLLllP6zegLqZkQD1XN9Hm9bzBZSgFR3QXTJ5jr6gcsn2htw
A9YWu1UIhf01BGbz1yK/Z1dTQqhMUqdFhhVYMV0RANoB2KsoPblFZoOQBiBb1PdZ
n0D3Eb1zWbFRbCWVUkpHeHb7mQZT/uY2hKIdo9pNs1QELc6tljiSVcZpsd2xqgS2
ZJs504aRFiiALaHjqDdXYPtjUrjeC/PQEb2NCm6eUVO1SYRYqQVdEtZAozGAE8Ra
eO0RydaeswDog02AUEPmltqiU6LSetg+sTN+crp54P/PRNR1Lq0QKrs0AVrYNVlo
ZmMv95IIlImnqONO9EieKWrpKfPzMUCbuenbq1cO/W+OZ0ws04VJZDAP/t72ENhw
r9UiWRSKXSxkSu2ItdfxzeHZbCG53NFFc8H7WRqTTGxBfFvYeWgBVmT+Lz4TArda
WvecYVwT3ZeqyY/BqyAUX4c6KzPQKdV61gqcedCX3atq5cipejAKouLOKpG7ubBF
O/OMhrmXHApOqJmBhj8S5OlykHucZqY0f8zJndfLWEGnN80/CJmyMJNb7WnGnGss
owNPP7jHD519leAjl2jwd0T3hrrB5324Xg3VGU8bjTe0MeclZczy2eHQ5EwJnE4w
HGcadHrx1tDFHqSq4noD/ajtlnTg8u/2Sd6wTcI9skiNsqAdhh7fTLZO/XfK7WAq
X4iqCfqrLs6cNr0cW4QBBWkBTYxMXO+gy10ZdQ5BmUPzBqzr6EZd3R6CwYzJxsJv
i5RrD9c5AgdgU6ALFXWfKCrVcVK/OSlgv1ZXXSQ81nDNW3ML29NgCA4tP2vCa2An
WWcqS9cV+yN0pUbMmuwngUqNC0GxrXUJwc8qgwt0pwhGRy8T3rDkUbiitHU7Jvgr
9rAlNFjExxjpdw3EJubeo49fC8JdvQbp0kx6YdFL592Y0gB4/0bPweK9qU741RYt
57hF/pxILeY4jV0x4Ch/PzRXPPNxVpWPzT2aLJ0hC7poNnkec0XJ3AGhG3vBKxFH
FWSBMsIiFDoFy6RFT3v355J04iPj1VMrEHrjgkvAFbERwBJe8Qu4XeDswYOUaCQU
otRXYvx628XU55cKtON9x9wsuLfb2E6JIqax67wXb3UQBNJilgVbry+fsBgoOnbV
uXMhZ2VxMG9Zl3VURnUY7R1rvh+JP3o7Sgi3ColQhKuRzvC4CyyMHPq6WIyELOeR
HPlzPOmFr/sj5/OMfuwz5kmGvG2AKMJoKXZ6iuxWN9oZ9XRxphegSESNJmZAc8Gz
42e5OBwjQLOBsY5ArJiqJp+K0fgHncOSKK9RB787nVkaDXJDyUQNQm1K1NTwKDuM
nKPNJ4TgsT7r8r0V+dDqEaY10aIcU419Q8/4XOGK0CgWktEuZRIRQzVnu6bYLGQ4
ftgiJyA9CZXll7p6tXoeHn1jbP/TLCafuk+rxDhArw/hlWUT5mJpxhKLqwOjGQQ9
50aPuKx4UXv4bBbzAqwpMlCuqsXps+yT6+EOlcvdoRkbNs0VZ8AN9FpylxhRP6t0
dt+N+6T+ayvRZaOTlm4+4d4mLF4EMkP/ByAIs2Qowvk3i3MMuKcOYrKWM97ZukPF
Du2h9TbLc3e5sd+K3F5yLRk63N4xesxRYxwbz2GPNhNibweF2EM/4mdxFHCzaPlR
BXlt1hLqcyA1EJwrMUKm/XfDYCqOeqX89q7d8V2Z/qAhlmsgpEuNTvB+UJfvpEbK
i+gg/IQltX4qjwuO6nC1si+6kIH7uZ2GyE7Sqdp/+AjmF1NWRzEyZR+yJdYVfTu+
QRBPwoAhqL0ZB95bVw+KXt5zgaNGq5Kva8rhErdak4oQxA0sOwuqyYBHxpUWtmsj
kREE6lhV3pRFDoZmq8CCobUFSX7YJ1dWWauAcA0YXKJlOvaxdvELq/fV/tfNFI/M
4kHwX7eNhkIUN33+EHnadR87uQBepwK9N4Iqm1LlJGQfIXLyt8jWee6umJzdlZsk
wdgEd/lalaBM1WVW0ifMhf54rbTK9adgtwzajBn2ZpYOxXe0LQ6+Hi9RJJnws0v9
iKZACmkE2G5oCZSy+gQJZ631cc4ACWqrACPoCV2yVNe2VS8qaS7YCyknyCM/zR1N
xQ2wkJEoIPqBabNxx5Fkh6tDXzC06XOLXpYIkMDnCMkl39RbAvzZGuZor1x4UFz+
J/A8njrC+N8N/EPmHy3Qr8h1EV8nSLZ3h1M5hgGWdSkjewXpu5kprzf/mcVwyrAZ
IlkMB0PvN4DK49F5aqF0EmiX0igLGUd1ec1e2/uixyg7+kV9tX70gNb/Oyiu9J7B
3sEGqTBguepYiyZktj98GL7u+ygknXlATncnGVf5szzP8psafqJ3kHQ5vx3Zdwbp
ZPn2Lod3AbkIBS5xfItchCZMzatupGMjK8aWTp/oKGQZhHz1aL3236+MTLTRJyG5
t4o7Y9fdRv2EVPviuiHAGtad3gtmVECvXUUYub3pN9MPaYl6ztbc0tIGfHHLZ9bk
GoYPdwmqiSo54ZGjJRBCYO79QDB1r3loePqkmXrufRxQ9Jv8Jk5XwSrv62HrW76c
BZOZPZGNWyz6SkgQFPRhUTVdTDBAOAO2ff7qSOuO9WAcT7i6r+ExxPMoKMAw41zo
M4CWhWAohXhy6LwiWHHcwPHjcLTXG7WLjf6QKWdIEL5Ia9FKTCKhAG+4Z2/ZxI29
znSnthCBKoQLdZHrdrYHBYpZNCLFypE9AKd7QGIcnIhWbNEoHCjeah/Piu9oAY0N
iaQr+Fy8TEmKe+T9qudPt43Yiv7ANqEWMZgHX162jVIONdoQ48z1YevtDihaf7++
PUBpEo40ZxYLPTQ1OGEsAbmYpHmyj2JhqLmmGW0ik/+BsstxM3OnOws/6/X9IgL5
uqEgvy9dA0CkQdJU0k755pcsB3SFE9z03jDuf81S2xMev7jPPbZqt6lBM9EBB4FH
OUJLUPX+khtONl3vXFxH+NGGuM4jtnAvS7rtfPDd4iFliWLhWxC+Ze2fzn/ZjwC4
DWd4ouSPuzW54jWrsQzHVhOJnUtxZ9eUn+LkXfj7WEl8F35y7K8j8Okv3O5o9dSX
/jLO85sC5yfk6RhX859usjsxZm7mkg8dBd9HzcpfJUgYkO6KmiyVzwlOxkqJXp73
+Fx7I8G8F7k4cijQfiWwnDNRONM6oei6RV26N8StlKg9Ngv4JjhNyrxF55DspdTW
7jq5FukxVf49Q1Ax44lVb996ryOUf8tJAD+TpOPRySwRO7zGQRlm9MBCXy29icyW
YIez9qDULqfSromQcxznN9sCb571vimQMkdJYTR1Yc5313VdXLR68Wzd3ENIoXk1
5m+P7hv3gKv4wVOpxPlz+r2gxD867CbF4JSvtiX0lMQ6Y5iB4Qo8TcVTmf08Sigy
wI/z9Fo68MqiATANwxowovaS3d77WHJjR8kob+GpddxZ3LctL2x+MG3uQRLiJAUt
FPWEGWlSH6EEgi7R1JZp91b2fUTVtwf6AejenxLuayHGb27Xc11RUuclx8+Jbq5d
W+CCElKN5RV9usTY7+hc2sp0hNytNLGXv3A4ilJLN+b+I0V0ApNo4xfjq0348Hvd
yZlHLiTNOVqyqs/ss1DfPEFn+34vWaDQ4uTGIG4m9R7UENOTu9yocgoIAgWDaLqK
EA9GhsbWD20hzPysITEPd2+MGdwnwidjwspvDR5nsk8lcZ122NHbsfHnkTGzhFAE
kL7qzIGpk60Q1DGFpUsmazrhdw7XmM4HQEQg/uUoiWxockSE1lHTHeL3/5NWrAQE
7KxeOeWyd8hj1D+7om4FPc8Fqfa8mJqgYkWRouxEyB242mxxCWu7BhD2ouyeRKmT
raMNCv9/gk7vfCNyg2kcvn7+ujRPfZ5nT8btzX3rle0RsMxtHTMIwYtUWwSIbYfg
uuBfXqhZG9f/axQznph73X+KcvnEr270Rpwad8VPQlKG76XZi677E0yWXXJTI9jj
88Qv2GUkmCRuwOT+qhNCW8o4svK5NfMnK/nmFmN+0b/unAounxtWx3a7YmME6hZ8
AlnzJmYLWeGYY7D4PKRtEdnMwqts1FaHKEU7uNswrglQQoWWVY/gNX07K0mEiaog
japykirO3u7klETCaugNuUXaeWktoFYJOu2T258Oc/ia4O8EKS1nTlSsksuaW97F
GhE6+zdi2qJ9g7oFA27FisI5HnL7qiYzKQDvyFFRPcWKPnsosZtRHy0zgzAKoEwE
RvkCnlBlzKGA0S+dZr6IusUWD5XD3IgVrQ+EgQ5ulSMq2x34wwz6p5kgyk3dnzm1
Hw+oHCafNKxXurOQwG+kTrA8mfNIYcGSXA4XBNNco7CMZgiLrPS9YiIzv5ELsuA1
M4jONmONgiBwDB2nLp6Q+lUuJuupeDKtVc8QFfJgpTmal9MoyuOe9K8Z2mNdWw29
FW6PEhc13AVeDN39s8WyZYSqOJEj+CXRcnbV0jF+DWptjNuTO9SrfuJAZymggO4j
y7Txc4Ku3k1P0xX5dtoyt4MUlUi4T3dt2HryDhV9PzJ+zbdUFx9EIfoqHEUxHPbr
O8W+Q9YKh729fW06LKg4Dqfhm6fU4mAuHNbx+gc+3ErPUD1kzz/41DCkDHlk8o9e
S7qTgAX2fBqVCC2OCBZrL60u+4wvLNcCA0/g0DNU+AgBLF5xqlN+sCneDkWhS9DM
Fxf3NVOioQ4JMpsa0vreufbIqzEFd/X9GOuU2PMZlPE3uHaMJ7Ys75/dwd8K2Y4r
6cmSIbtKaGjKFQDkOTCZhu1Ui2Mr4Hfunvk/DU2/+Za9NzwV39crEt+iIQUp7Ty4
J3G7sT1brbC0Z5+I9n+xUhRfPjQbVyczUWhOhVTubt3N2SC95Ny4ZA2C5ISqmuTJ
Ot+G8abFqc8syKExy8jh31hl4W+Q8LokxwQetAR6Z0Oj/V/UlRjgAV1uKSec2kFs
TvxIgfmHI+igQeIbaHnwmbw38KQkW1N8Zu5yNVEvLD3iwhmnK7nhzO9XhAU6DNXq
fghlis2n9RD0RGnza+nJFGayMH4oHUeJyRW/gZ70LC+FQBfdDXZ/Ci1ylfuv/nFY
2Bg/957KOtbZbUIWHPdhBV4MAHSirjsB0y8ZZ8zwa4Wq7wW3M99vJjQUSJSZOVI2
tilNI5fZAE/RZc6qtgMD5/tMyRzQLZUHFNUT8KEXtSc17E3LEnVQxV5yQMsrNb21
Y1SkyA23reFwjgFJCwW9yr9wEDavl2bd94+kKuF+ITV2yFQI8w6woxL0aks3htLR
JkdMEsEOnyJ6i9UxnsDgkr1AvFWmO79Yh9YvmkYisQ2vzgefrVnVX9K3Kkf3jv3f
w6rSAJHOwP7iGr5AgK36O33G42FZSRLzTytPVI3n3dMgGpboQ3gOhm0wKV94jE4l
l+w2XGeuI8izAvdSwO0o5NeEt215Evr/YhHN96b40bRbsTKXJF4g2ZNYziyRcEjK
Rz+XBZ+zmFSgR3HcJZfo5MNHgG3ESSrTljMlYPUGhSGx/GYG3ETfeFuW02gSbSUu
FbAUtpPW+99uKttwYDPX4JZN/sz4cUdvHXjcAhlk/vWbCagMyC2muAP90C/NmTJU
pIDwdBOo0fRZyss1G+lhdmr4kWVasNfiNGi/4lWmopCLc6Xh2s7zEzIPpY2Q9FHX
RRWcNETOEi5U52bi0a7K9EdNg+CpI1Cn3d+lGp4B1aPLfBzv1EMh1BLxpUuHoDgv
trt9q9d9vyrVWz3hljr/ExF14Ebd0mYbUxmQA5OwNm7+vvhRLLoL0D3W0k/wzZFG
QnVWI9xDphduHQMPmdCzjxdKwdgo7en5JT/Lfnhuix4UWl5sKwNAuF/HduNxaSwQ
PVUzaQkUduNVR8HUQAmF52tO28wknJ2LvigElB2v7PCreCcJTRjJlI+y4EUok9vL
JM70vEBA+U59FPyluwk3HhcAJ4a1RJp9ObZvr5Jgif9aSCox5jZrosahMQqWLx1/
Y1CcnVG1hz0EF58xOt+mtJBDp6kMXprikNgqBOwyNgIm1IA63gGhtNfGlN2e6jD7
hGZC1NsEm7/pEkUnXahBgtisJe5g43UK96WWSR1Vo3dZwb4pSErAt6lXtrdJX+N6
DdG9QiZIwwi9/bhmPyUUc3p/C92a6sRTgUChqtK+8hQjA97lwSf6eUMm+D4SUSpU
Io99Phu9g4TKQT7ps1TXmQFj1RMNjIzVJcbKWg+MwObAe5Za3D/zwQ6Fz5wKU0qW
OwMOQHJN9Yw6iitmcfe4f2zftpwMkOTrvPE+vzky9/aAoG3eVVkNz2IejCL2ytWS
vYwqpZTvSz2aUZ1YWHQx37yWQbExIP1hfkjvEkLwjB3poom/YNEF82TCtiSpcWEa
JRVvS12Lti4dQfbAUPBzwXY43fNWvVvYPE89BVRtcSA8onwmvlau+/68IocKUrWB
LbOVbZA0ji5Ae92JebM6soqIpW0A7/h8acTkSEvkZkDpRkdZj8xUAy7AWNIeTT1b
PtR8UCNCO14eb+k2kmB4bG0MYEPXrk/+AHdkNe2nOAI810wLRFvPv8JIA0Y3OZBH
8CSRGPkB6pmC2GbKh/dIXCkz5d2abIjMGrkQbpdzO/npK4Sl6EvLtJlxQ1gwerm8
Jya6YrBqEzhMFDHVIWwUaGtwvRiA6VO2c3sayuqhbawqZlZiE+Zhs7Lktc8xHAPK
FPxmQBfHaueD5NF50zlQsU/NJrBKpAqfmAvhkxpRFMp1H03gpyheIlr9CreOTPve
ygwVt+9LBtS8OiBCgl9Dx75uE0iww0ZfVKbhqDzGb6w2njkzINYBUKGYMYciDjRn
jy5RCimPtStRn4y6NkGW0hq+U5PruZl4daEOYEyKPwJQ8iABqxQNM7z3AbJ1f5PI
1APck20IXeiiEc8l+vfZ4YcjGMK8eOhEoG6mmvLE5FcPYZ0fbhW6nI2qQ2jMEyXl
lVlXL6miYEPk4y6g00/mQZNc+euySR/X8GVgcIkCToJDCf1Ddl2PcwL+V/G44L2E
tlWCti1id0oVgL3BrFGxwVdZBsBY3uSjeMj0qG+tDmm+sB0Qpk+ZS/EfV5iUkr+O
/lKl6+AqmQnlmLZxXAotoReKTtyA1Di9RXwAY/PxGZUJXXlZ8IJ7JBlr18zOOL9G
rAKSc+RSqoIkxL9B5Z0PMGYBqtkzRfFgjZ+b9ECnbxO1FG4eOjL7q/+I8gWbfNvS
jIChVAfey1pUJ74tWmpQ4BaSydGuMaGvtOsRBv6TYnXIdmDa4TJIFe+4+f9/NZnJ
PAxGM5ucGIAW6CxOQzr82Qhy3kQxvWjOQptVnnwulLX4otYhpcvTesReRnxQ0vm2
VAmL+WqGo1MtNf7ouODgG+2nijwi0p0h8wJ2RfNPbSru25O5II0tLCJdTib51idd
zrO8n17lGNbK8uzpq8f7tFji+BFPcF8TiygRINdLRQluflVZ1qFqqKic1F1TBnsy
a4plxoFaU+Avr8Lm/zmEwoMFcFRHIIXk++FeyIBf2pj03oIbBmUIoUqvLUXvmzxt
pJF8PVeLvhcqn2hA5y1D1zSZrzS7nZz96GKelcHUwIcRa4v+CMJaM1dLzFzUFvJz
7yX6g9Y+XezDuHqUzkp/jhRLxHEXzAFDJfxWjrGB7JjXkiiw1K2ixABkULCFcBE3
jPUj9IEE4JCUTagFkQNwhmTGy3TIVOY4YTqR5utuFVMpf8EhoRDWwSiztAhOWSea
PhEYiKK+w0gZc2/nBSq7fHjqJYPCxs4CgZyWguRLw8deW9WOMcZqzMbCYM0Lkbv3
NWgHlTwazA1HsSGtzN6++pzx2PMtkxoKc06iEHen127eudvWxUG8wHc+8coovJnN
aQiFGCM0rE2HlWZiLVE5hpsEGRHES1cicllFHaRSMSTKzwJcQ/NSPv9Jr/NHLPFu
Zyma5wHK48n/J29S8cUSfiNrP4ZSDvM59QT7xFvbeXn5aRp6ZBc8XTMhczzr0WTo
hcpwTQXfY1fx4gLVCFeacrz9AqYPfNb4QweEy34szuOkoTqPjE0Q7qoqSekZ05W+
yUWvuzBi1GhbcRCbUe6RKbFNmGnyknIHk3tymr7cqmEGru4sppKkl7Ltvsp4I5eF
fVrtUT0dBmoUyG/XZ2cXk21fYZ1XinTz7qh5+b08XOpGcircHnGqqz8f46I1wGRQ
sIe+RTwBkSkFt8SGvA1n/F7KWf9TcryKPhfCj58Y7ghHh22UlKQeDkvn1H4ch4Na
Gpr1D806k2psq8HHIxAgSQbAU3HRLImG3oXXrBgZDiZF9BMyipbPSd3q57qraA9K
MvCECT11F0SRg7MD6grHc/XZWWv2AWiAdoSmWwx8m3uG3ona2cSQh0knIrjY6opC
uwX7qsiOyZHPKenU4MnJDtUaq6t7bUEXM9s0PaMwGcg/svVbwt5xuh1Xzl3OXYpm
d0fQJUUgAKZO6++J9AGPD97IoFv06fdOZd4/9C9Xvqv1XeCP3LspCQJYXfabyetB
qK95BZuayUbm4+wpeARxRMBU5E11l22mpTzjtPi1e90s234KErB8YDEXD/x7MHQx
6ssIFjisn5eXLg4XNqNGTDypGFRsdATm0Z8mM33Zqlwo/xlPXFWqnIy5/MXo0E5Z
J0ivmEtLeEMCUjzJ4oFVABVyx2c7ZcFLGzYaXfYqOAOAVbXM2Xro+wc49TeO8EUK
RpHcqVhV8crYi7z0beedYKqB+YTitu2CwDjt1WG7t9wLU9kmLFQKDRPmYO2JIAeO
FZS2jiRJmGslBfizHdSq0I/coV0qbMIQ1+uqK6Mq5cOIQReGIYqZC9gBwZXi/tHi
/PVvZcGakAdtypNYw88CwB+iegX352HI/sw/rbYsn41q32K2f8tmlC50U3iJaGlS
9eY9S5Cvp0NscfwMnjv1TDHfPWOq24sE5X4re8OEsA8xnDA+Guhtf0E7v6XVD3GQ
fgeYI03gCMHOBCjpUomdSggFJ7FEJEhOKFS8Wy6Yo4R7Ff3WxePxc/nZDCH8qV0S
Zyl84qfOH3YjeG+NaBaszJqIK8GwJ+OakjGASEEi62JkpDZf7VayJOdYNpKCLD50
5HdC5XA0GJqN8LbZoPJRWFNK6B+CIQMMU2mT8n7ghVj7JYV/2ysutFd22Qtybm89
q/eecdIyltuHzCpCuJ6cgxDA5SR9sm4bCm+tRbDDj+bDgEeSZPHyuQH+57OGBK1v
dc2Obsf2dxHIzpttXTMJH9qWrKOl8GKZbt/jlYy1bxQi/LBaLrbh9U/uWJpa5t4Y
icgGM5zHKmPBbCKLvgCXXBX4yhlAMLH1HvmwdKQpcSWTkaY9WjOlhAth7ebx1HFh
WHj78zryQrLFMf8pU2DvLMOym1Lgpa43MDd6pXc149Yfk+O5nxDDAfLSP3YEhkPu
T50fhL5U3cTktlzfZiROUetz6aIJmEOJ/MbFWUjeHnTpUFp0/bP4fTvhJ+ZTKVSW
5evVrnhSJZqsnG8gvER2dUDm2P5KvP65sJWLGhOcnapJVXrExMMJ+q5Ae4QgW2uy
4MLYFefdJwQComfLQBsuTjwDLkZQkuy4NKeobDfloKZb7BD8JGP2wv3EbjsqPvor
UtDvoKlSaA1Prwco3HYy3j1KpKmlUcz+WjwzoP4BYYJJEK2qipfHCsaIZ7VRPCdC
XvdReCNyl86VndVGfFZhnG8ur6IKB6r+zY8cuCN9T5LZLDS6uO7Pfh1o9J3v6Ix2
c2F/uM/Zlj4FnKjhGUoM2Q4//RISjs2qGjnLlH5xtTCJwqiNdkukYrw6fM832/KO
1OHm9l8G4vCyTHLUNqFszcODZDtL6pxhxN6RiwZzwIkhMogMS3LIjKJ6OYOfUD+a
nb+iQLMckeX38ZXQcuFggMSfhS8p6Yj9z8MegyHNbbnwy6pUCoOAj6g7iFACPAJH
4EmyXwwoIJaMv8/RKKisc4qxtd96jWodh3f31uqJfJncUrlkA4ZyXZYe1P1fQe5C
/vTOJpfA7TIVXdyRjCXA1rNi85OrvlqkLigedR9uBB9A/G9USfiegrjCJ16NhTdj
OMkb6Z1oDsM5nXnSTYbk5wdtqu6AQuE3ofC36uu4IepxbZkqyxixNKkVMni3/SpA
hu50xqwLv84T2+BR/rwcRTbY6W8sT75Co+Wa35RvkRmi9PnBdRxhHwE0GNnFjVo0
y2eRjl+uCr8O/GFZGxscxKWcBzNKBhq+MssersiEoJuEO0ALywu7Xv6IkykY1KTe
0RmWO56MQq67z40daUjsnYnj9TQhjb9VWQeu8Vqm6xqIF14m6UI96CeD6WuJGxG+
zycidM2OP1L4k0GwdDEzA/M/A2RJXNIqEZRHpqTr0oP1Mg2W98rwL0kYg1QC0zeS
b2a4VgmmcpxlsnXUbvKRuh0cuOAxGOidRLVjx3RSYNSKKkE+6V2rrFQhKxdIOgfi
e2qN+douwnM2eombFb0cPdL5uMN9fQ6clHs30OiCq2wSc101tv9AvDXOpw9EXa3l
Tci2sjKEpP/LGzuSXsUsjy0PY33PPnQWwlZzFAJdqxF8sR0mjffO5NbY6UFBlAzs
dn5j6iKk7vJ7Af6sTO5OUwMdXzwbas11DeihoYA33jVzdhHinesiY+BITNaY2pkE
R0KEdUrNM7Gl3YOvF+WHaU4+CGUQazbiDZy+ydwUt3PKmByxXHZWSSZOSDgjsXTM
ombzkZ0b909uynXqkyUFmOWLlhhm4zM6iZ03860fgAiUzz0WPa+8weh06m2b2isy
x2PXoxM2otE7OzSRCiZufwPFDamdDBlj8vGKUacnRBhZJMsiUAlHyQg14BKT75SL
D4VR0ZkYS4RZ4apBszXBcunQ5Tsn3EWubD38/uGJB23oieIrTcFHawW78fgQ8yFw
L8+94z6zTESBZ89KZrhhk8G7QRIGFRUtu18GE5e9iWZqE74Y3qQCpr3JP0pJ6d3M
BMm74nxY1nlTxSxSlbuUXhTESSO5yozJzoSCuG84uLmTZum5cFVElf+q990nZ1aZ
SKZFTHUDANhoorkzIO0yhY343I5no2dT9Dq6Ps++pTyhiVOK9moBtxCVuhlxJmnO
MD44pIMboPbutLhIEzlPHX6xfArG9XT+TkKHzXATzxQPgIx7xQmZV723IxdpNm3a
c3EJ2PI6ksMerUDnuwdvhV3db443IaWlW8Sc2FSC7r5jbzP3XoTOkBiCw1Qvis3Y
uWoA5FBGLmPTPq7ck41lWt41A0vvhZ9nW9+82L2ZaQQxsvtLbLTA0w6+u7dgjJqi
dVyWCe0kiaOuPwd+EQiMD3OE9RlvUb6Ggofl9TaKCy+5RQyCyUIo91M7eEuyymsy
k/2hwMZYOAsaCZGuD3iZVCOh4b76YEMOzSI/Qs4bVOAEzpzNNwn+oFmxxrO3jNG4
AYgV7aEdFpYIUnn1DkNW3VUlLxmh0G9dVB+GKeit4nfIsjb9eA30G15hmyf/v07G
Zu0zNiqCRnrFcbCtvbxBBT4AnBtggt9O1a1re5Kz7o8V2FhDn0EzNTHW+osdAnlR
7EFCsgNUohACyjD7jBLFub54QT65TIUUSikoDhzN0/JqaVe0d34cM1BnbH2rojwP
oYGx43efnXXIrU1z0GjhwcLYtcTj+KmF8fq72/KfLrQ9JajxEva2b19cDxbf2WAu
8AqRcH0O+hhtcWn4idv0RBOZs3MWZdALTp8SRWNgwD+G0mv5wz4MQXs8s2YHSqqQ
W4zyhheNKAjamnn7gRvx1GRpejEuf9QEsjLv47QVc5gioLIeUBy/WQLH47ZfTeat
O3mwnESMNY5bCEtyj3FK8stJeHBC3apzQIlabbOQBXv67kUE1IUTbmgpOIHTB+vk
Sk48vkzd9o9CeKz40alXaFVFirkcrdqE9ki+yDCfwkqHYTyIjljKhAGCKyU94byc
Nz4SSampmoPtX8lp3GcCdw2uLFvm5Xr4rUOpwFysbZYsH4e8+9zlBxwip9sI2X2o
waR/gyJC1i4pV1hiXPwxbwTXz2RiZ12jqHsKYB299hlYBd0CxiM7kjAIxyFP3cmC
+gTA/tMlwz7XBTDU10X2AiZwPBt4vr62vFWxfp6KOoF8N55htVJcR/CS8xhVPpOB
RWp01vmQicRU51zb+Y8FiRtjuYQzdNBnieMHE4X1jbdaztjHTfknqnstkg3xMhyi
BQ1aSlpflcIi5lGlCwg9YbDwI2SSbmtsZQ8vdyxAYLvyMcDTSstnmnBNznXVi5v9
Pz2ATzrq1ySlte5VCvOX8a8Mq4GSP0L8jMGspq9sIPQH+6L3ZwXsVdQ6a61fE2L7
yM0qMqog0DoUb0cDGZuMSvh8nrYS51DVPBi47wWAsCA6wWZElOJEptMVnSJYCc/b
V6xiHX0lESnhJ4tiG9yRVZTbgGGx/i1wVLEmBbJYN2D3JTB5TLMSanLxqJdxabaG
Ve1XykVZ7Kmnzd8G+qIOxUIIruj6Jg5imZoml8Mw7N1oq/qS/CRXPhPLy636Enw4
fHqivIR00j8597RC/QRogSJS1R8JTh/wOGmD3uwST+4ecXjILd/W0JZPJwSn5Qfl
/ld0WiPdr45RSb2aKfSoMAgSHMZNKKeZVfMe08p9aTRQrtNtr+qi88tZ4WVyJ7bI
cjJe+TxBozevh4FicBpLmQbdj4nHDutc557XFOOHT++1M/WEB2rDb/mgVElI072D
XVi74rYsoqNjsanDxqZGG7HKZKHSVFKneOfc0OD1pYG38d+kXqvHcOKx43p1UzaM
uR5Xy0UKDNMxmiHsVaE7o/Y+ewxBPteDSw1At0+iMRgahBKRn4sICWKn2mvew9hy
8P9pYULIdNe02WqoADle/kHkSeeo+amJG7fT0hDkQN0uD5GphO8EBr8nGKQLt3aA
xklgscYEqSa+1xjpEDhq7R9DjNRJkKjcSt4MJ3ka7yxhARM2LVoBXiH0JNZXgiD2
y+iQEJppQe9NjHyyzV/59TVP1WMeYlsiHkeF5/XtdEoS/e5Jr+TmVikkjfK1/lAm
P4w9KGcddrXXzO+yYgw3nc9rvj3QQwWNzhlWbFs3WnCnzqox82wCd53RyKPOyqlj
hEnL4Y1buapgC+D5bT7RJRiQQfQ226rqoBBqSO7Ui5NVIsLEWt4tIzCT4NFjnTlq
To3efaljFPujigIMagRJtEctA+UrVO6evgn9jeL/irmvNVwNd2B4mnvDO1OQq3+Y
xS7rRxgOC6X9yTnqvbbah6pH0mZLr0+eBl2ty/V0LQz3Vw23Rg9kL5z7CxxhyPRu
h1bpvp6kGhTHq/o3jvWRFGK6VDiKPZ6jml+lRNIObqYEn2b0M4RPMEv4RZELTb4R
/1F0gaK9pvotuZPCLqFwcXSGL0OCEtqJv0zKsdsP1fGhrEiXmWGsbod/GOlj6Jh/
HsP/FfwWZDHfyzy5XONqPMIM14tDkjVZseipZZbMdobNjBK3Da0Pu+HBRkJzgtLt
6Cd+q6qousvcfetcbak8BRI4MnZrpMM2GhnUk+2IlXbgPRi547Nav07rAUjyLejc
NDmhuQlVRD72RS1GjqdVaNdkmm7B21okMpBrMcDoKrMCAS3hNQUUghn598UIth9p
08BTdVhd66u0MvQ7VRNSy2KKpU39vbMt2w20fb8GlMQ/5BIeTNJtHLAXz1ycXgxn
dF8W3CGnmI4ul5hFPQdxSL3A5Y9HSp/AOseUPV5VSUacPwXxTKH0erk1NzSn657k
UvfQeZLlajtA2xfB+4me/Lgs2l+4BnTEsE8DFqDiUzBZMGjNzbdVKT/rMwoDAsF9
A+2aOvuRMo7q4d+8FmJWuLUwXT6lkMKi/zJ2W1740d69yWcczyOcs4vQJ2AX6Dm1
mDmZrhw5C/8ob9AGJ96uwiC3fRfDFQfq6qeUjcEgo6lQQmEmcloXB7bhpZnLoOJ9
f3A8CXDue4oPrgLpWr7kJxQHCEXtKOrq2dG9f+m06FcCCtOvbxtHs243GwhJIDkb
Z/yqFcBEzzropo/wfy2m7CsNa9TvUWw8JCaAvuTuLE9saijjfbqJ7srCzU/N9GfK
hmO402HK4EkITFXFBX93ei4NPCECeoJQdW9dxO/EVjiCsAspkVes/qhtcE+5bF2n
Asj9Zcm6vgXficMvQ7r7Ulkl9V6Tw0Lzgqm26c6GSiTTn770y+ygobb8VdeQBVhG
zqbP+CGeF2Z/4049H4xoq0rg6OeINNXoOqvedetUa5YMfm1yALQ/W5fmPeVB0xOG
KyVG5CsJWvE84Qjuq8VJ4KSxQVQDrraiP0Vqnc+nTTI2DrQdAcDJN3nR3jwwXpqv
9kaRHtg804ek3v0FNHjyomvupVFYwgZ4VVhRIc4Z8Yjw47eLxO3hl5H0Olf4sA2B
jZZj9HC5kKVaLDbUmkQvu2fMsLVNiFrjBA4ETtV7pbcU1AmwjNS/Bz9816yOBTD4
qVUajcHsQ3Ws0LLZfX3VF9HrD5mu31BPx2CWvCWczJB+mIaTpLbCDXciIYo0sGLg
upL/kBOoVqd4bd2vVT8+/KcoT+SkSBgKFq1/zTg5FQAVb4eVSVXD5dHn/OE1Xj2W
R4BzJPN2NqTUvUxPGbEexS2MluN3y3LlB8d2jTocyXzRK8qDfmihmDMDuvTTaRpo
M0Unc73KR4F/gOxgM+LEdBbXgLVK5CbgLiGE8pl6H7q5osNb3SS4XcoMnt956+w7
qfu7tgV4YJVnTuj2SZwrTIPecgzZdf2HEnJz799TZAR3Qzq1U0FMi6GMM/lbkmmU
ytlqrUgNaNJnBa2wYpnoaZ0hpgIxdsy/a0px6yAxY7taeA4aN+Wd71Q1EJnCNJbV
n5pK6tZ+cIcOPxevNBEWxZeLoR1+w/2jdVavdSLdv1fsO0ccGzFEnT9lJ8gIllGU
3ecUg4rG/JtLVjfq2EFEhvJO3PsfyK4uzuWsr3PWfxqV1eX4ylMEFEJ0eaKhyxai
kdenoViJhOzHIru1QrKqbLOZuhfiGk1z1We5Sd9HZfAGIZXfJxxYn6a2KyyqX8jN
7URuaAHkg+5Lqn4lba353JAaQ3EiX5HDVDQuh4N4mxd1JjPYfO0OCpdEQxK6uWZf
QJ/9K2NJHAOPeZYvVGA29v1xqrjQoX1ilPlceO9+9vqPW/bTA5hPRgKIm//qiQPk
0HUMt8/24rLQdNzNZ7qttA+2PKdEsXUJSK57In5alx6gSln+HwJgi+SIPmOxsmpF
zizoxnvm9EZ39kUR0nqygQcn5J8RIvB41ZzkW5lRyh/qOqy9YcjgcL9MNoUIQzSp
uiLK4vn0CjyAzk2E6tOQwjrv/392dbJZyUy3K+TQahuOAqlPz7ZlwIkEjtEsfEoq
wQ7Mwxx2kN3uP4zribormFFzGrHHnCzhWzs0GyGlCax3NKsyYQzxQacgHXqUc/py
7vA9glY8HshTK9cNujF+qJrn78boY+o4mL6sRsYS4VZZjigkw6bSOCahxaq97VO6
364uzi3c3hWCUbsfm+N2Oh3RVAXQI6xSuuR3kXE3W21yJ6j4xA3no41k05Gz01BF
v2r6T2bWh8gY361monSiEbHR2HFaZXFY9BAJFy4AFBSltHgZAOp2VWeI2CQlc+T2
GxwmXNKESnW+LYyrtUgoX92I6d0AQxRz3cnyVhbOwz7lqGEzg1fTtyuu8dVPjvUj
P2e0pwP+YlxMwYXnYApLMl1r2w9976YgRHe8iZ8kLZ63ld7ytaBAcg8QDJfazopf
1pXk9pimHou7UhL2Bfa7CTYPrENao27qZ2EaWye/XIS/EiliRt+QkTrL8u/2vsZi
BMcQXa/XK+qmftyUj4qk09n9ugT7twttS9DF7W9SqCo+c471QteLQ7w1HRTeZyb1
vBwWW6U8LaENSEx9z2BiNkau20YDTALZIBmmQTpxI9NxCNU/fcu4h7r2K0Vg08Ur
r82uOhfUZhC8eXVw1ltqzTAg4BvJhHhYOhfwn0e4vdeBq3ej8G5+Hn8r2H2WXDsv
YCplT0TpqI+D54uLOFS1Qc48afVCc3guqpecdNmE/3hR8gdxoMvFu0X7Evt+XUl4
NSlem4I0fXS/E5iNxnGJXqTztROy27D2N8Wu8quHR1yAxhQvJs3xlig4kgKjjBCK
fbOh4WeN1jntCSEPfI7coWVPtSlz1SXQI/2QBkp1BxbFHR1PeRttJEHcxXu2NJ61
r4EaO3/cDbrW+s2MVYuG9BYyaq3OssQrMjraejNy1zcOsFkH4VjfFnNSM2x/+wuU
jAHEA9mgOeHWErTV0LWX415uToZr4tmU9ckeermJaAwtGQvrrgLBReC1E54m9Z4n
myMMAP1lMpBpN5G+fDaAe9xoUCoxT3Y0SD4/rsaV0krn0fbPjyIHuS4sHg0TXEFn
7fwI/iWZ81+eXHg1p+I4TJ0k2kEu75AwkZExG3QTneQUhra4ixJnZavNjlchtW0e
loqAY83QYVskgXrQD0JI8egMIVgYYDXBE5uKMmzKOZXc0DqPAYq86NGJ82sKU2EO
LtUylv38wKjbXdUstok4m9mbZ2ElTCaSyhbEzewsfXSkiGKW0k+ZH3Kxsr2qdr2N
IhzTPNH9b2o6rYkZ+2HO5b90hB8khmuhVntyw9HfGu9De6v73021AnpyWlv06phB
7EUvMmtNR4a/RueBtJjy+4/MNlpRFkUvXh9shgcelGaZ63F/2N29VrwtL3XFkJFg
Q9tf5AdCkgmUVMODzTfJZEBHBHyMff3kHrRZ/8B3H2OHbz+CzKMbQzQapTuP9pBi
n+rUL8aBMgmTNmQufz4danhDRXoi2PNvdeW4BekqkuGYEDgTUV/kAL0eht7XYeTt
PdCbCsvrZZ7wiGkAXiGiY5PaQ/82lKd3peZqvNLHjG0NLox3cdTgR7d2D/BHIp54
W4t+i/Ixe2Os8NbRLhJhzwbko5fzq1HkXwul+02AVShCVBFvymyXe5SZzcLBslJF
yMGLh4wvNgxsgtFZALTb9YsCNxMyGCfQ1+SWN56lHqEQ2v1g3J36gFiWQFkneS3A
lkAimpYk3s/NDqMgYbmFSHxsvs7YxmrZZ4uIJ9NSTabbCd6j19/2Nr0u+gjtRGAB
qFTFKg+0ljGbGwmdp2+5wO9Y9GyrY7h49BoL7+3mK6GDuUjDf6WpMhRPc9NYsVTp
Hev4oMDPv8y/S95vbq6A+KbYtmzZDyZEyZntoxnSht4tuhDk0MXOflFWivZMHafW
neVr7qP3cK1/WtMUQVJjjtoVAd6oy54a06tKQXZUkPJyiIDfWLYd2ST5P7Tge9he
IkeN83LAs5bNoO6g8Z24Z0KyJ1H2uQ4Q7VaH9VwhjcRrTqKJVGRHy42Tv7+CH2Xr
z3k0W4ins7hGxNayRX574jdAox/geC/65j3ewFWZnJTojKxDKsHUiRz1dxRT9qoI
t6Nqd04jDGKzIjG/uXMcC33wiWL++cpfgVWgu9mxFd9aCPsxmSp2Im5bUOUm9n4U
gaD4tlbwHq7WxIFHxXo900xaO6f3asj2islhBZYexxkoPLYv4+StoMEpPTxSj9XM
kC8LvDGdC5nh6l8VfsnzSWl0ESOJPRjDhskNm9xmYSA+ClvePS3/9MPxYo8alEbO
MLT1mWEw2JPQKcKb91ICl5ripY1XrYL9DeUDHW4Ghb5F/xXdyZ1ZwYd5ND9MvAuX
vj/Zg3Bvx5OR8GuGek6lclh7N0aJth1sNWkw6jtkU+ZzgU0ASU8tU1mYX9EAZrRQ
OyxtIxIlAehm1ej73FaNltW/pYaM4bTM1brNsCUfXxvsxBa+SgyTX3SIdeAvTQWd
52YG5bbMalt2mAXkaiymsT2h4Q9ZMK7qoUALLygcp8wRIB86gjcFICXRZsXzOhZQ
XCplrXvYnhcQ83flHkolxt4uhPhU914Nz+RmamRRe9GC9JkscbFXpYUAdsxT2Uda
yZwupXmTKTBs5LuAbmTwXZHS7uyBWlb0DfnsLQq3j6j4zumFwt4b3rJwWjp5VUwy
WLrmrrSraDr8DBW2ROmgyqhgrZPtvLzeBnpEV8C4wTOWBlt+y5o3+tyYqT6q4qJb
QDNRue7oCNtRchgkKKLH9KpFK80Y5zKvWYrW2dRU10g76aEap84N7a+eZ6Nfpujt
EmR9XGNy7YaslL+zY+mTK9ztfxMTp60ai3sPiDr75ESShndANOs5JaJrn/vaflpI
zAcL2ahwkT4tRljaVx+MYgfl7B86288Oe2LKv8DtCmAA8MLKHR4G77tit9PVcm2o
LVPxwS0FsykD2B9IY2IFXAuNkD1BQng3Sbw/FbdPkmVqos/NB1cDhKkxIeQnSQ5f
r0xoonHb6G8bTkIC4sAvIqMmYBx4cndh/Mv5+GwjsBvMylzsfGaqeKTNFdDVCXiR
AdwYAeAb58rWQqtFWXnKP+OzqXzc/Bdp/xQRtN15X3+ddOZHoji/a4E5C3MKhPK2
u9EGzVhwtO/86R+Odp+qxjJUACP/uPDhRBoLrOj5ez3Qp7pRoEMkArtbKEVtgaWo
FI2ho4V9xxVD5n05a46zxPLgy14XB3/FJQJ7Oi6VsH/2FYJYHuKoujrA27pVUek5
yyTnGfyyR1ZDrJPiHhrX41G+zozu16iXlZB//FMlBqnt4EGVVpYGdDeAW3UuKd46
iOdeM5/woJ5jW/htgORbPco9j6oq/NVgrxF5j7bZzfRTL5StbH28K9Orz8YxmDAU
Bg1mP3tuKSVtE9itI4KkXP8o5IotjM+TdZ3XwOOs7LU20Sqkz908uJpjMz7bhNyO
ikliTItGf98fVKulsFqPNHmPBvGVjxJa2GLP5z3fQn+3vr9E2VV97nqTLEGjvuUX
kB0bVxzAodIfUpnvAtqa2Xben4bwW+hBQ4CGHsVqv+T9ulpJWSLDXUZKdn/GjSri
958D7LKiSki+J4WhGo1ocTFIjERn9VZ1fvUfSuwroV4d9PFWBI0ErRWls3POHQDO
yytL/IVFybpFtgNup8z85kSYISgek+fjIR8W9iPN5Qm27JbHHiTSvXLmXHSWqCcC
TBmZcvCbUsB0KaZPaKjeiO0lVsoKtegkBCSszsT1axmNqAPHFNzvYU5eijlOna4H
IQJcGbJIu5MeVkmGT2gIx2E3r6hOdedS7DdOVJXWRpzEQ4IBJMcKwKmESIJ9+5Jx
JQGmdOjpa3YSwBlYAhzghf9pZrGctdwlwJs3Iybzq3fvs4gFDwRgOSn5XwNiwl5o
+uN2/en7GGe6ABvSeMbx2LPx2WU5GYpNYzfuDrSYAceEJfkx2efOKvCQthLL4cT8
XD+t/lgHndGpZvZMDjvt+1w3BBOJud3aW2RTcxcQ/qSOz1MvS4odOQZEpxTtxWr0
IUnhU5yVowMp9ea4W4vv/rPsuAzb6eloIKChLARnP8PUo2VMtTOuJpdboO03moOi
8k/KKUIF7cgGv6+acSCbeOsQuXUkwYdkcwzHI9C6aZ53oE8khZlnMAF2OhDKJZl/
JvK6Ovkmwl9SS0JifnLaxjANvKkJdAY+4JYSO0SAEUr/bvRwrOVVBYFIKfZI5zKi
kYykROWK34xjH/Hs8d3AuVmd+yRXKZrGXDQpb2Ny4e6HwfU99UYOx5dMrrUSShCc
rrrNOcfKOCzQTZ62KQj7vJS21CoJt5vkFYBNAxDLxg/quthpNeR1zAMwIhxCKHyT
g9RYz1zh3fi/mfSI4TD+Fw7dv7H3sFWTMJrIMe7KK8WKT4jzvGhFVlm1YQXAV2JM
tO+odUtvtJXZlVFmUSLjOyfe8kpGyNlWEKkeL8E80c24lynV7462efrI9GT8tx/S
io7bFZGsvnrVTXH7XgDNmMsqeJtpfuFYe931bZmwKTImVCRpH7S9CxsyrV6TriHO
0AN/IVeHadFpOyI19ZL7EPr7jEnH2Gyu8mNf/LcPvFIbb9oGhXohjYfudusM6jJ0
vRutK0Frgdcb9chfAsObgERpmJnRWUrzBSJWNhGrA9wqvKQvD30n4PxybACKa5el
2QPXdLFYHMonCXm+Wubhg7Fy/5xHYCOK+ZfNtB4KfG++5lI1md/aMwaX8NH1xZzZ
uT34UsVMLO8g/ykuoV8yR5DH+ZmBb0O25y3hipE4dqKiacqlLJL7dV//RXlgwlo5
EiCevy3KtHkTGT6nc19ukEOhQOIVgKP02XLRpaLnBqFFouTyBJmT36oLt48sWQ1U
YzA3xHlOrjfgvcWlBz4hcAPypsyzxpcM+LMS1YBQco7vtNtlBXtwKQcPjzc0XkZx
D6HysnV8NaO7oMPeZ2j7Fqqe4s3alPEn81+a/d6JdeqvBc9mOMBHd8MGAk7R68zA
ORIMVKJiCFqmt0jJthKzBg8Sy1K+LryLbgwK4E7uCiGIY/qklZ2XYqde3yP6Qt18
szmfXrtZ7DDaXhwP2iYS4k5SCclOw7GapQQLc9gj+EnZvFGar/Bc9SoqsCsuIVUU
BjNV4YlbPIMWbc33oH8YF3VKTg2fHw79nXBRk89pBdecDLHXy42H2ZkG9KMpcXeh
l7Mai7ZtiQzemea4pr/jLoPslatUz3XiifibkuukAv+YOBr23qjYpk2aDkvBuyql
AoZCN+w2lj75ljQjjttyc8cuocc4b6xO4jGljw15AUoKt5aVFBhP+0619GUuuy8C
dPJKqvXWxj2q85h4s/emFuqR2H8n5Z13zrq+P9TAV+4DbnEXUU4jbUNIAGF+7m2W
bufL7hOOOXgLtyFWCncmKluwp9lEmjazYaJ+xVckFI+/MtilQa5oaM/3bMGHo0Ma
cpziuua998ZDwKlWy7PhV9vLedtIv2AX8fEZuyzVAwK2M4V0+lEavkLVgfsb0nA+
WyCYp/4pPHmVc5F6l10fP+/QWcc5+7M5mDUzuh3GLv8fTJNRClQ4ZTK610TE9iS6
2WeCIZHWfy+QIuZt/U0pZtI8/SMlftCs/BIMWJ7LQ//meSaUX34wCz3zcxmyJcV4
9SJG6xcYmW4VRyVSfaMDgmeDmI29ebGKvBcH8oeONvYtrgTSyYvdFvVFu7sZ1axY
fbWFh36dj6cKDFWz1iKjUWqdiWzN1V75OwcttSE3laVGd6QW4YVVBz2GpsSHcP2s
UxHJ7ebUtyIT3Si4Zqg5UbXRxh5/SzTp2gqpqKyuiGHOwFoeuJG+vtDXW29QepXb
WIqSKdEj7zvRjbznc/6palcLoMpJh2zSSBshnTmtawr7he09jjdZIVt6LEyyTDID
9d2IKASG04/jDCSwtJvNAZTcVozRYyR+mFGek/GfUTOrYrV7XAMTGLrQQPjwuH6n
brwly6SYAO8yU/RNMoWLdsTNJSqRUkEo29qohygBERPYlWghn4Kms+bUfm1E4p7W
KGj0mOr5BazB9Ld37ELOYve0gqQ29mj8abux2FyS5F5couexxDZg+/7lX0CaDEeh
FrSGC2yZ/HUxadkjehQ7hK4YIYzul8eZ0VeNizdZzHFfPsE5r6W7hpCExxq+klye
AE8PgglA/sVQOzUYGeKOkL5ZEefUDwGeOKMxwVEoR01Bw92kIdowO17FpXBfFLy4
IpCtkx2duRBvKqaTBi+4gHE+hZkNn8NdfxZD84BbTFEqPD6okEDYthwsawhafmvG
bVBinsvUtJ6pq/Vi8AMvu/75GzpDq8hOnyMKv0gL2+YO4xlAVqtItTKM9wNA3wC+
qWkA3DdheZvd6kwT7F9q3ZoSlBf0mo6mBBB1wGaCiHM7GrDTfJMJ6eYJBxPmdbcX
Cqr9hWocJdhOX8PZUhOgeIcj2G9Y/a0CBj6w+bjaZVMT6L3aeBxYKPg6eucxuryy
0DKLEHMSw99xQ+jjMwXwdCfL2vg1wPAYyATvsg4xfVE2jffmwSy8IiGjT3lZvxZo
Kcn+rcopmz9sMKL9XvhU2pLwbeMdH+BXayydUd7gUkMJcyxB+ZEfd9xqAnI88AQq
sWisd693M6KDLuea+VhgmNCU8M6O0A0x896zAG7h5Dn6sxlYSYSePWv08mG0gLHA
Xtj38q6Sqd8yzsGnClt7USIO1Kwq0etIMHey6pX6earhM/F4tSWBzR/G50+eZXK3
O89o68sE0Gq29vcvEsVW/nOiDayy+VU1IUA+IdZh0D3LLCNOWh8QOIWUAs+7SX4+
0RproxzlHb/xV/IyVsqYnuyNjQ7B0/cr9nWKjL6Ob0brvPlB8GGgU87TiC4r8QlL
uJDYJw3VMA2F4z4FDmXa/a5+vuT33ECLdC0X/Zv+WC3Bo+la1OfAF44YpeIPxZIj
BPx0DAmiAtDwy+X6/IOK4V9HsnIrovE4HvhaDzgiU3Io8DX16nc6ggP8AsGILAlY
go+e6ycLTOOuwkwjNleR5xNU1ZkThIRY288CxWgBvyr+k72PH/xiY8J0TItjoLU+
p/7pDJDnvIelwANQAVJc2aOC1bIkYy3ebgLc0SKAHX+d9SMwi2GLbhWX6sKcoYe1
YDGWpLJ58dXnakTXZvL+E52D5QlxC+sBPrYJYg+m9TPf6A/LqgQZOEh1FKXINq6D
fmD2yE9H5wqx2Fbviu+3BA2ES1ZT1gedusHjhHTKLTsSBFxNPWSanG+JGNClIVdJ
3XbutVP7/DyfNmtuotv+DQCn3zoFSDMoJxmY4m4GWc7fQKyIScbGxXYucnS/7rjC
QT5YuPrZvUjXXLiCQf9ip9fTi55Ukyu6UzEf5ixLe2QjNSUCBA8T9tiyxUScyh4Q
dd77YqUyeOMIpzfHneymS1uFhZXoeyKWoKdwsMTKnEL+I91k2WzYnFEuEg0PPfcX
19Af7s3BxqCOOj2jQ9N8RhZggiE3rQn9eRIJXTZ3QhjOvOc0qVvBa45g5N6W6bNl
nsHRu/fskRjmpWOmSfPtitWQl/CBjqS5kJZDmJXBqzmjBvK8UzeGLgcJ5Ja6Bese
28Hl/quNeKQbzabIzwTPMisGpZ5/dvQOCEo7LBjt6oQiv56KzMGP5SfDcTqajoJh
KMh19NzGNcfmdfnT5Ufk+QayQTBzvLdrWCcw/6ScTtEaDnfQYsgc+KlBzno4+0CA
u5Joaa2Rta1DB/nJizu6qayOV2+EFYM6wHWY7PgErb49vxRGiObevhtqEE9UbG/y
ymUiat2VsPzW9rZho/GgeV8T/Kb6h8pMOq8SNh1h3KgzVX8KU+MyAlPKuJmswdtk
UN7GZAA4CUNVpYF52zFe3iQeswNWYmtQSEc6FPoDRUEA9F0+wf3FMrqdExnsoXca
xUYaRVVvaOAZdBCGbZD8LmTuUmN0zp14WY7HRCy+9icwUtKu8+2O04Zg8oJVPT4A
ptaa6LB87YEj6RmYWlwPmWNeuhVTJizMlwclbDt2e4GG6WhnDWzqDrp/O6cIS5zC
De6I2DNSLvA6E7UWDxGWVzDBt74nM1MzWIHtBLp7642mMOw9H+BcPp3aO1765gsc
8isXn7vN9AVvIGXXByO0wUHaMQl+DY6NehPk9ys3wUvSbF/4kr0TVw4SJnp0IqoP
ZDipiUdojzILmdMZtLc7qgI7SIoLjOXNnDZyQRjRN7oq+Sxue39NzqGLTqkfAls/
VL1oUhVotMssiw0AFmORzGf7vkztxrP+F9E7InvJs4mwg5e8D0F/XyZRACCEPkni
+nSBbI41ndYVSzELp9ZjvlE1Fw1z68c5tL+xtTVckLmPrRY1cUJGdqCnDRuZkpEG
OAZuGRFEV5oFPaO6Z/XaWTB6VBYazQZHhGbObeonEvnKj0udYNXGWi/y9dawwdC6
89NaxXnXzXJylSScpwPOuEbRjLkFvDh07LonIkvJzCO6tUSZjiO/vSQRRFKVjn/h
mSgM4T5kHZkk7puST4HnllEp/NdKgjdvKE8iEfQqTyHNURH0BF/gXkPeQoiI+yyD
PBtYNrIwOlr+v7zVjmDV7dC+M335MRp+WTNZyM8S0QN7MTi6qRnF808L1Bd9kGtu
3qZnXsmePfW5GFKnA5lhgQ8Q5l0L6hHl6gs//e6bvuqYQe2LUt7BKidYkdxRJ1rr
WBx492Yu3GzSJqQeVUtJBZUVN+XxCWzCX7Dll155fo/0TYPTcgNN+RD2UMKznMkj
zcEg76buhoih7HVz3R30nOqT/5wyFrEJ9xV6LuvNGGP6xldNQIljJ3oFgUZeSpwW
KxKox5o9AXyTpC6awZm5leaGZbVCK6xR9VwpPnw3KPxxXBzTx7HLhvz3u+svHaRA
5jPIDPVqn5R1EcNM92yPIraZRJlujeOfPrX6rNKX84Wyrmu+gGHtLCX43cEV+qJy
nE5cagvDUVmVQcQehbCBIaS3OFF2vyOwPMD9Us9CWqCmCXgqN2uR69IHoWMr8VKR
rkeKceFpOxIBE3w3NJ0VXPzYy1mNtN3Oe3N+zHCJ/c4t2ObfOnFbKYlKWrrkxi0R
S39ZLR+hmSVLopeoTHyDQI4C4QTRG3l2QRmXgty0Zj6dSsXyGnq4b5Luugv3AEU5
GF6rBzBzMSFJrLiwOjIrhRphtuLtkDP6aGcwR4PzF17vO90mu18858Sc1oswNFyD
ubWm68IovDtonyoVxXcuv4fVXucwM3OEGPPYoE+Pb7JHdutQAsgcmlplcGBrUbzt
Mcg+VKErEKhLPLUcjqHAH1oLV1kmWbnFEXiJWjiFPLvyG02/bJo6SxbiBkaaqxYH
l7voOUCBJyo4qbMWHC3gjza3vzdoSigwmlGmAthe65PdoLq8ub7fipTNdEXjFYml
wr6XZBksIRJmHF0qNgfVMBS5PAv42ME5BfgE75yRIuFHhWmPJXHFngqbSyv/zN8f
R2QelFNYAWcVa2rPB762Dz55qdXdfU9jeQFXfXXZRORJrJiYd/UcxdVfB8b11JVq
CAxKuBUmFCS/KVW2IZbN4pIK0tgzR/Kgj6ssJ2BIazAVPxqTeNQ+K1P7g3k50xoQ
I7PNC6dtmYA4KQx19C9IkbTwCJ5zeiAOaHklT7dxYdUZIH3sDCXv87SWKanHT6E4
p71qtL/dFMr2bgSuuYTw/QKJsrGeJIjKSwfhPe4TFp7/9xeNao241uOYkb6eOlM6
feV4BNY07Wl4En3b7xptacQBMD+8K3HJQ4eLOFtmwkghi2tb7YNfPDLVpC6t1Bdj
VZBYcOCTP/vIwTqQunClHWfiBVkqJggzLm3Q0kn99lz4XmfINwGU+dxPfZujeOOf
pPKxVA4mLQ9NyCHar00QN5KbXTTQcJ9yQexqR587okH5lU3JbsPi1pKSo8sZ26Zo
ym/NJLwPzJUETDRMJGUfaE3+D2JXkYsMdiBEArQrrGuyhfWT3FDHiWAkqUE8AQsR
jqEDOI+iQ7HoapVbGObhU+ylJkZ9iwDV5F/fJlA1DJiwnB5qBgP4IAn1JnHUmzq5
21bZASIUb79lBQlqsWwz+RPjkGo73O7tEVQQnOAlH6PdUsLSNM9Y83KAtORuS3kx
jBm3zXhxSnwFLcexcBL0bjCzVfg4O/cM68qYKAZx+cIYPws0v3NPwjQ+IKCI4Fon
I86wMSGsb0agthCPGdCRpcmHPEOoiAiDcbtY2RlcFs1Ba1q+jFhlPEzPi27jsAho
P85sfRt5b6zCvTjeJ/beM/ePoyYWcshmvu4q79f02SKTqyYVKgP/nOzYSdxQtQxI
LCuR1pCRA5CzCoADNrx/2UzZWJ4KST6iTzNBvvDeboVZze9SNZWlYlMMpA8OL3qy
QcG0/DiaGwcqFlk8GzldR9yc0ZZbzBdJucVvYV+zVOalPgzM4kQQ4eEfpKjc9I9c
Pj/lYy1r8rYmO4KnZvccM5GvIB3ksGAGPYcGUx2uEFcxxr6tJ/zMr5uajsqbjIgM
bwI9f9+HIAKP3CIihIam46iGlvkMi3hAom6tbwHEr8cI0fIIkw3qdEDSiTWgz+LC
tcfMYbLg+ASlrG/Wg7qFYve5FfrnQpA+s2MPn91TPU24cIqWIjdwujH2B6ZHYFSo
0EJ/0bni3wR9XhvnQL5JHQZ1wEW+8WGKMRRd/YkeW47OyeY37TfzFI6sdeZ8o51j
hG2v6rmlF0fvNXaMu0aLgmgWTlPKw0+cr6Ug8qDYE7HaZU0h5pGfJIzXUn00I2KB
X2QOKr19G0J3DXRQeYkM/39zxiePMk0nRrFOUh8zPBFlb+u3Zg/heAOVxY2JN/Eh
Dd/2a0dDyU/EFhEYHRCHoT/TQXPjiW0oj/Lfvv4ttXYPzFE39jsZzEgGouyNDSfC
cjZv0esSN84Fv1cEfX2RM7T1gwDkzcWs9nsgIOv1ONdrDidx1YksAv94vZaiKeId
0mySPwZ7Rk6FHWaAOrkSEdUrd4Jfq/FMlXqEYKrYLqN9aUIQmqnTx9gGohqzZPNb
qa72+ajasBoc7Z0Dk/tzD5osf7ci+R/3du1KmEWnQaJFG2OVuXoxrXm+rlUuoYm6
aEm/gFUANAmHAH4fYQWSbnJ8ipk3L1dDH6MyKEQPPjRnGnkiMQzCrzZiMRXvI2Py
BYleOVFZaHD1PWO00xzHIQe6j6Bjj6a4JGl1AZWIxNvGe1RVei/kSw22XrCiRAyd
hc0o2ACHTwj8vmPZT8oEg1PHilYyZuE8bqgk8wrFMXmkYWADTeSei9cZAZycmNGd
rit62ofsB9J0V2SU1rroWbP91Kr8tDr5w6roOR+9ncTojWOnCuxoR4+EfEmVierj
jAc9TsR7uF3im2l/731h/QVr6hMihT/Y0+dSVQgfmc+qXXkCNPXpjU0YgI+QS7Fv
1QcDi28sU4vCiFj57x6UxTw7S411QTGq9iVuMZArx+ryzqM8FigFSH+A/pJHxY/E
pLluniRDrYwEIR7xgwAiyszb7EifR7Qozvl6P4fgTBB2kc0M3eA7x0Vk7MRj+SBn
kZwrn0J3uVqX7mxzgu/dtz/BTDD3Cjbgus2ItHUWzXD370Mff5s7UvxIUuHjvVUa
XoxMEG9XxfYhBcBhZPLX/58dg9ZT2x6OxLj4TA25W3HYPIW0TZEY+BI0L4xzF66c
1H1rjeH9Hv+g/yEgIO0zeqKqIvSiW0V/sMz4WmO7q8FKrkhODXoslt1U8sttiAhV
FrFXlXWQjhlDr2iwu7yjzC/0ZPQW3I1sZpGPPdIyJspcAAU/7H8a/cXfTM8Kd0KQ
uYLRS6rtkb9VLD6xlom0qVVphYZNUjx0QzvXqdPNoD7WbnGwMQ3Gm9df+srGheod
3atLvywuZ8OdjvjPmqk2iiNKMBXxNfCAUM/kcT3vl5tGS7lgxNK95LK+cCBMs9Jd
0/WRmgTI5rMxIOC8YT4xwXVXrTKEnjb/FRSk91lvWrJrbneaqHlWKDs6PKab1ztj
hgZggw6xlJisGjWynjIYQYBb2sHx9rp2Scv6DhfwQHeHv+OyxjWTTqYb83htmMln
6yvPiK2pL7UbgdTOLEIkoDCXGluylFx5zFAiYUNSmTycioU01XYljGJgeSjB/tVH
FwAPqbnsG9evAsAvBQuuKIBbe1qXlAkIFqh9GhSCBUZpHV7Jrzw15TDZgdwL1Dfh
+TIIpuNgdeau1tUXbFNJb4jnBZlf/oNfXxOBgK0VWYk+SHJpXc1ygQmPGlE0yB+N
L8TG/3yOCzm7X+pIiwKF2SC0qIY/3J5YJfpioxdLuXDkDX8O2I6KB4HccAGBLKRA
24cPbzdHBVKeQVr86CAJsb4J+0zO94ZSCs2FZXcfO3jZezekNJxCBx8pEDY/5xjW
XTothryj6xF4hjODVsVpMESTdWpZPyzplIy+VvA1k3yviNRYNsLwUbxREKdtCkIU
uABM1nCko/NpAJWN10Q207bSM3qy2sKyErplqh69mSeuZ3VMrfhjopBDQwLFbogJ
0Uwk60jLIdTzFVnwYd5UThyFRafL986fESzIgKgKzo9a2aepCmaz2m1A05vw6gFO
P3EPXHGRYfwckolUbsDQs5fy2iRIQZ9cJOAJZAvp4MaRSxv2EGYmOeGRERTavlVG
Jq5IGxmfY+/CkYRRCiHUprjt88v1cyRgArGoqdCRtscl1XMF/oVK30fgFSdyGC6Z
q5jXoZ5iNM+XLPSVRIrHqS3kXlQekkkiHh75aGu/klen/D52svG9i311MW4wbyvw
dEs36BEyukrhTCHrhO9OePkbx3tJ7is7s0uXllHwVse5bR7BJ9bzY1BXmbBZxXog
IQ//ZykSt2f/toF0nI6mi7kdeePISUSUi2t0/d6zivFmjLHMo5IUvJwwYUMsnZub
S/aAltGWyLF3BNVgRtPrwSOUPQgvvtF4fso1C9MjtR2ig5rSXtzE2vo8gfNkPswR
i9lz/b02vt03ALf417cwokhsKLYB8Gp1SwWWCkigigHCwZIpkH3vOoWYhrEUv/F2
WzC/cfe8r06vs/NlvAYkqW7dPDoSHBlQElGbcGBxrlQRcZuH60J2Jw86+ZN5Vrvl
5CWBdusQ/ih71oqr2r+veJY9EuzyT/slrzRZvVlBN9JpYQSQ2rJ8x6f3xRcTxm/k
bvcev5eKZ6gZJbMOe5+NCsL3Dx75v269qRHuj+HOk/zlbUfUTQxdroogxtB/xkNB
qHOPBVomJxnPnbuxYzuV9phZY1HZkYPqH/HzwV0VyoPG5oHWh2w5MdUjLCa+kMbE
jA2svy5MQOGev+V5NUyw0Z4wile8E76y6ccDFqaHH/YLi0AGBGwtWobrGVYEOocK
bDLJgJg4F4+BvbNIkSSUmjJN2aNVbfW4iXSk2VwHxCMDmMHgnLmfBwShIAi4U4+Y
byVpeX4lvsZcLzZZbF438QUINqOyqmBl03XGOTccv4+zul7Ni6YpaZvNxzwA0TXp
grGA9xtWBzPrf4nBj469H9mw1kiBYle7CALfiCjJmM2MDv+BOgWmg0kv1Sto3Yxf
mELKqKB7Ee523HVGXJbYLJu8VjrLILVe8RxF1NYZkMGkJ5+09O8+VcUBR3spe3Qn
Y8l6KwMgu4qV5Ke+6RuOA6zmNKf8qSCfsAiVwZ7fo2OFAYk9Qdp2pN0wo3xsOrvE
aRSfxpmFEMdjygYE3LMmLt5OcpvaWiCMwNHFLz5T7/1lFBPqH481sEHVFOFMPMXz
FVU6Btvt5jrNffYTdU3vkrH6zUGBJTvtYtg1AhTSkhTqhmPa2fje343nYXIIWXFv
o+vHYTF7XoS4gaNxwSxF4XMxz1DHgrzsUVwHSRriocGCzLserW/LJ1urnfnL8QZs
kN68lF8tbDT0Pk9Yz7HXzkLGrrh34fD20OPVl31MrauVOkIrpXkv9hVHL7v/nS7+
gmwAVdp7YhFU5XWbpI3JEwfmcmrL0VEhiqAcPwVdUvcRD1CiDDbJhyZOzqQGoQ8M
IbTtx74TDrFO2JcMQcJJrEDfhoqTxP5MS6271032dJNK+6RW8EawcmphidDjHv8j
EtIEYlUMSfwcS2Wit1Wr3/+6Y5hRNlfxcNIWmEXtPrTM2Q3CLyVYtQm8hYZf4FFV
zdVnExVXAALB7EkYiHBityppeBOWk/ElQ+ALizwivlStN5GP9vXr/PSz9U+hvXSL
CqU8Nc/Ka46HTg5TeGjQfZirAqNy5SKdoDhuGaYWxeTcM/18MWEarwDGKhSIFiTE
wUUmhGY11wu6C/q1IGTQaU4wOOo3TTp54v9gQ/n+EhuXFfXllJdebA+AZeyk8GM4
zW2E8R+zhCWRdEALtmlkf+AmPtVBmdZ/wRtKsNZkjgFn/M+tyj0D6QsRmlvpYM/5
ZZ3g7K0KR4/AjgE8OBXRVwk7UsprZL/4QaRyXokJEo9PZvZJx5XZZQdEejJ6KURf
AF81jryTM4++HUyzWnY8CzsgYfiEI0xdvip2zrb1mao32SCqPKLAssYIybq21LDE
pDqaCto5gPYmliMKSCQ/6lsXTgroiEizu5SuWGkNWs1j3zIVCwsEjmdBwrutCPsd
EFpPg+/mwsXA9dP/rhDlGBuwJhxfeHRLeInKkAo+IPg+OpywZer8lEZ1e+TKhTma
SN69irJEd0SKxERPNDA3+7D4K+4hVOEzRDF02g1mBrYGo3luLaHZ9FSQusocHbU5
LScBwaVKB90i8oQEkPntTDPcKNLfz/DZk1UIQ5EDvrQnbgsrXGVMPSGgsV5vTi23
8ZCc+AVZe0jsfiWPMSYiM3Ct4Mbe9fVmzOrFRva+7rf+h23cDcJLiCqjjCZeYX5F
J1PgBqxSpnCFz+H2+Cizkifw+d32VEicwWwaXo2E2epkPygTpQi2c6qkT/d1tQ3P
AcU0k6dWbM2aBue7vTOkLgoJuxzbFAZsyyfxiJS8h1wxRzX8AIxzFCsj/h6/fSz6
2CFitwFZqJNsNsxA/J05VGPSevjKB5PmbMpYRBptCTfeLleLCIw4Uj2e06ECGqae
bk5SZYMLZot0sC1Jra77vbX5ppacSBUx3nFef9YlGjCFQrb0iGUObq6ogHASbdNt
2C/b0jxgSj6WrPU1vcMeoJIg4wZ6ziSlL7T12Qoc7m8jNv+B8uUGZDcdz0FkTxHm
Hv511ul7DMVZGf1WbYytN+f3fMJg6D94vTjkDwWRDliuyQ+N0SB1XYbzX8LsZmnb
uZWopkSmOrYVoXoBo+7ATXzdhcAgUwLx5vLWh/Y0sIl6pz4z3ujVxmT1eNi8tV4w
qjtqHSwWn3aPJXgMufbCd8xmE3U1KZ51KGsSnkaai4t6tCI+RpSCpSJ7eAcgQYo6
Uw9obbehLTPwNZO4cMp8lGJ79WHvaqob6iojOFXSAPs8bgirtEYSTTp+5ki37PVM
oOWq1o23u+kGwFOAMYbNwZqK7kuEbce8LztlfOwoAdCDewAZuurIcJCMccCYVF6x
nvUtl+ZdmTGAoDXPTKAC0emUZ96TGWk4WnSZnAe5tywj1I6Owd7Jztfdf0N/7xcj
rly1gS9ryVp+QefrfFjkAIXWnMGThI7wKqrQhQnGi8sPI86p/rt3vdIsjGfJxaMy
69c5qTcK5OKGyttDhBX0SN/o7fRS0GEAwAZuUaUPqFfYLVAD1d1PKv76NHgBYGMh
wlH1yrKaR2/Tu/YfTSnszhCu2wBn7Whvr2BF/nu5Zc74dNguVyHIGlIuAWN7aR1y
J+tSHmNqvobiGcYAZ4M6Aem4361lJz5uJ01UA6co7HU34aP3sicDZbnexR+PrIwi
dM81tSd1sKiBqfgB5kkblb/TgUlWz2WJZYaD5Z6xVW6cFHlPvN3o28Mmn1b3557B
a943lLfDIayAftftsTjBWSkwk5rvH5J2ySRJWcP3C/NIBOCZ2c8Uc4ImvQtR3Vw5
3ZytHsVh3JJr4vTBiaRK+zUkhrw/MExg+h6Zs6CP4T11/hqokCijnpLo6xTSQtwk
6RXXvnmuMuUc+gkK44sU9igtTegOzY7R2+StvHnoTzs9oVEk/EFUp5c//BmMFrIQ
cjz7LjoYQjkIFIGjQdEN2tF53cAJzD+5hkrNvXHTySCeKrtpO+6ypwBv0tidHn+z
6Z7RPSsl1nhj8pOO0cT44H2KJKPdB5hEICMS446lQj0FOyXnMQESsGsRUpjDF9+m
pm32mk+qqrPLT0qREHNT0nSQ9eaSZv/rOKOpsaoW/pp5SwImlj1Esnb5zf5KWv4+
hIMOgyBExdWx/8VmyXMG8eGNPcxz6Zg8NaFUHwfsOM0nsHYSxkbazdwmCKhV7pe/
yPadoUR883uu+KYgvlK//4bFoouWlxiNgKdnby6ijl9afn1zecPvzqpwPJWxIMPx
bir+I8D1KyHK2dak5agqctUetFcBYQL09AwVF+PPUIvbDFKDqfnwfuFq3PMTHnMb
RGaGlnyy5pJ4es2rNUwgJnyw17gqyJ/mzi6kNwjhnGkyLPVSHkM52bl7NXf/BfX7
ZTirz9hlDt4E/0bkNsHBvnCNApeX1jCqF95Qf05QbhW/sl/5pMNtGPgNB/nW5VSL
oX7d15Xy84dgrj6dkujnFS6Sl7t+NCPbXjrEvS8vj5zm6JB3D2ntDR2vV3oXkd4y
fVquSAHgpu6r68UOrrMgRATT1/fPp1eGPjJiA1AC+t2VgjkCfPsQpZjsia8d1Tuc
ebtRH0v8RMDgeI+AyzjBSWRuuXQll6oe7JWW1GBSaFNI8RLJIpkbUttALZxBje3O
9F0kQFkiywDBkUNR7YbEIZiJjncw5x2AjN5MHrLiVKYvcUqWyPaulMr3OBRmh8s0
CdMr7dTF8q4yY3xH24gZxcbubpKRUrfjA59FaVXTt7rLTBUbpz4wbvSJMpXjXoaw
kXmfqoKTaf7fKpwmkCJ0hu7PpdmK/J8VYLx1Gsy6qrcb7SzdI+TYnG5DClPG6OQY
x5FwsJQ0GeoInQ6BSODxPOVfypax9bOsr4PF5voZ9lH5tug9XHb3Nr8exKQM6+d7
RI4nfT0cvrjXK2J2D8GvwPyHsHPpdfXLWA1BFpiihDaqZV4nMydYZ2bDOMARo/NF
7keegDUZ6joc88GYSew2IahZfGEjyzTLpfzVI82eE6Nkmb+YxzB61xbhasehs9rg
rkJlIw6mojqT/dqGYVp6YSAgIghE/rRvVPPcZ6NF9eDrcQ5gAkonV8FIKgUBfeWq
obF798b2yb3te+Fb3lFsqWv4lgM/3qRaIy0IyTc7m+sMRNOy+83WUWJI0vm7hcMf
9R+S5Ql1R+bLCxdTE9dwdk1rT1cF5rlAEtDUYjd/LRqE4Pwc6xmCrSmRmwRasRUJ
0An3GIar5PHAqcqS2BTHD8qCBLBX+vaSPS4+OKxjoE3qsWmOeUyCjffmzRSqf+lu
oDp7ftNzLRmGfhnencIlZ+JdqtIhlS6XMOM3xJwy6OfzNUIM11Gwf+gN9GFZKgPa
I/C+SlS/pBWQHwRyZBmuDqBYx8EdbkXEc7B7y9w3gQTf+fDrWZhtsdQqn+Fwv8AP
LNSYqFf827knAj4MRVYPwTdhuUJ3j4nFtBd7KDIVcASZdVa6ckenfQDR79Iiuylp
Z6VZyW4s1cw3vZbOFbqgrPbjAEN+GFlnf9WyUMsiKKXwQhiulp9sk1RWOfDLQGT4
05Ur7+fR4nBwc1UZKHpzlq/6zQVT5PnJZRTyTawqgSLC2SeTfrB6DdwR2TBz/Ze8
d+1eqgJM0xFpi2dbN7VC8qTZ+f1EeaH7GYGlvsht9+XiKyzK7bDVtjebFFIFTE4f
LyynVYAKkCA+L+TX6/ZMS3vbBejsT1NPlAtspOTfUw77hCLgwjjeiZRbF7U9n32j
Q/TdS3zHF+OtaXC65NfxiI2GyCJIUmEqTJnmN+PclaJy8EhzsnCWhNcLHShD6asz
9Q0joopIRn6sSRjG37vo/KPVNYWZ03+viRy1pyvxWZquKc3a9+dDGol+a7TRJmib
T0reHinGIiZ13lEuIUCQlioGJdFzmjgOhyZjyZFa4SijAh2jYVOAXa6iscAaP7ij
3ZG8bgIH1uLeRLfBy+d9zD27T+WBkoFow292VtBsSdcypNWLsPOhJn2QphpGFgzg
vGHdtFGmrKffX5qBScchgm4OLoi50yl7QEK91/1Kh+ws7k98l5vOiFLUHmJhDaC1
X0s9XCexer7cocyytlmKFZZmC1j6YbGmXLjLw3BdU4xfXMsuEjKIZRkKvgW4G5dk
eKy9DJ5aAKyx/g5EIxqroKciJry8ct2UUT69GRtjBMjc5sMPuKci9LBllb+9xS36
oXBy867JeRKchNJ8B86u2S22ref8sMOXl7uhIWRfHVKE+J67NF40Y01G3K0RPMYf
lDZi01fOgAGU/wvU4FO/HCXTmDnmMJx22zZ4s+f3YsVg3L7cuzopATqPJs5TNhYp
uTVyNVZKKOMkLlUS8KZmty5v9bgi/Hm2D8Gy8NrZBGrDYknHpZycKYn3AUrCjrI6
VBz3xKtNPLkzvo/ypGcdXDLcuKm5etMMoOX9nVu3tH6B2yCu9oLiMH5fsF3FdPfv
O+xegvLa4uZDyvSPGZKnt/6DkE8hPXZCliK0ZMFvXYy9mCzJHeJ535VGB75qmQM+
WqIsqks/zzQ3yDYGkUVMBHvrXP4OgMHFYV4HzA6wq/DJzrg/LQBwNknhf2y8p1au
3Z98Ge/dnBDYK09RDyur39zFqZNJmNzEwXSfc94+NWNmhzh8N8KInqgo15dYxWc3
bVX7ewCpY7lv+d1s6/wSEOXMlFhLP/jRQGLnMB5bwh7yrLfKBW+MFUemxiqyi4BG
AtSjxyDS3knpc5YFmZlXrwDi8nEXEGB38jsyHQF38wpfeXm22T5fRRq5gCyKqfU0
AYuQbYZnAFV4xT69FLPE5dpfxsqt1zbBNoaauUjQgbBJ1Qs9T1ohNC3POe4dOOu3
GcyvLZxqEQSoPwOUDMu2r6TIH9Xnu7kfQWrwgEN68tTMTemIyv2fZP8Y/qIsobJh
D9xZEWZ+XPcx7w+FcQuzbFURENli4sKcDxtQKWDM03R+o0potydbhLmfEGKuG/fI
h1pxx+BWpuZg0ZBmikxXPWFaZY7AJ01RjMKUyMO/PL0fRMa+GI2cdgcKsefYVIqg
1Iz4Hf4aIvDT4o6VvpGBAIlY6rD6amEguTT+cKozgOfBDp9gbidIj/lBoLDp31mc
DGHQ7sqCxHaWQMhWw9Qxto7HFrxt+GVWAP7T5rIYWJ4ICHIVrjMswtcs7EadKtGJ
dD2J2KblfhWe4aYpn+xIpKPLH4b9P4Mx5TifPLQTV48DpfPOozTH0HW/suYV99on
GSvA4sWe5OmlxCAX6htrcJ2zX9QX8gleFeWsur6sVMPNX74XllIj0skk1siDVaTn
n8hjow66I8V9FsV8Yhk2o2DRWmo1EtRl0vx95LCihGKey4IkWsXmktT065i3n4DR
TfrkEEQSLNv/C5TDt1VIMnIY5pPUItUHy9BfBwpmF7LuZBK/4d29vsiEzO/zb61I
no3tpuTT9ng3E5wmp7RBtOkb1ecv70sFMqxPgiA4V8ecMd4UCFkVf8GZVCwu6y8c
NzS1f5rJ2ibb3zT9L+ZIS1TGmmkZLU9JbMc8iJgOSHjdtMBZNsiHIGhO9sm7AmEW
8GI4p8N/zyKkjoBJLJHBXC0WEui6WEtz6int/Z8XM84SPwNtK3tq3g4pMaw/AATo
ezj3qYFkAA1ksId18kkanDyKSe6BtTniICws7ix1dleiM9wRfnvtqh+osO89YbCr
FCY3zcKPjJ6Q3V/yAquIj9P5x64Mm9tZIC6d6m9MxGnbXCEh4rvcxtQQkbguWEcu
/44op8Wop2O1oYQyUxzvVp587HQrqtpmkvHIqj9PIZBWpFasyxKAGX8LsqZ8mDQV
d4C7VirXS0+rg2PAqSwbJOhaUNqVkNm7fkGDyek2o+MXQ0r3NTcQdHl7Ncs+zZpn
dZ6syHMprIIixdSRIYFZry/XuNNK+ElHq321yF6Go7XJWbvrr1+eP0cAw54seHAW
RVZzG02/PL6avbFVxAcgUBBsNhvE5QJBJHBpsmzeRgUHwgqE5kQ7UcBHH0LSstth
LlJtxdfqcGEk0MGxmvED4vgEdZ7gBnwN3VWsaZGI6FnAYE9hivGp5TcM1I843yFM
LXNX3Mlxr5Gd1GYtqOEhTn9esUxueU4Ooydt4wZzM7ayqFtKEXAM54eZqy52xq/6
iXI/M8ZAwWmmMVy+fizes1MzJXYG3DVnvjfYyeU8axDWcJzmLh/gg06Ktsv0l4Xx
8aVroVGh2GYYcvq5rl7S1hZbtpxKs/ZtO/szaXGKQy5IVC+ar6P7GSBB0ZlCgPEy
LvoWZsMuscnQwpASD6WXyn9wZJ1GpBkfLYiR1DLAvm7Pu0GpWqxcJm4YiTO/QhG/
dOQ2b0ddOmvVSU8aWp+a+7sIVF3Stbl/DPjD77ClF+6uoVYoW568TvyHTICNSsvT
BefbH7CZubj6NSxSaEl2WteNTmINQn3tGG/dnSzm/GFUjAknlLTPof1InzccfUB9
CQakg7Um1qbsGPCmyDHUOkOGTmPN2qR3JCuHV8dqJ8gxZNKa4TqGApj0cyLy+1Ff
nOCE11gz1lxaSp1np6DSL89+Bvvsg/y9MGGXZ/SjMqLP6My7kOJ+qaqaCI6I4Lz1
R/ldYm4VyRRMl2/xZS+X75r1wasYlKKeNpqbbLPFwLo46Syv21gWLIqr/nSJcoo8
2Pj06AjcA60li9IlveLxgYD2kH3gnBOqhKTUltwvcdza1heqPFXuOvm7v/yU1zrx
Tvnv6XwaCR/UrOahNgh1o2wZY/CK24XeFFNKqqpMX49pvM0fxg2HjKHCIDnfV3t2
DUJ0BaQ8QfrISjNhhTtu7J2tMIGITWbCL/Qj2oHFuMg1+c5mbiLv3fIzSMkjJdi9
rMMB7ojUeS0v1kKyqZd1lQl9KlQBEQtl2kTtJia7rfOGFHEOZZf8cmD6yba+3+oq
GUukOIBsfFY4KLQWRCjJodIzzsUrb2dqYxQnIv+NyVPakjFYnqaYtsuB/Gz/fxiq
NcjWbJA7LK6Ygh58125UscfmV4cIEJ60eILeZ8hyVuMe/dzX3K5sOGucejsMmUS9
2HYPUIMXLoEF5vZmDjE/LROQ2MVzjq1bqG/KNQivGntl28C9dJ2POnmUjK4ykDIW
9dxs9v8uV9CH8NpK5/qAFP8fSNaCkyZswjRNn4RSXeD47nIFb7hjTgVK0cKSvcWS
VY87bYme3rUJ4kT1a5Zf3dADwAvDInGcqBOlnGQ0myvhGfIHRgVZvoZ4qnhoEBpf
GM7HyEOh7/0prtMQo4sIWs4Do6nAmRLZLZKwZBWGMkYgVceRK342oicQup3d2qHU
vHsx6/EuA6UZO9246uEnw/hL0Tg4VtvnCGUciaAcq+58vnghb4PwMNXlf3J+WiH2
QV4eTA6Z/A/UkuGrZrgkeMjHw1Qvst6wapF+IaLSvWFk4dDL21z0G/hmmtEImG2g
OEXsVTU/07o65053G3V5F3TyXkshSSOmgA47OlS2VZCTO3fJAEAl7ckM4u+Esu2C
xqInJe+zTWbpW5urJ9un7MS4cHGUsLrQf6Mx0ZVWBbKCs97JR3OfNXeik4E1JcCU
vAVUMKwwwvo6pP3bUMZFGBKzmtlqFZtF2RsFcGPkoInFfvqvpf8Jcm0CbGhQGva9
zHxwwIE+3Ku0NbUkTFVExzbNmvF18m70zRSaWljTcKF9JgpuPJvjm7Ycw+zEUMEH
t9RhiK0rAaLr2De17d2qsuYTw/d/esFIc0XGfBdUGMklLhyCUMPvkHQwQguOQ6ye
wu80PpVw+vFAqMD3AOcW36DEi1LwFLgQxzbGnBf0/ZT/h4+mAsDzpkjW+9NIBWM0
LbHz+cunm1dMsK6B2AOCXMZRpyXlJpf6hhMGrYTD7vmffqNFIBbthDZovlqIQ9du
oUmBLM8sQ4gSQ1WUtouXrf8qiiMgLmJf5/5hTB5Bu12pbv5+QSpBq/eQFbsPBXnI
z6rGo4S6cxk3g2qQ3UiYLaBbBZli8Acmolhd16wLVA7RMWnjdhZoQmpAVg0bgT/1
9sXKd4mZgO4p5o0qrzpTTTtijt9d8G3Xgs1R2eNycEGegIBRofgbxk2T7EHMyzG6
APqI4NOYS0m3TC9xG/boU/OEiXeyxUmCGQjaUohDZbDE3nAOEoYa3Nm7yXJqXEvZ
gGyfII5ISIbwGNCznMSqktM9ANtWWx0zV0EPU31Sd15B2rAA2crWJ4PpZG9lICUj
2NjNCFwbvwlLdcWhqgcj9Yu+FQWPM2K2V6gBVQouR6A9YKpVlsx9HBjY1U3Ts4QT
fOcBvlqTkd4+zMCun1XJMmTXi/fUZmlnD1j60jLH5jU9UyPeJOYIbD+9xsUf+4AR
lsr50WgWNciGnmELilZ9xyM6Ea7SU1JbCCR7KMUAoT9fFv45MbEdybwbKpXr1Lvf
HqFpW/FnNGsyzzKxnhDZM9z2kago3govVMOjC9eZNCk7LxHSRM6YJ1VWL9WS0n8m
TUnuW6FJpGNT5axFj6b4el4xgKWHobg/n2GyJxlHe6jEBhZvC29hQW8ZmT/2nvHG
3dw+vf2/IxTCcVjlYJ+FDXWffHjCrA03PWLfKMCD0ziPZk2BIYvReaLWX6rl7RdL
W16qugp9Km9Yl/9L37psyWoWfqDdKgXRmUuVsPVuk1PJyhltKUpSfovR+1mrlihw
U0ZtF8qZ+w5pOh6shb+ju4Hp5r3xeT1cqjJjukf+2mm24sjqmxh2ocbv+k+qWGSA
u+tpGBYo2U5xLOSzd596Beozkb0sIbufjq1MDDMVDvpxryVbpGpbYjC1m+RHDZ7L
DZSsLUDaQ/5kyaVxrd/p+ZpCq/ZLDpm78hcu/I9G+gjgQv79Wm1+J5PnVTn3/RWE
eTO5H7k/kGTFioyu2XPP/1EglMWU5sV+cEn3SU881oQawrzvvE5sy2CQqDEYL8ul
X1UmDJ7ikIuXVARHTbr+UzHr5zK8GggKUhAqbdTBRS22Rl9O/FZxG9meNpdAER37
NN4iwbk5iBCsx+SN5NQWlJnya9o8xitLrOPterPV5wJgsYudvMKn+IFRMf7igPxh
3X+DTed2dqRWS8Ac9Y1jCNAIfmRRl2H4eVXassRapFqhUPNbjrtxFogfO0trMR5L
1UuVRC1RBogLl85epMiWDXffmZECXOr4R+THqtzb3ZxVHvWEW6XZtJzg9qrH5uZU
5r3lT0BPZlJS1ozFoqUAXV3O7JWttlfS+rYorlj24YmLBUgoH7TEsErUdS67UVXR
REIGWOc1iIpm4vK7Hvva4IPq2f1zSMIYipgrCQ0T4WZoIygo9RKTpTElnqGcPOTt
+Wqzqra0kpNfODcxMPohLZzx8uJOL1+IMSp7lbYGqXZovWE5iuF6/N5AsrIVNbo6
fphxFfxP5CnWsu76xX8fGGOHVUm9Pvqm5/kRn8xW6Av87L8xN29SBMn1VBV56aZk
HGKSqySBnVRLPv+hBO8HnIHLrAbI70+Lf5QkjDic5jwx7c9J59xX4aLCcI/4ygBy
DmJxL+j1L1J6JhQ29hsWaMksJVF0xz8/cMN37YytoHAknQF2YTfnrDezKXS+cAcq
VrCB+/zMeCCgG7HC8+wUtLrCApWkkZiOguA1tKlYeq2h8CjA+lWg1frVtRy+RpZx
DWHpxIh+KvTXx8a3el/+R3dDsmbBQtPx+/venWVJlwIKF26bOYuARaJ0E/mp3k8j
ytuA9+ydnI8FHu+mjbu/XK7zqzDxbxHdMDd/GqUxzmtTm/iA8t4ZQqQcLGxRydUk
7qUaVnTBAOT3DxlJkpKRrjlqU2HHYBWV/omiaGTZCyhftJhLYcmp5eVlkL+gRGAI
OCIEbpir6qxceMgyYsLBJL/117jHGyIApgSwC3G8nLK1BWif+5cPX6DhAxfo9NCr
ZC/w3Qp3UwfzakpR8iUT/FwcpTCrD1yzaARccb6T6JMBf119zM7vkDjfPCiCEoOk
o4gIbdCzlgsyceHnFjxsQWyCDu+k6EPXzSRFR+7xzdz9zzdxcqyxhCz4HSjndQYX
Yqb42Bj/dGGqFvK/zTFTsD7LwTeHqt13b/f2kBAoAW+sE1SK0DQ/m/4/wlKhAfN7
9HHYEvVT/rAzyzuzq9j1DUzoaoqYcQG1W1snPt1Ix3O8+VaCP4Ywh74XhuW9k62C
19sZlOX/8WAO/ujWnRIL1ytjncHgHAR3szhzFJLYOrv/zaMKE7Olh6QD4jM/T48/
bSlb8IZQTke42uNdO8xNDZ68POrIFyDGyhhtLE2wD/mmM6YpYq5r3mLMv4SaZOBy
XtgrLHKEznwRqTfZS2MWWJJtCtPDG1+fBZqgJ1U8CDnegn1TgQRi84lasI6FI2/0
sO6a5dJET8RI1DtEOSYo2mzxlCg1BSBj+JAmGatxYwO+YgnO059fapAwm6ADYpgH
b4ShWk0dW36NDL8kl4zw+9MJBmeVDe8XW3pXI7KzwYOn/NRO/94ZEWukIJ8jzI3W
84l0YzpsVqpaue/yPpjy/VzeZbomIiGVN+FqOAo7Mqy7gZ7Gu/9UVVSOsvmOtSQg
WW2lGPrU+QsrdmoKRXRWHiDShVGQluYrt4uDRtJmVtZ0txtmk49d5gTF3JheUWQx
faeY/DwB4c7ked3NuZ2lJJU2UfyCoiGbhdbAqhNxVr5NhJF48Ci8m7tQ02EJ50Tm
yptg5vAOi3KsjJM2PBYptatr/6f2N4azy9oro1CaUPdkCALhAxLcPzsxynkf2nal
JMu0vuXOQQcrgvmWAHohROcrbieV21W8khNxsuWLfSyFK97TpAyh/VMd5fuonsif
3AnC792Lfobvdk19Q3c+wuTga+JGeiw13dcOFvmrUBgbc2AdTalG7oZPgnC20RzN
rSCv1TI322/0NzEkWvt982A+ZEnc6SMP+YwOpO24Pj9zkJS6K4BD8BSKtl7lQt0B
5PandTsYx+5Qadsjq0s7hh6HWQslXdnWZoAyr9Vl76AOuaQJoZiHbebaS+OQBwoi
dgBNjaIBquo463IvR+C988l1+R32pJXjZ+zM+AB4s8NV1t1mT7psEGi+HxMOTDow
itIQIWx0EFgp3C4KOruwPcvIR3RjVUDQhRCJM5EjsaScf+0SxydNx5IN2EaHp5wn
PVaHwQohbOFID61bYo0yKVAe8T55a/h/srFmX/JxlxlEuAjfL9l46kUEJXPmnBuS
3uA/Rx2+dm3S7WUOa9U/CAGTRpCJv1f/Z4pkoxvkTCRZz9Nf+krN/I5VY97B+WZ3
mrAoI3iYaDD1Mng+ft6OSodYBBFDwg4lQBdk3kCZDBoN13FebroaY3VelkKpImgv
qX2HOlHXPSqg3AlEAdfoNcddRvc3WKPbV+GPE8a5ZOnCekPnDyOwXyHFnDW23Usr
CoMlvpdXc/GS+VW62eiL98ChRSb6oJ9j1vI8EFUQaoR9EtbrA6VaG9/08sQJSWYx
NGg51W9JgCAmlh0WMCUj9hYZEpziWFG/Bp7eQ5fWJl6BwQtgPN3LS5G6k9PudKDW
BB5kFJKVWhCmdxPmmppsZ0G0FknpuB36gizF70/wrFHi3JQr+vQz5Mzothg0m/NS
BqRANBs7D+1HV7N+LMFMRlqWvv5uCZ2PYJ8n/wSM/KLGRedm9sLMi+Sioq7S9BZd
RHWbwYYzN6GvrF37Q/Rlp1AmtRyUN5rQ2kKx3HvvI6i3iSwkefBr8Ui7NqpI+Jwn
nXjdxsRUSLIrqpLbqtU5I4QuW73a6nSS6bb4ZkUJ8Q6yS0GXXdEU9ojYpPiYbWP1
oKcRDI8Am2YCdcA03g62D1f95JsQj0s4+FP7prjknYSHo3roMs6zAVA7G3bWrDD8
va2AX9mi5kvrrJZoOrRG2WvzrtYlaDp3g23x8nh6jipLTrHX8x9SqclpZgV+73wK
vDoS9P5dHi2FkxnSms3rTDzDDk6tBly3cJb6Mx0LMIaSTgoUcIglOFajRnZ80l0n
SuJUREJgz9zq10C7JlVW8dve+GsrGAKtG1kEg8Irtr5lX9QJ7/q22nCYNBvtdBpl
Totdar1HV9hKHi1LJUNGGE/57xcQflkrsHGvy6+lWld16XPdYm0PdbZ8seNC7rkd
1FJDE6QMMp6cQh6xBSj2qdavRSd6mkOM6jJExWzzjm+J8InzJJ5W3CR7XFxP0GaU
H3PBFNvf1tWssMcAqbDSefY8iENHhg7OpO7w6JxmXhrF5j2yjNMuW42Wkb/qsZy2
4oSeJ/BxwUaO3x2zIYv0sc7/kFDqdhAIrDBN9UrlzWuIkgB50Ynu9Fdd/dNHoIKV
kdT36Ig2nUDZFxooUH9PVuFqr27TJMdBZucNBdcY7uVh2Nn7mj9YbDH9cC1+AFox
aIx/Byn6DAJbjAemfxBtH7qc8iudMfDjDaTkhyFr2wv/c1IbH4vthDol1FLpwDAa
6REwCjQV+2ikrc2VoB3oKnFUVyv6LzhYxgWFmdPxf4lQFhfeEvMHOxfUwkKJfPaG
CArRU1IE+l3DUEXSPv5LnyllpG3wg/Qv2vyAb7KGP1+8rTrAaaQvYId3nHBFXd4o
h4text8XBNEhx5nNuWRjiCme1YhrQqYdSTvYO7vlKeoE6MFdwuEVkeYeukU17xwL
goheLwjia0RWVrYGeubhoyfCrc9Vc9yKPy+6MKlEEyZXJsGG38/ezgjyk47/qGI6
YE9X2SP2YsqE8yuwJBVrKkzW2OU/5n/97ny5unrIAz3d666sr7X2HWhrfTp8OoXq
zC006oga/SQQ4NEtQu2gYTQtYrKKtPdcquK5ZDcCPs4GNqZtIJG3Z+Rx5Pb/URMa
CEpDYqej+u/buNp76LF6GbeXReL3c6p1yEwn7iaBaznmMfbgAe4Z4am39KnHQj7g
P4nsM0+5TfIP9fqKXJnHv+65UN2eU5JXJvInPh79Ph8OT8KeJTim3MYsVG4IUBar
NBWdWHoG9Vy4AW+rWfIKCjhbVqCyPWk6LqX09iJxaGMKWOUWNbSoDJi5uBw+nduC
BVJnNawiKdfSm6ISh9VbKdOrnRJmGG1nl0XYh4YltZcEAkq6D8ETJfHXIcCAsmzG
VWx+oB5eHqP7GWRAoRrq0m0Bw/WZ5IjfX7fLpUIXg2es9Z/4Q303a6ZxWxp7+5qK
hvq4f1ejQVSCZjtn+BEpApaloRFcLxzzaEdOk6PllxPVvqICLXkFSqqAbgF/3x8N
WIbhociwW95Deh1NGck0RL1BfQEDeAiGbwyAT9nrdphcZIHkVydL6TEYr3Oby0js
wJXBruKm1vSbDIX/85jS13WGfrTcCqBysoOD9rNsc4Wyph0T+Jhx43fZNO9hRft7
wBetFRh43OQuJb7lIeJF95bKl0pw5muqeaV51lmM4hpao7OSScXryFS8UCydImVp
yoXcG8kqXwmbMUUg/zsMHGXlQHXAI2AMNran1kF4/5VsmkOvk4Y6hjOoJ23ZE6DJ
Ztnrnj8ZtQJB8ViwrdnHibmoJjiTiBVwMWLTV4YVPSUORRAU86IJOcr07Ihs1eux
TUCw99lEIPr/yUBz89lgWb+TgCV525C+x8jC00a8HMulaI5a1gNrxGvdjOB/qqAS
kdTTei/4xVDe41iJo5UPmWL4doa0ToJO12eMUnjOfhBam4xTuZO8lFgz6ebyyXI9
DmFsLS3NlFUZJruFinbt92Cy2Sup/WJ982xYDPb4Hxd6PuzIx6n0+dFFhzz/tDbR
KnTIA9XgVY7nAFwUkisDZ4DmCHiTLzMhaVNyiyLwPqf9DPh3kM3WzPhfHZfwh/11
9l7dZ929gtGTu5TFyyhNEXMnQL+a8qLF9hJYZwfo4bdhyzvquCfxgxX5CEqSTJ1K
mqhZHF5+MA6Kp1hKvfN+KD7VAVvZOmdNUXUtuN6sVGQaiJ+oyGAFgBYgPv54BnJW
4OOtkiKl2B6qXPVt1gnJl3+dA8fJeVNJE0ZW+exzpy/Cx/b3oiGktpIX1xEx6Ww2
xX+Cs9FI8dxsEsLG4rLIsHgcJlvrIfU8ByCjayvcSx8QinS6I4BjnfSKXiN5Dm0U
yUx0/iYfNSXVSqTMjVtXkkHxPbn5K/Gl9uPPpgpzvU8l2Sw8Td04fcvNuXFmYCqV
Yk0fMPvuxqYv7kqAFpvWtQERt6ryRlgXNYczaxuxqp5Qdrss+0YbdVWFpdRczt2y
geKjjAPisjnAoOS0vrfdAv/awtSZ1bekwdVlax0o3dZ55quhmaSBn2voIm9gJeD1
AOZdBtgBpRQbTamm2irY8A5tDnMgs1yqXdTyrn0TqD712aW9xRq8cF1iT8B2DOCN
KQYYvcvX/F6+SI5naMsgjT3imOK/i9RYQTmaZNLJavnYWexJ3opfaduguWMf+67O
9dvA5bQ/PCEIMIgzvTc5S5uHKeZ8CprGDYgt9nBbvFvMaKHQYTxM4b9PUPoGEoHm
5V1KMMyuV8WYhsX5upM8ddkbuSOyvLem9EpGaK2JYowSb/qcJ8+JA52RQR4h7So5
AbPBRoICtqa3LSoDLa73KW41ak2Qxpj/Y8dZSfszBRnE/mwj6sjAxgfqCu2m9gaM
xFxNrASFRL3aXOmhOyRrHtoDTS7bDnrjwsJhPx4A68CUy6i4PuY1/GUaTF5CQnTc
vtMD9Yko8Y5cx1kv4D9Pfb1jR6k29G6q+mvHFi/9aemtUa/u2utz8dmixu0GyS4q
7SoAWKmfamW1cxJzdRsHsw3/kByQp9DV0nZZraRhvut6fUF/ge/c/BFr1//xcWVm
WM/p4mcuAHM2HwajGFELbVmnW1a85N8vmTodxo/kfmxhloNwe8W1B/HtP6ogtM4H
ucyQ4hMPM5LrTWtxs3+SkuSvvC+v4zAhqimvVaU1rFp4SQxly6VjRacwHbTvFck4
nidCa/Fh/SV0KzGMmUoBlJjdVAgvgVOFfGVn28d7jmCJvEWY/Q5gJxniwXwgSJpT
dXFEq3EnaV5j5ILSo3jkzRY3xEUl6CfbTVyHtGTvvz2vZ3GwuIroxsoqUVxZmRsa
3K0jC3/LxFxCDdLq3t5ys+hfHqtF2BkS+DWaIanvrvwwRKsU1IAcc/KvfbL99rft
2S4YOpuOvDqsOT1Ib+8nolydCGbVdj2gy2RfIN/OsFFZWnGnRduneVDM3f6cR0fW
Smxk5LPulztN6qZWkIavsZpHvMCTBO1/6eTgmrTrArEdelIDc9F+dKogYRgP+ApY
KFmTUQZasUWLTZOjXz4NXodFX8jKV2YYou0ypAjLK7Bav9kHfBdZZ6Ajz4sc0Le0
CtBmFQiEJ34zkJ9VQGN6Ac2DrfYY+SO+iwTuHaGTAHStOz3/f2+o+XrVtYGgxRRn
kBk2BXzsz6FBVdU2PT015G1vuDzrkoeGIKNEUJEgwosU3ilAC0w7dLn3eo0x6lml
5JNktd+YqQN6UbrUq2z9t07StzuhqNOCV2h36sMz31571mhI846KXiulX1BzqNZk
qJMNtWsn/9iFiETTTsyi7J2x33O6Lw02UJfYNLX8g9V93odmITCmMC3llSJfBkl4
jHOt0lrhXKRjERg0aRBu3MrKtr9cBl+6MlppGxHtj/tti+5Sm/I19DtGHk1wiGGe
jdpd3ka7CIvNAqZ7X0cIdO1OiH+ZJVkCPhHMXiI9NDpYDpZ3Qeu3GddLL/HXKnpp
qa28QtWiaSJZ5gsXdSN1ghuJOtxLSNbhVM3gGB5SnfAxEKVPl1CcT1wS/Jj3eEv3
rc+fG9kAbHhfY9QNUMHq6FV+dUsggIsJPyO0mywWP01YHPqeNc1sYcZ9dpTC5qQ3
lfIkAvaEc++Ykj61XTUeFn6GlAbCSivlTOBl1RLCJJhES3AYLdTwkmMWXqZwaYXo
KzNZP5lt9CsevV2TytL8JrSd034re43c1wBjSMFOF0ME74sj+8o1xBsVvXbL04y4
rklhK4GYpDPVJx2YFv/uDcMYaifZ8+uR3gCwmzVOYl7L8Hfo8D6egsa5464hsbmW
KdKShEQp7cUb/akInotymLJtFHNPCRK3TlVziXfY2N4NXRIRdplWItcZNDMixRxp
4bi33IVphLSlt3+eLnJifOk9QX9xOEtTtIkPgHO/o78CUpd4oFEdtpuwzZpsqawK
WUGqLV3LZkjHU+y7jqCZ2LYn0CfUyq+6257Jzyc7rY6B2s6cyEu8KzcE/8SxbfB1
Yb6fYLLOrL9/30f6T5sIfq4GQXZvrdgrZeA0iUViMSrmy9chHYbEbGtPwAotEIc4
O/BoIk+PAeFdTkZk9NY3l+I20wAew3+k0ufK8wmqy4aBHUguXcd4VTm/nhvONVXv
JEhdKW70CyyLUsRS1i/9zeCL1GSeX6jKbwLRTp92sx4v749XTp2oHOty1N+Sn3nu
YG7Wan2fCYdr1IpckE42bL+wZR8NpisVi/1MKvOCQPTagtuaiUku2JwC1fp/633m
vKr1OcOdHff3XAqd/qsdvE3wm0ckZQ0VmQ2wXaqWOnHhwfX1g9OWqn8f+5uAGfCJ
wNrk7/aiaWN2rOd02G4HTWJB2xz7TGUQUE+TUecpL5fJZPQFkYyQD9bH6Ihk+Qgq
OtwbD9qRfdYrZEuHW/bHKwoiD9X7xbh59cT1p7sI2JMMfVQ6eLM72SS17OD8WVIJ
pK5XYwqm52hRU59nZrcztEMtx117/AnLRH07Sr65ZBQzpIjk6TgguVWT9fCM5iX8
W6evG8uaWxyA+J1mYuGNqWNnWRhCXRvy77wnHOhFFTEdJDlQCam7szmnmSb5tEdm
QSMTecSVvjw6rgjT8sMM2sR3x88BrUlAeLRpCto5c/1T0T0bLG84tVANK/l64YVQ
EA3jTw+n7LSi7mVo5QGDWIRk6kCtFW24y9mnO6T4vsP+DxMiKrqZEUERSV462x0x
xWBIk3zX5P8OKYkdzt9rz9++nq8wggkeJC4vpyrXzQqdIMBVOm9J3Ua2gsJIReMM
TVQ5lqbFYNTDo8Hpb1lnruKxqpRuJ66w8RSFa/Weaze1DcKnsGJ+SxEpes8/MNm1
vLLFqc1hyZ6k31JyA6wBXs4/kJ37s87pgGTrkb+xFKJyg1bjN1vTTVkIuyAbMPq0
8MQ+wTO/SY+oJgeyGuqBX4Q7qhfKxZyuVB437F9rCpxlG7Nm1P0YSPw2OXkF/oVm
rdGKUjCA3qERkcKOGv11B8fwfy0K9227Hbdb5Z8OWZ5ykVVcX3ElASsTjFJcyqlO
QBx84kqmeI0saWBtfZALyiPl+YN4lGzZ2TZFqxUFVugzn4I4BRcV42urFpnWxpbU
ob64498CrnOFgqO4+wErDE9EcL5S3KoVT9kAWKsetApFmwyQFkWC0vdvQkrO632k
n769FLoHVfRcDRWre42LDiN9cidUBJeTwOYbJkT4OJX3Ow/TAGZT7BtAH2UQuiiv
2/Q+h6As5soaoSDZkZt4qSE8P1a+DRonaKMNX3hD/331CaHjO0ghfXFQkVp1EBV8
VQ+5eRGHgu9S8+CaQr9H1g3te8R8Q4jBX0aja82UAOfNUoCkmImCFbb5HBCWQEwK
dZCLk2usO4M7GpyQxgHjuK+7t+G8LvCw6nLm8e+r57YPtOBXYb4s2HzQNFV92HLa
X0AFLEB94x/WegHttLSLYugnNZXhZXLpq7OVpyKblllQpzoIDChEu0x+oyI3q4FS
9ciOEn76KYJeb9Oz2UjnatNempxyn62w71dwHFtgwhueOf6QPhFeA8mvmiNd372s
Afg4RBF5Znszan2xBvdCFUzcoVoAYE2qLVDhUFPdhCr7R7UVSrvwR0D5xWeCLpsk
H1ftTonvVvGQfcc4M7aDQweV/h4WYWxfAovLw0XswH6evkFHcozHLS23tpkTmh/3
WBNMWyj/L6WfWOXXKjiFCpIami1wuTd9HsiZ4RdGV6hbjCxsCI+l7L31VFtY35rQ
+JxRzD9sVi3FqS3oGyiIfVpCzoXR03cmP5TJAYV6Y8lN9novPM+fEdc9RqfL/qmo
S/byHAyV5tkKzVga+PbtQ/E91o05Lun5B4CNVfsP+k4o/6VbcCH+xh6bgD5m+mwr
onYxdhV9lR9+VVm90S9Yci8v856psGO1uRR+BpXO1pNl/H8lMNsdb6KquoeFYQci
GJ5jTjAjBy99vwnVNMj6wkmkVa4sE1bLny81TajgzaZ1iROG/lTVDTszeNDissv1
ztOVrNRDtda2lzyq6p6+t/7Ix9v1Bq4kTFeroHz+Qjxq0Xc6xd2R9Z9zisPrftVE
Uqno2CIBRP8iH5lr0stgI3pJQlO1w432Pk/7BTiVRSiuExJM995CEK+DWJHoRNR9
3aXIFLgIzvUQpLT6qci1utl1ayFweij2Rup/3m5HCQEjEs3fg6PKHM5HZSR2KCNN
AJ8OIu4qNk3ImaAzLtBf8ikykupP1Xl47oM7LU9VNYoUSrZHYfjeOPvONsycLEAo
WrubHSiGKg85dp862t3UnwgNX5C48gcyr/Ywo2N38ExeACjHQaiOJp2kHbg0BBi3
n/dQPNV2IH9kEGcFE0Kjk4QQWcGeoj3tuLlGcYYAeHBuNjf4TXSBmE7WSukRyxne
hepBkQLpDdg2Q4sMm4IEcmfDJR8CaTAjsYE1XftdycOA/omO+HvAOdSjGk4rNaNn
6qhVXEHJdCVLCMjmC2mU+V9euejhaOBf/TB5DC3R0UMXGy5e7bf2GRcJ2rqo+yJE
5OUP8odyXrAb0fwoMUTwHnjTWM88Guc9WMzROZEehcTMHhGoIQAisGBoZiSVCwX4
3x/MeeiUAQedPBm2nQww1rJssxjWyS0WmrjbY2cJnoKgG5M1ZzNOuxLdCKxEojKv
iY5ynXnRJ2DLh8Nslo+bWtOe/gpp697uxlKrk4k9EFetHs9ztYnMLoOmUiILSMVw
pbJpaOZ5dyzz/AddKdQ0eIa1OIq5DzUqGsK+BBK6OzhaMrIOWLz/fbFECJJsr2yj
j1g3411igKW1uw0WnVVowkFA9no6SdPCeXHyQvYwXIrpWPAfxs6pLB7i/RYNzd3n
y7RhJNyUrD5u7ooyFxshtsZx+5iOU8QQTpgEvpOOl6Mn7MufBdWU2xrttRt3g3hz
Yi5QVk893FTe/KcXVU8HX5Z+Oj8cgNJd705Fiw6opVj6EPkvgZ3ldNoxekqbxu3r
9tsPbrcXqzPTforYrKDEiWkh7Zu1avQO7kFpkCgHy4Sh7QmDbvm1NOx85/zQY20A
MenbTUPWl5fyXONtYmfnCWWUlfj1scVgd1NAE6y4sbmtxbTUMAtygJqDe+v+3QxV
0MZY/tENdQ38EViVE8kM6BmvDg3s6d6nH45hvcMfOmqpuNozF6OzjBenBbBbKjO3
tEpMEjLanpaaXI+JUkBX2GgLNV3dP7632g1pQNYpIn5NmNy7ySLqV2ykC/juQyh5
lkeqJiDFxPgATSIgRDeY0lrScDWp3x/s5NZm4C3ArvK3/knFmOwskzLcVzZgbnk4
roJCK30nnIBnyLS1AW9P9xo5+UwG7nDeU5KrLkTc3H7t+MJ4Q8yVfUCCvBNLwTHs
8jkYIra8NHV6Uw5fXXMzHnRTC7YNQmysD1iCyuTfUII3oRMhwKcKRG5tdEmHCmdk
MZVm1GoVnoxdbVM6D7lIqw7Ji1it4IyQ7DOPrG0r+6UgUIP2lRq5bxnXmPWCqw3l
mbrwOD+IRIqxooKzpRSEwbZFXYY0wmOwwzZGxD2+sZKZ+PsADLPIMl00PLJcS3pU
+lfZk6DhB983kkA9PTaqnrOZL58YtWJlUHEDdndKJU5U9s9joXBDMPL74yKidxR5
QR2J8hwnPNXvhxtHXL0cndFXppcjLnkwZgG2540c+42frq4c7S/4BW5qoXZUACH3
dVQzleCW/WhPOFne4tOthQl9tNUfqG+00qI9SCNqEQBx6j09v1zo2YInK+u3By+j
uoJzgEMVmdSKDTVni16azC70Asuh7Y3e3WdN1AJ27fNUOHw8HYKNB030A2SWQpMx
smA0NTXXW5DbHb0+JTWIEsMK4qed8K8z8xWPYaBIy9kYa2uVw4e4AgUilIDHZROW
RCl4E1znguS1+yksw+UePMf2T+aTyZPpaDQeetqJC5S6+iEI/miqvj/b1WQR86Us
2hIOSRlk7RalkEiB/wDVgUH+rZ7h4sFBd7SHS6E350pKMgo2SnNyMGMogCwdEqEg
RDdvk5gUfMoyCRSLjxe629cANgJ1VVtCuohmJbCvZtVJAh68MJ2ZrzD9rQJLJbLh
7JXmkpRKmz7THuiGcToBZdUbd1mdlPf3WXaqWmOKrhpFCAk/CPUPW7i7Hn6wk7mg
pk8NK/jMRTg2r8eHd05ldphq44lTO4Um6MgeqGLyjh5S1ivrMpigz201DkjKbcdX
3wmh3BhGYX2PxlsP9kapeKijhgHQoGyDI02TTRm+Z2Bl+2VyafF82LzxJOLWfX4w
yw6bVWm+ahAsYj+QL0h9IlD28xpgrecfhbjjyFteAKsXQJ2zLZwtXICMbjcohpkt
uHikzR7WnLJ9IE+sa1lEUQJRkf1Deve6p8r3/x+rnTnojr0pBYjyzBVv1NxfZnSB
230osq4uIBU3OlT5aB5DpwxwGyhbNIr1Azf7Hlb0x5nUvdkYTf+0RJD1KxLyTjTy
aD7J50ZLhjH0qeetKpTrv1pWtlfuw9WTYxNFjXytkzjPf4xonVjzTzu+5v3bh2bv
9w1YUS45Wmc419Lxdk4WaufNiDYIz1Q17kxjnccd0Jne6dESkImxudJqMJCSuQgI
EJg3Bzcr8f6mSeCStATXvgQq1/byz+7r3Nj1jczv4YBKbB+9NnFKgH2Nhermrsja
a6wqCc8Zu+MhpkTq/EfVYaZ1N+MgV5RSxaLEVr/dQqHyAYmQFwzHi3eBxTLuwN4S
GhxZsLffg6j16o1RZeqeMzVrRc1RvFIWVeyUUBm62DeIQ+chtWGWhrq0qOmCa2Qg
zHK27SZy2d3m431mjNfcRvaJQ4l9OH4yFtxwUJQc0ENBKmsrJWkMgDMS8GjKjHDw
E+apaMUM+xIjI4sbsOSB5gaigfEeQSQijd6/hH1xZGXx8aH3VGl/F8zEbjDeJ5qL
C9cfbV62PDuYgFo/QCwCzhU8V7RGfVQ8H+TPzr1POPlDOYuFtcJwyj+Nvyif+Zsq
1QcNkwAxANfoKFIs5dsDxN/zQpD80H+zSHH8e4kl5HQb1O79XoHsYFWcmMoafOPh
s9M6d+er9GdJYVTeGlectczHrV527rL3MldgcmXIUM7KdK/WXhp/jDcvQ0b3zj3P
ennsoNYFdIRBUbT0tvxsIcYgy7QsS3MTVmZZoKYorEBtw8JFnAr/DOIhmDUYsgI7
rQDBcoJFjA4M80gh0tPA4WQv76LPtnQjkquQWgpmXDIutyQJZolZcQKrFPi9C7pd
JtNyfZeg+cGHO4PIt3hR4bRAKdC/kK53J7IaBH8qn/8xVELWNhvtcf6hqotf9Kf9
K7Y0K0tivdPESjgmjSIPsnybnLpCuKhF9IE0dG2ebdTHHhgEjwMGNirDTf0kg0Eu
BAfLw6UrrbxYoI3iueLWEuwp+81KotnXzgikaforo6kzvaFTXB/+0/hXFF8Ra6AR
Zusi1gmn4thnsPlY9VFTRYi5KoXKVnaopl493lX4H4weL8RznZTzY370TaZy8UWt
yVfw7i71Z6pAqjnlpIhzujg0q2D7f+/nF3Un9/Q61FBQ9u41fckVIXHZQq7qnm4s
dBZAUJrjsN7Y430BOP5C9jCYjj4clgDPwG5FsEjQ7wV2SnWQrseQ9I2ZzSsH5S9z
B/w7Bk6jOatt/NV5pHbRNlDICUWk0ImoYBJZH0ha0zh5bRXcNf8EANpqm2MM4xd/
ki4+YKBEgT5wSKgn0Ii+eEPrmbz5ZHGCOcsmoAIqQCqKo4AYy00b2LZwK70MaZjm
nZAF14BiBr1Od5R5Fq9a6HIMvOYbdsjEv8gLiY8+d/RWrl1G6Scfq8YsdJZjNlSk
7Y/ojlhrTEoipSSbkLtJ4BSYEzL7P0NhXEsuw7kLI8lHweM+fMgMCUQpxjRY4URc
Yz3tmPc3/8JR7ShgKn7nzlc6FSnkYZ/41t3A2cbsKeJ9ekvmf0ca/jagFMzLVLI+
ehHi3ypMCV2q+HsVFLQVBqh/W+ZS7jS58sIk3iOHotXvnTAHji6xTipI+cscEPs4
MIDbTLRr8i0v1UJ0+1GoIKK/vfUovO+T3jSMnOV9BHWLoXD39zHVQ564IeiCLTbS
7oe1LYxdWLi/5k7Cnq+xfYoXzvtmS68UZqYq8xCVnjHBrz5OhKN9iUtzxMT7AJ94
bu+pPqHrZUXT/SiAgVygLtbQ1LbWyinAeGjAgIXWTAgrN5ikmRohfzB59rxOoKog
PrgpsdUxSUe8Cv5WHwd+6GXwBoZms/2pYkAVGJ7MlQ6aymw39Y6GKHhHxV8PF+VJ
Qb49yC0KeacIbv6w66a62/RZU6Wq5a3mvMT4+vBBp49kKvlx9YtDVfxmuLRFUGl/
gSvXZq7b/KOT8XJ/IY6cuuf34/X6Pgf8wNGd509m8TFUWL5LZHI843K3bSVesG4r
FGrzvyhn5SqZ+FtR9Xlk1kjl0VmuCnqFBxfERdwasFmcURsvENTd/O0yBZdv7KWB
aJRn0+7wURWtemDeefMJwRiChr3UHijoDywHEadr2IHYGR6HJ+76h1y1dt60QAGK
u3jVt1tXU3/aCkB+SKArZdKDtmp2ldT15LS1EL4TlsyYP5QpHYNn5rIjEcf+SzYM
PzOa/Lm/FGwV3/Or3rr7CNTGP0ZqqpMCYIRzyt0ZZx4UXes7y7upiHYu4BSw0Y7J
i9B3m4aSJt63t0ybGHSaO8CLnCq2f5ybKIoQBsLHVLbsFUeLLVVRqMsvU7fTYWTp
ASnAv0Piy/0+7AERat57AAxWMvCtbbr3oMzSpO7SiVrnjQkQ7/GHEgfg7pfMe/UV
Hm6AzwRBJKBUnCk18vCsibX12Ljar6y+yMoUhxq5oI9Zv7IJVR5CfPtF4O27b2ei
maIDU639IFBoCrOPVF1Yf4VHUutRo1bPrDJ8wcKnsDKMCSS7KbnRSIJff4pG5amU
yiF7t1eB32HP52d2ydQOZl3z4k5i2C369RcCGL0kej6k4x0dcJwT5WHZXugkao7b
KsC20RHPdTGr+/ha6KI0WLdmLEg4oZKNM5eHZavwET2XoKLgXTiQ39SL/Q3yGEGf
c/AOl5QdnM6zW/37vOeVXp3k04kDGfWw3m2nrarGczWj0LkxKS6ULy0rqAGIabAr
zqJkoqhdU/hQ4xypdv6MdjL8QQq8k0etJRCtrY+A+QBm+zL0lNR45ir21UnnCkcn
I/jijbVUswUz1afX8eO48r+r6tpx84UJCADLDZOfbc5LqWZflWFYHtC7SA7LTur5
eueVxuyq8ufZzg0oVBvMpfanf/H8KoaIJ4oqT75pXa/iV6RSNSikZia4KOQGgFHT
QHQ3hABCwMg22scnaVumoXWGMOKPhPrTE+wMicT0Da0dMTr/n8DbjHkGPVwQkZtK
JKhFA5DA0Nvycrw7m+ag5XpTn1ZVMdS+cutdLMPrMaDuyaZh3KAbuFngitclOfsD
e6fMmS3It8qUytIzPU6Mz/Ll/2Om8aLDVLOg0DzyPBvJud7l0FTPreX9vargjKtL
VahprKD3mM0b7IZhAP+Pk2x2qgO1txAeAblVZjJY1Yu1zQ9w14AcMeA6txZbJcK/
bqzWeJpISl4b9xDrwX59Z/4iZUwD4PQhBixmIp8H1fms0zSB00WElZ8H3Pw4C2iQ
Z8JR+ipS5d87dtYAM1XeL4+1fqDCsv9YQ6rE9BpemefSJgpXRq6O0f5tnQTSdalK
WCAWgMgIsRxCdB61RZlLmzQGGov3UdFkSTgxLMeEmOOoVUfAO3ami2K2SPJ7f2Xk
3CTpaekZURY9xxppTecoH+lU23qvExEiKtTe9uSsz65seWeEkPPOmj/5ae7c0VHd
6/RIce1/lXzXU9UQOPYZsPEDqmmjfLnFX+MzeZjtWhweIBPIXXRY4aShM14W9F/3
JG+YMgxaz97HzOCCl9/jh8zS2z/W4HEL/yagJECgU2qqJhuZlJjprTIw93h0b6u/
J4E4833VQ8yb21oH0gq0Zx3bWtWqoXhHrbEXs4K1GQTKr9lUYzr3vBNNO5KGiEwm
ICdJyX4Bj7Hj7IKdR0izJGpyzhr1ieeR+m/xz3kTdsXdcLu/Ky3vBOMyI5Pk98W2
87Rd4q7clqxnrip4EL1BalExhePATMHYocIEE4LDOHZ9MZ276ro/cOejSKs17xPd
iVvyCZ+CnI5SK5+27LhTOA7gJLu0ZccmHPzWo5EYNY9QMA2cr1OPJwfFJUwsCXqg
T/webbQUsEFxZat/R8OKLDligu4IQD2ebmwHSvIjLhiOjQ0/E2zAh1jUOEnPC/B6
iQNYt04agN4bzLXZ/jXEE20C2DVnNplaSzXk/QEj2FOr8m5F5rOawLtQbkWYuHT2
j3a05cO5nTyjYALjAjkGoX1s3sUePChygBqGp5EXFVdySxvzZZ15kaLL7uq0ps16
e/yQfBlDjXvpvGJLKCKp5aAIObWpuxLnUjct6KlEQJPta7Y8TeorwA+pvhgvbh1T
p2YIcHqe8yhWnJXKbQ7MiLZu08UoF6afk3JtVOIYk9ykpouCnllDfXEshWYJk1WN
RAOQi0VBCSIBYzdIqmB7b1jVkAOMm95S9h5TvNAfZxewbN1WncADdTXbPsWvjJtS
K8Loz9DeVRft84B6snyg/Lu828+C9+j7o9wCvKb/AO/wHdHd86pcT1nO8GrZuLWC
FNf3L4/LSVun5Vvd7blIYBetgJWf1V0F/gR6NQYyvN5cFOk9qV1FCwp9xc5mO2bF
iz/FMYD4D0Z6qXUyEhc3Ie4fZW3vZAz0THmrPl+4Rp09SCmL8/QMU6dyDakro2DZ
FMKYHCC+Vf1+TxMXw3Gc1SZh/UuVdk0RLw0iwqCv0zA/bE67G390Lf922Fw5TVNU
2CO5eFZDNSB/akW+yQAyd1CKgEIQWlRWHk3rQGq8nGqTD1yZwG5AbM3yoPNFKkQB
6BOMcQhQILvripSyt700dLdLralYFc+eVV1ISr7AYOcxbPtlwNA3iabvGAAXd7RF
RgtFhMancG5SIl8kWbgrHlPG7zeplADVb4TPyKoHQ3QAXIzoCi6mDhPd7jikZIKg
eEVQptkIrvgaC0w7YLaiMtXcWkzSel7DyS6cfaIALvyM0fPOCRlGQzYVIM50XTx7
GF2mGuPcdUHYNRd3iL1rnICduywnejvVYn81FyFaGa6DP3EkXFUat6suU845AW/P
fWlpY8HkvKTwhMfxOJWKcAXKItT6lxLt9l8PYz/htBIRCjly4kU8FcnstllTTGqG
pj7pWk2p1VUAquCiGVGYRCiUFrEdNIFQm4ylmWGX5bnkA5rSOBAkRLOyqDB9gQmh
3xuQYYXgVjgvtWtuHHf/man6QNhvqtTBUpQ5PI0F4/pUKqEAfX8okRW3frUInzBm
Tloy5Tr2NxNGo7ZSTzX23jymHCBJY/n/VF3DWhmMMwzNVOZ8TobD25ph6oawwcEr
Zn+6PCYnUbFwesoLqK3a/gqORJkVoQFeKm1YXnvbWi9F0S2zVmSlr2I2rvGl9tF1
9UPspc1Pm15Lh5GKuZUAq2tO6tRvOmpvZb3yiYaE+KihBIPattr9koRIscfV62yM
ORkuPNPuDFW5ULFEzjVpEPg8zgA/bmCjBQPLYftCO3UBE4p77ADclJ2+E5bDCMWv
neg0wS5PpQ1WYqhEV8dPyF/bGyv+UbgTEuCSKwYDSYdrVCSbHBay+cX04fLAh03S
bRXuyeUTrGK+ppvk4ViEd+fEy1/iSTjRo8ZFC6E6c23coU5bFMUR29bo8NoHTLZC
L9ht28mLXHCZplp2LPd33+CMUCWO9VrhvF34+jlVBYRZW4pMmpB1VMxPJQyaguSn
E97lexvxLAFHtf97HPqyZEXvG5ZZd4JVBcTwOHpK+ZzLpksg2XfvyW88i2W2wc33
5q1UiJVxiiKJv2ZeAcYuXXbRa0ojj1K68p3iDe9i5VfEWKBskSbNuOvsbpfZJX7G
PUBWl+OsgZX7OIyetwe5NP8gcNE+YoLmLOr/NPelP4hPOO0fzE7MwBzYSanRuYyt
/CaD1JMvEu5Jw5jub2tIzpM9Y4NI1lStad730Jfx61gmLjJ26VPhnxfgKDE3q24I
096bzuJ2WgftgJTHbXgUhKxq/YKvbZTrHxX18DFKs2T+VLW55cgNqP16LtqL3+u+
NYryVzAbjDDuy/xE4g/28LPpL3cm6g4X4SNy0nWN7wizfZb25ychLlttRoKdJ0+Z
E9hUeUB8POWNVy2FQq8hG4pVgpE0FkHnXNUz45v8qfR5MU4r3whKY1fZNnUvCyTC
EtnkCiRFB7o3kxUmLS51Bf0Z49lJi/KUYLQaq2aU/zxQ6rP/gqcJbfyPnV8wAT68
iXVN2B4/q479qRhdBBVq/pQ27bCQ8F83f9X4JvikapViwrzZDAa8/ZakroaFJMKE
J07dmvfkWZ6xx4EsrmXMl0bZ5IFeBk6Zh+oVHVnhOOPUuSrl2EJnbPJ1rt2zt2x7
i237x8VCiZU7CsIvHgKV9Ggfm+zcvb7zMxKC8sXRpZvKfMiAOB60nFBKOp6TEuVh
bjNvkMpEd2uUHkKAgjF9B+1OuB7bCdJ/hFroAtRyRbYwlVIEx0dqDRtXfKqIg+ND
xWm5RDqLuMQmQlmDV81zkN1NWXg8V20tfb0z9t4v+KT9/qxhSPwr83AJgKAyxL72
9Bf36BD+F95rlNwKAyPiL7HV9wYqzasgswN/LcmE9v++VqzifVBsukgZ39L1YoxN
QSHYYHSwkGTKsjnaVD8JhAZ67jCSEICMWBcxd1YunIlgM1ut5D1fmTB6vJwICSEp
PuqOdCtdyJxYzHUPa7q9/T2C1JF1N9KCi8mbIZaECO68F2ee2ab3DFaULWPizYlU
TWcN1pHDcFdHxRWkFcgp3TIaHz7k9XhQ5D2NH4l0D4n7NYth7EXZNKAR8oW58AWR
JsbZEcOmGpzcjqHotLQgJ5pPOhYwNM7rgXVIIditDuE8YCEU0qDqnmAnxYqpd4vH
Q/StD2GhA/6YZkJ4XgLLNw08mwFvFPveglzntZMQ08slBACT7AwY/iUpWnNPbyEj
aFRdYgKNQioRR1C6pP8kBIDvMWoOUXM2JftLyjYnzb7jTCbroftAVTj1XNXb6bmx
M1zxNFAogEknSIfFgQafY3Vb3lM/jZzPGpYJ/Y26dSXAxyuV/HR8+GgpxCUq4Tbw
A5ugFtzpHj257OVXtx0J8kBggMbsV8pBmkfjWhS/BjGJZ+Z1gr+4Ymm+62DSLeBC
fMWNu3VuNZChFjH9QHwTpzZchaOMJKb9LdGruz8myVDBLVZUEPnJA0khUBiksos8
IgPmLGG9r4y7IMEY/6NdZmUMtPMVgCsQrlhc4d49FCdonvJ6k/SQ+gGa8J8brsbE
ZftIQT1mVygmdbDEbtCnzdSCVXQKkRHWavx3Fh255OgRtdxUts+WqqQEict5TDpO
O8YEgJYeCScPfFCT48JBgXLljkYvjiCtdn5ne8ClnGyEPwuAMVsZ6tG9MfqNqcTX
X1GS2hXw8mSTY89gIDc6NGRB8kOZWKFiPLx1t0Gse8BAG1wK5sqq04jpPaloTEy0
+Zgvh5eksNrfAiAVR/FfnCEssepDAJ8Shi4l6uxt3UlVTeuElub9GdUMb4bRysPW
IRBzawKnasoUtl7TERB/TMUaDnJTeQ9u9PehkzeK8Ust8ZCYxeqRqy8ijGHh3pYd
zQgfwm1DrorxtfPZgVQoxcBB1kv+aLAur0fxosrjFrqgXjHUZkiMXIBB8utomglx
4a+KWqeFDLXGvq+enekkuwm9ud7VeUJtZ0bK8JGDeEVIvNtUXqE8E1A2kkakO1SM
gbuOuRUn7tW+kevtzkoRMf6E33BjTe7DDDw0P4GvfbANLyor8ghDLJ6xDlPsvajV
kmUMMFtG9g7NY9crTBpIV47MNpa7u/CkiTv22QXPdHdVkZ/jLGUbBOBIeaTGjdmM
UYEMYgcntonw+WN2wtJGH8eFoyql/NvMPIgYRh3QJAx+qUEpi4Obv1Pd0ERHqUxg
beFBOezZSNdB8DvHbghGu442Fha6GFmg70bySBrmU4mRMG8FTIebg324den+B2we
N5LLps5Np+OPpnSmtArKILmnLthnCqX9W0WPKa8pW9gCGGA5LdRpW8Op7huTs9Xu
y0oQJ9O0+HC8SiGoZ3k3MM1OUbOMNg6SzKYwDVOegvsfD3Oi9O33OF+MeDOP8NSt
op7OiSAH1En/XQuvHMhbKfBC6sp0G3UiXDmvtLc48pTDkLtGXIp1ubKLpFSLxKzT
IITfu2BOwb2ENSDDF0GRLbgFV+Ux+ifYPzxPfmU+DSoCp9Nji7N71n3yTe4Um1lj
UGs0JcfUdxFbXZPi1KIS1ZNGyH9xuOQxRQbvm9/fDxszMCzPZfkf7hp2iw8fCQxy
Q9MCigO9uyhlmWEFDSqa03sFEdeZwPT0PJ/QFwNadcPkNbb+wcUym0ObUk+I+56v
NrftDGzQ586iUjrzLEQGMEOslREc6XrDAgA9Ob3NigY4iv57Kl0F2vo08/pAja/N
Qee8ZFXdXEe3baKr2wH00w1+eD5DphvCRSzJDXHYeu67HshFruybpaWhlfoiNGGa
rCnU0CdSPYz46j36ycXzehua/MZZN5QYnVJljmPGT3c8CDW43EuyKBtqq9GhGQfT
AmopHD1y1p/ljr/KFrY/ZcYl4TCRmE1NczCoRztNiNo1lH6TDt4yza1o0GI/VNoo
E8RzhrBJ9Yhj9QmCU5Y32koriefYVm5knmgTcsx+WbJvgKukf9StWlAbyaLdMcUF
TnEWIHZKOU+LwJ1LyOY46bmxrsE3GRvHbgsWFu884qhZat5Gvdi/iO1R9LSclYqQ
qYvhWZnSdXFUDOi8IOl8LdBvQhEnVlWup7DhRH1ek/c5qCA9oKNKpjMKUF+snWd1
xI8x4q10u54hzroWONko/8QiiobMi/NDsszy930I1T3J+MZo6DiaYbVlrhiWpdEn
m2f6FZ09+BQSE8hpW75B+2qBxcHEe4w2dlfNZpkxV8N4jW4BY61fnAd1EWouUNMn
K1nM65gNZCYelUMolqP0yd9Ye3zJb33X9tsGJFuYyASaSxdAv5sJUKZ/ZW64dRME
beSfS3N99W8sfxxqsbgvrCsTL/5LSmIyso0vzHaaze+iv76EmjR8u0ozgDRRa+nc
6R1cFnbYwfiYJGUyceXEwRtQJhwOR+RlRrXOaA95AOaKG77D7epUMCkFNsLxlbMH
NE96fQL2Q7HaDWdXrFd0+fYiRAQuLWlUmyRBs/v8YnJvFNky5TOpOXL1k8VBXOZF
rqkMI7J0MmI07wxuAAl0/ZbuHADF/lyhe0kNKlk7mAz84tUQdCkjO4Y/CvEb9Qqn
J9U2We+bzSnBbvS6rP7VQynFnszVCDGYpP/RYUXuYBi7eRqCCVK0i3Ev6Y8JKgpM
GTi0PEPdnrimG/1wdn9eGVQX0nLiuvNXDCajF6fwSammGTp9Gv4vBXJbroe41Fkw
m9uuPHIxtzKU43ImJcx5Y+/VE2UbUjFarbcSU/jyYcE7fvlxIxBa9BalFt+hSuUW
tFib1hQvkgONsNvldfy8Ek7d2ySC/sZ1SCxCB0Q8e+9ayBr6QSKC0OCV9m3K9Xvr
ggtIL85SnJ/aUqJPRUHK47cWl2eMwAKsFu8nUPT07XvGSkk/tKZERGjkKGyCGOt3
PtSf3r+bgKENJHK4GPScIOmLMVFgW3TL9aB/ECIKN3oBNNKBvOsKzfMOevP1zqkc
5CPCt0tvxk6PiUd2YPqHPHh7OPav8dYngb9VGDQ5q0285hxgjy31v8kIIXEqVHfL
XwcyY85Ua2Gamfugvc5bQ1r12desWimVfXsNK3OeCiQc71J7JEouMLLyawd3wFhi
0SKL/WW0PARUqKjJ1wR8Ri/emVWYinxn+D/wXKtiO2FrPzP4SzmJII/ZIfEZkqcS
0PcBo8x9f6/B2er3Ubgbnmht0vSLhWuxGo5Rf90M1Ulk1fStaBSdTMcjrc6W/YK7
8z4CWeM+V3N4bWA0zw9fJuHkGJYQ2PaSFQKD1DWzTivMVbjgMsieDVjkcNRalEP1
J3oykAkHiaRCFgtAYF1d7hskhNMF9yDb8ZUnAL42aV4dWQOc3VjRr9blL+s7K+aD
xbgsU0/QGmyhjkC94J0IvxoAVnCOFsiq35yWwH4mREjpvXDxx39TpXId/JIlQb2n
OSFtWk2WHOs2lcn2Zq/iN0ms2GZJOsClascunVHyeow1I3WD+eNypRCFohEdZD9Z
rnjIWRF7o8INDf5+jH7onRmu2lSwNsrP33VR/02XxSJfap3Wdhl1AVJYpBSA0uYP
JSKIg8v5ZmY4xSJaSyVQGQPdJXNCc4970VnMAul0PosYDVSaa5LLGHfzR1SEIeV7
6LDk5jwjXHpAKYbOAdo7sGuQCmKdEKO0veGIbP9fcW53S/0Lb0hIRGGRECBVR+DO
Oea95baT7JxWjabyMZWARgoXJAUXvnYTC5LSiHqYfIaj1GoQJkjPf3JHLZY7843P
q6/6xER0mA39tm9FlHrJgH5soAApBlmvpK5QrgCdZIPK237MbWQRH08mMvdSRPqu
FeiM2OEFmfWtYm7OUF2ROWF6p2TTF8//oPXr1TFKs37I/OhBvrPBX/74L3LXS3m2
/b3VpTJcs68/TY9bmh2RzZmHlAIia5frad64xpAQlFlvN+HvA4Tl7Ipp5dVs/Nbr
jDKWN0Z/AoOzrDWnmdkhAEGZbsuBMJrgZPTSlysWyTbrCnA2A+I0w94BenQCQDw0
i1UKhtpZtaSjBuSBc6iegFnXmKVdRPKiu+4auuROc/f+H6AcNB12a+yqkY9zYd6C
EENLa04bTPR+NQ8wEJz0BGyBuNyiJYzIo3Aj3FMliDW2we069VUoUbRg6QJgm7A1
0NafV8zAqlE16Vuv2mkGRdPMb0C3R04DhOPN8xJFU0rvug49hufUjewp4V71gsjP
rR8yHieddbcqSlVgGEjsjYkisImSjyiWm63GR3ncP2IJqu4gCCp+PP6bMY6MPnPJ
V/cy1cx6foLhwTKqEwUZPgG4Lift/D0LbHOlBRRZ230cKfKk35xb6xmtYymShwCl
kRLKxBO+xomiNNSjHUTXf+UUOKdF4zbMLQ3Y13zyzSZZZ2AiqdfDPiM26ffPmAI0
pmhPR9KujDdbCO+Rniszb6sB0eRG1n3E1YgGJvR3nDhWeWTHv7ygwF5P2aNV7Ho3
AwGvWqqyVj6zZQastePTcdd5i7kEDyARHIXvDTl+w39FQG+2Ro/dxGMCVCCi3ymV
oL3x45vbKSQcIR7q0oTdM8LahwGsDZ9aY55LzKj0Zh+pcocurdtefcC9TvqGmjgN
zpl22ZA+ys/VMSMEd15VV6kU9T/tTP7UcYU5nOxtN3ZDykXSFMFL+XZB7RuWbQI7
nxo36HlHzYqmtLpq3P78Oxzz3r4h9ROWbm+ioeIThQgxH6onDcyrcE/4hVsd5xa/
6SrowlWoAw4LNNg3SSjbL8mJW3L3yvCdZYSsuvqkutL1W+oHl82YRWdtP+kKlX7/
ZUfk31Pev/nHy6OERvyVa79500qWu0CXTiYusreNCys71+uXP+aA3qb7LoUL1fDq
egoxnlX8oehgYLs/mE6AWYYMogoxnqkhqX0/dis9oe0ic7g/CBk34Sa/wR9ntTBa
kCnQXheUNfH3QNXHd08ca0Whh2tU6qG1dwJzg9OP33txafWujlF0n6q3YkdIstzw
BjtgFMNv/mzlBd3+vTceoinqHS5IEy6e9DaAtU8rkA+x3SAcQHK+HZwRYFsq7uWs
kMn1qjtFAe5Sb/dXRNgsA3pVimJBfHW3MOYj9YR+jBibUylDUPks74p2PqJP+bFS
hzKDKyJu/D7pOz+QojRyt40lnQBEWrgTBpEfuEE94cdQRbHaZJncQVDk82SJ+jVq
25rbwUVtDZzs+vndhsMzL6QvbtVZZe0W3PCK2xJOFLthwxIafHm7IbDXcsXfFh3M
EM3902i0J7RHXooqn01RggYMwguAqjofNS8sFc9dThC97wyF70l0Aw1we+MPIa7L
ZLF3/0NynEc/rOYn+m6vVzmYNpYjFzvWZiK+Qc8pD3O+4gVGufN/8AyVcF/Kb8P1
41za871d9qZac0QAwtB6P/dY6zQbze3SxO6W08yVMfNeFh6SpKrfxVptihMfe+NS
5KPBXrZaKoxWCWK1eUWuo/cGJ9I/OLjWu22sjvzogFGT2KQ8UdUbIRqvYz8jrFmu
ADcBUHvN0zcjvAC5AMirSTkn5oDRz+6g9C7NRmXZPuIvOTehcaZ2ml57Ku1S4K2f
AUEo6p4vVHWI7asHp5ZuLBRtDuT38DLiCZQNP6h/qDuKJFH9jDCNa+m9y9C7AEFX
L0cq2Gsbvy/X1Y3da2w5EZnywLNAiVkpcNzqgWwdK5xcOQDo5ih7RKLNdVRLjCv3
Kxdae4ADS7dhxWe+JXWM8A8SqzCcGjpODlDb3gS81fw84tbUN59CnmUbqhcIBAXm
jnxJr0NP2K58dz/Q/3EYXsOmMEF5nli9EIAVOolDkMGJxeRqwkmwJhwk/fLnorr2
BT0heiKT1RO5a7QsW3CXREvwdKsy+sXZ/qsYcKas4wbyOrBnvK+QQGnSZqJZE1qF
4SipSIa/2PZUIEqDu5ZaPnB5exNMJQkzs0kou9qsHHb2spERlxRoFeIFBp/S6+Lf
rZWVI+oYEJ5YAw6nsovgsMTZFBAoBhN/+HNj7zbSkS3JZbTyan2sX8zLudahEkOv
C358Ji0jLusDOnN3CTjVtg9JHeFLHa6gufCRAljen2136TOT0MQn10kRbfn0xQWH
ULr8f8VxXT6yXgLv24hsGr0DH+MWWaFL4NrSdBs/lptuGPFTD1yU8oHR7NF1Lxxf
bW1QRsu6I4wMBnI69//+1jpYIsYrlVxk7Y7t/n+2FUdZnYf6QSOhQsZyWm5QJLC2
pt2R63EuTfALD3/6BWxvfAMgKaI1cXaR28jVdtqIC3pshfH7M+Z7Z4V7Ithy4TMp
j5DucIgSZce1yojWWUuDr9HHXSQzG5lTjST6xPB65FXMT90Er1JIJaE/+FNIxbBJ
e8PMqZ5NRA9KzKvo7tCS9K4y0qY36qLTf0pp2BqC6slbVYT42rWsFgLydZ03N1ko
7cOxuJeKGAcIjGZWGAQGUr/h5aACXxXpPYLW/WpmenTqFblPKPrgLCIx6nEfT+ac
Mv0PNzA13FoaabwdjFbb6ClW8gtgv9bGus/bQYPuosPz61lRBD/wtrcGhD/YfWpi
rikZw+03wNZ+YLdBVbIu4YtXvAW+UvQIVNap9xGCNORqnUalcJntcymVca8KhnBh
9k2MmQavvtve3EVm8aXPWV//M/yEWO0p2tHYY0DKFPsHjIeQjDaNgSrZHNHq/U9T
ITD80gdnap5EgsJgt2YoO723iFHbY8PzeU06+8eZzDNMvk+y/6QxEYAMsa6o5pYn
yKdnd792462dMjZDRLo5PjKheaSwP6fKJTEqxAgWueN+gNvBW6dvn9A3xLCqS7zv
cbGEO0z0bva9zUKqb+vvnaTYHNNJ0Zg8Xlbfzh+k73CRYKzJmhAmFrRG15/3r486
6qMThBH5fPwqlKXv5Sd7FNo6Uc2IYGKu1O0wpvYsXvX2kWDYFaiZ2dkmzmti7vwO
Dj1OQ3TYeVo2ANi2HrfAltcks1c20Fu1oZDI7vfyIxeYKtfZkGRAe3Iu1KdHOh4X
B55K5KGmSWZ8MsUVuskHCyyLnugNSAyh7FDGNSC5F0bV66wD2k3RWAjwollGfrzo
MNnDBuTjo8nhDvuSTZOCIyG/m0GOm8yvOCeZ+vkvkRzyqeKYbdBWvUqdZT5Z+zUi
8VbOij49jC6b1KidvLgvciQ1SjEIrRSNCxvsv4fBEv0sHPBWrnOt3hMxWFsP/ajE
J0FaLKtyWuJklvYXVzuEpy/jFQhSrIG11mea0mV3cctR4VtYmJaIN1IU+s82MvBi
PgFwn2EawmLe8LC0qcNhZFJyovvdToq6DtoouaHkw7dZxxuzX8It/hEc1pTrVnNq
49ON15YMEHRhgsVaNvoFQ7f21gR1/HltNnCD+myqCU76z2ZobC9uzoMtGZHNp1w5
ueoskyCQYF3+W1dk0Du5eUBgIyT7dixRMotsBEN/E/SkxGJiQZHEeHZbQmnralTl
QbMJc+3acSOyafVsYw1pp2I4lTGYKnrNQCYCFAz7jbWlMUqN45ME/ijJ/Lbs7TrC
xC10pkuFSrersySBQSRtNPV5WG+rAhUV2t+eQi88UPuH49fmMXWdkHs9Bz64oYzI
ll0h7o6lnLlFWiG99D3M/L12q7JthgDP3pQWsDbrOB91hofjNHJspy9eqbZMcIZz
kQJaM6HfWwfepLFtQsSD4+0nDtWehiOzTBLoaoLhsSCRca2cblyAdbyWKa5D7XAB
ooa5Q4080Pl1yBDIG5aHq2lMjU36DakT+vYAgOSVJmbeOGLPArl5UVjcLGur6Dgz
wt4S6PTjxulR4WUsNifW5xb3BGpt9KpCMk3vUHdRXTsHZeG3Y34nHeIsc5yEt4Tu
tee1UmlF45QrJf3b8WdsDpTZxKq+b5FpA9nf/IgOcqPk/aPz/VcVjKnNV5lKrM6+
qJW/vxIQiwdpGTw96FFe4dm+NRo3w9yZLBZ7dOUm+48RHH+6MF89OAXs0eZXgZq2
PizU45IcXAzFp/PfHNvWn27hNyvkWJPJyC5O9+pkHWJa95y7CfoirtZmn5XJfTwp
CXFAB9jUvIDpEBZfuoBNtf+EcL4HuwerSvGQ9gJzBGGS4t55UPKvRy5uxKy91Cn2
5KOcmo5NSaOnbj13/HulRzeVg7zeXNQW0ZMLlRQp6kj6iwZJ18tCAPFZg3hEiIub
62Tz4LP1GirVCZ1xFRP4A8aoRxFFkFl9GVL25RJ2dK4Ij0sEbOM/HvUnK97gdgav
GBC/z39xcoxPq/D9U4igf0Ygnc9v1r0JrnT7JHDawpKHG4+TAYyw+GQMIbvbABN2
0vjFxcHNMs19Yq9m+1Ip6aodzWJeFpALc2e9Rj2yui5zBxX9NFQ+TDve9kmGHqw6
nBPkHLTDej2T4jAaRi1YgZr4obYrV6oA0wbrLGqPfjLgnr2e3cgbqj6bGOIv5GJ4
5qBUVcZd7TJWQtv+8IdlitFgUVD9O8OXTFkn3/chr4C64NeQP0XiExIdgW9wyCBn
xSqIkoeceKhA3NtSYKlqMyJL+wU/yg8pV7gKWlFcHJZubY28v2Z3BIycZ8b7/JiJ
CuDc/ZuX0ian/5scm8fp4Z3rCI21ippxTSuD99kFZtlcNMQVLoh1KnMx6KgvPNJt
VqSuX/XVQbj7WtOU80QFjWhMMetKhJzUaEPjmhMgNwpydSuxxlgsjFr5Nrdy1k4v
yLmgt8mnfiWrVwz/iWTdxMZIO7RNePGo3syz5R+z+Kfw81ZtpdOxA/C+a70HU82R
rOtM3Lvp0cfA2HB+5AWsQkQPsvedof4P5DnJu4FP40yR6MqStYw1lEQogyT/8Uft
PXvsmEsH5CgLDfhlafJA+IjVlAJJ7fq6PWNfQN6AFC4mexSBr7IyyY20ddDyjgHv
CTXDSayAxbceQES6nBrWpKM4yEybVJW4xavOHvfalAY4jg96pNOEkjR+FnotBXzr
/fkdPYfNpBGlwh+wK37daPUSxmqrHp9b+M3bBVNuNXw/uFGv3vk2ZjKEX0fVgBpn
982xykYfs7D1GqwktdPHLIDW30PvVdhgkwjAxN8AeRjc6nJISfBCLmea0CI8Srpy
dFJDJapmxtHIjUs4TaSDzJprxOX0cDG7kMDiLz2oyVQL49o6meiptsoepPj4ypmC
khtK6rSYWzQeWjSH/TOHmb9QuA2kfYo/FMfooEeWWX57/gyNByud/QtQURyCNrxJ
7ZDnskLYAST3O5Tp2UB/dXWmdQLwR163CzoScelTaeinfLASWS6nkoxh364eWKSE
kYMr9S1kPc1c2vYAtnMQ60qDoAaEcDia4ukNcw2icOUJkIAdv2C5q5KhWHMt54/B
WbDkAFF3YcvZZz3UqWAsWMp3vbj8PMhlG3Au1CMLttc/7tDUdEQO38ZyvpdKdnij
IX1HzLezfIu8ou4CWi6GmJm+uZj2aKJjLkeJklNfMfg7UYVP24f7dXY1tn4PoQEJ
lNUbkiUNscLdz0Ggkts3878ApDNbKU2wSfiWU4/dAmvh3bHTQfaMv+GyuYjWm5sP
z1hlcNjynDxbWL85u67uJ5k6vkxW+giNitvJARRCapWS3FNQ7n2xcX2MMXu5Udom
EL2aN3m9zstbJk95irdSZZGuGuKb2AaIUBdLcb54+VNm4/TYCsnDVpsxiohHplnD
99rdajn6kir06Rli2/114FLw+G4jAYALpbwIzI3+5LJT1JwPrZAYgKT69iHUi5jT
0TyTZddxwB9H+R0h7R3relk6vQLcgz+DUiXye7TNZolxe8Rzvj/u4CJuoiFI6hzr
3ZsgwALO7F/JDDeX6o0ocWMzY8CTvYP0rWvy0np1EwhchyklJ5R1sl8XZJxK61sP
CjsczTvW+aMZ+ujv51LSe8mlgfYXfyxCnkZpdCYv5AKcv2fGryf89GgCIBSXwdQV
E/jo0/XGjC3YQh4LuRFcl2mtzKsHAEIwS7HLnH80mfUe7u5wzrOPvFLRejX3SX/g
L6sQxRhL2/JvJoWkE5wxpC3IDCRk6mFNt1tFExpkxm8lZOlTsGTerIJ3GLlWXqOs
jezvlTeTH2TDMRJva43v9FkUbONti8fOVkA77j0b5YpH6TvCe7KdODVJ5CvPuzva
aA6GcOoAr0eKOtdWwU98m/yXZlj9KIV/ervjSYjVxFOuail15m2eKNGbvOaq/EwZ
a/jddOCXcqNB4XruxYXLKi7v9iKM9c3YQsKQ5AhwP1seO2Ea0SJSzgbuX7vjQJho
STtutZ1134ipYVs0fE4LDR9/UoMJxfLTKmzzaSuCCZ2WJ4W4pBDumCqZVTBlFa22
C7JV0I3xa8gNU6V8LdVKUVQERO36uLCuCMFN3hIUz8nKNyGQY0XQTtu9lI1+kmZ+
J04ZQfQa+ERwXVE5Ndv3pQI8OxIOB6c1VfFHb8u4sJdLdX7qHGjO/bFSBJ0UAHcN
i7zTRrKBNr+LVkje6J883RIOBJ20ROe+Ooz155kL5mRFnRHUKr/FmPiZbHFt7xQi
bnNwFdSt3d8rpLTDT9hReREdwBO91nDnS+mgst5hP9ZMvPAeAI5Qkp+mylfu+Ro/
udj7bYyVb8aSVkpno6ku1emlJbx8kYwNjdrJS3pxC4oQRqlGI91Y1NrwjYR651Ct
h78Ffbpk5bkv+0Z1R5oLtdO35/OuZ9NvN3ww19GI4tfLg7a7Zks2fwC0rBgaILbr
B2eFUFoJC4L0GcrAFoEXC3P0/9sbnU4J36G3SAR6mdlCUpuPr0TSLHu9+N7AvwnC
0NPqWpViCqBZ1eAMXeIQQuKGz8ucp5bANXyXuqdXwVJMFbVnDphcBgtyW1IsNx8b
vhKh3iez1ceXXnQXKvB2nb5beDBFOkoCcUo8N5AIwZxt/xEgRq90a8AKAVFO9IYN
BmiIo0fDdgLUtAPmlbAbkDZwYNxQ0T9NvcxUytdGEC/5Gy0I9iuXjrwfO6VAJwNi
nFzsM7yCPAfrJEKoczpaID1RaYouyaiuh1LgtQC2v18YEulEO3lJi5sALvbhjWoB
xQU9/RelASNiLLb5BFMrc8XIFQM/MfiVStE79PgztDmfCV9iXIfGrRJmzPBYwXR5
o6rMfvDWvMqhYMEmeUCpros24/zhWVRjX+jt1pCmP3Crk+k9nrOXXFyFLGamscR3
lgQxF95682oBO4YwWF2P5893yfkqB6nolN/icWr0WNsAuhcn/SjooaRBhNah7IMJ
crtNFewoBmdU069cgSShTVa+kInEuQBo1H0Z3zEd7K1HhqsViU+qaw08fUZ72M2I
79OgIsT6FE28NzGchn2LaBo7qoRED9mEA6DOnMpMYUQI1I1BDnMJC4LDND2kI2YB
OIkykTDCCfaI/uo/oEozj9Enpf8ZEc+sirlao0sELr53yn736m2Bevpy5FD58Dom
wBnJoNIL0yBWO9HtKRURR3ln8IevIkWQ3orFA6qumXkbd0pbZTCXTqTWFu0F4fxz
0JP2slWxa5SJbrSXsVemLLmrY0/qm+Yi6CxwfOO03nqcyKUBTF1mRbuM+VhnKjay
QEscFElsIcFk5dyoIpDb67Ikk6vzedofvqjnAm+/z0P5J0tE6QpPVsRxjd9M8f7R
kkzco7pA1Vd6P3F4tbi4HytEtzgCEMe/zw028i3kX2C9RMZ+F6d64AdOqpWba7Us
mTLTkOqoCVBhlAooaTqmDNx71jIWgxj4++syRtIgdEsBxKCyL8vblNORz1fVlogV
H/TtTknFgMx5gM8qgT6MuOPToAnQEcQdY8UnzyA0rTYyyonLDkP5XjToHwonNN8s
k6Lpd0iD5N6ZT/Uy5TLS7QRr925AcMNmXrnVdJEo6Brj/njrRDd7slxwe5l0PAlq
wzuCRjeLQMgWTD+Eg6HrzatvcEt6hbKG5118YQuAwGnDlUGN3l+3Hedf3mytHxQi
d0MDvzIpb4zHWFP9nMKSnqvv6k4/WRQ3T58JpexwpYrS3bk/PLO6RcwGLkTgMwQt
fkRnFFvaw5tEvTdV2mCEvuCoQWqhxKpXlxoHemL9NmEOkR/nGjM1OuDQDIIIJRxL
x13iwap8idsJf09PRBjwgGbGezs8oaPWxY8Adurg17Cgr4v+clzOL/KI62yHt9vA
QXn2EwZVPztMMXPIrYrNzITSnt3OWfslXgG/uvqj7y89P1YvC6Fg64b0arLl90+q
gX8Ju2rwc2FVFUmzb9XogL1ToFtHdukmBGfJGxMUKv4vTQv/LlvXt2QBDlV0KuKA
BEtW/3IQ4SJn9jsjjOccHOWxdwv5hc6ZVdRLcFLPPsho7pITb0CbjQUmLzQMdePi
5mbYpimQPlE4mLDmch0BQPm7bAvLZWV9FgWx0n7h+ZcmnV6iaFlXhtRVS5dug1pc
VX5o4R+27/Uel6u6WG1/ezHbs69swqtFSqm8+PpCmoH1IV1sGRjmu13WLZueyN6b
uvK5o+CLa7aJhPuXpIjPRT0JUJLe+zcMgon4pcmEqicb4px9SWF6yumgU1f35JR3
ukgafDQLPkj2phCshqvvg+brOGeJNE6gUJUCSE6zOd9jNjxwhUGcnKiMdLqQ7/S2
NWo547HBvmZnGx1PzcBE3YaHQf20oTAzwaEcf15viGNcPxLuFOx1nV6BP0hPfZPT
IlflirTuth0JLvPSAGV4rjT8BSm1AHTZep4p6qtkcEBmbziylxxGA2kMK9GU6jQI
ega1M1pe60kV+cI5pUygz7SpNK+QwtppCypaEhqtUdpdf+/M4jotsphc53LRIJCq
WI17YnWeSPvWVMhz67izfu4s5x+mFWFrMO4rqG7e6CbGTCjffQLCkIAGuH/RCL/B
fxUQoFvutm5lEpu62sHhU4dRB5wH2s6GFVMhgUglUZ4R4JpbGJGKO8MU0NPxN+6e
X6gygytCB+k0egB6xks5Yvhl4TNYjYkRjdSHHXI/RXSt5Zv6lE4ZH2MAIMiFz8s7
yHbMKc5Qk/QBKs4c0A85UyYD1JNMWGWtHLRzkp1lntnG4b3AcLG3U1WEp2ISj5/u
LI6RjBVFcXIgtq7zcx+2JKgbHEeLHwJBxFPXz5c6rJy8kQ1qyapsmE9UGIGNN9aX
cb+DAZkC1POaJJm7WTGH3GqktUh3JRrLjpYUlU2mn6WOZ/q8/ZkKw7tK1/lOeqeW
98Dypzgcqvrk7qAWMNGH4aQnLR0gSOddZEBfhBJQc6JcKGodLjdsxJmvoSADYXFf
FQNhWG9BKRKC5wllvBplzOdKRy+Lfus4ZcJgwU2K36LrtsjXIMpEL7fcpXVo9+qa
3vx/bDPXCV4G7KOSdmheJOM6r7ZhojQO34cYKRkLXYX7dfOlV8GbtvzeCZLQrfy4
A1C07YpHNtNsSIRdlV15W6OZOJrHlPgqJt7VPKEeqvlebIPXCTJMdlnNlpy/iYv4
3jVfmdVlWy2/5592vjytTcIb7c/hxxVmS4FzVDOBomlEGDAkYvF88oQwOSgHqISR
9aLAhV8bWyJm5Ybx2bnZinM2ReMHsjv7SaAi5+/B43r5XoatSVVoJPMEV5nIaHmt
cLSIgwN8gXhS4Yx4sEffilYFGCTfZ3dkss2z7+tn+/XLQfi55hc6MxAdXQVgUDyH
3KZkyYQz6aRtVak6NDWmmrU0t5F9byQ4Ai1ka9f0zX/GZXomtgc2Yg1yNEPxMlQd
bQc8uwdSwGtGRccLzgXd3eHXpNJ0CiSHt0W6+r1shtTVdXfWZqNNzNHUtr3A5UY+
Cgue/rcAonAZybXeTGpdDEQ4uGgljpzzicrainc/Y4H4itpWGQEl5Y5h+nF3DPpG
rXUFN7OfAxCKNOTZRvxSzRm8GkeSq7ZWb/HyOUygTPdSaAMSfAVogIMW+F8mnrAO
lsTclWaNTCzh5TMcssJXq9UUJEseBjKomH4in6e6eoRSGbV1qYJRekDhC1aIV2DM
5OgBBkQtJSlzDfRZSrZ5JHHeBq5bFoQF8efmRaEfd3pBM/0cqgzYuLQPX9La2RHM
V8VEGVeLD+/NNQTZPHVYA45XA80gSmWDfcWPb1SDA/Cqb/jzjAvtHuvhvRasLd15
N0lgBkq5IAVa/H5CzJd49WxVibOaMX3K18YTLvfRRnl01iqpKjGZ2rZ1QxSRqE8r
ga2BZa5jZ7aEQZ9vbtCQqP5tx0ccNzPPqI4kQfHnIpgYKrt7+uS4CNVpwy9saPs9
2xd9/jqd7UYoy3SQk3BxGTk8EXZ8nOBbbAMRRMpmLTV/56Xc8JvtC08xNKjDVnid
/PE/JJbtDyj8zYqyVqrQZt6gVJ+iwn+ebY/OdbeEiT0PflAzIfCME9HnEs08gWK0
F+PvvnTJYPyH7rMRPSQH09wrbDragBSMlaX6mqcatxqOAHtNfYKZ55SiOJ7UVuSC
Ct8+5s2U0AKO34CjNML4C1m66Qld7eBOTzYLJo4cteCIDMi3cEd1RyUtCt7Kk1yb
TXGEN+O7dmu0XxntFIXYmkusc8s4BtlLZa3q2yhyyB4h0pEuxPmuIxCjuQMA1nRb
AEEKu9uhsxPSOGuussdxlG25XU95SjFb/6iXQmzUIhZgcbZp2bRZUJElVdhDLNfJ
2FmjRrzF2z7ZTZskmM6dDDOnRmjtGE8/WAHZW8Dvd2Feq/aOp7jphgFUWZS0CnA5
7i8kVPLQiaS9/iuFS5RzsDO9Z9ZX8EsGQV+T1qHrHfdtZny/kY58o37P/q3kHdVF
qS+5u63EeGkqgXg16ysJx3+BxB2Hm2oUKkYLtoYkO0L2YEvRGm+S9avKO2Ndo0NT
1CFWVmaq0dRZ76lDXjd19WFKSIijqQQArRtKbBcm/leLConXt4AW6ZcDaqZry3Ba
H6wXSoYetsDVfklaJhMBkwWIonSO9WsYzAhU382lAxCgZzB5XgUOYdDu1E7/xX7I
R6ksZd2hPFQn0jQCKfcnZG0KleND1sfa82Oz+bpXZBpwpUG8dUe6g7H0Gfp8SAeF
n7gsTiCgGurq/U3vLQQIQ06quSOMZ1RjfDyVSjgy/U9r9kCdSRulN9X4gXLtKnZB
HClQbu/beQ0EWYtjOMuDhLXjCGCVdh6rGPDdP/oFxOnJaSDJjL9fDTzub1SGbJ0/
dx1+oos5lMtqse4vxlvlW4+AkmV0ozZqehnQaIdZCHTlg0QPGMgqlMU/eEVNzrJ1
qgW01ETeILqbntCD5mk2H23kvN0yciZJFnfFlsDFRP/AV3qgIa/PCRfC+Ura9c29
px0yMj87kq7EHbChAebQojXNbeHrevs588v84mTrdwp8N9BC5AbA+8zYURKedbtI
2JqNb1/kXoDPwGFnFAJRtKXxcyQ6jD7rzVpn4SpL8dTqwFA3udYOP+/s9RMbUrhf
MwnubtyBXquGxBJbWfShvE644HoucwKx7PqE32eGZqH3q14ipuxfjqv6nF27rYS2
4uZ3LSnE2TOL/FhyuUWT+cFHGs107tNZi6uDLdTjG215Ntwy7/StISbbK721WhPU
90Z96HoicTZVwJ4Bzmjqyip6qsVrL2JpibMP8RNYNROgZ9Xzh+X+4tnB3RnNaKaU
ZYrAWaWhDhp9ykNZP9m02vvKuMBYA9WGXU/2tD5A5Ki75wz8wCesCyoNLdzC992H
/66sXIc/CU4MetJf5rlVxPi9bM1R4TlRNpJmCHpqZkDNixGnKSsiXT7n0pO0AydY
JftD78jtKkdcBUO7AZ+Hm9hQ0HpI2LlnISmNySWqlAthYDca+mOK7ElXJ6LIDKL2
3TXLsTjWJ6vFU9yWJZj9egIRiYX7GxwYQAisATzu6oPlCAXtt/G/GtDsSgKBQR5p
cRxbq52euegfx17wpLl0TBvCIvO6vllM8e7eL1HI1Z3//KhlN+uJiXkmv3w5hSqc
c2bbDVf8+5i/fAMFdAfmmk2YMTxEjp2ebS8jib53hGVxTEOlL/zdxbSQ8oyvPt9/
VV9IiKBi5P2ZKIKvmntAonyIRJ8O3R65HxiiYRrlt+7TvPXy696A4/NoX2l4GepU
ogy+mssAJ7Km/b9oCwoHTpZXkO7FIOLYo1gBsiv/uvaGCN/l4hmhKv7cXOs33Qd7
1h0jxaGrK21TSSv7X3a+72d4rHgTTB4TAzSeqWqKjdoMz7l3UfzFhrqHDm06Tl53
sAIIrs4Zgw8JztC63Xk17QaE8Bg5iJ9e9yA+8nzZT1TJ0mHqO/K4eumattLbolqT
uQU9+N3sX5vpqzZHL8hp2LCflWyTmO/IJdOAMJnQz5GkgoPqZsHk4SUo+Ev8ufUI
VM+/ZXsWQknYiWyqJd5SS6k3FTVxHZ9t5JXZ6wp+2srCNJET34zRM1OZkWfHeH35
iQqxP+MeisUwYmUzppz6UdCQNLRh9OX5I14m+iPKsMsosi/S+rP++JORyUO1sIj0
Q9FWqAhO9ePat4VTrHoABvTF6bUUUU007yZnxzJJa+VH9Uk8ivHJm7MbiKkW9PML
I3gcaMuTmx3dMcfBGm3Iu+px6nb/5MjLwjCOrqPK8yr8ftBOpcHv0afRPOhJqj4G
ABdiqcyKHjasdoJ5Nk/ED8xo47ykkpB7g1Kx3Akq/wkOnzeIUi7wkObid/XX79uA
9lMZpvLCu0LMF8y9oKtynMhFbPo3bAz1P9T1rcvCLbKhaPbjGQbTb5dJTTCeQjXn
alsdyn8w6u2vPCmE2+by/DKfx3mHtb/2EPWtDswVuHvCwKuaxeo8eOwTYlfMMaem
ZUEjWEuGx5rw9f9E4SdMQPX5w3/uYxtk6LIDV5GezaOyJNJPRJR03LYVI1Qeilbj
sJbkXNe2DHc+5dd3d+q2KrvZxUSfFwKuj9sSO+7Im/3Xekzp6alTDYR0h1qpzMbj
maJuIu0Z1+1PfGyMa71emQyHI0Li3fsKQh0Y9gDXgA9QJgLtoRBKl9UXH6kHgaw3
XhfIfXhRK0NkvVMuqd+qw17JcWGuYVerzXAzDzNGC4CLguiqv7NcDjbQqmv0zKx9
lLKztOCM+Fcirb9GMWUZy5Yf/yVytexFn6gau2rC8UB1ZHKKW5f7HtSWzI8oYwOH
/AetzZgK/2o9u/Yuxcz/xzLx/j+o8dY/QuFkJ49WMAbKtzUtihzFlMmZaCGB16Hg
tiZX6kWHLqM6c7YOjvPeXUpAciBQEqayUXiL/TYut0cU2yvi6KGZRx95pYasWAtM
CIBiux0pv8Kwyqz58JeCcAbXdvXXDZ7d5F4mMfKfssroZcyC4mZ5PEwcWdhiaVex
TVRIOURFbqb65u3fyGc+uqtQbrrLjODGg2ym3CSqPHvm/0n0HlufZw15kpD5a1fY
5Tp0mlXqHh0aUUmqhoDroc6TIawjBB2EMIpoBh0aQeA5+zfd+qdhTUn5PFDwsTO6
SwzGjI7I4KuX+LCmnaY2aR2l7XsCpei+mJjGmGalK4x37ZqBvcp7YkSIzlL/j/S5
ysRuF2jKCSDoMlvrZ3OUdsXs8Z5JUKXM3sa4eEGz8nosSc8KoDF9JUD2D27Y7dAT
G+Y/03x/goz/rMrk4r1rrclnqD99dy+rAEKhaLheoDiNoyKRCjWLphskdyEFDrr3
WghSgYN0XpO7Vpgm6suKwNXhLfglPXeWo0PYpU7nh3K4NGDXB5UOvmTdtwn/FUFt
UiXtTpNPyxzkXpNjhJWq+c4Ayl/7Odu+mMKGzN0bVL2MVWBso+Ea8cBxuT7kxi46
1OqBw57DzOm+dnWP/TtfFVAyd2XEx3PVC8ssgubyhA82gqQHJcL1V35WROV9MlGM
5aDZXEkaO2wbrByYJBP6taCjKzCUGuC2MwspKQcJmgrVgiCHQj4bjW8uRG41n4Vd
kS+no73Hm7PD4KATVNp//DgC4Fz1CsNIKzvoDvzI2mobwGWWyT5lsw+XUdqtlUNd
PQNwnVo+VVbxYLtMTOeAtONlC3AfM6uYaCruPvplA1Hm9nQjEP5zeaugGDxF1UX/
K9Uc5p19k007VQ2MFvhSiafDhZha0qOU1UEhAe9LC7UjFEXTXFyrm01WYJWDqfVk
u8k1WIzvzN/MD4i4SWR0Jamf/Hv1DU8wjmUYxxwTEtITK9pxqa35ZJ0t4ADqMfLS
rW6dKPKIhsK+SBMCjrY2BZk0r/1/WorB+0PvxlaaMiA1acG64aSsuXmEGg25GbNC
DFEAQdu/UZNH9o8X4S032crWqo+ZW+V5cn/pjXOTbNnJiSqiB74o5AbBT8/VAHkS
UFRbkTuSoJSiGlQxZXVj3Js5UL6yRO6wLDQ0MAvP4sVtO9UEidB5Oh252qS4E464
Ie4m775i4xwYktGQzNtee05gY/BM4tzn6eR5svcCGhUoPZsQq1N0RvRKZ3JWoQqU
NOlUkIFkiy0peFt4B2BOSJrZC8pVGpFujhy2pNs0fPGTrp9Kr8r1YLHFBbF97s0c
16w+f8zb6jI21R8Ws7oOdb0Zs5yME+YQm76EIjOmvacqL2QvB6XWgiUO7r18PX2K
0944k0/MeKU9hSL1GmjqJXPgHbV3+4XklE0fsO0qeAwmGrCj/IgiQ0nky6H/N+c7
K5EskAEM2TMd8dmB2HCIKIeqtdeS69HYyvZn50D11PdeCbinvy9IbpMLf+HXG7iU
M0Yo7Ua6Dn7V8pCUiiV1c49bi3ouoy+iBCCjsLVUt0K1QJIM+ZKbxYcj0ZpTH4jY
fuTjF5nuY03ekxczR+1+A3XqP0rxm4NWipZMTt/N7Mof3DpMICcIB14vQ0AX6Iqy
P2xAYNmFsJr3qXyUg475odY0SzqJbEbmx+yHvSPPZ7WI08usOc6iBc/gOiScD8do
5cGbL7fql8z/GZ+5FL4byPsCUafncV5STj2o1Y99NTaQOVyZQyMlBkrZBgBKK4pe
9dvxQ28z4u4IRK/NVMEOaRJtmLzLwJaRypggDLqrmRIVXg187AZ6gWcAQ3JcjufM
eVC5scgsLSLzoXh7Pl+1wSpoXIw9iQHecoX/eGsyXrfoci6ZcHF29Nal8MTsgJnC
DMU/5jOCvFATEWzB08XByLz88n7NF/iWXvsO6ZXuiQo0BzrLor9YE7Lg4qBuZOrd
5bHc6KOJ17gsugcty2c8tstHcFj3ulDs576AJ7i8b+rUeHDMKAxw8/9aE2+TEU2f
uZkvNvvdyZGg3VoEuSEkHEUKCadVbJ5iSAZyWfYYVe16tj2uUtFPGGzQwEIdZsGI
A1Bi78dIVqeMgHgWPSkG+1HbiA77A05xd7IFYOuLpH0tiSOKEj6k996lLr9hRUtb
ckwVQNaWvmMwgmnPtSlgsLH0dNuuQaR7suvnoBqVceKb+aLfB0/ILgjulw/7z2g9
K24n5DXksfRfiG1HxfQEnJgWKLhQnMB+KEd++WFRLe2/Rjgfsqgztoh5Dg9HZAUB
nGPwbqbsFfDvk7jMv0e3OX+Sc4Zfubndol8keriM8+1vUNB1w7PAchzmM2XaVm81
0DK596KaDgsD/2YFC9u5IhEXhOXxZbsiCZPt1hJQ4jfWFxlZmbRYBjBbpR43HO2H
cz1GWPL0XVzgNTV7SBXYfvLCVWi85F1+MceN7IMmMxGDo63Hlqx7nRTYtfwJUZ7x
gsu7QCXIH7G54Ydiws1cDjYKOBWteN1AWP3dlPm9wpzdf72+HFXHVDMANjh5ZRkF
LC40ubpWyRxxPIo3lUuYuYNpdOmI8SRYdQuTcnlXgxmZlzlhE3AV9I01Y8kBbFs8
cfnk7/ZNcgoUphYioPc5RhxUMctxTwuV8gvaBrTxsZvVM128y+Kr5oImqhqIIvG6
hgTVsaAJ0Z+Fe4bG8i875EHkNHP3TeheB82tNnx6nC+ocv98QypYskOtsUujVo7r
bfrjfPWFhxQynfvz+tWzBTRTGaxWhgNGMgTTCLI9U2y13b3DqUXcQX/iHdMkfxgl
1c0v6I5lUT0CO88GZQ1NjfEA4boDypicH6K1St810U7A7WJwK9hI+2eV74G8AQaI
/EpGVQWVf++CJ/bzzm1XDjR9KIEMPOW63z/LjK1rK5dVA7HcGKD8xVLkqWX6m34i
2SNf6ua6DtOUY4OxmmZzAfQizEGFf3LJiYEjW3Hp/0scE61k0iBEfj5nWKqa4knC
BPgRrHfvssbwmAYn/7Y1qR+tIV8Y9ufobcZXxsYcE/ffrY+qRD6mPmd9Vd2CUdLr
Kt8zQute0zeF+1NGh0hk3XlYq0NY/tkSzSthHGlNMpBcir6N8ePBLXVMfV1c+awH
2AlamnofGCFfDO3cLVn1ArYEU5W+wUDDmR8mx6Diz/tV1zoIS6kjpd+ip33CIW2y
5j0n/cVHmbWzN1JLeHnvzdY1lbiv2U09NqSziteXq9NvcIucnrqhQhcUhzBZA0nu
0cwvwac+Fq7FLpTTTVlnciX3D2WyaFZiEkhe9MPCqWGwLp8FRlW10vljuePp52dV
M03oxaBPafv+xdQo004g0LuUhGfzzfPJK7e5jVrvqPnSVlem9vuFXFg9Vrhay/hS
/+QPNeEMTCLDIgvUxQScULr2GJbYxQXSrBacMQJLw3BFG8ty2/t1TzBfzanW8dbv
rYHoKbAJvqfW2y5TTmqJs3S4f8/ptSYPmaY2KY/tUEzFg5xfI/JwNsoNJRD4g6QG
xm+LEJaXawyrIxWoUfE4mQh62o3l+xQZgha/RSARNCDdls9gcAQ/jW2T8jWJEfU2
UMSHlevGNAUl0XCtUPll2gy0OT1KQlKx0w9BAlVtgkqGZVzcJWcomnOvn/Ajt06l
peYYQ4ZafAvk04ZuCXLQlx1EQamrzMJeF8uR26VIkeGbibBOx4k275lZsDRthT37
KDUv6sE1JLRrq/4+ug7smZKwEl4l6o+Bzvawsk6jqehMtEzVXJp9exhXIPGsPeUo
rk+bM1Mi5XMqx86S6J1TJRSxvnYCDDCy5yPh2WDY1yeBkZhxYylfL2aUxa65sO5M
LT7eIM3MU28m0EJ6esrzNWdawf9msgy0lnVCwVoF9/mO8b4Ys2jXRhPdcZXJqz2V
zczTktuk8kLDAJGylVOUNKEL2lVyTPDL8Sckbq8Ufd+DTh/0RYTLHnOvVw/2MhAY
xxtMUzBsVgejkZkS6MMQGiz+P5vL9kNL+tS/dCqIMkoUtDaTEEfwd1rnY/gBrAdm
uREbyiK1v+thnA9TMF/a2Zyq4UzV36T+BJ1qK/7kj3YqzLGTItHKMqqFyP3sReAl
ocCB7DMa73qwj5UwscEGrsJ5HZbilKtrGFLYiBcT2lKWfF5Pf+FNZ7GAjkYLhiEw
rLvvyGEHX6utsOgnpawK0dYwz+7unJYHvG0AK8wLcSiM/QkE9/quEkN7yLtCFmrr
MsFG6Fqbpfd5m/A54/vcILYjf3WuTK6ObgOa7uCriOXgtUYG9zt89qrUcO4yHupC
BWbldiQ+qomQtKNf1I1s5d+9SP82icd9fSyaQ2wt6yJlt+SVuByX9ysOywrddQVF
ArxTHfWEjWUHdbLUMVPAJUTu5jcJ35ye3xYgbKXneb4u0iBI6tqvopadGniXzBjj
PualCa0lSPKerJSbsfgcfYpod9arKiBw6yLo5sq0i8BdJujEoiIa6CLoQObnoVyV
0mlQVlL5zaRIbjoDOkK20GIqLmzA1wl2n8isXADE9ZJmLV3jBxE828Tlpbb/r7Zm
1Frg6phDMJwFR9dzsXqY5BN8Zn0uPUYaBcB6n79rRW39g9iBVP/q8yKwgpH3tqGv
QmXeXKEjbEhJIa992bMaQxwQRPW1AeeOKqWBx2ma28SU+d5Z5GUm6kJi3aph8oPS
1r8KiBr9HzyLMobyV4YjJ9mWFbUKQsdaU2S8EEMRSqf+rfj5Zp6fos58kmIoIDeX
HjCmPxNJAzTG6YHpYCfcZ3pAfuRmr5EW8lhAnCAGI95dOWubQTP9bjNpwEwSdwjZ
uLkK/smLCPpzY28N3aEC1L/earjGR/+icHgVZJr/FdurFfYXc3oV9xSsIF5pMNTp
54Xws5cO1NXoTvvq+I5wkW57gQLPt0Jg54Uth4gXB+oxhEj6B6yGRAVqIHQuzLf3
xX2ynW3VeqKq6GuCfNto3HCimpmpHQ5j+yz16BG/d+YZTssO4ZnxsgSQ53Le+3E+
tCCbxraEJn2BtjSlJ/zEPWNZYtnVMB28TdFvR0lWI/GprTgUqL/a7GbUf9QFZTfl
BQVQspAGpaz2/+FZ4Xxo3a2A5Qg+DT5lAm2g3PuR1uE37KIiI/UMBsQsRq+LGzpB
+2H+riVuozNI1+KfhFK/yew1O2nmsg4DuPRFNRjsgcINBgNq3W9U4E7RAw2r95fD
Y05Cu17wubyaIYqSY8NvFbLOLbizODKFuvQq1yjdV6dLSP2pzXYBuQFYjlecCTVl
xHIhw/Npb1h2a6zKPC8oIQYMxl7Ozy/RurlxLaSrLqgydwORJNXF6BgISUmLYgr6
CVprqG5xtkX1AIdWiOZsvHYTeUlv4Cn3GO9OR1nKdHjiI+QzDrm5zw10DYbCm5DV
nPeHiBPuMvkdJmLLsiAR8ZKGUGR7KkzZf2m4duEkM6aKlEhSW7sxy8aqUeoY7YrO
PWJLmrcLVRWF37Doj8hGSkjf6CgGZCcLIHIiDYUrZ9j8IJx1tsCPTvJpykmTQEM8
yKjRiLy59mdc0u+Rm9UDPS3pyADauSMDVqzeubPrP9VUuO6Y+4LhGPzZ3NVphG/7
RSJf/Duxi1C6jfDu8m9sshp05a+tQrrkA8q7wrGF0/iABVN74hdBMyDVkq32jez0
62ZAL8oVtp7unIP9mLEsLfFas5vj8/WEEb5wulFSFb+2P3Mrkq5G9LTnxHDKbIZx
3N1Tnq01UfM4ACJS3ALEXpuBeNhsEzEisSAJE0pkUsi8fNL/mZEt3B4jiNC6qIGI
IVh0Hw9lYYxVyp0+wv/vWsQqFyaCqmWCh03F5tmUKayswR6qTJp4XIrL6DsBGAY2
5zfOHwwAHbmjs9X9w6H5vAgsmhTpCpo2j6gMgZIxmzWJm/QLW6TJhX4m6y6UD8jP
puNoY2/o7LkIJ8fgQ2A2g32gv4/SnTZY1FdyBqePyFphaQDUvoDxJUvtIOd6BWpW
ZvpfxWmZgEZ0BCbWTBccB+98dbDVChyc4iFiOva4bOvcmHqZpqELxbf2JDanUe3D
lmFGKFge+kcYG2nRj8Qdj4po+L9TYIQHPWNqDeZa3NeGlC+6mySvpzg9RJcMvpd+
BCEeTP7GbzgK707Xf92cHWKVWFfCJ1oDLnedvFYClctd4hrjxUxExQmmp07sSGdb
RPgrgUGuouNQZk55pUKAHnbf5Lyccu+hUsOk/f6oL88Oiv9XZ1tVx6sDJv87jBy/
6qGcIPJ8cMOXPl3z2Kx/i5lzpjtMDk4m3JhxbXe7Db5OKKG0/PMYeAoo2xXqapcz
/QcjmWu+iBQ88q2sVD60urnypzKBJutGjukEtaFFxZvW8KpRV2jFeYC/K0Elrzjq
oaryh4DLg7XoIB3lym1LUS0dcmPnbkf/tRujssVJf0VPw4BW4cEP+UfnJjt1l6Lw
okH2wIgDf+Ou8aIYdQzH1xsrJEdcesXwi99eQSccoa4QJdlzLwtwo0Xvp6VyY+R0
jMZyE0Tzv6+rWx2fE6/+z5HDmC5P6irKUfd3GoLagDigYb59QJNJXA0AsFxI0FDS
OKj9AKnGeCbsc0fGtZjFUk9Uy0ZqvA/DQY3Irv7iZNQe9XiTWIDeVTCdgt5IXDIc
naN+bYjEzhia0UoOU5n7ekmP1IsyCfylu3L6vQheZn9k1YhJ3CwOfj9/YJcrWDqe
7S+ZHekj00U8E2xBz06yyG/kEtKtN0SzTUTwdYZpuYWgpuVpnOvYy/9OIlNjhStY
kdbaGj3PtlvFKutA0mccpRu4qExWhCzuRByxE9KLq0hRx991UT2mVJkc551fEDZr
z3+JZZHEipBglzBHUSuCjG4wektGyq0SuZV9dfrcCZNzjZOrgMEaGVB5qvCG1UPz
Jfh63VKwt5/jsH7UC4uXlpgrsBqGpigv3eOYnCg9Ex5z8j4eu6DU1yB6guZV7f/I
ClIxwIzyY8hQ/pYiGVzCJQcwhAA08BPpq8u4TrFyg4QD8TpmaQx2uzl3SH9EgVv4
lqF6TXMNh/HHefkiXa4nvgh8q4jQioXpaGwPvY2XzocLSEpnuVDEMWWAmkqah6hs
K9NdrQcJMoQJVc7bO8eY1p4gH7PStd0zVqYQkaYsrU2/2WseO5/iR9I2RXn8nVpM
tS2IuVZf7Sk3zUnGvj1FiBV4L3MU46SH1iMgM9SO2w6Lsyq0nwrMhE3IBCD+RH0L
gArYR/pr4oTKehhi9RLJWwSwDuqXYoQSVW2+mPxXPaW7+VjIKz8gg3nLyuuUi43J
BQw3TTQmYca8YSzGX7FzJmTx8Fewx3AqWfo34cZEHvfStIELG10GE2BzX2IcdACZ
cyx8SJzyka5hCiZeyxOGOuEhTOcMYmEx3xp2nlj3CkJNl2Frv+jTWX3xOZhQ0HvP
QxA6ywBPHqWyG/+edcb34CUU0PVotFo3nCHC2+otdddZmriZp/EqxbbKjBsWdbir
qfPEdWVNr//EnAdwNkLY4jciLQ5Ai+E+JliUCfGoFQyj2puDYUXJj/COW9Tx95HK
t3WbbJz8bI2mJF8KQJJhnzSA0BofDu8Aast3Rk5BlDwPAf8yh3mfSVfTBWv6OB7o
clKxRiKP6G6xmOVuKrLJVIfWkfB5k7AAZkIcSwVGitLmDBFlR77lB+USTBpeT19t
jpzFiBv7d2zxmGfdJIqJj0dQz3vjF11IxcN0Fvr2rhOVqooft8q4C5RSA43drWQF
MGTRMQsLfqfGAbnURMEiFWl5bOYHGRiO11dJwqLbETJn66gfFq9RLo7Ocv8FyutN
B/JTMq3f8P+lNGuo2z/5FXCnmEajEanMA6Q1vUgX+VE9/Iq/bGJqIGg8mN4B1Ucw
Bj5B7ldB6h//cAVr3OiJGwOgPDoJjLl045Em+S+//iycF+IYhR3Qzm2JmM/uA6lw
2fbvUvEfVhCn08zyfkqot4/wu2X0tSeUYH3UnUs64wMB1ViBCCVSmbyqY841GHyf
gAWT+jFGBhbeoEvmvPV5ABp66VJ2cgmniDpigdQOP32kHeivuBGOyDAmZP6rAT3b
S+A8sBj8mxOBBMWIC6kdmjwAMY0dXPak+bCt/sJGIRFvfuqndmR0gPK6wwA18zO3
nkQ5WDeIcOlaHTyXBlf2ChTDpADcXi4AebZPb5K/bmT9W/uQrFEVK+8Nm/1Nc1D7
1dMOfEw5JdAQv7F8yq/BPKFDHMW7FfQPxwqu3UHlHsOcMwISd4b8E8TynfftboFJ
nqOGUwK+I4V99Dw8hpWHnPX/EtGSiu/hJYbJeTp3CE0c2V9cTt74Xz3Bks6Qx1SY
0TS64apDT3VaN5sZ4qzk1GfqONDLGXjr6dzcxy7Glm2TKznKH0tJdr33IlAfVWe+
lBh66UIfQe4WXrJ3WAs3YPiTXA1ZEvEwLwEqHxkkGW9XopzBTSrq8lM8VqybR3gW
jUiT6VTOqjZQLk06pEdPpxMHrTS5WgfVqYVRSijHSGkXfB1W5ej4oOX5/N9PMdKp
ewN+Uih2P4XNPlhVsvCuohHmhzsb7Ktn3ADzxtty2VYGFQ/lrUNHLFtsFgp0cKK0
OObAVqwwONOYoZ6NW+nO0+wZuWuzUe2ouY79Ka6ruEKWCPlPJqOGw3KbJU3pPXwD
RemkMTLrW984VhjH4WNoM4kuFH3TzarVQyBul29O6PMI3vwcdcELKj+TI89mN18G
AGjc5nK2jvUzlcT0Ej5nOklV7QmsH33qrUiKcOd2ErZfP39z5bQpOdhIQ78diMT7
4mDOvQOaoUcpsL4vOHbYL5fxlipN1VVj+VAdM8dj1HNrjsov2BFfbIP3cELUES6K
mizhaYZXqfhHSBTjkBmbbZTw8LykHWx+78y+SFl97dh3y43oMpQlTBhWo4PfQrQ5
HsTw3cIagQUPsu91AGKFhYYzwzv8mH+zetOIFU/vW5ZR0fBehHY8LIDHWmMMj1ty
gPL0MgvJ6PVYSVUTpFxK/x5pmv+TasmErmhaPA7Wa1dXwt9VkiGOjLo0XT8SX2Ps
dAz892hQmpxpAL2fyDgULfxmW9o2Kx30M/oBG9gsoZBnM8ywcqpHVBHslWfrwp6p
Jk55wTrG+j5ioFFb1Oc7hIgkCefW1Wm8zv02FbJySe5UnkxyO8f7sMKyyB1sOJ9l
TRNs60F2Y68ythwdHS4kIiVofHkGSNHnowMCU5sHVcU3u0Wmy+lj+VM9j7JxHMlw
HHL6KwtXckJo08XfOSULoEjzIHGHmoz4MhAxDJjB34DveJhdrBNATM2tzsCuJvIR
nYZF7jBm9rahWFWrtyoEysbEq4JvZxoUEgQ+ZD5ZJ3XiKgtCVCa7FMCDeZJvqdDV
EvdxbfIkICzlyqHfhKgKY9dX1JDvaaq++jrod2kwE/L+mgMYchrrEJEjYjJDfUup
KdwQRq58KZ5X/LvP/y2hC0L8cOMcjWKMDFRuGwwN4LLQY4F5MkMdoiYh3QFCwnYi
NrwLfsmnltDteCfzWpBxBWDhlZrI9CiPKmuna/LoXCayid7aU7ElKkbopDecIcyt
F18hb+vyqg0uzMMdIO9UxqeXQALJfXlQsIDGjE1ZfXQ9QPCNCq0RXAmKkw4eband
9HUs9Z8OYcgm7kEb7L6O5ILCE6ufmSA7v5Zy0DNzY8POYirWd2eQTgui0PzoFPcQ
zzGsgRzPsCLFoAnwUQfITsdU9MMdHTaXObzv4etwPM6clM66i5GZX5Vzyj1BiRmW
sxAdYb7rXMo2sgiLtZGeYaUZiE9B3BmBF4IikfpNMPn89/Bp4nCBWeDe/3XntpAJ
9t1ClbsXb4S9FgkASkH1/2ev8zKGA02aKcWzFY0UCetufazStkIuU+pZSKL45yrR
JStpZ4INyuP8lf1UsOchtPSW5jk52xRUGt+J1oih+/N5qt3JOShH28hkctIpDcPD
M6vyzTsHUtHW44G0xUyU0V1kN2DrNEk62aKqFJJiC0HTTL5jcfN36NCEH/xjZ4P+
wNMVVV79mBVThW5+Z4w6Ej7JFAZjOZAETv4dvbr4PfgzRuDenO0+uYYhynMHtnyN
KndLukwSDz8BG8ZrGuEeuSoJEfzK/rUbZgWvpMo8ZfbjhQ7TgrVlsujqR6aj9Vek
O68xg6VCCIkY5hNr94WDo7A4kY3jTRBVV+0IEhHZZkkvdq65GIRpwY0pn9yuaKeI
Q3boAyMYRuwB10Hi+aVTwzjhPQPaN1Ynjq73kSI+5ahyrt9T+gaN3AqeFRfYTSSb
j6qNlhMfRNg7G8UFjMvZkZQIEtploYtv0FZV5zqUxZXWRPZzslxg3qBE1ZkW0ohJ
yQTwv+GwSqfyqnC1bNpLcOgGDnxyKEAdCZ8fz1YNZtBhgMB5+h2Eb6/0RF+yr69D
zI1SO4HO2OEmtm55K99wrt9a7TfysLXjuWVPE7jJhJ7LRNJDmyJJoHRAmiY1q/ud
DOdu/CeNC++t44L72hCIeA9zqSzMLGN6jYafsETKPczgsmdgSbRIiK9IzxlOgX3b
g6C+Y4P0Q1nO2FerpoYKSK3vkS8LbeRxXdzYAEhhU/kyrlOzYDwUvsQD41vQNhfr
y4AlPjixqEmeHHepAz2AhxgIJ/ddXjnpiggwdaw4JtdZvDDrOJE8I/UmxqSEf/nG
w0jX0yXn9ULN5xQnlvSwUWh+J0OS/cSvkU16nHSVtIb8YMUYskrI1U4KDZb/NxB0
WpQGVEfhtozMN9Z9SWeCmsG3Tkn82bzOe1dUbVJlrWNxhgjEWhwX42mdPe3d4jo6
c02cwa9CPcI2sehHDxesaXZWjcj7xo0AFvvhrGlWx9H/OBNsZE3OUZZO7wpfJ7Yc
SWGZMspB8K/tlxPXPVdE012EUetyYL0pzp28aSI2//taTgNFJRjpl3Luf6Mlq62k
FOe/Tk/YJghX/YVCiuGIeXsHzQnEdZqspSEpm1Xmh1JEu5ZKYe/7cCw674db6aG2
kAHomXFB3tqiepQ383D3LDkePqqlff5hXhghtWUAP/kdN7VnJwDVh7Bp736lfM6u
uZINhALcNq5Whpm7Z5iyhqKL1cnU/zt8bd4aSm5N9oHMiTneLdOlFMOxkpEUsTE/
hImf0KtUL04OVWcpopsEzcZb0jWNgnieh/HORYHS+pXZ2LgrD5dkcEzRvXXCRkRO
rzh+H+yX9RADF/I807nAKC/fLvddbX0McvbmB+24COePOhJL5whcsGIMN0ejgUjE
5um06iWADN4OMsHlWx4vSMdebro9YWb0XREvJSHBKZ2xoQo7Tgw8ke6Z6Ce9jSZ8
UQr0NdkHSEegpb+w2s5VFN/+H8NHk1qGfO7OqgFBa2Oq81mWUvNMp0r2Mx7hYOYz
TDtKyUI2qOIab7lhc0CN0zcH5ItBUDvJMvLuIcrBqHNZ5XneFPc5PZ/fuauxo8K2
1mWBANZubGkcYUDW945ZrYLFe56HDIGfp1SP7nEp42LG00JQk37DpMVcM4CbZyZA
Iv4PxKfI4dR6t52UjUyUubbNwn5roDXW9iPJEzTjYIkNnNPlNrxX2txU0KRpycTR
6GMo1ENeVtH21BbyxjmtpFTGTbzAOoAcC+S7S30Dt5LIqbgZMtJdQacNMpEM1I2/
XD9csfD6WNalmvZN8F2D6UX4aaq32lfgw9M15GDjNtd4kZy8LDi+YrWQ/UCzbk/p
s+aKNCl9hsS0++QvcmFjaQ==
`pragma protect end_protected

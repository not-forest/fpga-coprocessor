// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
U5BsuL0/EcPk/1FlJQLedOkF8aUKXK9INDyrsLdWHxdhf8Rf3oCKpUmDa394Do6t10IFj5sBUipi
duuLqtZqABDAL5FPUjB0ifRXy+z6+Znp5HE4pv4rk9Fno83k0aYRDBPfIjvKz8njpqX4WsOmDBAr
nQ9nd3n2Y3IEw6ZF3COHYWzNcRaSjkX7YCWXHWXt4CdOsUPsgTiBymeGcY4WJpUO6e0+GiNENfj1
xPA8lOQLuOFk/HwXJOeRle/E9EXnR6dREiZXWl+A70bk6UpVnEgoYUH9ipTbcAEna2uBe2kdka+g
i719K/seNxvFaxJdLOuut7epufw1c4u7Q3F8Zw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 9216)
QEPijhLwW9WAttohO1/tztFdLwGa4n5Jh8xVwDpjbc2TqgiyMH87Yr7ZHGXMxb3gTjBuJ2304Wtd
rTYUY7+0UPJ/FsLz2CkxRL4yw5mNjCnmqjeeETw+x+iHz5sQ42ZRf0uZz1u3bf6D9IUZhWUcSGNa
BfiY1KcMQ55DJSl62s1HDEhdaAXMGdOkaLMpKgdQ/xL9TD5P6y2kCt8lqzzmOYvbHEQyjsMJPmDR
2u6HEmnuL2hKpU2/lucMyB8sE/ZMhs2CcCDE8+Q0VqX8iFxhhwNjS4tXLZ+JBmWFhhcamK3cnzVu
lJYQTFD7hVhY5QsYSbVPhtBnNJs4+BaCa0FCSquvtByOi2Yrr3nWgZxictw0VIEpCVXNW4WoeVwi
vjlXJTmrLuGhkOG7Sz/KuY7EW3CzBT86jxE42on4tj5V6+XbDfJBt9syr9VXNkE0b050f2Vi0XTG
3QEsD09imiJYQ+Hr4GiAmKR7UaaJ1HjCM3aLfK3CF6XV6sd7P9iC0bdLk6QtU6IZtUKiGvcI69Iv
HugpdX2Dq9CPz6sQjWfWwf1V+xZdWxZlrJee3szpWHWweA9HJjGRbS3YAvVMAh9j3fcGm0KixtnO
PVYiqfLqKjZ5FSSOLcIgPH1iDBTXlxofXIvKP5g6i2TwE6OcTEE11dJ8Ia2pnbr/cK6qn9n4lVwM
hp/mY2m/HW5zYlq4pDXwMnMgrHjOkHrWk0DzklK21jxw/NA38DgtNmVDkGyeDOq02Oz/oMonEphW
CVw+E/JQ6AH46dTBff+/ard5YA5JO3Uj7a6mG7pGurXkclv2xOe3hXEgx5i1XLouMf6fGDHr8N73
l7AABEVq2EUYN9aq2uxVXvyCdqiwfuMJevsr1B0IkHrOqX5veXYuoqchDkpIyRtNJ2CcQvp36B+y
LsywoOo5SW0EXvNYYsEeAJrFIHwpHwvahrLzScAYReyNa2eZjdqJYbV5qbb1DzG6CA/33uIP6H16
3APESkJoAqAuf2ZMoO/s8rbzfUu7/2v1pNxSccpQ32aF9oqx+BLHvVyk/xWV9P1GLCrWEBWOT6yR
sd47ezj8LajYYnKgzpEYTapC+z0VKPXGtjamZcYm0MyAbjJKRoXXZ8xsikLWeCb/zVGAiPdFZ31H
Va16/HJOlQJto83XG6NCZa0b1rSII2dgV0r+J1ZdiLofqwXf/oifn6kZUJFqYD8P5xSjaNgxJpmB
rKEN0VXb59TFrUhGG0gQZmYjTKEXUrYdG3cvAhs0SpKlw7OtO4kV3WMISQK+nKJCYfC1VoN7Rzra
ObegSXOOONpZEdrqVzwkrfgLT1bPD4rQ9P2M/OjJLpqDQIpk0wyn8SpgzYSNuU6oyT1o3MrkqMny
Vr1Sg1u7LlB0Xe6plOCqFYIu39vRMX0CjLguQHJgsKSqDgRfksgtcfhzCZJ5d51yrMYAMPOiFwha
NYqjTcznpcZkVJ9gfmPrXhL9B956QwvRF0Sup0u1vZ8CNJmOjIs9ElTFED3tAVfRSdbNQ5uYvl3/
/yEDzwgrKdMnHAdhQd/vfkkBB1jpG8Umg3LaQ8bJswxWtXFpj63dW/Wvi0q/CYoy9++wzGhbeJdF
l0V9ehiCbyyqIXpW9UHTXGX9E8SPRXa0OfURs7jCxRWHiLNO4tbNhRoN4XzzEQFo+gHbnzP9dUw/
vUmxRL8y8fe3kev4e82O3PL2+o/tk5ez5y5Hr3hsfkjnJcuqGi004ycwRox0BmgHWxWftXjO0JEX
yHM1wGnLnrSQx0A5NyT4TqGa9+lqQMZutZ4r+k93kPuPcJJ2UyKbkCvjb0gbrCQcdzWBcI/Dv6lQ
m5E8baCqzR0oQZP4rJGTTXlYbZtHTLDIFTvOFinEf2hpdME3XioN2A3XrV1VC6a7dX/lObLjQwyA
TgbvCo1S2x0wEjv4X1cDsqvZaMHctET0MYuz1T3CXNZReZsuA/a8sMcAa3h+NvsbAkyEJZQzSUr0
lnrgkILiWMMSKg44exSMDWmcpFQuy+vn7pgJE1/HsRrTOtbSf00slpLomTdrz1blFYvn6uMYlZ3y
DRIDiB5WLiZ74hSaTt2cfAkdaq2nxjQQweFVin1fjw+9MKnm1RKChxCrUOjjn+7Br0+vNJlTgz7y
bGbz+6oc9hEOc3tEevKYkLhVxvyqUzrHDcx105dXeRUGWkQ0RD6aTAD175JV6ZlCLiAOm3l3mmBP
pmaJ5cFV9XgYAdu/7ZhUkduoeF7TQOx5hgS8tttsS1Rpy/g7V4QURrt0YdXTJCae1IyKBkFNjNJo
KBY1j+JlIBMl8/YC+X2asWENnCTKks6KyJEJ1uMUZhBGd6Aj91qlm0m9wlClnI6/MUOLUUdGlO37
nlE9RdPKj1f/1H8b5zIs4tVrFe7+N0LEqH76oUc52+17eB7aYeLjWTUCu+BeRiI6TtlsTRbMHVl5
tvGOiTZyen6IxUM9j0sAnk83PrHcHIAN6l1KGwtMe1vtAj1MAVerbIOBMWEEGhj5Tp9j+XgJtx9u
+j7xyyFIy7tN+UHnvY0jWZS3q85rq7xQwYT+Df4+U0vI720pv9AFVFBZ/UoazRCclRNoRbMyouOx
Zo1mgA9r80jyN8j9QRyZIPTky46Kp0l50MWVnNvs5YD759hCfEUTTbz75scNWHMbDybyiTDRnew9
1yM9hbVUEsyyC5BJeLtb3vXrTKOumjEhTyOVHra/27NkNn5k66Z9BQirn8On+ZHD+caP2Gkmi1Pu
thAGvQ+T57ve2mFtTu6+CJWSYhfChVvDRmWVllkbCO/KnPRMXPbAQxFaG1jVMbOtdI9/S2bvaPpj
RBUVQTVJz5DABSfC7F1a3KfXcwgkq3PpfzUV4vZR0W/oieL6tURXejNSoZW6bJpU8M9fYjt2FbSc
kyiU9eTXtO2edXIqPpV6AlQKsieaYuyxU4LkRvwT2X3eVR1s0mH0kcdvNwzs+xH24rrjOtZpFcSJ
gKt+rMhp1puGuwdJMZR3C+diitysWlNf8BLSQZj7J3Nkur1gtwSX2a+Rg5NVazx7e2sBDMcqcXwX
cQ8tmMhgoHhfqER9e/sA0wu6yIt0tueJvVk9C2SYzZhK0GQ9/es61dNzEqMJDwIyqQOZdNA/e6+r
tnItBinH1T+feB2BlTK+ghRa/Wfy8ZpAxhihDBjaalFsVrqiqPjhiWtxr9tatBywZWW59+B95trs
aWPd65JNOuEX7BAWp1scSqnuHUWH3a2ejW7H6eh2Qc1Nq0Q5LMIW/c+YbgFUbSqbe736vjzomf9f
xmv61iJYbj9rUyZ88h8xj+p9st0uaPyaYDLzYBYE1M6WAKfEH7AKi23DjxCzQctqZV753FzpLver
0FcGne9jK/Z9wh9QoYHjg5l56MRFdvYiNGFddkssfUbnc5iS7FwUZi/sRoOAcyuDcUnIgcD3OViR
zINDU5Y4L/k/5U5z/IJQ0kGL5NBpcIhOH6EwuMZGqChzYxXgNjM1XYr63AHUa2Zp7NwEAQlZ49K1
HoN84JImzYhCCtEeP9fek3z3/BwQct3gBP175XVqsEhNycBtyRkcBSnA0EizGw7L62f2tIq2wdGK
uNq7iHCAl5evosbq+GZm3TIn86WthLrfBsEhY3MytS7Z6AaY7n2j7xNjzFyniX0cnvnBMyYj82Yp
bDHzSWq6OlAlNFSc9GPHNN2SYaKQue2kDmyHdcje/aOrXPRs9FEwBSICrFHFIhBbvTMoCEDfwVXz
awB4r2ta6HtXAT8jrSWhtMWROj8MbdP6bvk/wqyfejL3J3vXQllX91tw6HweXANdi70C2naClFyI
tD6tojbSfr+IdxEGa+xw4+1/Cq6v//qz5YSjrqUkFndNVTGXKp9409emzQxMZ9TncSNqwJs/MBpM
uMu8OWdXqDIGOn7I8+1cL0Xbk8MgouhmmWyVwrJJ0OvXyu30L15Xi+fcJMA3e6bX6+PQVQSJKkXi
sU7xOZDErWc2auLOGSOr8MIRjEK7y7d0DgFvbLSDK+VPCAgJzdSscOyBPwx5z+Dm0kfzez24g3K0
A2xum97txUv/Xcc1HTSUIDPoumcGMEWqbnZJcv08rvawD6V0i3iUvFCd4F2G9ihqsY8y+bzKDhtV
DB6ATot5N73CpeGyThGCEuZNDWYNRSpSvkLLefpwd/kTooogUOwGPbM23cHsA+fs61eHSNOyTpM+
CYQ4aj/tldnnGlCd8KXI7qWqO/NvFUJeGA9gSn5fRSh9of7N4Q5EUW2sRDwmv2VFz3QMwmWFrKeU
W3rl4uFE55ae8tG53V9pW2azvMCUwIvIosUsPi29gH0PHxjsA/thaNBlvxg+DHqG9k/sBwL8IjCt
oCIEyiTFjQT6aMVBkfOwMlWCuZTTskbUqSHo6M+JAkigTEap0FHo3fZdngvB2UolHMsgQHLeOoPf
tbgjr6GGCsI6lVSQyjrq4RkxTpB9D3E4VoBs4ZBSdO/wgRVTG1B/y3N2SKj4/PSDW//sIQaqYKoT
xotf5hapoZmfh1zgknZ5hTSCMbe7H8nWrrpIbyr2OK8Jdi4Wh/pa1LRVKf+UCi0xrxA8G96BfMhu
8NGpOUY/1xusRUufKrdCsj7e1ZaMXKdy2+RsDQxTBB6tpjs7jcTjqwg0jT8sKeHgLRyj7gwaz0m1
DC3Ng8rFLOY+hA2uvmVV88zgeByB2S2DaHyeHPLJxx+HArhGK2+G4bZp6MkBFeq4da9WdlN0yOAn
MOwGYQv2yyJfHmA1c2D4R7ED4WP1csj004lpbCxUDKYsSzvfi+JBE6ak9Nh43jxpMEh8L7nZHJQO
bh3LZpSFua+e0hO7KfWap5/+Qw6hjJ302f0urzvTsSdt6A44xS7bYlY9ENaSIfhxfpfsT3nHN9Sx
3cdUv8jqqIbuvpICQFJ6njOD/3gxb2F+vcjqY4e9tK7EBMUoYd5YMOU4EPPVnaBwbX4cyDKnOnTU
Ysy6Wotk2YWx8Cls9N4Q3xuDhpslk9UdzdTCLdLH9YW7AHuWDVMsPlU+vOATN/e1m29KRdzrqA+l
nplumIibLVjEtsQeZvD8iZvU1/eNKcEfbXKU7UWdhZkXmQfJJ+J8wCMFdUXCPpYl7PSkQMtCdwfm
Jc0WwL2ZBZ8/36FE4Fxci7aym6o2vzWdUfawkLTUiYbymKJMMXWkwHPMbEiAza9osrHY15nlhtb6
eobPU44QARg43EX9pY5G50KdW2kgcAblsKGhQK8euHwmYNplJD3e+pEhVCQ4fa25mDQf+0ND6WVS
bWeVs2q/ag8+fHW7xZbm/4sZE5tFg8AAyUoXVH/mjm7icfqqzQ9iAS2lQUIpkBVgLMykenAV3PJ9
gvW/W2t0dPsQ3+hDxinyQukjUW5POMdDaDmaIywrWa6YQ2hdNZ7QfJX+4KaY2w9TsXrvPWM3TlVH
uLeqU3MKXzMrvDkuHKhA889DnhwJ1JUQh+cmmIdY1y1450AJcnST6jDXT5fiiXgK09pSb4s7fd/M
fXJIUv4/Yy56Xwu2+XkYpI4uclhP5iRRJ7CG+pY+XC5crxy8MaOi7p2m8XT0wuBECD5+Q7wdvZEp
EvV0nsvaZY5VwlgPjIe4jabpKPgqUIToaJ/8Oleo1wEb9OFGIY+DPGrdHgJ0ah5ABUWS7+d/oW1T
aE9HU7whT1GR27XY3cddZ9Hcx1KQcUPP3MGH3UcaHf56tdZm2zUqqGJ9A2jHAo5GghpDiWf2ezxk
qJ6vrPI/TqQhHAsPPEMQDXtBl4qvXLvF2ZnqwTIUgEZR5Y7bOPb7IyweL40o471cN+VmG1QAqSvC
9G/iXmBgOq+am5YXjDwf9YBGYsgbhi3xQP610nLSBwSDE5ylunus6jg/Yg324wv61yRtCfyvferB
qjLVhnTduuG4hNN5TehryQ8OzIIN71PcvV883GXVQEEmVgkgaAzwso85Lg+i79xf5m+w6o+zs6bC
yJ1mHLw+cwCgr9uZiZ+/h4THdD/FQbi0G7fcr2OC6JAZvFHatzXzjWNjL2MoWD6IULdUqf29murp
5JrjM/4fJI4vOzmor2wznhsD5XZRe4wBRj32r4+C1uQYyR2okFo8mkyp10lcq5Z27pkFYUvpS0bk
j1gfMdGD6plKGV1h+pkrqeKB9Gv/dD1n2R7BVK8Ja8TGPVIBxPDEtBtAAPFwLjemFH70QqI4v08r
j1rPpZFqe+44za1p0ExMX40Qq4DsT5xafV7a4H7JxYPZHgUFOdR2EF99lHdECkuGWoTIEJ6UcxoL
evsQt4/OfGFifl4A+OKfytgkId8ZBi0xhaKzEjWRmWqlgQcktETihNu/1tyP02+ARAXNBlW7tnz6
jO1QRc2AOR8XygYoWidMsYQTuLxlyKhvvf5Sn3hdcNBApZuPXHyuB2sDSPSrZDDemhEEhc4Do4A0
gLdPmOzP/Xt5VWVUS9CeFBn1b3jnfcJwvazPzxs8Ro1+yUnr88obzcEMonHXCgVvBp3pgoeyFkMJ
TO6AZAjSD6/QQhqYEqG3QW8Z2kdhHmoIBvUDrZlAG3tw2/SkQ6tzvEKbeCMqc6u1llp9fxI+45PU
0IbxyWi3z8byLo7kKvT0TAXekTf8KmKCBiU+ekr0RIf1I47fkxC1BV6Wp5T6lwp5UQgF/gz5snHB
XdFafBGeOsQUABHxbAcdrMlmDMGP6epKizyk+yYreZICURpZnf/gWXIEUi1cL+HTIr2B2RpKNN86
O5sYgy/BUZHyoOik12QE5q8zg4YqbUc/4UUsg4/ClY+9EeyrVMtA0TeaJRPogLCb/pfTXP2kculS
VKwrThyNp3PVvzBEhOSVv/4+gkFt4KB9tSp0+Vx5Py/NADdwTkIpr1VKA1hQCi9lxSHPgYRgB4b3
orBK/MbgVt8cORqC6Z0UUVkfyMmX0hM0kB6qBqE9v3B7Ewp0WepnFKfvo/S9DZZWqRVHthhyHss9
fj0h5JDRbvkLWkisU8jS/i9WI/krzb0BTUu73BjmfWGjh/KcD/vdGRLLHsjoxtH3xioVpSes90ZN
NFlpdbiXqAa88kmcBJ/SvBvlzkLM6LkCrFEr9/2mv8DNqA3f2mTRdQNJlLZkvqoWvkZ2hO58TO9n
PD0S/cM7WB01Py0nYY5ecDEhNNrd08YcEx0OtN3xJyuXDAkuIKkbsyaYTbxOC3lKYKGesj1kbRLi
ldyI5wZS4iHjJydTXCnw6b/i+k3a+9xa/e7enCt1jEiggcXA+As8j36+EbhZ2ldN4yZc/NFzf8Br
2gvWOKazm6CL/p+NzvsjVuR+Idv2VnSEax+zMgK2BzayLOkblnBSvWSQgN62dlkROPHgzMH3dfhA
MJMWcCeZKz9qLjg1mx4k7oQvOxVtB9Mbw3BR31kLAovtH9cNCQsVIRUmJoW7uVn+QndLgZtGTlH7
XNELp3XkSlsKsbga/dkMUKfyWOAVNt8tK5/45bN8nvp89tF839LvJfwNWecupLIvCDmpuH8mEsHq
yk6f6ngngowfFiyx5Vdx/izkYQRh4A6J12Czbnpa0LmqX3WjVTcTWjEvJpaTr6xhgXrEYIlbNhEN
Sp8ll8V+ka6FQu966mU61uUVgeHSKZtygOhIeG2bMQIEVVpHpYewlNvwGkhnX8UMJukSqofrB/d7
JPLzhXRfPThcTFMfSL0tcf8ylCx72vyd9vZIhxXu53nRHpifZ7i186nZ5sSlTIFtoT5/6kX09tEP
JanBbqpswZ3m3hArjwMuHJOiUToyFjBFra0PrAnWkVVBfrnxiSfpZhTprO0q/riABmDqMRLe1T/p
26ju0vb348CqBA/zPdbergHDyVQwp524xZALaSuq7ke2UztPEtJmA+no1XnOvASeu5F4bas30BKt
fNlEVSPlXYap3Fh97dTrfJjibgFe3pIRjCOcc1nDwv8zGfcPlJmDe9oWsqQdMVzfHVgWQcx/p42H
th2xu/yQSSUTo0yeArFtTpejo0LG3t9pX1/kqxKp1E6qvQ7JZHBOviHngj0j0wjb5FFVYLRJm6mQ
F4UVLzdG9rGHS7Cy0YEyv+l0k21ET2jyvCsI1dInx8FslUOuaWJJ1hrYrWwxuZSThw+nrSiPRkhk
2xRl3acvpwt/bKDyvwERBtAWjliz2fGY6bmeWB2YeU9PsNgJbFc+1WisDlqv3C9X7o68+GEFe0r7
ZTcCQCjDEHAjsBwgo9IPPjQPn2wScv6xNgUT7DgEXOBsijNlDr4HUngSdUe1UspGfc74tWb96PFm
1PVWUwZfDz2BOdkM8lYwQmcZr9HUuZWrEJneVQecfFwKmEstD3ZMtDQiPu5x5ZMB4HPNI9enBGOS
CrCZKEq6Bye6KwXRT0I9xp9kEXIVS5/gHKDa5/7dAj4BVR2w/Ts10B6c6ligxdiimNNDpTU5TFwR
fDb0l41LlXNY+S+zyD4suaKi6pUDXKKL4/eifdVkVI19D80Xi1qcN2dOOAl+8XjhEU98n5fbcBhO
OCkaRLezvRjVrqGbvBQgr3aDFSZSiZ9xEtmik0ckHG20cgreCKLRi8oaD4fLFrx/pjjMegdthFPp
30isiad3NsR8FJuEfDQUcmpjkA6k9wfJ80MJNL9udt+c5UYdueU8uwaR4pufZMEse+XLpGu1cecK
uOw2bo4eRpxIe+jHhnpZQ1ZQlW+8FdprA0zU5AOEaTdimwo5XfiamQJyxREVigUCOug6SimS1xs1
sx7SmTLPIc4ds8R0W9V8BBL+VAwz4sf7SLvJ6pZIXBl04cMh9IrrQxPiyrTAlW5HaS0DjEg7CbLg
uQI1KpGrNbbhLpPCp6lgUOIhQ4s/ecp4OROW7wOt2MoEJeHmrGFGUbPiTLbxj7LX82K5I8eLox7X
WLzKrMjQdsw/R8/MgDIN23P7KlnFb6B6s4kENho1EZVWFDowHIx9c2eG9sbXt7onFKK2Ue1leGYc
UR5fOwrqYZpVaUmTsbBlSUBObvDwPi+JCMjCM68BtEz4gm0HWxCZ9BsCgRBpSqFpFlS8BKS9zwnu
nqtt3S2nlyIo9puh2BKkK/+xzy/+zTSyhoBG1R/tIN9j+2Zosx5M3kmeUhBOLoIJ6C6RcYvMuvkK
p6AckJm3N0JInYi4PKpORylhLPy0/36hKxsoAWGFfDG/mIHRStThiVojgEJJDtR8KQWovYDBgGyw
I0ED45knyyx3z60oNgF+o+fP/bLNafdFOIB1o6tMvtyIXQ9HpuhcsuLdjO9pQL+igBIjXGYrfFC3
CdHKdtO6LiSoIKEMRkQNbNV0BRMbDeRPYnLfMWivk05q/NMqBLd22OZgYPRJwK8Ik1sfqrz9gjAa
EcoYUsoKWULuZK9mW41kAYk2TjTzShn2ST/OIWRSuKUWGKZc+28hMSe74ZCldiRaNTZ7TIL27aTj
pd3Pr27A4rHiGZecD7QiuQVG3BHk4wsP9dkB5hftTbxq3YJu3sa/mLNymfIjGb5IVDEhqzW0sZ8Y
P5kVQ/dSPVHZWLWc/c4M3aavggoyIAtMsDRMcOYDs/qIAI7kqGJMynopeSil+AeKMB/wzjuN995N
iz4qGCkJFZ5nXvtAAN8SRi4ZWnbC3A24Pca1N9JXIQAgSlQcBHuqeGDcF5Xzk3zbYbUpBBNNXShz
I80Ux8XPYufNePnYOIsj7SdnClk9ufwav2/9L8JjBYfw9PCYVCAMwmWZsPLZP5+OJy2HWJ7rYvfJ
sG0OmPg7Wak/a6ijkHGXRKXDbeGXMtQJuhdeT2Btnme+YKynTq7Ty3fTKSl7W7O8uP8VyytWav6a
PAo0ar3Ev6kXZ66T5VAcFYv3Lzi/Pd+qjStGcS8fmpOtLIv3zslHyTq9C0MO4Ogb/bL2kwUoU3Xa
JSmdOnnVRhGFXcSnnljX6V3F7oRBFHIAZWXxHxwTDiP4hM9NtczvN6sIC7KOzSsWQ+8Mcxu4n9fD
q6DHwK0vv2iQBskqg5U504tezhZjAo3MtpfLDoOrGF1ch9KMI9rCdLC+ANLZUNnuZqC8fA1Ki3xI
yJhSUMJfw+cRHOKrlrcnZXoHOsiA5+uhlGQT3xKfs6jUZYJ5VOeqOwL16b5qn6zRzdpFVLy1u93H
wcBIljINlJkrFYM2y3humd147ptq39qypBvFziMPb246sPXHzF/oEvUoeJDJV2EPOpHwkTKlWRXg
VDxvX3xEgkBTRhkVXBAXIupCVEqiMMQsyZWUnB62TbFah7lfwJ1+FLRNFtzuVL1XKgMwHLlwLhcG
yGTvUv2NGf/1rki/89ceuLDVZ9E25x/MXB4E2UoiG5A9Csr93QLqTgF+X/e2QDdCW0z3zExWoFSj
og7ulg7ICn83e28Z7sKHv5dfDBBRcUI7MTnK7deJzJuLtV+FbtjvDNfsmcpcWRw/e7JXUwGnCcF6
qDdpigd3cp5Y8mrS68iHqWLHBpgM0Ga+RlFxBiNiDMJ3f2lWdLy5U+t3MwN8HZZgW6kAsNIrxsN/
JIgLFK4PGYeGq9tPIC5FAtvno3AIAmHpOhqbGRxGHv4HCYjhAMnVmGgxFcslZh9Nr++sFBvA4BHk
WmNA7DZmwZOB/GFwZFeyC8bvEhEnTxwcKENOOjcP8k2pusxcvo+k1YXqK47bUzfel3aYjGYHUrO4
j1C8Vfyv4EruC5dj6usTNGYuuo144B4PVwd0H/FSLu9rC080Es4znh1XJGk14hND4vHsMKrhM4kF
nDp5P/ssVxwappq+UgX8TZ6jxdlXbP2ySq93XnEjq2D/zDAunFx48EylA/U+40542JX0zSZIJqfm
MHPDQrbYGECsMxwAxnM3KS5XZhJ1alri7f/WLqzOUAkR539xJYvPUzpYa0nPXzLEtVPD0hjUTacD
HXgi10KP+K+ltNrd+TCuKOW6XK5JNrA9GFHNb5mHa6OCvOlsNxDBuUSVP3knJm/FKc41Iz9ldYSL
HInp5JNQ+qW9LeshBSmFllUcW6FYvvTibCXPnzGGuOUrrMyDLAcA1sqN9+AeLsI4mYcm3esemj+h
NF04f0EqMp8GL/LqzlXBYLtVjES5OWfh6TOzj7mOylqnEXwyLTBkFa5FCcVWGb02pV/ogYzQMPMj
SEiW/+NpvF2ju8OSn0WqT4hHFl+6CmcT15IdGNZ0O2cNY4Yg2uxfnTx7KxeqBPXH3/ZGROWbYh5O
wTMPEZ965cT1URCoc32c2otVpdDofSfGobyx/eIQlqYnzlEr7uBhP1TycXqf2qljIsLfj5brdUDc
uLCpN3GLbNsBnxcuuRBJ/W7A3uG4kH9EEOJ7yMmEVBWs0WIV9+WymDa1X6ENXFsC9v6/8YbtY+9U
q90WnrLqyZv63FRiA7vS6xN5HloivkHqzyy7BLCRZu8ZFuKOeRk++h1PtRF9oKR8mUTCMPrMvnpn
NEhdYEzL5oe0YH57qvz8fGQuIJPdm5h5tMIH1XmqCqFjkZjoA/pGk7QqIY9JWzUdXleWyPtBvlnG
LXfjZKUlJ8OYD5Wo1ln2p81tpCRSLC9F4G9ne2R4tmD3E8D892yVaUe/riw3GjPtxggnMHp7T8Zk
HUPNCyFLMFWPUyMEZ//CByOlGpO8U+EUs/pQ7m7ZS67BLBelcKTPRmFaT+qMLvnOquBJdplOfFEQ
CVteM+oyc7wgebaiTsTNZvim/K2Zr+OY7qesuGl1gGC8Y28BOIL1LZtXM+d5uR88lM1JIcItfkxt
5fW0+/ncwyfh5GjXme/N8gnlgMogJDGpXJIBgXe2vrFluFgpTZ6/7YT8o6AM0PBCAKC+b9Wd0+oD
9X/HesG6LLP19BFkv+CKdGfTWB11IXWjkCeTOEWD89yHEk/SnPsOj5XXmkrU1Anh60YRzCnk55IS
6mqQccnNX2LspQdBl6EXxRiWgsHSaG5QdeJQScvAsdAJEPBm4awlwlQG0ZrQyjEvjWV0YxJ4Zsc2
qjh8oqhauvgidcQlnCSZLrmfmHp9hUQQlpws3JDthxZKiNIasWxFB2fzyriz2ylkM8RRO7EGb0Vp
w9kisrL04LVPAQb8WW2o4X/RTXz6T6grdYah7kMG4TWPxc/A0Fg/3JMKK/lyvjzyllyLReMmgUzu
xWxRdZXxpvN0ejd3w/SF2Mfw4gY+US35g5kuQR2LfWjT1zB8syug3zg4v2QbSDGZ5uWxWlIaP9BX
pZuG9H9xkh3Z5dtPtfL2+wkGE1gAvNDKRTXtLkb6YDoTn1tTY4GQYy1RUg05omm0bxPhzdW9P/9O
lqwY5BEZghh8zWsDv4y55YZpFwNK+GvhsEDrZhngWQyDtSNB/vLriTWGTJab3Jb4FhzuqdOjPz+A
Ah9VRFdfc3DLQiMWD+rCTLrrA5Gfv+xbseCVaoTkbe5PDtoeUT94
`pragma protect end_protected

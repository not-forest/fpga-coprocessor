// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
3PoZKWgb+oLiMTs0A39lzyuXL0hIBeleTb7sP7uLfiRV1eXmn/iz8qIOsXma417g
xi0XQa48LBe91ZzNrkfcZfE7U66aBf3kko81XT8uxg8w4rMo9xUtkBJmE2KO1h/M
QeITQiUE46r6rS3STreqJS/T7owI+SLJ8O3sOmRdfo8=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 6736 )
`pragma protect data_block
qd58eULePy7iXR4Y6vv+UoOc+JXrcXwBK/lQMBXypYegS2qlQOlnPF2CzL0wnhJw
HaqXrmVOUXsHdeoVEVFjkNX2VP1mF1r7FxlfEEjc9VV9L1apoqr4hBqfiuAsJzeU
MLXxQftp+UCSSxJY2xA3m47NoJZXrrnl9ELgQwvYlwco7vPNSdV7S42YAepA9d9d
T0S6feQoxnA/IVk98F2gFkMce+0gvVcLr3ls7jC89e+14PsHM7Iymq3IgmIXLL3b
LPNi3My2zQMvECdnLjmLSEqP8HDcZnfE2LNeQ1ntPWgim0EuBQosj39JuJwc4SSf
BD8lPnuO7s4GG4lUUQ2iiQjuQU0HwOCukkr0IQSO4hWTEnZqnB2YoDMkpaP01krN
fE1KwM8nfvGfJ4SetfNZToxejc3LJor21WWhmiAQXVar14XsOFpMBVK6PeaEXs7l
hSbKV7XYrZEIJ4VfvT01xlK7nNfOV7bTNxTaibViCg4w5d5fzCCVFY64unFw4B2U
2hreQ6QaXXVEddb+6WYcXPFer+DwXQaZ4z29ZY6Zbh4G4YVZ6aLtQO0N2Culw3X/
OrU0woFnh5v5hGEmC5Dtb3n1+pcKX4eMOLSUMhLJKP0NBRUi6T4s7DI87N1byZzA
RkdZwEXAJfIKiOLvclBHg0XiH1YttIfUNwzN/gtjMNyiKAiB9qN+YF2pVOjqETZd
IIss7YcVlykIDpTgRym866B0rHF/Tew3LFgNT3OLSpSedYJfqxaou4k+YClppcxo
F+/V7x2+aWm85cJNsruACq5nBxjCSnvaj+IECrx9824FLebGLJh7SxQMpcekKSiP
uOaINquAnHTQExyOuE1nwujuovBg4EwvAOQF+wR7oEU1zAdY0c2284SIzC+Up7qk
yDhUCfR3jp7QZ2CLRA4+8hzceilpmabqrGq6MdbLUb5pFADOWFOkSdVChL/4KkZE
HETZ0Yxq7ET1j2a8VhkrrChJvJGALAsguefo7DZttvQ0OlX2PzwPKqhlukXaxDiq
Pxvrm+RKzAR5zgshCZ/srE98RlIUmqFLd+iq40+3KSsBjGSoe7zPb27XoYPGs6/3
OL1J2UxjcV8CD0e2j/5Z8i5lv1osvpQDnKYTn2qLFb70SI+bIwaWm2JP7cvyU9QM
GU/5UYlM3ex4EGmUP7J+s+puTyHdG/fTs2Z0nVE9LIJu0MF9Dd22Ei+csTL78RFR
74sNYqHJpEwD8Iaw1g7uFNy9QQhfLRNwNgTzbR/GNSPPwIbLPMajuSh/eLyT4iO7
ekkzSl+GMG7D32cg6v/c37Hooe2hj6rAuUX7+VndImdzG/O9K3RK+mpsWGxH+Wil
KBqXhT6t9csr7SE8tJRSFtx0V0pQ9E1Hzm6Q61G+plcKgiW0ivVMrM5WJmEjSuro
qRtsgWyKeFDDXk5GS7j7RDgTuiGM0Mf/hn2/KqWhCufUNAaItxhAPq/MrGP8BqoY
FoQlgDhDAe7Mnb/X7hUWU6Dc5yrPdkN+7qFsdo4hGuUm+rZUHg4YIP4U1veBpgFo
T5Sya6EEDskCHn05K6bN67tK3QRyYqf5m9C7IUKh2fWPLp6ocZ9v7WwynZNa2sEX
nx621pxl5scnNqjrhVtSTERGHWa7lDAIEHbGoTz32Dq16Da3ETQXwzyN4AHVSJxO
4aCmtrx+ljceNmsCSeuZUPyjCDA2tcWOe9UnPIS6EvDpQWLKWYwCz+OvBy97M4ag
wq2znvvOmlL6a7WARaoVIMUqRsD1VM/lIPS8qWAiGwHfYzFydjyBltdLltmWahpE
fJIhl4q8hFpzvoTi1ICZNcvUvJJNcLkXB7YyDqpAnQbHPT29350ZRUNGB5yQ0EX3
6PJbRx/q7yXVg1j8DTTE6oPeOoh/upwNAImkVm+2ULAo4TUfBdBmXSxSneTkk0eK
J5s5T/3IXnJAmHNl28gwUtf0gwG+BUtF768W/GSY8rl7v1REF/Ow4XoMWL+tqdu7
sJkKJ5GzqQkU4wWcCC66PEOk3skji5hUAvceqcRbs02HWvuTBN4HVx6RArcXbPEv
Tqpa+kezXjB4ozMlC8Bs21cLe4CxyLeO+M/1VA3TS9Rb3cDKHJ1eGDl3ySFRr+cX
4fwg4Sd2N5XCG/atLJXzWfFK/zLRvy0vWxiEfwcf1a5WHhBbrOROMOLhAhFaoogk
p116b/IhND9T91ZA/3g/23GFJSd2t6XLKXybX+pnsbap45Rp1zNONBiAhythA6M7
kRnQA9pxKLkH5TXwbgWjznqDLaPa0wXwIvEwRF4KPrF0oKLc5HYKPovac5NilJ+c
2s7BfoiYDhWriwtjZSWkHVkLaqq5Q6eHq6IUeNB8LyOkYzdg/eKSaOfAqwBKWCTz
+rs+quX28yMePJBdxfz7UH54k7bom/Eu4GLzRk1OE/YIH9cxKx2OmV586FsSI11D
RQNxdVSxHfOtbDh/06bOn68XSiImNcupXVTEqKWrg42NHjV4lunrsAVRGHMk9/Dk
khKc6Vb6O9BLEAvYtwjdbZOcaPx71mW6x3nkNYCLhby/+1NvGOfDfDfmqJPNQEWc
oWMwjNUR5KbdofPCAaO51cnBg4J6xTPg+TCC0jWNoBYp/xUem79CINXAMzVp0u0L
g54rUgt7hLCzxQQS2zjqbcpBTwDIBaeX2zZJ9emIARNSvEqj3X0PSZCMnLpONPJq
r9V8ENeOwLX4sdeQmPaKo/0L4cTVkAwZj3fP+wcSIt1HrI60iLvkjcSiQVYfPnpV
pEGRdXD4KnthZZAkd3bTLDh6RKh0z1IZgR2coW2GI5kXJZQ7U9gwbXp3VWW8InxO
k74b0vbTgd4zgqlXsfr7z8t2S/+IsVVR0NUJXKYV1s/OSlsYlD5JZ6YxZnq+Mfsd
Y34IC2yH/x1WrsXqJJbaXtPTkxkeC3sna/nFtF7wXygYCdbf7F97vAmhmgnrVVGs
ajDSk0nd45mkojYQrBWNS/Cyzy0H1drdsXVgBEmT4JvX7igKlUiwqe/lFco5f3uA
Dz1zj3QPH87DMpNQZLiB+u8KFLjVmJ5pkCMNdRv9LchYkCWPfVV14p4jHnXczVFD
GnYvUTjXgvAbqW4I5FBX/e7CqcV7Q6tNI2zIBqLs/Dwr/awrNl5CoPSSBL+ojRHe
7drMjakVjOtB3hkJw2m1J8SX70SSzvMJ01ygwJYNHdlhYi34ZoUshPF+7HKGjr3C
IIOzFVCmoR5tFJtK/YrgbPi58jfU1PncGnXNPYZFTD/HUnnOz98p+suJYRwr1tPw
3liYbbYnFiCaF9O0wuS+EecOjmUadlJwpu4OUZcFxkUqKkfbevUW+PNjZsect/ci
vVw/ukh9pv9D/rpjZ2k2jpblobRJk2CyGTLdH9vZtzQbFp6JMLCZymRZLbgeMhvG
/ScB2TeApXdSZXDQVDvMtKNJ8ZgNu8cgWiOU1mzAIOBMDrUvL/JXQ7nor+wY3bzQ
JOu88uh/mXZxmZVEuy2Ik5B72xdmBSmhwp34OsHZeNNvyTWYDnIRAiHEEbXKhHFZ
4DHIWRXfroWtUIj+Np0uReg2OLrnk8v7dP+p0pcgh5s5aAqWJMOhPxeLluZ3O+Vn
GC5mrtJcNlpNSMXeNUXoZIiVNXyE2+N5EuCr+dovJ+YD6Ktoz7UubIzViRzlvPrg
Nf1umiGGg9XnNcispfkLjdjUO2hc7W8i0pOL5mkh/czwGAoiyUAssqT+pHqLZOlg
DHX87Qsm36NVEe0y4Ntzj78Q15l5ctaAUCcO7yY6drDQI0AXSgQO5AYHNsLaO4Q/
hue/oWnu5cMZq780Old1Wm9E0jMCME/6SUYfmeGOSe4ZvvS+Vwr+GMPawvoTNtM0
ZwKwjDGPB6i0947L4I48wfB5GOxuULsWv1GIqxHtqX+XzVcVy8eMj6sBJw/YTvfR
VmgjYyr/pQJgFv7+lNzLekTeuKpdjJQMFdN4OVtXn06fNewQSMZG0wNSCuIiJAed
NmecFWIN66r1187Um224CT8CtGKo37QPpz5GjpXh4lVnZPmwqrQ/SsglBIs4Cppg
CxmqjzNZB9Izj1Zw0VgtJGZusdFTzrAgZ2VQaxlqbNx6D5ISQHcHFMRGIMmQ8+XH
NekTX8d6Y09aFH3Ol9V9ywf3tM4MnPIHsdFV/YeLD2rxkcYwPoCc9X7mwgmDx2R1
/6Zg0tOHbGff+cZU7Fr9nSPrHhtE4Fi+gXvnIDP8HhbubVVKZqe9sNzR3PUgJ3vh
MzTGNHWwfLIli8vdzHUTF0WIbQOZ/j6syQg0IGXL1EyEaLvARe3OdVxLi3MqdTTa
diXT0TlobbrM56rdIronbe1LlU3kddQ/SKApunfaQ5Z6ETR5uTLNRg+5xGaBXbGB
C2rcWA6P2CQA0f2vTaMAjmPSI72nt4y/Jwbyqvfi0wot6Pcv1wCmBcacyAQAG2yi
cg2sQA7O9QilfdnUEII5ObSjHIRlCorL8lTOgZy1eww0og6fTAs2Ls+lpcnFucpf
3LEZ0082Ftu5YER2qIK9zfHU4aaeGjVMer5d58ZzMEzRZRmeQQvcTgU0cik78EOt
rPKB1I0Za8Y3mEVtjKC5oVwR/D+gFoAWqRqINKpvfzoWgnaGqgY4rOQVWKsFAIQH
TVcvniP5xqKKjfiSIXByL5hZoDeWwADSUFwKUzB39/PyjIXb7RKTUiN8ogaJtV+5
HhFkmrSjlWDhswQ6Q7PHNEE/mfxusMwt3lPru1kDFKtX0H0nnp1xNZyh+h2rPqD9
qobnuZlCkVDxgDIimuQXi20JjZSh5pplamrn5c5hrjf6MrcvXPdkoMx5BNVrmgQW
MCsKS9OOfkgJ2gsiQzGiRY21YJEMbtVhMm2RZGRnptrfQRjmK+IbX+JslpMN2kGl
nE7B67uQPOJLqE369GuT5DiZ70cGOAjHfEeanocD0JTzShsune6xVJdO1aalE87h
9osYRhaZZZu07cerZESM5shD+tQIzmixegrR3HEb3PgS+fLz7qdMT+lCMPSablPM
RNgd3eYWrJ3fvl4GqhYJ8oIUSXh+iKZwfnAre0or9tb2v92Q35InmANCRvRDvC+o
QKnkPU7j5ljFQBxrYKU5zRxtiCNOb3GfthSY4ZT8v5QBxVscYyFQagJ3MzKDRlGG
tLvZuYFWuUQRZIEmCR6D2+pXqpe+mOg+gE9NWkNcCeuZ8/lM7ajqoL4uPJwMTCyf
x8uH+pnYy5xbnBelY7Dzl95mB+YDvhYxP7L3vcHBYgAiwFMbBqy9tRJH7h7PcS6M
KYbMNEGmSTRwocAotLujRCFT6fWl7q7mvbp3hTV8gfcm1LSk62t2sLtd5qOA1Tq8
guigEaZDeyTiYuyJ1+wGTIfPJldsKssLZm738cdEqck7GpR5NNZpPU9qwqxyS2CK
JTK9WtIiUn1Zh6QvYk8jcJhcXrPjrlY74IsCTklmILu+S7pcpje+FJ0skRtfCt0g
nTtJ85V0bW8JzQ/C4eAh8SDyHfuhC1tLW3X61qTu/wqnFeVDc9rzf67h4NHlcGYW
4d8agujNp62gAc8TzodEcj5yLkTWPkPzKV61x2vWSHBO/Nl/Cep1U0KT0YXc1Wyb
43nXQgFrfzWXNHPFHDfiNUKID7us6F4llixa7KnHXdoB/6BZpY/gEwKVWwxTrOqr
vl3WPi3teTxr7mpcjp0SXols21MNgY/hcl7DEWR8YfBly3j68OdTgpe6nDnoE3pC
vBOUJQ+9IGAHoXExF6Bv0YMglTR3kqpa0EENb7psy81wt/pgFQmnVD2d5BAoG3aK
sv2PA5fKwuGmSjFaowT7SORqFh0k2oKjXjPs3VExCTN6GKmD/HzZ5FGZvxG95OKt
rsvzeqSFFbs63+0sV5+nu6uEDIErBZifm6DuCgkcj4x7/4tWyZLbwNgY03TkGKfa
84LtbtkXGSltJtnktoqswdODiW7JZ24YuNJF57ygQuVXTCPb2BxYJYe/66ZGoxsx
vcZus9Nc0dNPdfSsjqpyd8kpX3CKPGvNwANsyQUO533OzyZlGVJ1P7bWroohLVdo
i9NnH8Ju2VUD5jgcbxkioekgGz9rdogQ2Dwt4oq7aarjJ6dSntjUOkxEwBP76RK0
PYUZ6phunBWgwlXihU5ac9mj0FWZpsVkfuZFPdbSC8ex8eVG7J4E2ii9niMRhF5f
BN6R88B2zxx8oYk7TUkmz7fivMkwQ0yiFbk2rbxOzbMrQvjYRKmzYwzfsM7XCDLU
bIZFcj0nkixTDJ5sxYf9E+Ju+a5R+JomhpczK9dFkQK+9ThTl78iUfyNjsotRuUr
CembEINfvURV1rVf97kc79+HrBLVmUqM/mWANxKYYxuFsG8oGreKIg2FbhGaP5Ro
4vSD1eCW8iUYq9We2OpYhoHcBxNUerRQf8dmuutnHAVGBqTMFGYeS8ey97LCfPvi
ws+hdtwbjHKtjvnNVkCCut7YMMox0oWyNuiNm3T3LUA0ykAeJxA2vJkp+ZVTvLjl
MfzFIK8yttkm2UMdtF65Kgba2SxJDI73WlKeltYXyi53mZuET+7f636IjKyJZf0A
JXg+oACvTT4oxwhzoikMbz/tdYtRTPVElEE2nuMNJ0xtQCkshvf5KBcM/+yg6iOH
yx5sNNLfKvK3+oF89DQxmRWVYoNq7DGAEYiu3nN9uFWbUPQFElMQZ7mNvgtQykue
7H3iakiSnUN6zur004quV7g/Em35QH5dRDa+I9sPV9c8BY7ywj07GZYb/bUpP8hC
pDw8AkvSLb4SRlz8iBwBxSLyUGic8avT8J6JVFd/OM8Wp/iK1vZ1Fu3URj57mzP5
jCIgW54JUnQYNExdfDwhU4lyWdkk+pFSzBNgR/Qm3d85YNv7lPVCER7EnG2vr1kp
B4MFbKHeb7tiPSpGywE+WTtpznwBZZS5i8EpeE1GEce8RbSEFXc7TnhEYPNXc4x4
Cs20XFQEtmgjwpdUF/WEtrMk+FvbTX25kO3GF06q61bc0fGG2MymoOXJkdM19Uuq
9IVcwZwo5NGmapewkbqOcAc+WWtCMzbWvmpw3vMtsuio6NyfGdNPIhh3hwEIj7E1
hZXC7Gu0hfc2W8XaAQeem9AAKOc0gc2MwqYKfMLEICHAs0i2asdD03S1WPcQe2Eq
KLPb5oaoLZbH0HsTbvO5vK6oBkyO3EC90pXB4jgax0J9EZ7WP0sP/v5gm2mga0b2
VpqxGpDQ1kzRHtr12kMKCnhpMX73tD9YtWhjkFgGK3GtW55ejHh9nBNtZXKshLvh
yglGRndiCWt474G8P0VUR5oBVeLCR+pCm6IziVGW5qVx8RfLidJAZl7ccLomoHkK
3tfECvPrTqb4x8l7vO1gifEaIsKiPVt8r+L2MHj2pDAXYENad6pOPrEgxMxfq6S/
jfv+ypPf6MFjgZAi+7w+PUqV9daRSa5FUw1A81nLYUNyycIPcYXVihoRV0PN9oo3
3r3H0ogL3eg629/B2Ha6acL4trl20WHofPiUlb+Ut/SvcUOr/m/D1CIsNW8Zba02
P2jQxrwf06pOarmSipyMVBrSApo2dVuN3yfZodC5OeW9Bi5V8RPcU/DD1HD80Vyo
Nt+iyiGcr6ubVwljs81tyseyJEptdE31WFOZag3knTl7Z0ocl4+oritfSc3Rh0Ip
iySALVp6tyZFU4hYLVcNn0eBHjQblszntZibvpq+0Tx+vET8Zc7p3CD/Xn1GMpV1
85v3/c44n9G+jnz2LR8HCmfA9od8aLJ88mkmFNTJ6NaKiSKW7HB2dtTkKrE8aBeu
YnUf8hD3UEaryUMV8KwFcvXKfkKW8IVgvDmV0AqlW4VsjOnGh/SmUpm+gSm9eT5k
qTCKCtgAdEy3tXtHFH8xZX0MutZSBP7WUcFfoRn8AxQawWbHG5cnoaIrqU+hlHE6
qqxOoAPUxUTD7RGNZat5ErKVDiSuawZqi6Mw7nbihN95/LXp2tfUeU1oJAO2QKF/
LdkK9htvbW+dfsHe5OI+U8pcBsu418omMMvTs0eBSsgyDeTQsarUtQAeuCNEEwtd
KPSSWQWjOMBvT5oK9wIZZ+mc5H3yV+R6kcslPwTwBjXwv2F3qd34LD1wyCkXtwo7
elSfHcvPZHdSCBWkx8zsY/4Ep5uLAWRZzzOo9DHusMMy4xDRQpmTDjel0Nn57lw/
QBYUUcBQbRLReqRapHYSiDctNmLorGuGG36rP8/0S0QDP/7y1FOvq/CZd7r3c0aN
587eAmhAHJMCMz9UyeQ7I5Sc29WLpIqGbU1U11t15SpvQBRVvaFmYWaqB8lnhJNR
0OH4zdoBK4D+8ppVdbsYqc2kxUd+kLxfyvvJagcG1IJoNDxKPD1atEEIKeDe3NZE
BC5pFhx9F+aQT6uoZNDbZa+08IH3jOk6r/ZTD2u6AjoaAzwchS+U5bw3Elc9OUMr
ZwWxMJerLevDjPCsdcyx72raIOHhqUV71ESqLzvYQkb7yrw/Pka+OoDBk7fR3Eu3
ZV7hiLgTDQAQOPbHr+MAp4K5hcjdQwn63ZS8gQ2T0m7UUgBbETmVfoJ5u85t8avr
qXj7d/bOepUpmVleMXL8YMfv4LgSpPr7/dqPixanMIDtyDskwfSfz+dGzFWom4C6
Z9r5lublDXAVEKY+mdPJ5eeYUoug7yEf4Tg6HrOCun+mkMV2IjhIlLeoO4Vkl9yd
0iby9m83aLC+g9pjJX3JYgH6zodylWVqoVOorazz5WlspkA8JBMju67E0F/Cotgr
ReXTsypRfe57tR3USV+WJEeR4Bff98gCaF0sYDyTLnzArInBm1Rhd+LBlnCaxySd
l/s+o3zbdhGOm5OoyKzfUkkEGbFMruR0+PZuWEPIBAefBZv1Xnd2VXs2+KVA8ECa
sO/NSkUbBKGe7RoW35gYYUL2UIg/VzwqK5QJYsJx9+zbAVbMU0iCYnHG06Dz7LqV
uJi5dj7laaky1/2GQ7e70fTXZORmH4e3A37CPaxZ2aMc2WLcsx9xIB+xUnvWCqWF
i5ovmkWYxeyXm+KEoZBx9g==

`pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
RrHuDEuCwNbJ9sTbUFOynuksWvqy6UA3LP3gnSOLLbABlbC0EE2QFa8fYa4laMiS
JTUnOdNdyjqPVuBsya6jt0lIk0VO+yXWZdz+w+78Oku0NKGP+lR30CtLh0Cy2ENn
kE6PatNvBbbukRBkc+dkFhGgGsDk8iE8Vn4yGASvRgM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 48720)
/I40G9txYb4ntc8F12oUs2d8oVNyDhs6gCipt85DAf1oQwJrQorPPEyXa484EdEx
59AiBNvWFq+DMT9zz6TcDMZXwaZcdX5Kdlb3/fC6c7/vlFKRLMb8G+qhQRZgTJrI
fSyJ2ITydJK5KktbA3fQhSkSzXzcCMesOqxrttqcbTN+pJEVUwqn90nqLq95ufOJ
PjX/ii4uP2/WVgoUf2wYH043DsfCEuLCb4j1tDTLl2F/h72EDUaCIlARp6tx0NH1
EJfOG49cOQQXE9F8oKOzgCk/Hv84zJBL+kiFPQbr7oh3fs8ZL/tTwCdWxQW+ImUr
GziDlGFp8MJeVbwmcGempMQ8J8ewAjk6mHG9RAy6HZZmrPStdJMA6O8pEDReP5Dx
u0e5+OYws2hvs+TwoRe6pUR5g7zSisRAsJ4Wp0tDVvG0UA+3sPSkPagQvxdAApnL
y3uF6p5tPwl6u0kqCRMuhe+0ntoqHlG508Unc8A7k6+fWLaysKLnDQRrXhp3iGXt
czqGVomoaL0n3n3CjaiJGSvOuNrxThLPeQn0burcAHuo9ZYR6diNf61OVt1xTumF
c5xTXQK3ab+u5CMcS6kat74NHpfZdxpN+CpinUjc39SedIJMt0ho29ToIlL/E9Q9
2tzkdtI1eiNtyjJoC0yy7Y6QWEm97g/ktWwXnEIQLrNgkliRa+wVL1e7N+kKEGky
igmnuzdfSegM6qmYkbvTofRmrokjNoNHTGlN6sgPqtjf3D7ZbAjxXn/M0PH4CEAs
fCFT5ikVewh2o9GtiXOX7rce+8R6WwLO4j5ARRkZcKN9x4pP3oiIkQluG7QbM0di
x7VQwXNtdMBJPARlYm+fgidXh9HGOEzyR+Ct05v7lYqLv/x13Y47ZyJBXyBLT659
YPZl92Zqxp6Cw8NK3oec0jwSsPdK65t1U/C90D2p6KF4JNbUjF+fE2+hWVIiOmOc
ALjdSq1gQOy/d+hdtnZgLN5XXdxZtKxqiLXzMLCbFpsa/coSHJx2YZLIwknhoX27
LNzOoPbNqIpvNuwq92/PHn92Q87IG3sFcbrIrucMRm6m9Lzq/UH/yqx1cdut2xB1
UhOAYHN8lJGBBihPIFjBv6RHTIZy2cs24GrQbAkSTBu63ZhUfJDi7vf2GC6mB8wn
FbTPvejkgZL3UNY0UaALUku5FyA7P6kjlaDz//q3UZ0k+oh0gm/XOFxFPO/fJ3w/
cE3UKG43FWNKyi3UfOTZQs5pVZc9GPn1GGMW1+yiYEM/Jd5E1KR/Z1CVn/DiRHIv
Kighd+5E4RdTPcktw1/2QrMU0ja10ZXvSivUMIrqKTzd5+JIdPSBQUzN9HJfWm8J
ZQBkOJ9Tgq0oOn2FevbXvTEEO5MApCyxc4lNj+tpK7zNJNq1Q2y8f9grIw+htDma
x4ir1fWdaR92AvGebLvjCNjq3rriz4lCcC6YPG4CBdQd+znEw0oCOfMxbc/FkJUK
pSZcm+fgzzlk3oZUMS//gN9sl7XPzGpe+LEQSTlRu2AwgGnH0BwS14KF2wtOaCDq
6fl2KcocVyRoxjGq9H0EfwkgpGkPdXcGrwjAM80fL7hTrKhHwNKr3RXbtLGN7Wn/
xKdMrtVeOSda+Fiy/g5o4M8de6oC00NnN/sB3ppf7+ID/UUly5tvzskrVdWZ84Hh
X+P9ojNL8kxFDZiUmn677ZzPFihXtUOXmHVHjhb0ymBLWYCKNtsTv5wHBKRD7Gym
OQ0pB70KPzAsTFLRWQuPOJmOBuXpnzCATE+6ZOrCNdg860TgwcicY63RPMp9YodT
arzaDpfHSuMxzup2DED44mulRF7LIKtlHjE579d4WD4zrDTeiuQpTEsTo06tIg73
J5Sj8LxvY78CTSsfnbLbnsX7pYLID34sl3bcHw+DUVkp8DNr4nWRodA8zec72awa
rdq5hkZ6dAv5Uz8l03tqvTmJwRJxxmaCRc5Fkac4zMTK6KIcuECxq9r1Qp/G0GCb
+ADJhoUAIBKxGUDZeV6tVrbdYaTnEnIlUlULCD69Y3GMOq0zAxk2E4dX8YoEmIsZ
TvuWEBKqqZyHU3eSulxDTt2FU81FWt2GNN/U2gkDkSzDhfzfshiI91yQlFt0PoPT
SfT9JPtYSD9cPt0lMOpFB9hwBCr6nTxCBrURxqzeySyiglrJSnOMYMcMS212FeUe
sX4dO87NZxv+dzqDNGf01DnGfXjX7FJBAWQ5md3FBJrpTINFtjMslXQajtkq0lv0
Wt+0i+gCfrfFi5mdBhAMg6TYIyxBxkrdk/UofP7CUHoeSz6yEMTJ2YaDYE2OlBU9
JenXJbDgo9e3MNwRBP82UDOySvDd2DJagxYzH2l6RYa1H3HOZrlzMDlFpTZlMthf
UGZrzEYPsp3OroMyZXRh0mR3pbKkDZRjCoFDZmM/vI8K2oQ/2zYXy8xfkA+4f8/K
Hnj+XZBtT3EiBvSz/ikjLbk3zzb4N4lmaNKsM4DEpmrVJiLLfGcqn92LL4GaIZFe
oBWrOPIKU/tqoMjnE3CWCkkhL6z0+rn/z57cBd2SeVuhe9JyQKbN+DHkYFCTP9ZL
RSrqx4WRLRhRDdreENh7wvUZ9UIK4Cz5MHMrc7t7QVmndC2fsDqT4F6HWgl9Y0iT
Fx0AUCkED2UD08w8Rvd2DmfH+H6sE6nJIRqCNAl+7AL9W9pOocok4YC4JoKL1vpC
GUfA9xewtRtSmN14m9Omc/QEPvWtuiYXc/ef0GjrouFkHtPqJxYdgepjAMBFWv4B
+nTNDizZWj4wEV8N9uvU1Ec35LdGgCn0yYf5GHyZqnb3hhpk/ods56CnCQ4UIOLh
qkf7nvqKp7L/NsdTh83Ow71fDY9W4sjbrpF7E8topp8Ri4plNBd2Uf4EbPBOK5wY
Ip/FZccqxPfv6HnJvpayNVruYKP20EHzlcDQmejjdUdMjL9Gatgw20o4N3gwiYFR
WhmTlEp9Vh0B3MPLjPqscoG8xr+TMQBo9uhTE1eDAgQU/vEzVJN7CO0SwxpailsL
D8z41RhcsFqMVIO5InyBQJ7/6egiI2N/dpRf02aXyEsH9Wn9lXt79c2OyqGDB2ro
8tOSHxb99nYyVn4uFMtkT17yTCwOVclURsWYSrk3ikIQkKP0qope/tGLdQxFdObE
igZC3C9RqM94P01Dh9Si6iE91x84UpdB2a8PWfnQjJTdH6euLETAWHUaRY/EnMKe
NC8kFwsDgGdOY34PczBKpbNUVtUFVBPqm0uj6ZztzpkV/Q0IDmQt5JroqOZeKuCb
BlOvqHxyzQp8rhl/itNpoQ0r+7ZFi2SKqebXA4g9SO7nvGqqvb2xmsmUFSscLbEK
f+V2+NHAdp80EvAmaYBe1IuCdY55v9h9VdMD6TOwgcFkRCmchb2KS8KV8YvbNfe3
h+h6dmC4YOUcjel4HNPnlbLQ4m8qd4nLsWn4sCFCwSHF221lOA9Mg2belKDYblI6
B+odZOskITozqtR/Q6l29ev6+pAy3u7FJa37N7NsH1kHKSyEdRkEn3MCWjDzGJX6
unq2zpeCo73eaVBtlQJB5cb0mjV2PBq7gTH58Go392+VyFi8k0+RWbjDjc9rXsid
rcnxd0eAKJMfjYoH8fViFHvaZMBiAo0rezKCH57Fm7Ux6y4+tkKv7DqwtSCfnCx+
Qk9cmQg/kWk/2D2E24M/suQ9jBHrJLi7kf9Nzp2eybrRefU/k65tjfwEin5FWn5G
/zeOKDgEblr5EK35e9CUiRi4Qso/6AqWvfnBNuq7QGwOdSlalAlTSL1+TtRCXV0s
+JZZ4DQzBAgnVSoZBYoFyiadSDqBMswaudp/XE3VgfrYjjXuArW/JSajjTElVR1g
4fKG8fBXx2IoTiZ+gQ+fGAH4CY4MJArYddNFyHi7oAbqTsZ3XDGJyPXY9zPuCBcq
gGvYlAQKCrWRmccaXCXuiOwgOGQYkK5/x+FHPmv16thQG7zQSjD/osGlZh+rfh3g
AaWp4bt4DXGJsGboN0j22mhEuzYg+jZ+NjWLPNDlCHCty9JZq8ItQeRYfjiz2yWd
e2WRtj0GiwZtOCKfRa7I2m3n310LNvDoHCPNsSmjNO0K6Y/L0Tlonz1rm5gyoVaz
9+9RpAMTsIL6lBAb113iGL3JOzimclnKdA4g+ju8nQLBImAz2N3iLI4b0PDeEzDi
UxxClIskB0HH8KmCTqcop6WjSiXz7efWRD2s5wzq348Vw2wHtCdfsFDZ+d4D1Zyy
S3HNMIyBqWcDChANDRaGAmVkXlOxDpQvlU4uS3INu9a/b5P31jMOHsaNh5s0FVy6
hLCXgaeFpbBenAaev7xvjGGlmLo9oYWBEYJ7J0Cj044A+suwXaWwDasXC91lYhLh
vgAT+UhynxgvrWWHbiQn0sdf2vnT60SfiWbopjw+pDbr8ysob62b6uH5fwiOlheE
kKIqacsY+c2Lx9bF95D35BuAe38ysHjwGuJen/Sbjlds9Sfwfc31juelSH/fob2C
Z243eWJwi8V1/FQJ/XCjKD89NxCAUbqNs0BFC2yRhcy5RLe6G+4QUl3JBE6gZelI
/NAh0pK+6WyL2AWNhFEESbY2+bP9kEfApOBXLM0x/65Zny59In51KP/dgzaDOBfF
sh6EiolHnwk1cd8YkGw7enjs3OlWxK/IfJ6pIMPfvvo75K22JdokPIq/cMjVqdYA
SGAGyLszVkIBO58VH9Ow91l/N6uxZGQRGG1M2baexyhcjK3C8v51O+6gKA17m/oX
2qh8MWCUWLasEJm1kaz5HwCp2Y9U//IjjmmLtWrXG+w3O5mgNizrrDH++Tw0pmhR
qGx+DIEjVFI4K4bz+wTjdoYUaTTOzSAy2rvd2V4em+N50tNlmavMUTfmqQTlsur7
skrW6n2DzbsjroUG6UXA/SOcfG/RDT0CVowkxx2LsOfqAdbOW35LhLk/7TiPtVkN
V15etKv+p5ZQuYJkqFHT0qySTMx0Oq/vsiA+7Mu0oJPETe7lngIe7cDTYGTp9dgM
4HcmkM137BKhLhsCV6f/ipseN7copZkAMCLX4J9o/71c9plnFVClDDJxZ7y1hCBF
ObwRfyEAemipgO+3UKKeZRy6LtgIzx9kHH8SItBLKXqmL9npD7p3OA+Dq8VYCmeh
IkGdMY0CpaeLH3hXLhnJYtZGYscxun7QXkVn5iV6D53GHMAmIkXMrdQMDtFp0neT
URB7A4UhbxUoOogMjnE/muEdPTkcDTDmgFGESNj/2XUd+issAX+fwQVKvW8cik89
OydpB2pQqXCNHUZHXuytQKH5bx2OCVMUI0CV26MSTYxgMO+4g/E3nd6MttEObAgl
ObOvHyHRWaMIGl+NTpehws225OwYIeuYtlJZTOHy7wr/DoREzsQ2fFPYWk1qaDGa
UfZKgsVgRmqKgwEClVHKv/UaG6sko7rrH2yFZxEGPQWkf7V7A7mCPIFjMvh1TaI9
p/GluNbonDnLEqhcBtklkVtIeQR/Cy67qsIoPflc3l5InL4Ep4IL137TKdH6llZ6
VTDTk8nxup48j45bJI6CoL46ac3SMTNERQ8XbD/CeYLHegNp79EGR+ukdciH9Nvs
3Qg8SVbGDQTsj5oroqr/rknaEGmLExVrtXnxj83FczRIVNmEaL0JiXkSUsOQaFHZ
hioCjxsT1qqYU00bHxbU0/4cTJRDWcn5oAJNVLgjdG+EdUQ9swnBOYCNfhFxkuCn
3gnDo6VaPkEWT3OmyVnGsfY9aXbTcDPqe92vrkI+bMojgUFUDmDLq6PQGiBzs8r7
Q6nCWFPKH2XLVUDayQVgVU9jPG6uWhKoEqi5+khlTj8I03JJsw7iEQPQ7at5xdK2
BrhtdLZIqBEb01QF2l1keYl3obMnwzKiZt1oPC17QtBAexUvdMIiI75bYM6ENv99
YGLZAPhqdd17vTNp/uboZtw7K3yAod6H8CHCS0DN4cpgKUC9bbHzF6kPREkYr6QO
MmIsOYvkl24YKnDM1e4Iurl/yDg3OTSbk4Mq7QLR18nOoStBldLDwhE5KwmDsLbz
O6nAWenQggagW2j6oVTNaUMnPjY83VXDE5YmT0/yewJtAiyyHTXmkEkT0cTP14m7
nk9yn0fhw2UBOGcKRozOg0WEV0XuJGvltTA+qG+rRn25SIRSnt5qFYPEs7fnXOPO
/kw9PwtMqGvuOuEcGNudsXiCBcV+TxbyS1AuKbf8QbDx18eybfNW3NAxu52OjbLB
q6VUj8/wwCHZ9RpcrUQGXGcBbPDJvdeaB4jtw8rUv0gkAxgMniCR0UWg7OvE+v4p
ans3N5IE4i84CHRelK7b6HToqrYk5Je854d0xd86ecOWYEiLVLJv7nXk5RaGgsH2
88hDItOrOoaNFfxhz4ulX+KDDvlM/bZsl4soYNGW71qu+dFRMFGOgTQ5NVfRZI6K
NI0p+m5Nj4PxCJgDZVrO2Sgs9JsTnS8UhXgG9k3IDWFSXIPLT8xssIbADBTgmH2z
7aViErg4GEXLC3TJT8Ek2GBLm8r5tunNrMxgP4SagNK2IBtX1cXh4W6ua7NPFQtx
q8QdHDINiaXkBnSXJpcd/uPTPsKUzcuEeSj4YQJ0YtKP6VkmLbUwwzKvXKaxzb0v
2YfJLeUROfOQ/pEGDOx/pHf8igRWfM57+SpnQQBKMWfsDW15Dz7kWrIm9DB2NwKW
qVgbKKyu1/Xj2fqc5hVTXZ6vgcqk10A670f78d/v8jUE/au+gtT6OpNA/UpzJhMQ
Qs2wXHsljI58ew+W2t5ek14pDYWxvVaYo6YZ6BZT2T6BaDwU+TrUF9cPNs9f1sAj
UbvIn57CMnAuaHiD8TQ4MgJO/8E1dEjDsbQWWgU2sE0wQGyT/3HvGgapg+hhF6eA
aQ130nw9RaEMXuT3l+dHNAdcEpJvTzPXXPZmYQdIDra+NJbYUHTc9w1dopE45cKv
OfropyLs/WWjgOB/TkC4y1i4K6/7ubVHyNc5CTgWS9dVjA2UtAoivQZ7KczVLGZA
Othvu9oxZ6VzBN3V9QXotSRgGG/umENGpLxeXGlLYbQbEGhwAU2dnjIsDjDzxCyX
EQGfaxIMOIrKs8hprPkdli+UjzU9o8pkwGLx4igPpZjuUG8ayknOMliJDNu4q/yj
XzRQu6fgaXKfgRbsheBkAGCyztc1l/QFCe2VQPPnWwgi5ZBa2nUOX3HVZ/0TMY0D
Em0Z/JcJ9wNn7rEh2TTR802we7mgqcwh97ItmteJ08A2K9iymqPquUDrF01zlaSi
ezZ0wBReuYHdAQKUe0Q5Do0D169jiPhu/j4MPWro2xQ9q5DuhcdeAr76DFvmNutQ
aDUQyH3mXfjzukhX2UN8HPQNS5as113k6GyG/mycQGGJ59SSl3xAI/lD2fmE9BVf
ETDLRPlTv4P0GmospkvsqZv3+iWUbeelnc5s5x0aDYfcUcih9oQh5oENde0ixRLx
Bn0zR5NYFsB2FtnfTt0XmSXBswD2NNbJr36y78UxIR8EiwT4V4JsKQrPgsFks6/P
ufLA35xkxi8fMkE7MpetudgwEZTPg6JnUBjyqXcggVABFr9rCUqmZ7DYRxMBpjwi
nZtYbVO8oCWJuFqXY4DoXiNPV6+g5PZbNLFpK9iQzmVysGT6DYw/6uVIaW96/5QW
B8Pv78RZpfUkC+AZHTqoaefl1+NEQ1DNwau142mkWWW04J8qYjI0J1F8zYtan8BX
mhaCGp/Ibpg0NglzV3wnmGeRwCJf6awnWxY/1BXNxYt6tSOYnX1GijPHo+9EXnw6
PRKypSDjPYmEXhn5/k+A8hCSmnc3fJ0o7H8zg5FOIqsYdiPA1tBzIiOQc3V36wwM
YjRBJEp7tRm1kkrJhhl0G8oZ6R96rP5hb4/gX9xc5f1SubRU1jjsK+NnmvU4s+V8
gFk2dstEgwhOkZgVd5w7xDAH2vWijq4jEbWj0/wxWRDkbax0lxKzw/t3UBZ9sbbX
28T6hbQv6Vwk5NHL/jqYsIHJ5Ylh0hPMlO8ForOfdyqVQSCjwiaIlZlbY95VftRB
eJP9e1/pOpdnx6/guImCQ/3zi/OM2v7qzcbZZodXQtFllr4/PnC76YTjNgsjwWxw
HwrPYVotpCeZ3t/0jVKiNgAI4h1G0xprcqhB7uHPtLN+SJecW9c5jU1Cofx0DY1t
LgfXc2Plb2bdnSSoOcbrDE8B8vOzbHUHsuTqChkY1mjWckHYHzad1tS9szfQ6rcz
2gMA0lUkSzi0ZvGWjHjbS9+9XisOU5tF8UBVIPTChF+SAEHFLdpD3b4kHdbUTKt1
uK4gCkoqnM6NdTdPpBKOYBR0dZ/zBILA1obiNCCb+0uske9uerM727En0WEuHeuz
HThN0Ks3z9+F6B+ITYz58FmVNewVaEDZIDNiiTWozSaXsBk7iDD8n5poQftstF14
Zzx+qipBKEnmnU6dTk98WdmWwSxPSgFxUTS5w7Q58nf6mJS84SOfyQN6VYkoTsAz
Rj/X3/AEgMtYOt+SnE81TxlpVJr12ma4h7EJIUKXUMmLbh8ISJrBQy1qpl6gfarO
SsbOSuYwlYhrKnbEH4cvooYHQUdO5bVZcNRudJJ3nLEH7WhRIrslKRzOBcFHN+lW
vrMeLBKzcSLO1WHM9D3/Y9wbZPE4Qr7bnZKkcnNPmvZPnJbnPZGYZseFrnRZ2zut
qMJTE4bxWTufKc7j8MYimqm3AZtGAy7XiuGfrhTExpA2/Bq46iGWdvaPqBRVXa6C
6/aZxH4/of2u0BU2WM+iTFKfempsOtD9ZVrrCRLDf3c73W7z40Z3PUES4fCC1Fg2
JthIXIWUEuzGfFv+LWKIXKj+X8PSt/pMuJU2cLFl8/85jiu2TIpod4bCgvwUdvLw
Gr+ZNoOuBYfU2OY1OCOCsHxGzrh5rqvX9Q1WE5RoC/ReA+hZlPrRwjI8Y7yhGtef
jEE7r2uGOs751LsQU1Uqb3qZjZZ8vgMADBNt98+2hmXWPXG8zhJ5AA22W93DYETh
SQTrDMkLBhSiBrvUr3o62rutbbCiCVdQgexBnA9FPUzOqsNs/91530bCnHCDC0nG
3eiytmrgEInohkox04QSCvqbBtn1aqqhw9kcNo2qoktVF/YEe7z682PgYwyJZskd
TATolATEm2PutHPKoSoJXZ0nat59FK77uCsxVXGpZ9gMTkSOGIHOTcT3gpUA6cEl
JOuQlkI1h8qgWVedK8hsIq9a8eHDdrh9uHiXMNmj6xg/tqyj4pAaX/ir4yeI+CW2
kb5fl9dvh+1pH8dqJ+o35b+Y5dyiMygCGYQl/12ep70v7LIuF9klnnVMKZ9Y+JUR
LktK0fVzhCWYVCLAyc8+G6ONA9wjb0J/WZhLvhB7TDtY62QX9C3ZrrZeoGO4EvPU
+p24d1UrMwbPD54wuiZsMpQYauhOAt+8It5W9ur7CCoiea/paMfzLp8jY1OQYpgZ
4hnabpx49BLRVcMkMu/KAD/dJgG64DPQW8QTd6brGP53JbInBfHtAqdpqEfzWXwu
rg2O/Y+HuWWxKb3V0ulaMu21GCH+kmxf6CJKuS1YTgEkX2xdc591yKqpfovtiXK2
z4QWcjUrUCbOBF/asdYAJ/LSp7Wlv5e5XRY2hxhag1zMWMVsnzYU2EWIgUy1AG11
NRu3w6wfZGbC0Gk7Jq2KeB7Y3o8KriKEhO8DcPNVZyjp7LaOpDASIl9AD+zXqsJz
gK/+6CI5XAlowh2sCkWusYxbHgAYBA98BECIcJ1sn9IQGo8El13AywjNPTF7eOQn
3BjZV+AaWLM/KGgcQkzIy476BcuZqtpJBmwz1QjZ5RzYYrKy9ccYwOvUTliVL5T/
aSGw3qBPASNDBoAtJk2QzCG3RylNBTKgcjdLudvfOXi40KsrqNhQOpYUmJ8Cazbh
cYujloFPgzgb++oebiRVIlzZShNmlG8omg7OR2cytNJtsENmHH6x7o1dGp8e0azY
17H/VB98W5Q8gRQ6NMNDQ7XqK9Itfjqj5W3O0MszVVnzYhCprFQdsXHQRQh3CebG
Fbt/QufHxtHnC+vk3+O7bLQigr2SYrTDCOoNPqXpVEqdN/x4jdUQbOvBcYoOPRfD
QCMNuoc9Pvk5kpPSbZbXC7i7LJWFH0UdytcKBb/s0p27kVVUGFRG+HbBZz2ZfjWn
Jm51mzOnraDiuw3H9b9xg+2s2AxuDlazsRc1m8RqQZYn5A6EFnWAZRtKwb/aVLiN
2a4EmLitM1edroRxpLO+J5a+fybZJr+zkF8CLTzhu8hWjTtTZTQ+m6RVHt7vtnHL
hkw/Bwfth0KYGbtm6m9vDLm/4jWaAw9piWviBVyYUzhXMq1ySqqaNoc3/T/cN0xd
mStN1p3rIupNcyA0rnmqjaFUAbNsMfOL6cfZ8MdYIbt/gxIkhsqRCMwDNdN82ACr
9K+NIP6eWUV4krQsKJhvRC36LSfgBxbjZXMLZdCXMa+0g86whaqB/XNeAmGbJ4ry
bfkWVDd2Mj1vMAxSe2QsadU02LY/pEOMMnxPtl5Gx/+Lf2Q+6bV4TnTpPXG4D4PP
U7pv4t3DYaFtJ9Y8cv5cJqrPoh5iASyUNmJghh5jH71+Nw95EUVoA+i8pamwhm5M
dhTHZAeKWpHJ6I7fNBfPkKpMJEHvjEBnsmHWszdOmWU7dZn3UCbdjynH2bCqUTmY
o3vUsLogzsBBzfzR+lWxg2U6RvURtsvybZQf1g4vbpNCEKkE70I3ZyUoI+mCWYw6
XxFpX8IOsO/LywR8U7iKq0ZyvCWQJfasxCa3zPscIblxmCc5jyGA9Muym9c93uVm
xTAxEe//MPnmy4YGbyNGEdX/xFNiA4hsA2sKOdb5i9Bl58HOa6iZafZmnxCyiJHz
UBFMB+5tFYcteEvv2bVj9NC5UAtPQXKAjcVXcitZBeWAHiKSZ1QGccCAHM26lBJp
9tKHQDxIRgeE1haX4C1OdbmVM+11nO2qsjOEvroML22CDic+0Nd4oS9vka8yxjMS
pfS6JdCGceJH/ZZs62nmYtwQECK2e+w02ZIE740wmCKjoJOTJOmF4fKV4+FfMl5f
FqisjMDmX1DcO9FtN2ZgOtbOhHiRCff0KJoNvjLvJLteGNjXs9KICe8ui4EN1rU7
kdz+lPCIjXU/qHGBlEHoREXpYjBPkVx0/u1yJVEEpw8BdkNH9JdBvd2/7ca/tS4V
5Tdbom920HMu6oxZC5OntZufAs473eW4r+XJ6mR6FtlGcCr38wWCuv1tDYL9kKQ1
YOqfRlQ0naV/8i2wRXaASthTxbue37Hxl5198+faajjrkGZs+qIKMbORz+nDY+2O
5vU81I3sNpECGsz4U/OY4PvpkJ/tiwp9F08ZO7SzM3QgGXchOitb8tQgemwCeL0n
FGlDqoTwA1AIptFepwgdAuM4lR+PKEFvok+Vry6fX0pt2vIWEskqBMcJoovbuXQN
s845cLKZ/SUImsEW0JwkY64H4amFw/IzTf7NXMp/UmM5B2f7GsAKFU4zJy3bz0V8
WTjMw0spTyHIPnnnmDPhkum3zWIDzbBF54qW/a1sYRL/TbrkP236rFNJcIa2KpsV
FM85avopW6U8V6c3N+I5riAhJPhKXumUWk+oRVdjHs5CNoplH56dBqKdACQFWUlJ
GfTN1SNCLE5HdvKk0GQoZwVl0qgtpqEyIQjCFgIZVMDkWu9BS7xHNv/3C/wvB0Mf
BR0Vu3NEo6LDxoj8fIulvoZhKCYiFga523RTX5T32grJSTH4z3wi2Sxb77vQz6Pb
5L1cuSPTE4fLBygvhCxJGQUc2I9mU36OiWZ1olvHvfgqvqr1l0F6v07k6IzQxhln
W1VkUXOO4nI+sWLqOjRx9D8fyfzAhBPpNsJGrFDff4zv8X4uz9a+4sev4/WB6Z6p
CXjbhH4kVh9yNe1vL5wKBCJk9raIhHKGraCZjTM/jeJhRXDLEAnToWeqdW39TqqD
S+TmcMQTfzwyHnn0m0iT1Z6xEXEQ+IgDv6CjsAZJwgeXc5Xk56YlqPGKs9BesgVD
T3WdP2mOUAkBKrgIOKn9pgNho7hdKvDQy73TFW43as4Cpf4j8LXMFMNV6/5KadyJ
xifpHtBmrRWqi8S9syCoyozQiQ9Lfx3c5BiJ5r53AgzmSDbmi8IeZaoCcXY9OuSp
zBOUAg8s2T05IUanCWa0wmQRXJWZRrH3gwochKX4aa8Y4PQH7w+pVrrRU7rfW0xw
6O7OZZrDd1TcWhJZBxqPOWjjG+oELRgKQCyt7qkSjylXer63BSi+xs/jkeye9l3P
/R9lfTyLUr4V7RoT6gilnfQ1m14cZ0Owm8HswwT0W6/xadVGjepvBXkYu4lgaTGG
3zXQCjs8DA1/CiRChneG7kTIzjWTHtEvzvSB8KU2FpuFqOxNF/Sx/QaQOpbs56n8
Xa2eD4pgaIwI1WSvcdJCfYP7fh/6uwBsyoZLP+/ipLRwGKfm0X0sUKiUHruXtdAW
5cB8fPlJv2Fw7TXqJrUg4aTcb148wtxRx4TIluUEQRECu/YJNy27EZrZkrkxt5bo
MKnVkqPSet4MSyOjnXyefe9wF+6Sj3SP/IQFa4x/7dd0Rh2OV+3QGufPAkpcf3uX
AoH3Ni0lXFf1N1TmpYVbc0oWmrfx47Z47v6xT7JpTjsjRFdh2sHCUvmrcftINxzW
RCe8dQbXPpYFqSoLyO9uRP3aZThUEBZz9MM+RdfaqQv8/5PGBz9YvWjtNmaUY6Qw
jiZNcCpBzPjaDgkyNqWHX9/47GXywZXwaYXHS2DbV/fv4O0gX2UV+sXLAnB82Cnj
tt3ZWnQh8LweGxBY+2X8QnOGGLtF4nfq9FPg/9ggdj+JGPJv9+aZwaWuEt2Y1X2j
/+7HZD28y4TRIm7u9LFzvt5/363ChqfWm4AkMnBo7yt3leEdjocPFSveBelXUpyJ
tIxdXQ64amPlLMDwPdDNGF17d0S2jCFwKaCn4S/hmX84ceMpizTZPrk9M/FKXP8n
h8/ZT74mGZnIJdHRjzoHIdjE3hKN0rKe8auTKEm0oxcHXweq3SeSVB+JzVtTMuA0
BYR+dwd0+LTBiR9z8a15PXDT5CUNQ8lzllOGOO2XZiMtwajDHb/hAkpM/rNwVTQo
KP56jSVQYufUWlmFaGvwNqS2hwIhErswM9p4J5NPAw/XTAxSKouebUSqfxmV62FS
EvfYKGftAIEd8KeijDP9NyhsKL9PqkXSWN5i5dJFgpapsrtYyd5pnQCpii2Tw/F6
2WsgwMaWrTKRmtTfrJ+BWLL8lP+Yu9RLOePHDmCn32aZY3ybptjHJ5SExI+nXqfz
yCH3VbOaFOPwKs2ahZ61OtyO1fx84BahDxPVgF/rMYttXR2FfMj4PSCYQNTSv8Lp
GytgTR0036sZV/F+AeHcnWdG06lNVpeTEqXCtIzhsaUDG0aZ1XinqztvKH7bwkS4
LdX3YjNJ1GYzD+RcmBpYrPkEpGgqRiUj7wuptSE4ZOIg55bWhmE1HkvBwBwcLrMq
4CrAWSaj6m3j06isoBGkWb5CMFDaHPCf4kv2aLF6fuuW+51TQkwgHKF19n6Z96iC
VLkRn46lo4XC/fzHRuSSnWJ5mIMeBS6SBZ8QvHWHoORFXDDJUD+eA2wf2kpSxPZ3
T2DMhjLuui1mskaf8HR1a+j8fJUq+2EZJt8jbg7NCzNSYU0QG5Mbpi5sok8Jk9xF
tJ2F9vxbvwlpm81uTV9jb2y35DXC91teFB2nxpZTOZ9/iGwtGe3s7rXEy1mv6NFf
6WVhBq923+YqBtshYQEl+u6/Vb7Smf6LSn8RId0KxRf5k4XH0TrXe9JlwCDzuZev
AgRraBgKKhJkEpiXyzlDAq4jY8lncc8lwUlhzJqNJb3w8si2vsMrcpMtXF3ecIhu
YtO6/u4/Lvmk2mEuRldyLXBpKXu7uHIfKNSuy6HyxDIUeufYwcuNuvyMLEmzSgzB
YZLQ+WnnFkkmqLpSUxCsZHu9C7426r3BvpGmNrWCG9JhxPEYb3UTWYX6gaUGgwzE
BbfP+EqGYKz+itwOcVJlBoa+ki/zt3Pv1ODvukuYy7oiKnpUG3jzz1wgpdpHImkD
modPLCK1d3LVxT/gcEUr5LICKPZ6aYbKIu71tq5JZ0B4242750Z/h7/nbAyQSYyU
+qrGYPvrZg5kIXbEb/tM/m0LfZAI9ewZdhbwlaf1tQHQJfAS2Qlv/0a+XlLRNOfU
R1jAryEACtzHtJ1AFntqwTMmZHDiJA7LICOlVKSHYHlJNnD/MmZqGi54MgxIBh15
hm6hc9my0aSGlHRj6dcp6mMSHLiY/vC9s08vbOSqwYCZVd90J4+X7YgZPWS5Gzsh
Xp+eAmkWNhVGpU6/YSxxox2yrEkOeR7F3phVPW8qvzHOhzBeorj1goG11jJvF0C0
zY9h3qy64AYjywIgEaqlMHtnJiMAEF1kpHg16gvhSc1mjt84zteJKFaK2vvMRUNF
hF9ZJ0Jmaum4ThPfSBIznfE9QajaymT1cVj7dnfW5BrQbpYA91/9CUUJrqAw6TKC
ZJirKwIVzAbRznXzk8RYUfoFAh1ik8IOn0W1x9fVBdrQCFAoc42h4PiLwQojJEsX
lxZnxvlSt3hBddANEiLcxeXxRTZwVHEutNBBDUtMSVqHjcpyROifhLMTPK7ZDR2I
Qtg6oEFaqW/Ep3TDO8NcCvOo/VBW6cAtQqNJsmVTRy93GqR23FK7LrLEL4uOG1nq
iY+fQeEKGL17B6B9R1jaiiR0YNfowa1UobO39WslArOvVJt8wgReOcG+FWwuIaz+
X/e4loT3F4hkxNdfQc0vuCnFUdx5feB/ycrwfA/fc9t8VelqvILkaO2ffxQs3HHS
30mol/Chdpl9hLp7HVoOYHc3/3/5xPVUXXjwK7uNxxEGacsJVZemxZUuWByF96ec
dGy29LWjJIgF+qsrr9pburcAZDcYGaTaPSgsC63MMPNFUZhrKsCauXZYJKXCtfWp
63v9JqZ7o1N1pZlBGZ3DMpaFC8HG/dbJFGl2xozA+y9uLJqwo5/R4oOnvfrjphxZ
28bhAqNk4beLMNLcXFQekqfs7Qzii2XQUP1dtrIfY+PHMDLs+W+6UQKLFLYybwU7
J3bz28ArC4olwvevnKaD5M5LKP1k8zV6l1dyM/mvdxBby+5SGIvIqWl028fyvnYG
5X77WHpQv3frOCq1l89mUZnmMmzwuU95xY7mAmPg2hTEqL45GNrzUPN4GXBRu1v/
p8OKA7seHFizasRQm3qcbyth/HQMnUkkZ8N6zHxoD6YIrYYT35M49YsxuAHRrujm
19HWoKzN7c3k3+d4e4k8MHZWYLWo5FZFRCSyD4r1CdxvzI+eRNjAIdi6kuN4C6BZ
BIhq9Pvtxz1g5bi9fRiESL6qLU2DvixnWHlg+LEKNq7eLif/BAYMefih8H2NYpW5
hCzUQxpdJgPbnBNZTsu/1lzM6fihDMzc3OC4/shmkZOtPBvWQAo7BbqK+SYPlJMx
Tyh2nb7CGa5TzWCVvSa5gt/MbZ3DVfVvaK+/gq4CO9jKnSWFW4K7sDuiQNIZmCdV
4jOMqHGOqUtfxM74t3OTSjY5SjprneEp+Z1T/+iKce27PPvYpWc0EgQW9PkMH0oC
Z8ZypLD29J7irlyCSlAMAczI8XjTeOxm5nhjtMLfnzZ+EFsUK6s0ZSgobnoACbOp
46IqCvXyfqXIuuyk3VuRfJRZU5GmOMi0fesi8BXLrOhm/4k5aSJ+aeJnJ/gUdxZO
uROVYj6dxKWU7A01pnta/qDbp/s6wawQr632Tbtg0bQGZa+pa8tR3svhLjgBT7Nd
SoEV1T3wxfAQX+Ugyhvo7LS6HDZx9IPNPk13GoONxElfCyZEwRIzIFDFh4SbMbq7
4ZvaNcWvdCmIYPQe2R0aLB4ducMH4SPUMqBdxV2liQ17EG0itlF/wAei4oBWtCAO
nDKop3U+EWv/RWb0C18DBIgAfwVzSiqpTQVotkF8YgnMpZDGiYBcumYTnm3OZso6
1gSj6/9zQc43KVSG3gDLxj4gnB9tdKlgU23YmPqSW9xVViId3tMqlMendsK8WzcI
xytdQw0odnipzfPPmYw0JwoKoPr4N2nYs4eYL/PQlWyieAjl1Aqd4xJHwKvaEfQ1
m4R/zhZBbzaamUWiZkF0km7Kkb07U14txpHy33G9LiKXzjDPzg2NEDeEZOGUrdhh
g8SHcr8qaBoPJzQruKGEn1FqvwUXTYejDB4paCWHFKgqNgbGJ54Q7QuVhKtJJnh2
5CLzpbdG9BxW1P3RIFCIog+OTVKO66ShC1ShFJKfI0gSCt7/GkVbZy4hqZcMIaRS
S9ffZ89Hr9WD9XZ95g7qaIH49JnuZxbvTST8hYBX2eRU34IFRx5VmJnKAH2GhF8v
7p4jtRHdzxsK4fOxy8bZlGInfwHjDvylmnPTVKdTD2a1nI63Xtq7TIZxVJFMK11e
wnvcaYvCYGtdVj7WlFI5df6LKqrxuKPSs8QrmZw3LTcbrmk/3M1IfwqTlYyQJp7s
2+2CZBQe1J9tLRgOKttWX/XmoO8Bz9SEE1HyqwgE+qNdI5FnpO/pUkSqP16EWkhV
yE769dQeo+SAJjokdrURc6xmg1hIEXDbrvn4pix/JzlBJAbZnzCxoNoNoKs9osSa
NcxgQp6pn70KC3ayXeyO0Uw2FkuWp0IngJCTfuPT69ahtc1q9gGocMvPZ98AK7+O
y23B0eJthX437+vRuvNA2+ohqZ8X0Ftul4dg0j7FG/kwWZ/d5nMsE4NT4i7Uin07
vx+ZZ1732HJu0KPQcmV6y689BhatGqOhqJuJZWB26UnCtQ0Aow3oqlS41sOW6d3T
xB93mqQz3e6BefGQJHcKkHy077iVcRDNX4sJSTptVIEiQeeDsYnGo87uFa03aKvC
N1O8q9LpiOK1nm1ogEDsu924xmdufEK0hqfhxabXPSE9gWlgdrGPqy21uhFFiklA
krlSfLu4WGq5XpLvKZJre4PGmaEcckgURC80ZSaqOaH3DzvsglRP8iANBmTu8vRI
/ONvl4BBirwxqz4EH+gcKtp4QBMYPWSp+uA9b4Gw6e9rewPozcqi/ZBktEl0IQTW
U0fvUz3FeUaHWqRHrCiVRlxeN07V+r0N1WcZsegcB8zXwmXFgrVA6T4/YaYyRg21
0C04PiAKRBawfzb9BC65kHPr7F2rNPwl6/9KbQSX/wBuPrWb0NrCXLoquu7YpTXP
pRHAbKq9ycxfGcdaMNvmz+HyqY0IA5T7rim1fxvii01VlgzKS1Z6euOzapnTQoOq
UgbwTxd7kp6o1A2OuFSqY1SKoK1ECj7MoN21IZMxYLkzUtH7a/8HR9YHN9sYAZ62
Zcnn+syrOKnw5pWnILjQdh0dvqfCy+NyoapMm5Z4hbwJrVBGodIrmBGN2DqdGdAV
AYOOWpue+AI8BAFcF0afHQHO7GzwuUxQI/gvHQMi6wM/S8IL7rOdjntePI5n68H7
wb4xkoDce5PKxTS8nn7HTKGdHQCE00hIE2SzRI6CocU8YH0bKHlVbvZ6dOG+K8z5
F+zzhRypQAUw30M2Dqz0wQvLlchR2LtreerNtTTKOZZGCBCmYxVyhyDR84uQuLJk
FaOgA+d7liVKPRtcjNgwfj3JIoY/9ZLr/NyqsoNcmonjiYZEzWQ/erbsi86//NA5
71yLJNzuCdIG/gqK9/pjE4wqYW5eUwWMi3PlmRlioclJ7yae51Eo0X0QFfMk2uzS
XCFu4SawmmF9AN7uOaH+IbpLo2Q2BAH6m4LAjTexruH9J++FirElfzd2riYrlfXG
vxMvJ5P5rzOp4By6FhbX0JwKvYPukdiKtJlFNz6V3oJkZHVVC4G02cO/PxZ/fWgp
qgqHo1yBpPtqBdxq7ZsWYxF11EgvTVjhbcET+K/ia8VN+fPqhpakG1wW6ScwlhSu
suKFunjV9V6bankD37c/UcV1ZVeW4Bx7EQwNZTGq9PeKUfC45s8ZIrznZW/cvWWA
TqnVLBR+fKF1t2ALsC29oMgsicdfN7Hhkr/eaSGUaWzhuehL0wIjS1tfo1V6DR+R
1ok3TPj34FqXoakz69AkVFgm6C8B1VMJGt5kaHD8/Nqo2u4QSg5qOl2eAdGudwEQ
woLsjxFcsqugSKIBaIff/LZlxLByzQ2Beo5EUbQ7R87+/z+hR6cuZq+QZd+hla+P
8SjZzFyOGfMIMZvALyviEdq9ydqnaBDAadtrST0/bhPpaiRY27BWPzI+rtEbkGPI
3kn2eaEJT1oeoN7SU20zJnuHwsHutYsiYAR7//Zqrvss2YrbYXs3WLUon1jIfLkx
sseE70poKcA4nafEGbciA97PCyLBDMURgIxEgu1uAGBzeIJeIUrR2lrAlwkDYBrj
Hty1rveYTY4J0WLiyw+bzK68hwlEsVWFtVRBF4lTxVpGLZsz7gs2kCEnp1qU8y1C
s/x4dxywLgS0JsNlnK9U/ou4cexJQbzl3Leq8YNbFC6GFlTkFLkN+NqT5e6KKDkv
NBJ7WaIpZ1u+8mLGzMe7g390rS1zUQCNtHvfiqt9Nj9dhHxWr5Y8q0HesZdXqj3p
5Om5Q1q+c+yw9C+yz/mQMK6Wb/DiJNAd0srAqyHwvcIVSS+jvQlePsEIpjfDK8g5
V/sJKXDJrp8Zm0DevJXzXEhQ5oAUud0bbok0SHvsCNpSe7eBGgkawcXO4cTQmF/q
Amh/LvZBOhB+6vDNznK/FlJaXJP2oomXF2SNFcAC9VohPMCjDhG5aVcDelZ+elzH
AECwxzB2IRoU9x8ZoGz32C2M8sISA0ckcSvI83M86BJy+VDbSSTOkyYrjmzpkE/k
reXew4SmjVuIAJVQmpSoR/+cSBueVDvGCeYBJl5Z8Op00+DZXpaMm8ZuUprzUmRQ
Cx1k/Yjvaa9wKfQ6K1dJ89Dn6STDQO02PyP/aIWhz3yU3zCYAh3DReXSV4x+5t+y
noBA982ul2SnlGBxKtM7JEL3H8UBRvsLrmwoRv4HJyNZ/JS5p6CxZm5Uc+KlQD0/
4H3xnLaG+xsp1GLeD9puKJFBSJGcqopsi9+oh7Ppg6aAyVGkzCvvuSwV90TWlhyl
KNbYQFSY5jW9T0eeaK3EboUbIVodJ6xBxgP8Q9hL1xO+5ELiSwuMkwBHD/mdTwPn
BqwZrlIgkcAKV4qW6ICHf9/oy4qdKRmblezECV5UUJZKDA34ZieEcNDolYo/P84t
5SgQwm9St/NcO2WXdIRMOngWqEkp63k3WvTJtYFLmz2RwJ4nZj+ffu8yyxDAYrvK
iYJq+bC5dM1zZlGIYKzzed+uzY7lftdE0p2ALwghEeUiGmgXEZNwAbgufRryNWnJ
IQps5mxswv+kIBooNJeXlIz4qUMTUxcS1RpqM8o6KzAWl0+czK+qZO+lMH7xDmv5
Kx0cc797+42GYGXjfToHUXmd7jvTegrt4IUaSJ0HTCz4yr7/6GSvVM6bIRzxC9GM
TjvT9PtIwxYXf8kl693PxbUYMtUMRE193IOVL/F/2i55Swe41sLna9TJkflSiHis
TXM4yfs6BqjxcFURXWaWiNTe1CS8hkkEYxT6JBPNnidzBln7n+dduw6wesawp+e2
0EzFMcPmROimkNmhCC5VWFX33hj8b4OmCAOIGA19z2PnFCPwb5wdARLypz7Tv9vN
H2uTuQUBq/WC0L9dBO13o90cLv/8F1QJoBIRaVGZq9sKml69nJ7cJDCWanmwGC34
fUCQel/dUblhR9v453dMvd5UZjf5cO8QU6PlcpVcYhI4cFm4UrwAZgmvOFrgtVqE
DnH6MKy4BYPcbDKNI37nVKoZuCWgVfsSWK2/BQr4tkPzp2qo8IogzXLAaFYz4nye
bHq+gxQOZ7CQjHN8HjLJeoz+ssAdnCYOXEYaT7zqejcblUM7AubTHzskaTRA1Grr
upAdkLqXPAsaHIXhTkm2rBt8kNVMp16R+63Yk+aW3mu0wclybwOoc9zUk6xGPv8b
oO0+My7zqRnRhvz4Qh46vw7vHUFObTzf2AvqRDfeJgmLjptzDD/AXuatQ3UgEUvG
2/R4yOhKI/ulAAr49njn2HE6uaNUJ15tIPFVO4tKl6ZOIMuE11MxZGtXLHQrGcZ3
sqLK2unurPsJrJS1sHwK1po/DUBSPKrLuCyeBVlCBOGIr9ZZv/WYMX/7Cn5DDLVH
vrAp4EMG94rkAT4imNSvfOFkHpiG5WE4FnUv4zy0sRiccZb0FEgFh71uH5R98+29
QHH/EVvREfPq+orZ5dlfWWXtuUtY0wHRJN3B2G1qY+agKagApg8O/LQVGecBR2T4
GRv7t2UaJtLwsUz/pn81GyuoZTJXlu/eangKDT7ZZJfP42XvCxcPWsPsdQ9o5EPa
Q/5ct3EO4fNG2pjmf/PEO20JeeG500vGWjlyf1lyot3cD5R45d7ooEEPJ2EXbtB2
IXxkFpMuGbKfYmJV6vjO5Kv7RQWLqACx2ki90qPx0bXeygBh113jK8q+oucOEgBT
kfiGutwdD9fs1zHvTOpq7owXUtuz0xMCXnF1XSZ51YSxUZqtXVdR8ayvUuyJ6saU
o2sU64ZlGIcHjBLpzj1Ft9uY79SsZgT8PKEviYKf6g4iczgjHWCstgQ/I68Op8NN
RoPHgjmBaSdU9zKeQPHWO30R57aBYCziBOTLUjNtAVk7Vk1NDnxW9ACOlMZXicbV
jIJ9uET3YZM6fjfig0KGmaUzj5quIQzsFsTsBuswe4CD1Ft/C4NwavY0N977ZmTz
kIfQ9+MUTrmNRuAi3xoFNEXb9Syqgp+kmRIGM3QvTstn9fZm4dzdAVtV4LKHg8by
86S4QNDXHc2k2k5WKQaApzpO99oi0EIQ808Zp72KWdcpBjTxTZnjhikjmZ1AJnxf
XAAaOxkTGLjZbprZ2ZZkpiZXxo++444avQYWuWM6F62qY08FnMBM9C00m4+ww5FG
qU9yf8yBC+tk9tQZ9CPa2cp9sUq96ya9ZnYefUhtzzVJGtD8XZop8r+8RLu56BbT
fnI8KpJxNDCIizLRkjvgDb4lQ8gtZjT9GivbgRfwiRLZIQ6k/jvKWGoqYlpwiSAK
kmzordf+42LvrpTJ/7oOm7rAxIuYS6R8+JGe66GNmIuwhqjLHPQdHlrEn5U9XeTC
yz/m4b6zPGfnQt2O6C97ORjwbSLwipYbHmZ09AlGcVlqzopjvHqKYwakCtcwklAc
7j/1H+A1P71o4hwhzkn0m2zNo0wRSgEZrbak2LfDN8QKmbGyEEspGwKBo02k/4l4
T3zGt/ATrx3uLsDVSLmZCMAnI+KSy/1Si/GfCpB51T/qXG5ZYnFJf+BtEdL09YvG
6k0ImzZ+GyHkLD1d3BsvIskaoxaHunPgPurfJ7IYBREbBbSaxl6ZQlVgl+pRZ8Xf
szK0gGy6VrA8+HZyD85HsCJL9SUgNIWtEboJXaFHUGMOKXBIAeX2oTLq2aK/x9oa
D9IbfpdZzGCxCXUTqdUvazemQOumIlCwIaC05HrzQtlMkB18Zcp6SUW7ebIT72xv
+0wu6W+x2XvdOor2upnz7CaJtE/DqyzZ7bAmEcxz5YahoWtTiQFbCBmRRc2OEgKD
f1AK8LRtxYR8pHqgnwEx8cDHbit5omQMn5KLp0OaCQWKKQTqFFoF7RESfRc519LX
h5z+cEpIJmT9FhUoVVOUM44AFmij8U5w6wbHisKxUsNDhgHg+NMX7AvT+raGH4a+
krJyQoizB2pAW6zPYitaErkRQ54uxXUAwyvlwgHN5QNhdEQV/uYmm49dodBydx4K
IU75Fo230cQ3taeY0Wr0WgZ7qq4PnNuqkouXirwfn0OoC+RgclNNvx2YAXUPbJad
DsONaLbiHnr1r9fZRqWrRySuEGKxfVlUdPZ3NgCKgMV9CKNHmHKdNSsYA99+0Gxw
4eAdwXZcn7LdfEjcBzPLKh7ipvyyXflvQAjZBkH9bIykH/aL36TW4+TztJyM7i8J
j9VrDhQ4y69oDvgahkEj1uKz/UGiBHJk8r4afBKEzMiNSqvSTsfDf8VSdVOjtx+7
D9H1d3syH5la69ajv0tuZbPOATquwa2DSZxUyZJuYYg/xaE1SkAYf4v5AMV7T6y5
Xai2wpbeaqpuOP8mUIvFHYX84W4AZEQp7COTw62QnuMJBWeI/ES/vtWXGDzf6LOW
nafseipYdXSCa+4Z8YQXkXaAkTQDx7HHRSy9O5Bcu6yY+LoHXVR1UcQPPN2iIB8z
yxuE6szNKvpE5EQc7G6NfBXa84RiTV3AwQakbJPHuTsrEyYSCXC384vUcq19kPqk
IvQtgTzMLUzTGz/crD1AWMPMa+C6uvtYwHhD+GSANNkzf3w58FToErY2EfiNjqmD
5SyiFwgl/Wyd2tf1vt3YgCoePGlyFUihSj5fFb2aBKwjX5uIgZSThorYFoWdnjZI
aYMYs2leu3g2EUAWIrp74z7CJR2ECEq45QRaYK7YRR8N7/HQ/ZJnltlNO21BMju7
+VK+zs2znGJG+hfNHIruDPO4HzljQGx/mZA9lQW0tSLihpOOrYMmxTQ4FS1BURLe
jAdGkpywflh4guz4j0S2aqDxDA1NnvBrkkA3lOAlJJn98fT62QRgznvucIa4+wCO
8z73sZhc/kD7WzSwPSbz0NvDaM1pLf8x8TFaaj4d4HDnGbunBEjem18slILfvzFs
+XM1rWF8/dt8VZw6XSnt61g5EelX77JMQmytUcWiZVBs49/xf3NaSdWhxnxF/z0M
W/MwCqbxJzCYRiFQGXjO/YG4yzMMaGcMCZ7OPVpqASA9d9/zQpb5XPcN7yuAbrni
RiDIGb/kHNDYngiIpOCTLRZUVmfXLb0NLpiRq8hD1ghQmb04laCnShQ906ILnWuG
IQX6mMEWxB3fNX/huxar2LlH14FMXpocto6KzrI5DPiuNNYWXe1YJQS8xVEY+eXX
orISp4eQdfFo6VTpXFvFPgc9324/63U8Abbqt5VBFSO9r6CavIvBwHUq7H8FOWPj
bTO69+x3fdw2iaBchZyegDd1oYmkO6wyZ4sD8TrFJrr7/Wu+EAL5XxAbQ9FQ/+Qg
aZIREGI212WEYg1gttmS2TmZ/MUnX/kSyTBz5bJdE9xhITIaLsasRTT9tZ+tsn89
GkyMtzgGrleDO4cdsOr907bnxp3ze1MfpNGqIPGLW0iayY4BXpgx4m4cPvLyygZz
X9Q962VNNH/nQR7U2xWO1niqUDueR6h4ifZaO3FVbF7vbl5OTKcDOHMvrJkFLbCT
S9gVo7/14wRMxDXC8Y3hPMXuZTlRsDkTX8DKz9HTmHLw+v+JeA72WUgC1a5t2Ie5
/BrHg0a7gFRbMAb7yOQ57CpIahl3bCwuTNE525Zp5oTrnzy0usoDYabSeL0KvUy5
4n92yR/Va2Pv5n9o8/5wbcIBu2Dhpms1VxhaC9VnMMHuBR05NPeHRhPilfyE5gJ1
2jlmzzE1yMsKhUXC55B9vHJQjv5AzQyGqVZgbSjNhJyzkzD3ijy9Y4HjsOaKMEpt
Fl3kEltObco5qPotVthzEMxsJ1z0fDKyBP/CSRmEnuSRKXMZodKjm5CgOBvT4ScJ
Wiypatwlex7+Qi0kiSJF9hPkiltHtwFM8FqQ3fskMDf0yQHlm8fwhDFdEO4XxBSb
npXrnlfd13+T9DmhfwIY5MYxZ2bIhsQGWdytoPo4hVBruT+ENp0Cqnl7+YfJedq2
JNi2rgIJ36q5PyIwvU0Coi+GktXEun4gtCL8kOOKO8b0fDBCtr/UFtd/zIkpSW82
tJciNfsIdGX+jyDRNoGLbgN09STTJZodL1bfMmZuqvNCV0f+470N7zh/kI/hbfSF
lZUM0N81oM+CF8RMmz16RYjjD7aQwz+qbnyQtFUFHW0oEiOqLzYGJ2ogTdsAvKxK
A2c2PWaWrN2NPq2/QOVi1eV2Cm+gF0NrMD5Zcv3mIfiJnlTiXocAb7JBzx2Bdx3Q
IWGgtTj+LA2GLRCjI7+AqDElAfIdhj9LfBsHiSpF3gJL//AtVJcaEIQDngQPabvE
NzGBDqPb651S1u5ghLk7Zkzd56KHrGGluTRWKCp70FaFw31Nnnc+Zfd9QzQ5yTn0
eKYxg9Pjep4vEnIX9lAD5y4HDj5zoCcw+n9iDmZ3G2wKk4Z64gTNKOlRVzRLq5Mv
P3ilJyLQda4iKj0CWzRX0YaTUzydUxSMf1DE8RSFg4YwJPgg5dJKBGqY6URlXDn/
yYDUNNz1c6K36OrKLk44vZd9dTIxMkwQxQmlV+Uhub0HqwI3jc7HSlWt5VtjyvBj
rQDsob1qZOlgQAgnIKLydyDmZpUVTm/Dyd8UPc5mIrphmC9uQMPopsmGe1Q/6v0U
7CGbHRhN5KokAn4kmxdxC9EfgwB08u49bNNPvvXHCgLsBQVwjDT9ndBEYfGe1tii
+BdjmCmRoiIIQiLRDCWgX7h4WHUkHtdV0zU/l9DPZ65GzkeujDG4mMMIr+HypShD
ao25fLGSWcV5K/4bFD0cIrr5AgMs5u8z1weYAeic4JgaAMFyR0d3abagB/vYES2i
AF9xaV0vJEBw6kTLbr8vZwZrATEZjN4vj2pMVr666yZnN/XGlU1C17tCBFEQAIjs
4PuStsmOxAercMkTPHT7KZeWFXKRMwqsroXk2GWfsUuJvmI3iW3n9Nj68YYF7UN9
EMG6ao+vVrfazJqOqTv8b2sKorRdUuTFy7ArpgaSuA1/skg/W1kFaZbQeJU7BaE1
i+xvu3NUsbxeDwKmZhDLlm/7t5GaEGttOwrP8EJiOr0ubAHB+baB0ly0vV+EgS7S
3w4iWMobOQ3Q/lsrV8pz4G9e08PtjOhXQs+hRPrQJ7M0LgVlXtXsSJRYNWxR12br
KrbKJKxGecN7ehpN9dN/LXiAr7ijOzJmEil9XW66hjmgZZPcEHml5o8I/C644jka
3z/3RgSVFl8BrZ0Z1b09icRwvsLLFDP2MfnlcXYPyyeHDM+jCMtxkRtSd/an/RBQ
Mv5XVxuQY5JGF50VwMjGCyTKmLyDKVjeRz2SLr/fS4K47mzOXa3r0fHY5rtkoZy0
e3KeX+EVfecmiimaY7S8E3GlSUYuhrLuRLUqBgkbXkZfpl6VVaaGw631flme6HzZ
ZV3kju9fM0sp8897uwM5pCmmKwu7KXAwpC9QnQh7I9MOqvhVL8H6e6i7Z2waXuIs
UdS8fHjZ2eiiS4pWxtb+XuLf0I1+Ro8kT5WnZ6c7dZoKpPusrqQEweqBkGeWMcN/
pvA181tvwg6btQ8mPfk9c5wCdkYYt7U5vs2bazHSGsiSz7eCtgj6qCAACMrfcLJn
9RDXEyv+lwOvYlybtPsA6P4UsRq2tpoF78xIzmPTq16nBBexiHBPRE6xWqloJrHb
EvRtxdhmYrxwtOlXzjCJm0HR0A4cp4uFLvR4ZjcoBcMk4NDDIV/UvjaD6gNKGpVC
cQIvhVddqZiEa79QDve03/itShZKzLoMQIh6dtWaEUvoVnOQeiGMkfVZndYsslNm
ufXj47fUZCkPTUb6ky4jKmkVIK37FDdQ3VvzN12MRHyxt8AGHjjdDZPeZubns9I9
3eK/WvrvFuKvtZUQhhm7dGr3PkHIZgN3wMLmHbXGia+wfOmtq2WTzalhT3ntBYph
FcmChturnGCzUt/HUX9pCF2hwrGSO9VTpxwQU/zThl2G61CE2tMYZSIJrYr/0a9I
vuVG9r+WlHafdBFeHAR7sAjoL8zDZhEmgxCi7BKQoKxldNIhjfiCyS6PsJn4xGHO
xGlmhyLAbPZFCVa3YLV+ZwYWld0DtWTaiG4Wwu9AO/cORZu4BBl+2bBLTj2049TP
NOh5vPO4UVK/IY3XeVlJc1nVkP0HsSL/LgIqroJV9RVEJWuezeI/OdbUAsQRuhQN
OHfuGmBkkKPIERns7Nmq7WsLaNwwboWS7Or0HJPCSaPRpCBt4e03VtZmejtcMj3i
RugW+z3rHDnRNMKsv/aRlGr+mcOBc130A+18Pm6FRUWtxDV7Op2fJkjZKgU6vgOJ
Ee3zO4T9DAGnEFmJ+9SKAmXuGgrZwbRxzxUp8lpIY3JSUtyPb2E2mb87I7Fuh9bX
1/yT+MyujrCLkDXbzPJLujqzVFff4SAMP2I4AiPHAOWhSZdZu0oSemmT+pEUQuuu
kjTXxo9+FfTeIOtG04kljmpUZnTr70c8puYr2yw/+Ph5+9071eLI2rxmhfcqd1WN
C0kRvs7sh9AJDv6ndht/jk/epZiyuGpczwkMtOGVAvh6uVtSWLermnJ5/60GXAxk
nmslNBgTdawnbGUCmKQUH84ds+RzaNK4XoDnFmwfF17KAU+LawGhQIJfdxoZ9Zhn
/noIERSLhczsEitW7kdfOqztt6lPdfOXgg1nUSMn3chpgXvnLCw2YZOqUhl9rlD2
px9Nu5cpMngu9jGMeB9T6hkatyHfFU7LXVNxWhUgIfe6WYOAbXdd8XQBCBSE71Ak
LovcX8d/aRgUCK0wS8igaJ/BWm6rT18m56NZrBYD0MQ7vlKcGEj1UD2+6Ye/hO1i
q9FjbOO2rOBeUi6WhZ5ySBK/t/m2hcywheCX3qVJOpGMWarj482+Sy4xS2Pevtoh
6hHeRMmzIhYMBXOYwJMLS7zPn3yNvRQee2wgJXKjLGefnkT/VU99y81rM+QewSmt
zbzJ00/2wSanILdlvnhvuzl7RSMu25vAOOD82HFSmFBHwKvaE0f0ZBY375auJt/y
8LEONSOEtb6Xd59qjC4yvsTdehEbHjCLOjt0Cpezn+71Azm7JKqLtbAlP+v7jjHo
Ik1kVGtqGuQOuRlbiqWEZSiTV827XFCiUH1T+nRrldFQf4WGznjhEuQgKhjhcAvp
Eh1rLNKhIKPAEWpufS0IW48ajLq1+lAv36YpswgG1S5hIthLQfnG++U1WysGQE4s
pzGRl1UeTlMkRnBr+UOLbGbZoyu2EBXkitMAl6l8z60kVb3IoagpSvZ9S4rgjwm4
ArNab7M5jE4wbxvjR0VDjgCSEcCyGUPJCQhlvcVM1Injo1FhoE5zcq7vYLh9KL9E
P/rEHtgrhtUcNZiSULPzvR9rPKdALvQSuOGfLjgg4VIC/rn9PsMIlRw5VI08wzkr
uPNTNOfC2I4puv+MYgaNQ6YvhV2OSL8yT8qg6NAacD5D2X7YKvSzKU7EJY3Fwpkq
o9Hv24Xa10HgAJ2UandZn4hsugdeY9ZyEPwHuffC5n0M/xxfjb2Ucvb5uXcjIh4l
8DEaui7gFxC6Ak1ZMsHRT9xVfxu5T7HEWXXuhM5kEDNG32Uv7bKHDDAKh1he+u0A
4bxnMpvpmQsqRnI433CFo3lKVIpTQ+s8Z9tOzgAIs41rjlGksJLdRyoTtmltPxQp
g8+MFxUxK83zZpVonWihmEGAlNQqlG8n3DXlkCsaSR72eUG5rwc89JpR1EH1NExD
iaJ896Lfz/pelpZW01dWNnkrqUdyiup9jYGm6Hu1grXxmec6LzxcRiHk8gtS1Lwt
4Dtm1cA6lWHt4/YkWpzkRx8hHhiQR8kJ7/d3qkoEQ5R9RtTx2zydjIESJTsv54ZE
Jzm7X7iCR2c7Sx4Dhd57doDF/AY8y9/j08jN1IuMQsRBoYIdLdH850bxPoRzaYVv
jDoPbyvQ3mS6Xj4XfQ6PJNAusfs8ImjwQD2DQaiPkx6lNufQIwEB31gyWU2drTa4
DeM13mbMHtVaBcNMkCv5GTh0EGOXI5eqY/5FX14/WjhVqgzLg9x8giQWp84K2MSE
uXEg3EcX7QynWkC5It0/guXB5wBo9oS9D9b/Lyyv9AcpoqlqizkDEhu1oOkSvRyC
xlFepHOk/l5cY4vvMoSlnHnBPlEX24IO6oU+CSR/M1fEIHLp6pvf/Q4LGnGk+0mo
Yu9o3MoGiOw84FDy5gPzMjQGwb10NaPIIGzMEQBoPy2F66hU6qT/4KSjOgHtomND
AlO2CTbSIr/bPLHuKbm2zGQY7MerA7FehSYxplg45GUdZ/JH1qi8JQMJsxd34ZKR
9P5rea+c+LtQ8n4Nv/cCn1HrSAo5XDxBycTxGuwyDtS/4yZ2w8cWgDt31UUgtST8
6ez78pdSFpR8+FdXF1dDW21u3nOY5N8WYPO6+ydW3mEb36mAmlvthQhA1O8WXOLG
69wpQi0HKFBul0cjlrqriSgWPTYYtSVGa/3quVthi7RrDlh3slIXvldIdgfk6rH4
Zy5R41Op/ILHMOgvWA+iHRhoHiZxwXi9aP+55Jmcz2AjKFmR9Lqj/MvAgmgjHGva
KibNMuU8eVskJi1w5uQjwENGCJN39HJLUjo5ySffOe6AsLr912hfTYPurNxRIofQ
i0ua82E1Z8Jkg3gaZQBaa4JrtuLX4AZwJDU125hALI6YmI162FfGaT+zctANbmZ7
YGg0iBXRRTX55KUliaemEQxRtUQR8pH2bpEe7wni/3J/KGcFaj7oSfY9pQoxX2xL
lpwBvW3beewPnNtyyFTrQOa/E0w9qQQBaNAJTbhvGsG5nZXDt6E8KOTy0ywt7gAL
PDHDlttXkUuN3yhbGnCvQXQrbvYw5ZkIf8gnkQYW2zdyEXAwizMF3r6ILOizOznI
HEBCk03eEuwvwQSLTm5B45vjSh251QCXLINiR9U/NrXI3oS90e+qUOiZzDnBG4JZ
bjlggfD/GMDyHY6j2FB07NAK18hszppfevFi1knuoTHBB+cnmFgSuPzpM7OQdcH2
UmyJNx8ng+m1hIo1KUH9QpV52JbN8JAYOMPbad30/NRTy91Ib105DCEsp8AGEdAi
FpnJUrTplHZM8DYKA1cSg5l38VP/XrzWDJDbUeG+MbRWwdju+eEmo7HaG/veozGR
VWqdN/BPiYTz9Dwpja8I+/WlSI3PNOkCci+Xa+1klA+/owATgc9CUVwqSiMmczF+
hNb7uVpA9nziZ7jQSUgAamvLtI+VhcWpmfbdY7xRAFb4S4Pgj5ccJntsJWecJJRB
XpYKQI821xK809m6lutl00YnRSqx6PszHz45YK7zq/rKpLBBeAs+NbrniaP9SKDp
4hNx88IiIzfVwrKR+ZK2ClNWivDJD2UX8/sxpDLu6fJg483W+BRSjHgQW/sDlX4z
GAMEJPKHrGWtPwGcHdxhVzcaF9WlsSLxUB+sQewMOibU/7qPvVNaB6MSDOGRqR8o
lsUQqS/E7mxyEw1EU6alyISeHHo93/dOcR5Gam0xbXWUFEhn/7zffBrn3R+aNyhO
Y5u5Z37jHU85e/YLwNxfPNsaQ69Uzhwbtw+vQXvrKxOFEsnGyyHAVmzLAz/zNDYU
ih/i34QVhk7ZeWAeiNM2BJeTvYXtEBO4WLLoAofW6M5JRjQCmEE9rcMwUNTfmeRn
1H1V/Xe2vJkrjDbVQ6kjtmuu371lpF3r+CbpDPJI30s8O5Ibz4Lxzh7Vlyi3dNG4
uVb/tcADQ15TPlcTttcPdkT+C09ep0mloylWHWixzI7rQEijs/C26tLd1FHAim++
gq0w8my3sGgrM74x2pjG0djRiFYK51bntyKa65Mzmz3qTotMmkRkFSbpcJmttps0
Nt0uU6qXRR6cdwYHk21H2IZBZM6LzdmHogcttUNo4PH/WFWzBCkjo3CRo09HCXh5
n++mSOa2G2kMsPWV66zfogxby+RamqvrP5eGfoaXKD0ba3dF+Hjl5oFGLpGKmYh+
0O6OK9fAn4nqIr1BpE8tQJqrc8edDehjk5iwGFZmzgSR1Jhs2MQ9IMOYv7Ggo0sz
w0zYERQmTp0ltiaYkN5J3uwMvUuTRaknafE6BGvlMu6qZ+qrdHhr/cX7MpIdPMrO
lYan8smKCmAkPTUGFMMiGV6smjj2cded8FJbg1V3C6UMYMbn3bopkn0sWeT3+wJ7
z00P/PsWb4goShQ+mdeQ893DK9u9DnpeudDec07QfyUYQIO6sCERV59uDS/wti88
0CQFBurWMSMS9o+Qo8025ynCcyUOv2Eh8NeAl4oX83V1P6bYshA8jNR33nSBMW1K
MuPv41zVIGXZI8/q71W4XOdws3TuGZ3PZx4EzgxPnau5GLukzvf2QdJ0Wx/Zjh+b
I7atbUBCB2xfAJS37bVzfm3vn7Bw9oYZm8EPSKEw9WPHj9F1EHQ54tJsQqz1+oP0
B0aFjMAmAn47c0kyei+p8eHW8v2Lt8WXB3cUXN9F/OiwKV5JE7UikBa/NCkx1pmZ
udW2PDG2rgDrs4OncE/F200VNNzGEFRQO3aIdGdAx+PnyNLOwF3RutPtI/v25Q/U
pBkhaMgU3s4mUakAHVBSELq9Ju9HBU65blirhVygXbFNL53yg0rWFzUGydY6iMLv
nPkXuNF++26O9pOHCfZXIe54yxZEXmj6aADh2t1Fl3gxaR0ie53ouGVLABawpcyN
DoZ3OAS70JpufSNShMMnAZ5ox9ADffnRVP+ke+zmqsdf4El+nqVnj/nldblEWh0u
rGslx3yvH7AyYC5xWuQrJTOa6LdPFr1FUpNJoUuu4a6tVpE1FuNnkC6TmRc39Hvy
5MZfdXhvU5L6VPQirTsUUEfHcY1TlSJW0O53aZHyMOSimzBH1dugFdrFJJHXgdIy
J4dchWAyk0oH1zZsBciS1mvrE87CKCfe5vu0W5pmYssT/l0zx/fOHetMHEWqtHHj
Aza9in8UWUgY+LpSpwo9BPUU6esNQiHfI/Y+kiS2CzvFWUy3IxINgEOKxU6T62Cf
hGaE87UirZKemyNX0+Ol9l7nC1UnHS2iRi51DeOKBwp49lam9HY85LUdpaOkgcUD
IO16Y0pQWqoWXwX0RhEYhfcoUZRkHxXg77K2sb0kwsmQ3Qg5xwYeoJEaQWObMJMw
AfvyMp3TjNH3Wqt27ObFGdTyyeSB49xHxae8CUEnK5oe9hjcUZAWntakZJoGpCBs
Rzn3vuVQ4cYqYxFTPygMZoHarjbKBI+VnJW5x0CQgQlrjg12+8r3d1cz7lxxmYvS
Mmddc2OQjqxnor51wiBgIo8/xi5FWQst7fwV48QTZwDOlgrRt1G+jnnGvAD6JInU
Bp0GTdA16oNV4zZ3eCthNtwwdtvzVlKt8mFYaTTXp20gnQj6FbRV6b2/I/jkEpca
3bPpCeIRDnep7fK+JBeLvuRl8W8nkTuHwBHcH0o8O77vT6d2j1GhjQDDJspWv8VZ
ZgTetrvWR27eDc8dPouOurCoGzpUAA3dzPa21Bkb8UF5pQngms6bqDsZxVLKAx70
aiF4m5XYoCgMhiotxJyJ6Cz//mzw/jgavsmdkaRbFHbbru8qZ5Uub6Avz6Bhca8/
dslCWIoOkcM5kDjpR2DMzQqzEmkrXAWqkNMvP/r5moePwHAcI3HSkqIGBrKDEir3
MMzW5QSLuKqsRSFXARx9IK3GntbOKM2XQXCqaZOsHqpDMu5p6+GNDyOsQLvdwIX7
dFIBWB5qLgjc1al7xvtEs+PQcUZfrD9etfuDgt3U6Aop0wd4OMZKKHxYmdP7a4R1
/GDVOnNk+1JwvAIOY6mdvVrsYfnpen7+pfqeKleJxAZrTv2pQUBKgNCesLqr/NcG
qzCVoo06gsAAcEWPJhwkZXZ6Hq5b7olbZZTI4QLJKKytnBy5dOsUij2X8VOVvnQI
25ZOiei8GaeAn5DER9ByaHo0DTk9vgCgO56pqY6brJI1s8Ftqu6OjbI7wviweZAB
u6d812luTOF7/GOFPiQh9Jx78O00wiiK/ehZ3vLifuI+o71Vk6hmSjmsqVbIj407
Soy/NHxQXPVYCerspp6LC393lPtfBrQN7GX6mGBKOEMBax88uGEm9SarcVLjmsR/
gK/L/rYFaKz0QfedNwuKHqK4Hn0LCLc0ScerfSWjpfQh2eM60kiz3WKzwS0I4B52
MXNuz/bfld9pS6GQ92c61/rd8XfBjDNWriKvbGBA57WKqNQRbwxAd2RCyYWlRHKR
cRgp4ffL6MXArkegFP5LBTq15Bzh3vm01TLpTwMYEiUCU02JkOPXSiQpAuWiw+NS
c+6dp13u8GqBliQkuJNbFvNiuS3K5Qm/ttH18jKbNNyu4KjnY3w8pNLDBPmlllns
9c34Y1TFDtHR1iG9ikYaRdEakPPyW4JcU7LBNNVwEl92O7F3j7Css9pcrp+x33Lo
UFCCPMfkWafAhHc8hBignDlJtwSerRSibF+/PgOb6M4K0vSkc0KrQ/XcC4lAXFCb
WWqYEKOrXjiKvxWBgW68mUKNkuL2lLCfosXzjBhI8izUfuxPZguv6/454Qmos+mt
G3l4Cw1wVmgPBmuYbnduwmpB/AB1Do+xNVDfaenZYsqy6eWlBvHosY+fxxnRLxm0
cAn9sG+MtC8cuphCVxlvGsU+JPZDeLNy4Rf10Tko6wQMm2t1wUYJlqfdhlFhIZVU
Ifaaj/mz2ZoqOBWLJRswy+E1P59KvYYwBF4vp/RIqYlFEHAebMkunRzmwiwEPmI5
4APx+1kSYdF0lQ2VI1q0YetaBpnedyBDH7LP0WUnoJIKw+tqYUij5UwLafFd8T2Q
wTqHUcm8kFWcQybo1ji4Y3ICEIWXfUXD61jUGNi0L0ZCTrtZ5aYLREdJpaOzEAOg
E4lt3E+EAoSnGedJtitRUPE2CCL6yWEgc0iDbD69AESODcllt7I4p4TBWP4jbvfx
QBqoJDH/ePup1jLvhSbEvC0D7gC8LpDCyFvULVjQYhdPQgzOH0n3pEXB4tm4CjU8
Q3vapBNfIVFYgElO29cbv6Kg+DDr1hP6+LuHQAaA3/aSPY/m7DyHKO3zhHrFiZQO
J9C6J7XMq+ZTJSF7k8CgbAo+Zvm5NsunvyLX1ktJHPZj5bgdPOr4+yI0ZfQfiOd8
gYQgkT73cZlOsKkJNbqrnWERe7MYjku6QOc5TVmwNkb8BNttQBa1KvNPzt0m+14f
PAJq4mzGJKTwyauanwUyX7Iql7qXeSucLoLuyCn/JPGU46V7PAfSoFMLOJGy9SJF
AaWsOv8XC4FYZmVa516n+qKuVfDfkmRKRW+w/6c/M0KvG892p7i7xtwMK8+hihTw
8NvPyOKAKNeTtn528o6GbJTqWxaci6MdMznloNdjZOPNihnVTx3XLaASl+Lzn8um
u6/QY9T0AhKJGfElvAnaNRQQQT2a59+xbfvys36eTApkORCPdHD9chfvRgwBwfZK
7L7Ba2ReukCMfRpJxHi3U6d3ZYMC/Qr32Le/d67IcC7qelQPQW+/iKPmdu/J3O7F
XytX60zA0lUVz5pXU/w+kpDajDhHh8+4nKdLB2Kl3cxf69/oLJteiw4uOJ12pl80
YX3VBe4mYc5Tsxr/QWU0c8/6SJL3yh7qA19yUCJY0iTD079et975EBZwNI/lyQaX
F/wbHh28vo3Ru9WZ7K8yHdrMXN2HLp+0/5gx6ySSKbwOzYySgxJQxv9w8hRu/9re
q/kXw2aoFMe2ziK4dFumbwtx5oUeqJRQG1ZZsdVl1yhsjloGwzClgX0x1isvOb/V
t0MrqBQBZKRNXIezPtPTst27W0BTheGEkCd62UT/narAPVk6U1zqhA6jPCTufQuX
k9xaoGrO/RJXUgsTuQS/0rQS8srjDB5hXbwH/5VYd5sAzVFqYhISWHi059pYEK7K
rFFcF9HMvIcW2G0G+tSrn4tsiFipN9KsqrqnRla47y4hdPuXEem1Re55hgsuqamC
H6yOcEUxEDUUnRgKLmWss3Y0RG6s8m0H3EAA/Re4f5CBi/gEUNvkGCxlVbvdjfOJ
yZwSqaEe7kad6w/hjeXAGR+4w0rrBt1mucodA818RuYyQhKl2CScB21fJoNm2a5F
nbtoK82zH0D5WN3VVUA4Odw9bARzExRLwm5bQs+Z+dPc2TGWtzXWH4E+5IimSJP7
nkAoqthTA6XoLWhA0PrTNH5cjOsPcpFY1fY0OQ70hvejdoayqABsXrpe7OVpilpb
3Hz+cwYztDBM4W/hF6i+kNRLB1mNQx9YTNg94ljPuaESP6P3+EOYYwCODTS43tZ7
JY93poJBD1skPgzy15/zBR/ICTKoTFN8AFOBEEFlT+KvbT5bPYSBrXUqBW/5Wa5A
0DssREfP64c9lohN93qAXcqZXnp03EAyhNMLWt0iL4/Azxh+aD8tws8zDiS8hSsN
Ls8jQdqJZ5RVD22giCe3jA5kK/WeMLPvRaBhJDAy2QMTjkR7gQuK2FFNjYKqziAr
1AebWtoclBGK5qwVYveQrk611+6RKCljSLYfb266D12y0+9D37G4DA0uTq+5JIEG
JCT0sIC0ZThUDYIaSgY7gQXrQg3IX/wpPb78XCled5EGLXxLJaUfOxBkvOhQpXoj
VMUePTLzAMCsmTgz7oLk6o+TxIcOnnEN3LPMQ/ZjA9W/uyqgodsMWvJQwbCL4fGF
f4dpyHqgISJdtZ5gc0ufKcdY3LInWPa8O88sWqdglOwweBorMXbRXC+Pbf1/wis/
GMPQ4AKJk86R7ZchvBNU33ka4FOnD2emkcty6fkUEBUuu0mWlPTSh4c3SO/Kh3Zd
hLQJALtnag50fJbRhvLltY2SoUKHjHki2aRVoQg0VzljvuQkSKmb5R1mDSxfDGlF
7r2yKo2d87VuHkX63sJ3GJ0jRyAyLHNPcJs8Hop+RARBUYyqOwqXAh1zXxbK2Irq
nmX7rfTqw9CitzARVarZJsPwe5j62dxPsU6pKRjeUx4eDKRsbkZZvkMgt6Y1uPzD
iq/cYYhmjZ3vDVmuDO+JTISMSiD4uFN4+kbCCNVjnGNhx91ecO2TWOyTa/BFlayf
6tgcD4CBfwI7ywnAn/rT8AI8eyyB4pg6RtpL5IkrZKcl8SKjAgQfqcnh8jO6NOp4
hwue6sNW0BngIy+rg6yuwqGG8bLY2EPUbUWVVSpvlY90DbJu5Ydgurhi935ZImd0
4szeqnhLUOOjm1h4OWPHU5u+DQr3OInpYNyp/JEw+9v6uJLqZCOwdq6XOG+5cbke
S77WiMofvb6A2wTnMhg/9oKdNGMWgkxn8zEdv1ddRbpvh8JduZbHa41XN/2ns6f9
PidYWwVdxYVyohsSGEYeXt6/B0trSKSPzvJFPkSWGsQ4MMsCQQqe/5EPYsedq7Kx
3vBmZxlmRzALTJS4N3n2yNharWXcfhm4f5V4h45cE33FvEuTnhVP5h97q9epImcX
ds6IVhdQ+HvtYNdf82FNTMq/hn5VJhSCErVtnOwaUCo5WRnvyv9MhpOSF+z5L3dg
T78JkmzfNsCjcwSdZ7GkX8Y84KawQTi+Jbbx+SB4diMaX7Kvfp8qI9aA+C9cRdm0
5xO9g2OGzVJiXYUDEQjJkowpo3nuRQOhcMJr9H6UHfy5JyvTISAY7/YAD8Icnr1T
rOnMQY2J/9ypdJh9+D1xXROFjO7R+XYAHy4SSyiSZ7qP+6JH7eSROWD6QOf5Beyn
bCdCgDHV1QactuaDT6b5ttHFxI4EQWuK2xDYRBudmtvFG72VxYC4Pv4rUEzwtGVK
TTEPgJ79Tig3EAcgLqUTd8awe4mZVALpo3kCV4Jki4bYNNb9n+wa0NgS2hKs1L2K
Os8g8+7YnsbrOC+cF9qkJIXymMw5kBE7JE2AlWtZfBujmG9Au+1iNzzITCK4Dtld
+mUYWz9YLSo7mmDDcfxmwzVoOBFR+mRY0k+//BD4151M6k5Zsvc/zHBlzkT9rSY4
QYf/La2ySTSUcHu9XFThZ/Z8Qh+oD9avQ0K20+zF3qSuSxSFVhxan9M51024Ozhv
LKZ1ecwAW2qYxIl6YB4K8G5U37xiItBw2TvKxj2quizBt0ESxOcNYbuNqbaiiecs
6I3I8/T5Is9bGOyZQkXhUXroGOUGpt4NZ+YpfdrOtu8MJpCL6jldhrozD6xSXVQK
zjKWL332OrRS7LeTy7X1ohu6SyXvyuZ/lH9CAxV2vQcGLCMA7uRGsvzYsG7dR9Nx
hB0LA9vHoMBKENQti7WChyNbXbdNreHmdGDlC1CZlKk/GDYNXLQ8SeMkhsfM5pAc
L8vEl5pxethPL9UcrMEHHIDOSLJW5lEg1ObiyFPBEBWeLWX56P0tQQZWpXK+mwA5
P0PfLs6+aAM5qYMwQeISVkBLMp5pdXi5r/98ccBbRl3UokKSQM/XcX8IBJxl0JXf
Shu8V1wokQlJY1l0MVAxXPU6YdYJNG1y+VrPmHyVsy0E437fXTx7jHj94XuCqfjY
RjD7ZcaettSCHqZQurbpEgMmPCf/8bCUe8g4jOeIt2kdEZWOMk9MhOWvewaonlOw
IpSRqzjG2v7Wl6uIcXEEOHw1B3nTP6qwFhJAn79p1KGvll5+5sOo0HxwqpSiYyOu
ZbsigcpOVTzh7PytV6Lrn7jiZP9brWm2Eo6VxrydS9Xw0BqfpiTielt4Zn0mzfeP
0SqTf/gw6U+VmTZQxhMC5rffK7JRGM3Mx9C+w+9eKfgCQobJZmPKTD6La8Pp46Pb
3xs8Abyp6xPgsMo6iBGi08MmHhuCQkBV2hGIYzeMnDvjTeYdIyxrg1XdZeeGlHCX
HVPE3LY2bGqq9+pBzG/lfLNOfd3fAh1OqZGtSwuv6s7EPqGDJxLHODU1QeO+mW2e
6iCNdmMJCxa5MZegV3weDOHfWJQq8ZZFQDOLXQOLTUA5hiMgQ6ztYmwRCXjwpY3f
6ZDJ4T8f6JcNe2JPGpG4CrF7hhivV21xXAOfQpmBvv7EyJAw0jO6c9aTC8cHMzdw
R6TBteVmTzLK56Yld50Dz5j9DN+QIMhBObxgTFd02gd3KjwiXKq94UnpEsgzxuLP
O9xTg6P9MDjmw8JyyMGnngi1lA37521BC9bk+DWka37joDQeyUX55YFEY6q+FhuS
U+mtxpsL0EcRaCbgBi9QhMVBgOSJKWqKqu7HXChIqZ6/98aLi2wZ6K8xn97Zcbye
+rUbuZGos3rQMCVp2Q9/YIZBepy3Q68LI6zD8XbbXvUJH4tqF0X9IZatkTaGkel/
n1pOTRGk2UrsEiJylSv4ky23eZOsIGXbpB8JFAF8UhMBknUY74kh+B/BWzTojhT1
9Tuj1JR+oADNxxB+umfJrwedEcBDeGP8ZWfZFRKhwzhobcy+CJBE+Lc3IsNhTBYt
Cg1JvCGdLfl0ggvgaOqR2L3aekaP2w+c6Y1M3VkpPpwUZyEv04H7EIYu6FylwgVH
cUtYJAPdHKLy1BW0RVBtfJ3xy7xSBBF7z0uIckA+lgQhuLOVwcQR68X8LJatoX+6
jw1Mi8olcJB4S5W54A6UcTU6lFYyITBJhA/KWo+O71It8h/RmWa+ZIACouA66JXj
hROcy60yPrHJSJLLs2AhsR4AcJtmfn9iWSwn+cjth2YX7G5mbTiWet5iwvdIU182
j55tQFqZ2QlGMp1s2MWLY3QqlpOV9PywW3ohIY59FujuFwojxIVewvEBgvJAK0WR
nvkk8lFvBDF/mMVADSukIdg8JrANApjEmDXfyOUnp71v3gc+NbPwrRYC0SKEX7hh
m4uBldCc2uIg9INg4xZ+GEY4CjJTjro7vT+Bbm9XiQMIIoMhIa7DCwe4gySOiGPX
rnZ64RLp7TYyI3Rw9O7cFJ6dWxkFpplDYEijdJ/Mr1Nqvagv3azCNpcvom9PxYNf
V0UKwclJ3m1GSU62M74Y8SFd/Hs9janC3+DUC5mVPuNSz+VXMbVDOvfhbup9mPM3
zUYpa/hKyml3Y2wLnb82pKGrsEU8Ppk/RHi5hhZJJ6ystl9PdbYIC981veqAVaMj
f6mzPPzo/fs4qOpWvNBcxzyOXPG4TTb0KvW5wYs13QqzVy1zeFYvExxdrzmwkpjJ
y/2o7DF9mJb6kcMejR3F9gE3g38gQMiSakuRCGRDvNSBz2SkBBygn+kZEBJR6ydZ
xQ4tlLN6hvUa/Yx408LwZ2eWoskgxZc9CNlEThfQlMU90IwVgMREBo7iQMghg8oK
sNRvfu2+nSHIqIj91EF1IVCXZA8EczXXhsJk2oRMMB8i+rC2uSoPXTZoDH6j/C/i
4y28h4i9SrYz0EZ+n4HVX2RRBQRa3WKRBQ2KswNjbgxUDtSIsOTgbEdA8YaLS8JV
kz1bRmnyfU9a3gGQKkrcevKDRv5/6CoeUfZ3qGcii7+Xhz/48VYe5/S/UyCnuGWd
3yEuFzemenB2s5/6fEVrVIfdNsAVRaHxAyNCIJCEOWvdcCSHaCZFOrgdTtmM61a4
afQ2OIUukzvcJiWD2sH/0PKJTDZ8ls6sicS/VnHcK9o+HyO4iVW19j/tSgyRlv4T
pfILszgVVB3qykhLa0oUUoElOEZGvCNwoZAcWWiTEzA7qQJOlAKCSe0TyzFOKAyK
8L32JysNs1u8yfxWpD5g0ilAlEVY3dRx4tjWUAqQcCZA2l/hTh0LzdXsFFP5vQYs
YpzzK6sde+sPfvx4LTl/EtKdbPg8aqxtAQEfal9ApBB19zb46Wm2jS7C8hQNtgNl
/C9MbPEkqcpw8A5zJguSbBu4QzSQffRjqp2s/bhusaOGog8RLWFEcCBYwE/1MaUH
8TJkltLO+v/yfWUhtuD7L0QnHqZyX8l0DjF1t5nXXYbgoqD7h1RovbhDHLmo1vRC
57tGBd+mRsMjJd/bSW/ZQiTDTkUHIGzpF2op9TOJIi7jKtwJElkdSk3t4ekyOSo2
opFrYpsx1xsEGhhZMEBYQyy+D92al/3q1nt/1gvachCvXtDOcXycEp+/cZMNx+wV
5o2Nr3sxD/WY8U7IYcY5DmU7oCfWV5FRT8fclpqcuviuv29pDHO68dzm/K+zhZmh
oF2KZyQ7RwOsgWSCxSyPgrGxhoPQQy1RLeP3LNNvyvWuZ07KLQhVz45aD2nUrJ8L
MQ+b3t6yAmx3g1dxiZpLcNqIAXkxiXJiMbhEVewDUELznA4NNot/o8rdkN7/baFk
gMUbgaEDomScJ7bL5km2knVgjLutOfx+yEdXpB9/AVRJtgd9b5RGqC+ClUy7GMww
LhkKFxeWU+PCHZuSvJI+YLXSte30bUK1q2mwT8HcA+sp5GN7uCJ/KJpQYKki5p+e
HlgaFyhtgjx7rhP3PIfLMCrZ7KaurBXoauYz1iByliFG0UoDRE4KkIBZlSrImIrF
oId055pdOalGFLXlcEhtGDKRzdiGphRYxKBbhKO/VO7ChZlJ8r/U6+INmCD39mvL
JgVxzsjNxmhNeN9A2pFeY6J1E8EE4vV0+4DtYK4Xutf+ztu6zYiVQ8ZXG5KXgYmN
sf7WO7K2r/5ITmZ/B0iTfDTB22rEVsz7wLFxyyN0Eo8u4Atnk2DsgI0YBVwFxnVA
ZMnMQfaBz4hAFAm9fc3uP1HzfCZFWCWV/S0tlNKcO+CpWnDBiEaw6APWLSHUQ2ov
8NdpsRv5IiFDT0gu5dXqiAPiG6XRIDpncj7Bc2qPDO7m8DEhZlCkmVdi6z4iGZJN
8pBHYoebAekbxbWSWLVaEOWxRv+9HkzSp75tQWUaitlDSQdKYKJku/9qr5K8j2On
x0sOuxNkXlc5HJjSkmEnPE11ILQ98Kf67IPJzEfuotth8qYQ63LCuSHjjJv9TeOD
gMIjX35W4gCylu14NiHruTb2++YV0hrevZAbslvNYAgc0LnuIQO6eUnAv/qi5N+i
t0qDDbo5673BMdL4lyN7Flb54R7MN1KnxUQvFknEldqK4mEJMWv3WXEV8dTWKvQx
PJWEPV2Hv0AxBp1PjRCiOwLPDMZbWJEq1AO3Z6vMG/zVC8m/FxauS5TwhqDLwg1n
8I+ICumv4ZCdhtwzTAPv621AnFcgAUGxUlIpwVoWcHX2YRvyCdacr/rLm+CSTNKD
Rt6Mns35fjdK0ygspTA1AD6yJ75nEL/6C6xeWP61kvEKssLOGO1x4VDOqx3BP0+N
wmvnIizxL/XoHE+V/VvldSstBsV3deoUH/Pd1ETrtkTch0mbV//3KVONWTpbNIgq
BtMZRtAYvp3mSK63hAyGBr6Pez7GZLep+tsv8fidad6/5tcPXYf9SZsAYenzHxfb
Q1o8hDCuG8SQ9aobdX6OlMMQ+u2WGbD18sFlQMhoj7jFWqENNENAfvusytutb9fb
vROVNgvAH9D6FQGQSqSitUq1jxf8rWl3M1i3XXjA6iTGrrGiQdkezUEk1ta1CCWF
fv/ZOaGFMzcQwEDcTCvwoZmutbMXdvn+4zZSUkqm60RLNp1QHmGULYb2+MwQZhz1
yQC612uEVZvi37WrHZyZ1bXdX8PMyeyUrezeINM7fbn9ubtRyu8HkpwCem1w4knv
qdA++77iNohLEkTSt4FEfJVDzzR5i3XDSU1TSzx82UksU3lUSrz83z+nNrzL+yih
rfrihoFiB15tR+AuGyB4H8i1rAfeWRe8y5CXMsF0AmH94e/a9oqfWUcIS5Bpb0G9
wyUhfTkJj+tqOJlFa0nw77LgWvfcslusic9ZfdiBXXtpeLrZS8dfqtUB2mx0b2oE
j/Do4NCbZ3yYk9+eQW8hcoKt1u4n+x0F9/UTu8aW5dyy3F1pDYVy3vbbGC0Awv3H
7JPMvfLLynlXFpxPjKw/GUMvzi2kkAtylHjNZ5k7KgwVCkGixJ1ShKHKIOjk6Hae
t/p5OgEFaHvnle6QZ7R/C9drWi9WsDfpVE1X8Wd5PFkTFrVGpLYxmWWOWy0dqalL
hsQTdowNtQRo514JU/1yGj9fIdSKh5cPQUjbvUM/fGAZSXaes/FbKFZ28FsK1eRA
yXpcnlzCJO5SmCdnWc3fk6eDY6mROssJSKjPWYd43uMwMkYJ65V2JijobbncfZ3Y
IGgzIiGCxfOIMcyKsD8UcZDGqrZfIkG6ge+xh9u2/3vuExE6Ix4q8HivTB0Ry/LQ
vcM4nXLJWmj/r/PlPEs94cobZYKbIRnbyLmzbpaGm6iOYLfnvMeqslf+FtHm1LqF
GpZgWogGOnnAlbLedeAUz7EkDpL9sXPTqH3GNmJYxh8SOpnO9q8A8Mu+wMOLJ26i
8fJdnd54vpvWZbUI78QyEuwSQvqUMasPryWd8AZHerkcx9CuVExTSUE5UoJrBitF
czEUGSYMcaRxTnBVMnzAoEJu8WRcMi3eRfki1Pk0EyXF7cx0MHvqu5CZ+SQekn3L
ePObaH6oBj6WkRpxfjurL4wSZEHi4Scv8O2CU53C6+568RRTxBDPTJQnZmBWp3vS
efmcW1YieJTVXWxAyvZhSAZsP41okbEHPYps5fresVrc5X/w5amUyIGWh0158VH0
ParKbi6IPqA5mVMf5ioQcyVGstmEXlCMJbCetBc2z6zMqD3O6b1vIZIdlioEN6N4
8Kf0Z0iXqY0Hr+EOnT+as18YPkIqBluOEjqrxFEfgYg/t1S10Cjdmi91drILi6jw
Y9ID95SRy9PoGyqvmpJ94HEJDAO2YtMYgSKOeJnPf6ut6ppWf3Ic4dURs8sAbVhe
9Or4Lox5VVvthnp0IEHqZ7OpgtvKXNf+5epaKz6qjARsbC44B3o1iLsH5Z6zgYWE
wIaW6xYWG2thgqDO+/ncEbqG+3eAqHltP4eHcxxruCJDdY1nee/YmR6fn80FzhQL
ZOpDGZeB4XGM30WYGGoyQa28vg0iU8RWElVd3hpEJfc/ZCQt3R1q+YwXRWigpm4S
ZyeAKOo843BJw3CvW9eFSmS66xjUSeF1KBAYOjXhevm6zU6C/7CSJkuQRnN53ArS
q90GtxvgnhCS8SpRQnCF0gRiJ2Sb1PRs/RYE2KuzVM5EipLwcUGbIbaYnwOYCVOZ
4AT1W1lRti+erIMtKh1UYC/JlCTHy189oZpcZ+lEXs1zVCBTxY2ctyTrvYqkZy13
x9MgtTtbQBoXpIf6A8Az3HERg1eUIG3dlzWe+Mg04Yn3gwQILI+Vi5ChL79dcYc6
N945l62t8X241l/J7KGV7ifkznNM48hZoVgiVcv7PZOVod3UNxcnkPgk/p2va5FF
c/pko29lrgIuECkApsE+ZrKPlCrG+sCCGxFNASgCoAJeShNSWfg5pYNmH3ECLYAD
gR/gtM/Ddm6/CHdLVam17h5TkcE8CEe+q7ly2HlHlOYCT5Nht+eOSpWYsI4Y7d2m
xEmPOHZTb5dmXCKeyyFWXxrMljGagSCJLQxD/+FHap2rEScyTeRuSW0hOwnVsEe7
eThjLj9vbCBsFSldCdzGsiFXWKs547T1BA0Q8ufsV8qxW32VtaaWlQ0nhM+0pbgG
gj4cJR7Rb8I562Ise2MaYYXE2pW6vT3nrRm4WXKRJeZACMiRgfPm/N2kmjQRQPMk
R1l5rZSWBW+z80WvWyD0NrCEGSOT+YjsPeSoH9e3P8g17xZfWa/evVUeQb4U1uG7
TDIxhS4CMcj/cLe9c6+vTWpj6NTN4P/McOmBy0gkOQ519Bx7Pyg+dku+prs2nq5c
rREWl201sgJ4K6wC6+QbOG7FjrqxyzzNKECLPpMC6VxEUDcSbaCjaOkLhUpj44Zo
po77ULh/NVoowIruLXWvChXR26H5sEc0t4msQjqmnx4Wf4eMzWumemvf1HRM2++k
+FuQfU7VSZuL3Z0BASKrwIPrMLBCG7c3JeDdRtWOAOQMajYQFA1Xf66c3vY6PPZp
tFtqSKY1m7WjfX3V40WfGXJrxVlV25sX1CuDInTTgyregkiEeFVJd6/Xzmexm9Zf
MfVnPT7dcLssoAWHAkeGLTF3D5ZZyxUlBkcFXtk8g5Cl95Z1H2862NjnBOdpwsI4
t2keSX63DleLN8Td10DaLNUCo/OeQxGla+Iy4LhIG2BZPI6qsoHhI4YoISge+mw5
XgLO8kWd6tb2MMm7bDWPmnMSpLUsA8jd3161AmhVqXObIpOtmDTngZh/AL6Zp4uP
vXYwSo4jRDSw7Rx3VE4G0dTCVBWoN+Lu2RPQ86KJXAUfdcVydTuReUBRt+cl24QT
wyagmyd8Iih+uyI3oO9ZHCVMY/SJz6O+iruM7FNNY61TbEhXDJzqrDAKirZqh8Br
7AKp3yw+I/W9TKCQ+4ubaGF7s2ug5e6JCJPk6YSeiOJ7UEl2tbnxesQ0HV+2TEqq
xIb7feRygRU1QuZ83IjMReZXO+5zaaUu2gTWwtSMnYw7epOoLC6dEu8tCBKOeBiT
Rz1XyVeI3Mi1yLics3WEDz8mXE55tbZMuP1Rnvt8Q+NfucJkimgBQACZMnNKaT1l
HkrIGpZKSGQ+RTLXtgOtr/u0ufnqJkDuW1oVMa+veN6PFECM52JWD2gG17PyGzRB
3xLN01HQKoMzQkm1Ewt2BrySqRnFVRnl4rCl5WX9JrSXzw0isS4ZEWQaovNQKUMx
h2T34kmcbVUTQ2txuXTFKw9cpmtM2y186Qy/Nk+1YTrVV9tO32xX7l1uUeyzJXKO
NMJKbLZSKRibkgDfW1oiFo0c5MErIML9QTrFfIAbywmnYBOfaZgjSr1DhKj9PL9d
Rw5O+4snkiqsRLyTdw14ByJJiIXGmrR4wts2OlD7ChfPnVAdKgqccqAN48wRjgO5
xYBgGn9fJB6zPSc8KSHlQSVM0NWKKwyM3F6jhum4BVSAFB4CFUfKDD4cNuc5g0AK
S7lnRo9v7ecq1ArhSOon89LW5pGOaVhTZpdgBuwwu6rf13rTVyufXBcC5DLpo/51
cP7bV83GmEZYQtk0DuIN2ZLoTTSZF9ckrBkUzJwyBgKw8cTzlXbsfX4DAB7gGJWJ
5F62isj/HY8hDG+MoFVc4o0tmwAxXiYVNcd0hATP2VG3ryXUH9WfdoPGXTpT1x2M
zFLdx0zhc/EiYn/uDCwRaBlynmHUmlfBc9UvCGiymPNicnDYcCNri65qKITwHOax
38Pwzj/4g2LASa2zLIDl4iVD9T6kmJK2wOxrEJ3QjYiOnjFoSscFDZ9KRPkJbwe9
nzXXbSSe98NorSH3jMxerFfDH5E90z2bAIPa9efz6uhq+PlM0o0xEDGVANUtlrSv
sUL1PhBUWjvfZJDbKAF2WhH9WTejUF9Svj62t+i5Yf9+2JuP3wMgFxICK2cx6bh3
fDNQSrouS5S+UiUAx5DhdG/YQiJcyTTFZCWjhx5LuqyzTrASyAO3AqTRWauhi3fI
R5WU57FEu72LxOpFdDkNsWd2+nU5SIGNZPvqq12YaAZPBh/fk0LOB0oVEKw3Rry8
YHyDuf1yV85EAJWORDlnPJnTblDkUhZWJsvES/ajWqCiLN8cBQQRsw3gpEU2Hvgk
PWks3rCo2G+evQ1RWWHwpmKYcJk1XNDAFhaZFNYi+DIg1R/StBwoia1rehuH8Lhz
qu9vNkp2O5t6kn43UT4AitVUKMWbIZhZmmazu55VQ+iclOis5Tvjds1omVOu6VAf
3z86ZbEKRB5KDVW24eaP8vL8VrkmdldMNp95yjKQrP4ruyyvYETcu6lxkDhWD2mP
pQw3mldHx99I/RFpPwBINJ/ZefqHI9thuN6um0LTj+YG7eKrnCVvMgIop3gsZPVM
mt8cJiHLfakiiCnFQ+Ud+TQ8BXvcNK68SaFF5sOrpNwPmJ6+SgA/S269KdL/7dLZ
IFJxjN9D7+FUeZgygHBlL5qwTDfVbLeeIrU+FNOfID5hsNmfNP/1nBKmTtodp1ZB
Mr3fBHPlAjVDZOHtPgn7/0S8ycp4/7jlgPD9zWOoSnmv9Tdu2AC8S2ux8vogaDAU
eo/iIqbvWBCLU4TdcXJK5ClL2M+1M8oiMUYgp9nxwW1WdDORJ+TUqMjvKQ27rb+g
Ar1pozD/P5D6kfHPOUzgo3HQ0+A0VtFnee8FbwfmCy35K3EeygFK/e+PrrCbRIMu
MfnJepJfzEkDnvc3XU9qkj9BbZU5AsAxUgaiKzXUrRarpsvy3RAcL6p2me06BG9a
7bRrZ0H9n4Rk8t+sC6vbY8CyS+/Si7EnMGvjvWuVluEv9MblquyL5E6Tkv5pS5Qn
XS/6Fv6aE1Pe0n9ov9Vsu1/bHJHJSVLUtetoLqfwth8ag65duIO9HjrCM1YwrPhO
ZVjxNudWtza0JZHixR5D1TpIu+IQ4eAHT4eYCCGVxNPopodnoGSG1EdqBIR8QLuk
PbhpDljxLhRegbJz/SXDpB5Oc2CnRx79G232OClThUcA0Q08R2FJfP2kY6HrFaTB
kY13d4rDZqBSIaVX6GnvDTp7T7LcOy0P3Mh9RtRxHFzpYjRM0brmh0gTffhHCm8T
b9WbNme5Pz17LGqVMOxiUkywHmHHDgL6zsrtx9lq9A8THsn0g3FgTZMseRysja79
GKruPZxyWi56IhWRchiNrYbxw5NU9eYL1VYFJO3R/PAU09AuiVOiDy7FdvbsaGSV
CbHnLbXTcArLuOwITPk+Wo1/iRELMpoPZFzvjY1zeU7bk56akN0P2BSztQFoRIV6
9X8hsEt4BH20uVB2qPBFXyv/HtilfgaoDPNDzb2DUK1fTHN0IDLP9/TzXR7au8fn
+us9dQ4krVEBIk3hhVDe4dNLVsPM+RQ0Ba7+iCzFQkEMWtjLkBLrCedpQXDHGYIN
1jHDEuDJ1zwiY+U1dtoWjrIckivRiTe1HcRGnQHWCYyvnkM2JCd7NgApuLBBDLiH
KC7jd22PdhfzlCf5PWhOl+e3tz32ZWZ9t1/snFF7Hi2ztchYhi34H0TgAHhbhR0Y
snbHUmjl3aItx9PKIHdJrYT51KhdyQqgVpJ0F4NKazzBteWCEwkJZIA4vRx9ln75
2xqgG5pBYbaxHkTROmeRRQFy/fTbxj2qNesk53DTPIac1ZMVyIOPqaSvLUfm8jsR
VxEXW5mwOoP5nRHoYKz5p0AJXAfPY+qs7PbSDYEPZmr33nu51d5iAIWWbaXJak0A
J2KJh7ASRChV+A3rSL/sCTu4sCH47uVQNLTRXGNgluWCl9JZ9I/nGTSWHPdyLKWA
67b6BmKvnzgaGh+BLtdwKlRXLW+yN16iZ7qjXhaghsdOrLUqHhXV3MLS2x2BrOu2
IL2VXHludOojuhyHaOFxO/zinbJlkEFw98NblAxp0yNIS/0S3xT3U2Nr6rahsqfL
lllhLg8qC54PzsS1HH2/PHLMdacaaYmi0MvlnMJ2i9+5wA9+yQJt0+Y83FF4dSA0
EvH9tFCJEkAjA3O9WgsEhooWP5o4ZuwQJ7xt1/M18Rt+CCwuQH2bhiiB91t74rf/
0n1AWeEhujOaj/7KoadMBcnYoIO8N5azXWquf+0oU86mAC0mWqiahCy4PuBxIvHk
iJGWLbPGLKfS/pvuuAhEYGgy0aEQ2tlDLcbzOz9TaNPZMx2272MpVuzvPrGxeVAr
cFW26DpOxYy9csTxjwGtcr6OGX9C7daLO3MNC3u0oinrEsDdLR7d5AkBEWDS6NiL
yGfbSI1kcDqWKqi4Sc115k5bzeoM5dPdg62c4T2rvN6J452vk01MC09+T6utEwJP
ZueQgLDLzXPix7ieaW/D3/XJGeVBd5UuLAoWWV/uOsJT6YPT2sprSJT6iSO8S+yT
fp2WYRI0fvckk5syINhhQC8za7YcMUpErSQ9ny70VIs25QsJ38T0b9WPW+xrL09g
MsRFigimMi3p0EBBMwBn3i09fRIxhHVIzZgrmVf0arwEGr9ZRp30ct/TzT3rE6xe
I3IwaXCafKy/QcBnJ56PT2Biqv2V1ud6Pb8H1cXxltWlRo6VqOK27C5Hn5VBJKRp
26DX/TVLuPSzHyyLKsE2AgTUU71qGU5VT7+jHcTNdozMdyD5BunyFm/pBnMGBHRB
1zYj5eL9z4dANVnj5D6gKOjyuqvl5iQx/56RYGRfZ9SApE9mHKqpo5ewffC+hItA
tuJQEtCSx9RciFNMMpt7KqUvpxtVWe22QdAwVGR8qvBe+9qJ/syC4QC7+J6P+hgp
kTEK9oEubXOhlCe9HSQPtWpKlpXkwtu+tOdVr4gdOZBD0E9YaPFCJ8xOdPc6n2vf
TlUkcZCE+z8i6iaFfUgEr2hUjyH/t/KrB86NNmEVZPZeV+31lkZE1EoGSc6tJ2ew
lvqzx7u9TfeD5MvzatGgZEsB1bBi2wUVlm/tv9B06a79yVBRkJDdyWmv5KKUAbLT
mrpY5+ged/PPPnb8A9UW2BPsR0dZFU8Vb+NEWt4iw+wr2qTrxFVszA6UxXImxoUX
IIKF82yRzata4frJuA31HFkUXfFvMTQxzZgfjiyYL+xvMyJOzfXVgG7CBv+dqdKM
TABQlOMzdhvEp2/gJOIhpCNaG14FK8JOyLfu50aP2gM1Xv5DuJdzf9MM4krE5mJ1
31ydoKwFPSSixLGjYc258FN7GoegGM8kr73MByaG649LAUGK8MnCeag9yJReINtc
xTW7fYzTSYDKeE4l2kaJHWkMGlC6hxPlSPA/BnWNtnIJuOS/YpQKCBjMhtsEztEV
fsZ7dpyz6o29QXUdQYH9gk7ThzcZKsfZ6ydU37kIcpMKairDIARLY2lzckDWsRAC
GIyKJGC39sI4mf/WFi2FxswosKrNpjWvcqL5qBhKJ+DEnby3jdfwmSdw+v9CpOge
qmpYuKC9i8+ejMhuIK51EsX+0gTTYNiTo8dvyeEI7gCAXuGOViUQL4LjCqxYxkZa
kDGCizXI+UOu9OR5QNdktlPHOgYbVAGSfHZT1WK1nutRXnMmW/Uql/klTO2KvBjX
aeh8v/24G6hWWUWRoQIVrr+NU3FQ07fI9x+DBeiKhwVTdjZ6rBmDJxzo9lrkCvF9
PpfDrFLbOLLWvV0Inz8VN3sp5IL/vx2cw7yOaR7Sx9n8CO4MiSOJJ/JdTwZ/NJjW
nX8VDh1p8Eqm4mWhbxijlQJDIPwIj1E/IQkwnbqcb7qKUva83PNd5HOvsqdMT7w3
ArF12k2H95xDcekoJBlbdEwuFnfGLW+Cozc8BC+a+Lj7Bl4IXLvgo8WmFU7SG0xS
t1p8MXpa8B/SnpzdbqA18l26MT17OY+S9D2gah+DBVC5GRwFF5KNKvrx9jlWsS2Q
okGkgbCuKMF6qZgsIirMOl/iEsgqDavNjRvhfqwXniTA7LnKCr8AGowwaLRmlAmC
N54a7xbKHEmPgICFYDfDXVXvsdYCUhaBRaHYIArnA91yMmhzonvE0s1MeJbIpOB5
Dk4Y7+itDE6N0VhVOAyNJrCufEScEI3jaF17pZ751L1bgTze4Po+tXbxSfpnYUXA
mwLzAxIiCWnEgb3HulCXUXJCzvJZxmrUHMqNO/PEtRqdYsz2ukHKJiYS8Ov4gjZf
SNqNiJ6KaKac/FIATeD/emBlzUMV3fjjXwh3y6aUXpA2y49bQ/YCR1xZ3DOZq9ky
W00/AmQbXyuYmn/o6xuDXGBC5SD9Q0IJ6ZzIcb3ImX1i77Aa2RiECdQ9uwViPkRO
K7rYn7W5d2npRxHnULGFHyAxVLc7Ty6VDWgg6zqWY8nk1Zro9ar9RQPKp2n4vIsr
yjGZrnI5e7Kdy1wLOGTUqpjzm7htNRFHX7mUXuhQsj1jgKyT4VuSRXGDst1hqYsP
bUzInbr55n91wCF4K5OQ5VClC2ayNPdFYvkwR0dm+Q3lcTheO9QKe/YQkuvarsVs
F79Z8/emgK02/vYylIgoI5texvEcftiMB7BI++qlHRuItRQhp+D4pvBHXNsnVWA1
af0b5PJZax0Q/oUH05bk0noTfn9cAEM2d4Mn0rvS0Q8aq5k7ar4vqsbkS8xhMSCH
LPQ9DPkx9ZoaUwCIVQAyFuGAUVl6McucLhDoXsEtVWb4fPRmGF9PHOneIuDf+gyR
ihdvigFVMRjUIqnSPu/826vyMwqgDpre928or/XfvXpY5nT3pbLWCQIVEkf9mldW
m19pUPo/xaoCMn9PDqKHF0g3x2an9gJbSjP+KK20bicBfrWmFJR4c8J+f5UH6aaP
1221n1/lgN5gVKJGzs4y3VtnU1QKX4x2JKhj3KPBgYbF5Eou96m2yRstXfWKPtFl
SS3C471sgQeOrfG/spFEhEmyA/hbYEq3dsfXSww4gk3vxNa0txLra7pXYU1WCRS+
PkRQnZM70tnQpaIceyhknJnbLIaCQHJP5htQ+1s1s3iVoj6CG40gbpsoaeX4g+yz
xA8JwQ+le9sL0r9B67u4Dw9jRcN2dxphqqx1ERJBbzeP4iZo2O67km3H1eqqiMVV
FN21iPk/yOxJXRG/h7zsWeRwfa7Se+hgM/g9EKM+Usbcxo1gMMmOcb+pgMVRJzsg
RrYWG+hNwMEA9gRlCKcr0BiqsbEe/hv9HS+aNHsBDZ/xJFa3g11wP+ws4t+D13gJ
jy6kCrBu+pAMaNQVJd2nlwaMgQvh7kpjFJ2+uL/JSjY7oadySzyYre2TgntueV+q
H8dukuG/w26+b69POnOxS1QEDa0NOpmFqpxlHbXJZZvNOxWn6DIzh+EKynqUvAHN
POAlX1j+qhOsx+uyL6j3f4nvk66yM5C/B3AXdm1sLIT9cyhRu9VVfb+hTX49CM3J
+SJRasuU2XaZIveq1MwHLGuNAe+Y3PwyVzMl/x8ISC/pseGAG4FNQsN0cDXlM84W
3tMUj+4tGxDl1kvy6OWVa6Xz9h6KEzg/G4sSJUExlA0Vfq8YP9UhNkhb+PzMYcmf
eMg+VnrXTGvgFohhWVCPwlvbNOzwgG5pPlgJL7G/ELueSkmX/pE2ya2tD7fQ7wUX
6d2fyPXI5jZMr25dSHg2D2wGL1NHDOHRHokekhx28+2YK1xMTRPYij/33JVV+Xy5
0BbnsXTImUfROlc0X0EhKxBxLGjbcBDB0R0oiq6JJHhiRUp10ZcYvbT3T7Kn6JPA
FO1JinSIP4THkaLBkFE83jLjyxw3dwTwI2EaZFERYPpGV8uAeyZ6cp16LnLMQylA
W32SogK0ruU4G2aGiSJEIcgB5BWfDTJpanFKN099XKil/gzG8/0Mn33PytWfGWxv
iipS2IVPB/wyN6Awinc9kILKM1Yx9ZHGdGt9+cVCvX8ZRK7gIWr8mh0BeGzjZ4zy
sMyT8pDmVjtS3AYhf/FWs4BjP+hG64Pu3Zg4Km9viuW9eguLW8ZTaYNPGotTj/U2
Z9LhkW+KEiUS27SP6zTAFUF5nUqc6GfWO0qxt1O7ofL9dIQgyqTGtqRsT3WR4dTK
VjeXaW4MLQc8S9+mxVTKIiyvGQHZ1MCpSe+BMDxDWQPvD//d4868ifBvb4YLveva
p7CG4ZyEBH7ur0gOXLAPx4hocNawgrZTs/dHDffiK8vn9dvl7dJMcuLnDaQ63RP/
IqvqYXQoOvnc+BgGtV4sY8ukVRiTE1mGZIRN0CAVhkTPWTJ4J6ADrOAaQ3N/sGYV
uHpxOSmyoI4WFOyMo2bY4SNAPLiXU4At9gB+s7Qs08Swi1vkZo0gPkS9vKCQ5UZh
ff1U6a3hSNm4TVx+rXyvcnaapWrsr2uikvVaDARlUudmmkHOEUD1ivbm3qVVWzHj
nhqXt83Kw0BvJ9DYSOTMr82xBup9bPqCAgbdItlFYV2YMy9WItmicHBdIeDwsqQ/
EgUgkXWUE9m2/zAKx4ymlNm5rsbpF370j7bbUnEn0lGw1iWigU6x6tF6bzWeLmvJ
pqQek+3zixHOh/Ddrsyo+qiOuUJfEnkfQ8h3umzHUkXphlY6fYOqMBp4kgENo9D0
an5u8q6iS8nGlrC6FUl4CcJC4A52G6fPYrnjQTv3ipaCZE2F4YuZpxN3RigaPiWE
RJV8ucl54FfMvWe9rECisIn2X2RfW1bzlBghTQKncwf4YmwmOSJlUrzShfkd5X7V
XFKdISKxUTLLWmm2ZppGcOsRrOa4M0j4Xzsew6PQvVEiTXfEku0LIx8NmjLphM+w
Nw2kah2dmPfP4otrBrvHQlCXR9+pCnVAlx7dTiXqNnuBt5p+NeTqbmLbNOwnbmWT
OpDf5m+0iSgZOhq3GvHgeiGwBE8+7sDJn99aftwogUxRJiAyD467Rg2zWgYSltGo
FPz70gjfEIRAbvwhi8UterQt6/Ge7ZqsrcOvpQgyvqK4CUEjrWWEwYFdxL4u1TuS
DE/dOhPhhAWey8Af+OgoYfYNLkIa5c9NuRBBlIBA9je9aCZPfTlxD8kmqyKzZUP8
B3Qpf7afJ9K/dZ+++slWmuTbtkojd23Jrf4CdGorbMnPcCtafhQCw5hGFFg9qvmM
6wImZ6SJIjFwmiRG+qNaXGJ+i91S2vS6ZtklQrlpl4KaDNtSUa0VIqYHjHhVBQmk
UPcIxAJXsOTmyyWtb1cUhinF86gPhl4zU7xKHu6K0Klz/CMwrqKUtqo7nGepgMsU
igEO1SzJ9CA7mIj7qORHS+LcvpHIIF5EEc5wvbbuEVQNvnxqF/xixcekln4oxqqz
Y4rr6IU7W+ZMFhPV1nNIViwxDGUHIGZifFepZzEgaEpoUiDJ+oU57Vf/w9cRa8Fw
+kwLFdbl86Ro1S8GqC8wYoL/zc1VTYgo4KEsgga1ZyodLBqkurR0dHbpVNAg+2bs
MMo/pAXTmBvTSYBsvJ9SpeDbRCg7QA9Akv/Vl4Nq1Ofdd7eubSSkOZku4eIvxhw+
8ypxJGnv13Eoh/1isfKYsBqENm7c7LgOI7Vq99YuZ34lwgZrDgYwxowVFK/BD2Fy
SsxUlPNToyIE8eo2QB/wR5iGsOe4i+vIKM721BWEzk5ax380KthtugTV+9UG2H0R
1cVh+balDRcq6RmsrYVmDVrsuWE2GaOkXOI4A3WBOcg4VTYlg9ri5Ydz5xGN79nV
vqlu5d/tGma8qwJRAP3NSJIZZOkogQITH8D3hxO20oEmGK7SH8fG9F3WICi8NhsT
2lHadwEZ0oAsBRKcYAgV2rf0YRWAtsVieRfuyhiLA4RGlhl15/t/3C1eHylw9+H+
6cwIC/vlt6IOLerlGeaVvPtLb0y2jtQ1g3MChTYCRLVx9+y2BW6/om5eR3zRdRlo
Qj8kJi5xZWeOHEW9VSgfNWMuirs9ok9BQxzhZLuvUyqYHhiUUndq1yyjwq8kQJwZ
AdfjildvnWFhMI7Dt087WEpbWDrMpjHpuYALHlTFxRRpIOnrVYnH11KLUZAMEifS
N4PXCRx7bXhLAOnL3K2dAj/KUXoTSmiWm1VZpp7G+EELspIVyrEwQ2fnDNXX1L2T
NIQwYe05ZjvdzsdueSFA7+kFvrqCySFdY7o3kGOTxbly8wlfx/K9J9kpYL56zvNh
SbOAkojSXx/G0mbwP0Gg2LC0c1NkmOr9dFiNaX0z9q9l9wNfAo34riFXuM/EVS96
+dBavkJ2n+b/jFA7gp8oIWnvFnXACb0n0sk0IMb2ypru/4YNQiK++utJojcFsOi7
gErV+ue7LxxJBRrqVsrJmjFc6Y3L1wl0OcWeimEtG5bkWngsR0Gm4Jv18G4BFrkI
l73ASBByzwjNCb56plG5lFj21/ustkLvBtrAyvw7Nvf2nqgytAhTI1cBfgw6ej52
RIHLS7b0wW1PMf0TJrzkx7dtYNzlr0CXwvnlsNwWUDLOOVLsaQqgEE3eJRvN0onx
cSJIATFsAOGxJknqevklhm1mLGsEVBeBzQT417nYcMPO1xhSgqjhkLK0Q4+uRXKT
UfLEmvLNXwziM4/QhhYQCFN/3U7NNaj5jLWQNUSZjc2s68yDwSVIa2ll0zr5Ko30
Gj5aYWBOwI+79KR+IH+Gxul5dbBtu00l++AuPvREiiCoao3vNOceTGRm6Lc7SFmD
PWPeH1fzHN4Z9ERZXpTlWKggcFV9MwLZEVWs2wSW/vjJszvDYTePu1MxjTdKw9OW
HAo65hQR2JvUby9wan4N+n1QWSZkwEF1fXxBo3Av0Ug3sm+W4PC6qAg4V22liX5/
t6y/NcjLKSPrnvskjTzXxAiUa1JWJvcyKUCKZutlqE8J5vHOYQBcW47ixXgmAZI9
DR8JlN8qYuAoPMIW81L0VJyjNLJ5nUl4uddunwKoLMinQoh5iCf++89Wq4wfXgot
jRvdxGpQ95OPdIz13fUsFydE4jDtUgHkVKG2bGPuZmM8LtsaFnbOh2hn4KLQ43fJ
LREEn9Hbc3KmBqTE2w0VjkXrkDmRL7EEBdH2emBl29ujoEFueFdLNoME8QWBIyQ0
5DXFSqLlEaih7XT5qIgVzT5+q2yScbsA2oSBFPj30na2Gr4ToAQFEwEiw5DO4LmE
zQF53aobvkUiTY9HxIJr75p3nQAVVA77qHvCzNd/4+qrUtnPx+ZLzdyk7v2EheQX
m2/Q+nVNpYhTJDRWmcN2LIW/eaaAvn9F7hKnSD84qWqHOzQX2NarjjpmqG0GhFkk
RBI0j9u8MqP3/zzAsrwYF+LwIJlukQQ4cKGnL9xRbCjjLqNSRYrOVL7JQt6NFk2h
EPAJYY1kWHJ+mI+LUvoRldI/guYOXYm90cRatXU2fQLGknwyptZa4B4QbRtZIRF9
YKDfUjLF053HuLdq1EgOg+I4MViQOVLbZjklHJX5Cx2dbatwpFoX0/Agwrdkw8qa
fWnA6ifuclVcZjHzd6w88Aoy8AWbgKJl1GytpuMnZtKWCNi3GtS4X6oQFZzCBLC7
nwDoSC9SMSdXFPByQe1j2TsoG2H40Pzd424fkFx0pMdzbJEAjVZxf+aU2caezrmQ
bg1019Y9DG/3TvdR5yhjooj38TA/3q1SUtaKrRvdv2xCFOSO42fwlfoa+u7+mQuf
gTUuAM8NCwp+iqVNXbGOPCSUkWnzfJfSpbCmQQ9kHim50D5utb/9eMEVpyooS3oa
0P9tvxgOhwXW4miWeUKGAf232j4OXoNan+ClvmNIWI+56XGyPDJmv3UrOnXGOHHj
TnSt7QEFmR4drwOx6wcAmj07ymgD3M4YBeXmMz99KmQVrNUl7u6rsNt6uMF5s3d6
oBUIm1zDdBMMcw9M3C9KRY6Tr/zXYZq1kCkYoDCSTMtAqz3b9D1XexlAAgPaLIKG
XAYRLDleuR/VHy35SCwDWzbNGxJPLuWkf4N2+EPh02Jb12Ho8wPDcd7okTbij27O
5NfSgoyIK4O3EvZHCx09SADX+7qsVf92S7qfNyYG7KhK6rWzRWFDHK7kERfn1y5J
+m+oBz9zK0dM2Ii2sZcFv8MFVRlg5rKwAVuqhqMjpzwB8zEpQY59eHyLda8N1L8W
8xxgBWT0zTRdXOwsaKpleCqRtPmntxg6x2rIVFeXMtQCteRR3ANR4URNUg4q6Jk+
EmmRoVP2B6wZOaG6nE5emnZqO2vXkl7sXpoOYgkoV0RUDI19tHaFNc3WQ4DC8Ytx
tXRblmAOVgwYzgqY/nZLrhfW+VCZAKD61afNAfaULZmcaR54a4eZhfngQJWhMN18
y33FYmaP6yE/OPtsiZI+KmngF4J+FUGf+RzVQOneZs6a3zPy7r/1b1JNg3yV+L/p
cVOK3WorJAU/vy+69rPGSk8C5fzrNAjR61zRYtsPqFsqbb3RHV4VSlkTkGTxsDfv
fCBDKcv5gRAnVZLVV8s3GiPSX6T9qGTQPDdTR/kJUtgt+FzKmsiP4IUSIrvAWPI8
1HErDS5rVkY1im3VUgC12zq0j5u1AEyX/cRrtz/3J0Ba4paQD88zjL2/rRKchgrS
PCiVaaV/CizgarDsvj/2CXjyYEiE/NBuMYBUceSOtsB0ldsd8NEyxKp5qNIgy7lM
WxY9dtzFlJjI2r33mKPxol/gu+aRUUePQ5mT58h7yacMquWDElSypStZy4cz2yex
lE73LINqi+bYJI/RI1248HL4yg7fQFbqBURBPseCb+jXz9YKK91F26BmZoj5rCvo
TSGFqei7doi0iF6Os3EDpWUjn0EhZGkuw6EwaOC0bxEOeT7MX/wutvJazziuec/Y
kjbi4XKM3XJva3dIAgkNsAKKZoePvkh5rG+2XSuTOmCKAqRI3fJhNFAium19RWGl
MtdPC10gUGuBdaSQYgYpL4CGZoKPwFdDzIp9MuiHuyzJF/i1JdZzEQDXxobAJ7pU
8DYw4G+oF+Q3/6uxE3y9FJy35htFQkdRwIEzoUqzfhwNebubKPkbZVPRlxdmXQyK
vxVXKc8Um8Mjcp8gm8DlmBusN2kaAz9YQ+MxnieFCXqH6fJpPI3c4ZsCSDHG+yNe
XuPLMF3TUDUNcosEUHjMyFOq3pxs+X6QcJvHKKuRDQUCqEPcnFyKvCtmN5X+WDSL
sgxhNLdXKRYDFwhK6m5+gkpjbRbZZojbeyuPwcoSFPPFLZhrE4YwZgpVqF/4yqd6
N1uN5P4bKaCEh7mHGFjPGHxTSe74UxRHHflPALvcGN+ca69EZuZ2rfSfZkKaFOKg
EE+Bu7sT5u74OSwKygjKPJrH8wQCmovoMG7RV9UHDFMsPjuqSfWjlAN9znh1idEy
YjEIDzNjWWSQUubV/zZxo2fEg4pC8qMY8OIhufNAEy52Uz6v5I+iat2ZcSZo6GYs
AANZBQ6OvBhyIj9ZtX3lZvNm0ybHbOj4KngH5IsCLSQLwZ49FpGWcxuo5/3QbsRx
IlSMfs9ixCV/TjkVLMLhd3B95vNdJ09MgKQbrQ2iZS5HWx9ECzP5X+H2W0xeX/RR
GkovBnVM0RILU+BaPnhr4lHkwTluDSM68daSDB9NBy4av+zNHm0P6gJR6DF5b2mo
I/MgxV14iy84RDQpI5uxekmrPbjHfnv6LRYiWam0A+tLLR0rrz07o9ilS/UFdG4y
Xo3YFyH87Dyh17iisy9z7hrbcfJ6j7hcqfBncLiXrzRZUMml2S7eq96zGK3lVQvl
6eN0/khhHFSyZaUWz8BH8jr1vmFds2OE36wCsFrDkBjc/FnbrrgNN8VpobC/xkwi
x8TFhiSFG1pZ31rwGNFtGkOq8LoalimJibR8H5VS77XxEL5DomFj0Y8iva2Lw9Pj
+xmdWj6kqGQA5WYihDFpUhEXKxTkBy7Z6w+dW0wGqRdhT7f06Cf0oQH/T3X0Uje6
gScBbab4TwyxgUbiwQs75UynSNv1Q2ohT0YC8qlXmG6OaLbi75slj7TKT0oWugJR
xngxUwFedjXmShKzqjJJrEJPM8KA/kwfw0xcQK9hjq5loAbpwqOXMKiwRQaylnu7
mY8oQHtPEn+EnqLE7CypwDsWl3I5ZKLpjgGEoaVJ+g8PrlYm92hlT3fclmg8VTS5
mDpsKK5PXvkutH9CYjlaLxOPy2idqBQ5FYWBOcyI0Z+GdNsngi6r99qiobo0DEEY
nUFPp8ZwdSTaEVfHjkLZxq+NLAwMUjJmVAb+5/4pAjnJyKHUtX+y4sJrCVbMYIeg
V2199t/ysmQvdf4aKS22ajgDxJgtxjQf4Z7rUtGsiNiJnThqi3pqX4G8Z8mGBVBT
dEl0nfemKFNuwrSV35t1bk886i46gyOIx++ahs4nMo8hlmK/fJhcJR1x5fOMuwHf
chyBVj30Ryy+0mqEnmZRQjBdbshUVIMrfi0Osp/nIrmxZMHR8zfCsawSlfMhWvxI
OFi4I5rzh7flNAr3+EhxhB7BIRj57pJCu9+hNzEjkdeOySIaYy1cZwbRzsV40GHE
jJDBylBuKkjgtX+H/7Nk1LbtgF0LdgVYNUXw1iPOOsUsjPwro0f10+2b2Xt7AzjH
L6T19h3DQiiWproOtGHVn2F9dX+GzEUARSc3wrvNCJLAiS559riuchLxarRIqMia
TbWOvV0PKATvQUCtg2TSu67WD15ab4p0gumZ9gqi+4MRa3/ywQAwSjGsS57hLvml
R7cveBk1PeTuGIaq1ZqaLKFr7vurlTpgJ7Jh7W5RaQ5XMZoqqIJEUYeyUxd8Mj9c
FboUQbuirRM838Wx8++Am2QltWrey3bjtCLXmh3zi9EXWMYQokawcxu+PjRHAFZE
Vt70UDC6rRBYLDgmU/ZYuUMNwkVfsavUd/0cNucZ9ApWuFoBgDO6DpB4kqckbYrK
MS/k7JRgRs3TsyK/7zh50RAA2+DoHSqXqQH1sTWOnZFkRPnhJSvxD2Emn3briyhq
BUQW0+lyfMyYO+pZhx/CO+mS5F2dyfFEZxGc1IEBK2RAe7Vy1pNoNOJLpbDgN/4T
90YY9cTtXFUyaDKOl8FDeUrwv+teJ+6sh/R6a7dPZXB7ToVYQD/nOBoN79MwLyPc
cOedlEZrGGZpzUUC3SWun7d/doJX0iiCJkcNGBsq+cGGtrj4eJQ5UjkCu/66SbMr
by97ewsO5m+bCHPhpd20KSk2HGav7iAbcPSCwVBEKt6issfXMjvSJeRgg8yrgBUe
F/G64a3DzZrkv/XL1xgsZepbwiv3iEb91giioommoh9l9QU89ytgNcHXg5AK3KhC
bRv2p2MLxjdcDBmTOrWASawElOvuibw7MgT2XgZnBURno8jTzbdHoUgN3SCrV3fr
ex8PWzGlQ8ChZMmMM6ARqKsB9h0yPFvA2V2FTs8ifdx8vf2IjGNPPLYzcUKeAkti
63Hfr3zHaw6hFlWcYiyRVfQcxAFYGghClfOvQmCMccFtKTohMaUxx0S7izlzF7xb
vPnL14BpLQTeU82i61zpIhysUqgIFIcGKcm/dktzPb6TcZ2K0YUz+xzd1RfTIfrL
Uuizd92v0WhYPHfsaY6UXAd/Dw1WjszjgbiZ6dp1+pbRXWbOlwEeNk40oBgqDT8a
RzybY0lBfTlUxstVZ7W92fVHyhGs9ysZi1Uxzj6PaDtusMzEwd8JBuUd7LgX/GsB
bhDRo2k7dmbvo/aTWxe7kDP6FUQSihAduqxx5lxPCoKIZnQ3jAT1bSvZaBfIEKmh
XwWKhgNximw0oskQqMfp4SEWjF+1qV0ZUFyDXdpxcbwBFapNuuTT2/UxcpmzwHEq
thlHag2q08nWQ3ciGaRVTmClqoeXIhmGnTTNYaXyxTYWgo3CsBwYjWnDrNTS1eJw
1xMg5dyGKsWOlMu6hd/7GJem/AvVokpXRjQhXyD8Oyb/NIQUqu0ZdJXymy42Ebg4
aqHTpb/uqimpV/BTI7OFztnNgD9vbXgcF5cMatm6/OCxXa9cCu/JmuberiACYXzA
NyrsXJImHZ13g+l6pJDAEMZhNb8748PwW9gj4Ol9UrKI+Qk0VT+uJlnSHNv3+ayr
euTM4HyvSFwotcCf6yNdAfFoDrTKQdJya1TfPLnOLLyUKzTr3zs/DtqkhO3Nb2yb
qMzmWcxGXH9KJsTLFKlKPZF+X9UdCRuhI87QkAow+37us0/ewa89qYjmSUp5jxNo
qpQ3N0YchGutdTwk4Xqlx8/Mq6LdVS/NMAQR+bu6klVvSfqIFctxVMtXYWu0kRbo
AY5ElZDcvsWDU5nA6yjLhYETIvfhKQKq/FPPks9crJBp5UPlXcpoQ3NEcyChoilC
xE9o6NwMWftHyuaYx2HRGHNxzPME7AAtQ0380peDAytPmkMWQK+bM7vR9x2mpEIH
bf0GFXHSy6jmvfs3G5noQgTxIFuJUafiScWB73YizJ1zTcNjc5Hju+vOU98ddecc
K8FFtFk9H98n8fgUxMAVjltsLbVLkKt349BQznLRxGw18V8c5zAJPX1klNtdOGEg
t7kWK8EmaU9BWrLLuz7jIvQNoxE/ocIN7gHt8+Tt2PXq5Eoft2clP9E/sVrGcLlF
BTl4C8wSy2nVaKibS5eVK2CfijSMNoGcdbF6Lp/MxHw4ahpcRy/7xPKqrDNGNbJj
IT7gcULUqrG2xYjij56Nm4yZoEuhXyn+sbDB3dZOtyqcfDlZglXp3U2YdSuqLln/
CpwjAjc6bJ7ULztIm3JMaguDVlRr2e0oJITMhV5t0t5mHn9cbKXM0RsZzYrcOGmx
0ixJccfLds9kpuwGZm0Izmlipy3OMQlsdpvnXPdI/oeqI173m8yZGgnKaR1ijnrD
TUBspLawaWZm5mnrPj2egSmHeGxdF9oDSb4AMD1GCgd9dryHfH5fyJw+HO0s+HgZ
2fnC8Lo6gAFHZa5vTLUulBPC32rZ5I8Lkix64dIfzUAKKtQzyMsSeWsA+Um6PG0K
8eZQWXtUW3Ox4AXnvlV8aasl3jc+BE8itP6GRVBOCPoHEYFxkgCKFhuKgLiu+E+J
4m6jFV7V9rup+GaYzxC2hp0vQ+5G/9907oKC3uGO275RZZTC9H147A2xXQ7ZT17r
FSXLBH0t5ICh5LgKb0bPBgv4IWdCTyHOQiWTI481gg/h4KuHxeLEQhBJqyDk6N7N
2JdqjjBcCsbxQRJJb7L04gEFfc6Ec1BLwxZsXJUprr+CyNAr+WFVAlUs8HcXy/7G
75oVuyGyq1AxKDFPF281zr8/WcGusRpPEFiCLWwiuKo3kdUjuctbzfik9NOB5Ve2
Q2d0ZGpjY7Y5OF9u7uxX32gOn/RRfHsdOYsDIU/Gh3KFnuCYPop2HJJQolFrNZcq
b5DyGxMZ7LvY0hYG7Lyl9g83m80pQwJhMN7E4gQ5ZJq3bHA1LmQHEL4Zdd11q2by
+Zw0l+HNY3VH5rySFQ5Sr6z/M/H5LpnYMeG0Wlvh/VTS3aPXB37jHRwBTP7kr2zy
+/72jGb/WOvazFteE+Aihj6EL0qCcuaEuM+8EtjKEhWjgxoCjidZjWl8tPXo3FpP
eLSwgdkzIZ8YCn3MQ+JL8eMkonKgQIh47uTFbl2yZLQGhHzbxK+YFTSytLNB9Ht0
V7VjBxM1bkLKrQIDPQu8+ysfa/okRK+PMpIreVGQb4PkGnbGtrFbNbuCtKGF1bGC
HRY+rKaS/6thKdukQO0FUhY/G1qCVfk4xvArI5J2pjPlt3jKrOnMH5VDd9peHx0H
ZNLZrnGedupMKpgsSkLT/k4fouqzDPO/unhcbj036z2IuL5MHpP1mzX2KrMekjDN
XE+C5qBr7w6q0SUuOG9MT/qsAqsgO+ElRXaPjjNZWp1HdXDgV+Gv/EvlrfwxR4fv
ORj7Ui1nq7yn+XRzz/oTPu+8rqJC+jeGgiq79muF1Vuvmbe9HGNvbDMLCiR3IqGL
a4Yc9BJ8rD+URQPH23MrjHbiwWAMLXiqewTCHEl+dgNrA37rzETQQvlhuxoyvekG
SxMHm1AEhsa0VUpfkbpg16fKQhM569C8N+et9pbR3PNVSA3yuR3CmYnJt0GFtRFi
YmwgP201GEB8q8B34ZZASSDapdPTk8TAnFilPDPG4TcCaLgu+LRy9x3A+EHILwdc
/7aLn62cIPOlBM9wHR4y+8JCaJ0692cJOJGK0GuTyUeYt8UQ//kmytJpYgW+iUXP
myJPjVI4/Hvsr5Ulh7qKwegMM6D1HPHNm5pdZNDxpl/AQZp7ffrWrBC81uT64KAH
I4p2wQ3hHZnRiFM4jUGTZa/w8hMlVtHHVX3VWaY+tDh1f/MXMfrjrcUdjJs12Pkp
hFkmzMYSwQNuQO0MdIRBb1U6LdzmzzNzKc+pIh5K5NrHkNE1H2RmdlW6/HCKtr7v
mPiJ928bV78Mw3KU842UbKDly3SgBLR/rmB0uwwFBTT/VqM3eNNPB/m/PpnzDXJa
92ZE6ezQMXJpYAbOuB0QDTEkMfhJ2oaPMgp00SpU4VMt9DXPQ0UaYio4WMERdV8K
DnTqqTPYinvTmfUorY6mfhjF4duzJSeWk/gJYwaQHTv2ayw4Bjj7RWpIsPndwWVG
fHl6ODa/9Yq1urCPbG9Y4F6Vztm4NBJg+0jDeSUKQ+VWqujeFJzOSDvCH038msPM
PyUSxuwlAv1FFfav8TpKl9HBx3dWzvI3FxPKs10JHvOqcLNJ9dSK38p0I2tWqMRE
praijWDgXQ7ZPusJUBe8T+Eo8Puz20/epVIlGQeGWsi8aAdDSPJjmDgJeh8vxezM
ZxTdmuBjgjb/7jHQmcgEId5FBRhDCb9sdfiKwBw0tzJWrhlTCoQRuTJFUnobs9A8
PqwyqkIAY6uITiABQOcegop2GaS2pEBTlnbE29ojJ9qtKlZLyIHNlCkRh7SN5NSQ
6hSkjk8Kdl5BI93BI9Gts/tFiVa7y0MCiKXISW3zkMOoxI6DtUSD8F0iy6guJLeA
xAE8rhXzJ8pi8z6WRjtq+7jfdlzi3JFZxnLTVs4Sr+/4EQTdsSh4DjQWUk+Z6zfw
sjgn2u7/Fv/34DoPENpPGibxkDfbJQ3CH5v8vZEMr4/+4Be9Wu7Qb9/CWGsJeyqp
Tag8vWM+Qql2az41t5HDn/4k+xpaHbUoedvdhrWsrx5dvfYIwBCfIDFJICsMIurV
Kyi4sYqRKaFeL8PJBYrfLQuc2KOc00ni1choQyGF6S0bf//EFP48T93qlb9pXlfz
yFmgE2kpOkSMyvmN9sEOhSv4ZvFsL/cNbUn5tPt3y0v1qcJ1ID5eNWzNS7zavpFS
qpPCIUVG5WhKBbWMHQGRLV56/Dn/swf3pPbPJelOv2XsASkmOZmFktIdVh87DgEP
IhEwGrWiflVdjRbAaY7CB3An+c3VHH5emc90envbYIE30VOfTjqWrUwjX+FWgHdV
QwL0wGYQCrFw7mcpAY5BFvt+Pxn+D78PmSJYHxEEJD4w5nlSW05rKox1DoysUyNh
oJhNZKJNWc9p3hHRhLLM9PT8HM0glcoE3aUk5wgYX/Ls4ak5CKWIiYPFtwceR7Ju
iTZ8mjq1uK/+73MfRI1LXP+w2b44UvwTSDb7Ehmhl79iHI/dIKpIAUX5/HsPW7r4
cw6KnRYlPw0g8c8UMhEtVaeEdQlsYwlGPCOus6TIj2LzGWsMFzzIQVTQ4/0CamwK
4NrL3jAhU2UCzEqhZIj6Zvqh6uwh12OQ1/WYqrGBQlXOYAs3Bo676oJYAzLLSMk6
soPl/nWxKxv5YqU2KjWRr8I9vRHDe9jHIw/yfB3CjwGJkDgZACdtB4t0yPTTgp0Y
sI9qGQdAfnT5+fMkPp174mJoQbbX8lG2JALx6eZjRoZ0JbR/qQOqbkBw9KMF0V2x
mqoT8d1qlYbsIRD1WAw2AwIvStCyN0xpC4bINr5ow64fwbHTlfrFiTKwjE+YTisS
8gJf6LaNxQApKAQgYGReul+lTZjyoQTh0wvzcO48dxfwucWnKC1kT82A6cbOLCtd
BTdSzpqNhQQi5kq/l5PVpaO/T24p0uO/n31XtkG3UQD5Zu3rBVEbELkdI9rg4hcs
Y/dajOt7fnNRCSjYyQpcTQ2l7XbhuBHTL8F5frPSWZ/HcKbCnPH9aSN84+WnY1VI
Q7hX5ty18I2d/1IkOkgZVbSo2DisiTtN2XZnAw1mQPMEG6131Co+0Ijpl9b1kd4l
GfIX5Lr/BEalUUCHMq9tt7pFOrXMs2fbZp1F6m7LSPNjRSryLSmYAoiH9ZxxU6J4
99jdvWlN8fYIUSqiQdTjKe8tpUj2moiuPCd08QJaRAtEKOiufI7W6UMrvyY1mjO0
aKWcHfTye/PKOq+3bAuAXdKdSvnNit5hs0WFE3TgPCZZNqefFquyD/mny+2O8aRK
XRs6tIara9H4Tsyb6nvybbKZsqIdjqZp2Q8XAn86GpuanSlaGD+9mrUmPhJVakRy
EtAWtxDdFlcpKXLADpw9suKQs6TVMccWPIYhmm+9x1pGqVRPLrNqFlwhtbiYVRhw
OR6WZeDk9mf0H81+l2hJqkteqaQgAtx01fYq7qp9xGOQH/Bv7WNVhj4ZwKD0HLuo
eGxkjgqEEBvpC92ILgrArsQsxtKCSUFvSjRVh2PWAV28KABiEPxONAR8dfxzYViU
a85mSpqKbcwvaNJnCEevajgZQj2SucXODusGXJlDYJM3Jx+qMuxlM9Te/D4Z8Ht/
N+XIaIH3ouwwG3vDiyuc9JQMZIjnPrXBriyp19m0HmXps+pnE7Zco3t5bmt6E+U8
TiWMvngLL4pOk7TkW1fm0gou9T7goRljFgRTWw1IKky7aFF+UuD8J4xACLoL4NLi
co/q/HyZ9LlFTmzc3uVj1ehBCo4titgycE/oi3gnmys6rUbuZTzLNNMIi2nHSgUY
o21Bl26kvRQ6Fht1+lSe/ll0Vs1N3ohbs+vgME+654IF4BR0MxbHxJiQSg9N1UZm
oeLZIhlb1B1CFkEkG2WBUkapnsJ0Ul/iVtaG2fhEB+z5YWGVZdiLxTRUUharEiHW
qmcmr7kzk/c59JdBb3lKuEYMBYZjPMr9e3ycvGE+v2KEie+jycO6qufy5t6FBcBD
EK3QldXHhQ8QkuSE5ubyM7FAV8Iq/0lAdUzpN9/AAWW/dOory1zfV2fkgOUQSFJX
+ZBP6G9ZwuJZjBmkJNX/dvsQVboeMjzYHBL12TrvgLDZVis5bDT3PIaFFOIRlrvW
mUXQUpk06RDwIn/At9a5jekAaxqfFhpqmnzNBkBbEpYQsaG0tlhfuTEsh01IaGvN
N+zkSGSpDwfpb9RoZTDbrwkBmcKb9aAxoGGY7o0aIJwUBia9r/NmKQyglJ9dbF/+
33Bl0yHh+Q0vr4el9Wa45E3CtJ+/NGnHi4lJ0RqjnCNWgt+IRdzcc1s7yI40WYYF
WWnmSsLpQmjTi6itOEgadz/ixtnqlLqEJgnYsj/fqHksDpDTdixlv70LyfmDVHaY
bzmutU689X3ZavgUj2QQH5h3ZHw9P4CvIAwNspYn1OZqJfAR8jpUKPeOv+ZKeJk8
bTlmdSuPPPa/YxhWgQVnYE0FwYukSm6IpWSxAS4/paDlpDqz3Lg9IvTpTOYG+iH3
8ZhWHJOZddIsz5oE16WKtfZduSqQeh1mnOlZmnz/1JlhkM8ierBLoiGGF3dVvun3
PvbetUicqSMLpTSLyTYy0z10JeUvX3GraeTFhcYA4ugK7o/ATDRAFpuddm17zrF8
vt1U7eyUPJCkiT4BV1bGNWiiF4eEPEfO9yS+6+9n0so9R5FyE4ndoi2blIGDQiuV
PbqLf5L4dYizX46GgFhFm6xioVQKTb6qeUfw/JPlZIq7QfFqAuUJaOwUO6Hxp6Zb
pUImjtOSoSne/rplp79hE2mCbjD40kPDz4YR23i6IUl8Cpga2VXnflP0YVxOcpUf
huFRzPRMBCrZhplDQk33dvnzRpgUOHAQ+bOcgiCDZUX/jPEUZK+A8KGK4NzT2Pp6
gNaONQzwDhXrZwUlXdVUL+2QSw3HtvrDUzSuy9Q5P4WY6qdUj2DstXeJf338R3Ae
PvWQpFpPDT5smeW7faS9PXsYt6coE8NL6bbfc0tFQYujjoC3Q8bADW2jxdjErc5d
wK4MNu9DHJnClLAyW8wFHWl66kDWOPTG9AIhZ9YLGN6HJP1maNBQmRJBdlTffmEg
KoMS5kUbwjf0izaIzufBoq6kQmJjWSCDthwxQ/j5a9TuRn2KDMOatDApQFHuffbu
zXP4POksXotZPsz9BwhirtScf5kPzR+vnD40kMhShuZnIc5TpHUdUGSs8pux3Q8g
0ziT/wgf1VzGNCTq6PsSr+vV2mGCFki67W9kL0RUHGUU0/zOoXwodYtuL9RVLn7g
KtJbs5lInESiD7DpFJC4GEOm4uuJ+vMmR6y5TZTpkxoRE8AUA5VeFcmRkpirZ5iy
DHhvGZQsTjR9HiTaWIPmA6UjdCXZE3Q4fig7tjGlw9LClYV41KG4pOW19SLcNQRu
6hFebfkKu+p9NmCTvzdjKMb2Ul00HHNMLQWyQUHWNnE50I8RoWAaxk87n9SoQlFM
mJourrfN3VmzOnFc0WLsNUSi5HXZ0cnvm0yBfcvilN6sstDIgM7bmXBYGK7YrklX
weVVs+m8skpOVvvFXIb4IfLQPDqNWPifM9CGESWppa3VkhVfzwH3Pw1YIaOGay5O
5hVMcIkdmMQ+DGTY16HcN2vr2IhaK8/9LaIfaS/m5RAuzWlUGn1C6naFWDPdbLWG
/IRjzIO6IevxLYYz+ovggU3k8F30oYzLcq6t6bkXQ87M+z1HrkJkqEaaqKGAK7xF
MeNTYy4Oo0XZywlLzzqv1PsM/GJbcNZQM5pU+N9Q//GGPjgBBOaA5oWj2lcBIEDX
0wSGV3yV3UHwV2a97Hj7Ayc9/JtH5gTXIGHRINNZ8hYI/Sgqjx61DsExIx7GDCdx
i33sPpfsL4CKNAb312nJb5b9SoOZ8dzymT/WEpqvJIFo8lbeFjlIJjScNITkruHz
0s5I61pJx5O+lEJorR/glN8vgmkVGIJ+a8+tWRB1zFIxe8Y3dJpMvQ/N8u4Q+n4x
0g15xR8++pYvzl2oLPxEdd7zJeY/kPqK/wnqrS4KRbUoGDRUOri1QZO4uR8aUBhj
AZ61CxeYHSWCTaTQW16QR34tSoijhgzrq/aKKlCN2U+BBlB/Oh5kUe221kCu4ADH
DsEejBTxb0pLhaPaZqsYt9mF60onfwYj7M2ZcohGuiQSqYmaSJvPkke5tjCbXzPp
8NFjbd1GAJG6Yu22tBfGX4oaPbWdFjmkKoIm+lbfoKoRSe01v1XJTNLs8J5YOrGr
CV/tTdl6EfINqeegCsdzIE+EYpiHSFQhgrSPgdvjEUtcFq3yubM87lwi4NtH4IIu
`pragma protect end_protected

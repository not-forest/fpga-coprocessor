`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lR7JxiLrSoqRLbdgnHkACmNEhjQa41ql1T8+bDH5mQKczYtNII0pWiEvxzNmJrSl
jS2GkzpTkAOxShGLLdZRWbIt86bedU8B0K9GNK+7dU5PJqX3/g9sc82XEO9/6PM6
VmHzwKG4c1IEPZln+NpSbSqbb22wyxBo+6wfNNlKkcI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 52432)
xFCdoY4JVT8tz6C/YyfaDs8oUc6tdAmgoasr0qdF29rrYtaipncNqnhFOH2QaWAk
5S27UCM9QDduMkP6A0mN12usWVEIZg8kNprEcYNLFP0Atgm418UY4nsfY+1CxQl6
eEu08GOVlYc41LifkHg4KnEkvA4d5PFnaJGMxJcqwHLiAF2rq33toEQ0L+sj/JbN
MI0vAoEBRLiFV9Md45Jq8QFgja2V6lmd+oqvYNmVsCft3+QVvUczPZY1gkqmbTnv
Z9Vc3EZUS/aq1sKqC0aceZV75rVVWb0KluUUVIYQw0wm5/RQjFgSfGcjrWj8PDJ1
HZFxQcxZo1h5uJJNe2nUG1vH+wf+gWNv/UO2DU/RUNljpY1NR2uWt9quGIYpqrJw
r3i2G/AHJ5jb6QoBzL7Fo5v1bjbwTGDiBYoL8iIZPqxxXJ1pZsJNLq4GScjw2wHL
H+FFADhRo/sbQsoZepcCv1Ct0l6eybFMERc1bQOdwfZDFJfLL3yGTeJ7Mm2XsgEP
vLvhERZAuxpmaVpb03a1tPLlOB09yDzAWXJII4/7FSonj5XeAb2xqyFS2ndahWa2
0DqW1JTVLDzNHRd2VNc8tTcZUIb0fl1/Er7HImXjQSwExI3IjWrJLIhN1nZGhpkv
mFnJ2/NHM/LnkuHWbGcoTVsltFyltVswcLMfCky8iOfR7x3RZk0q4YhoJ8N5K8zq
3fbZErDaBttj46d1VqqLXCCYO7ZP9a6B9fGyD2BP1nJvRASCZ5idXY25v827V7vq
OKExqDXN8VpkI7kxkpGlbGXsri5cTamT3Y+NReAlYXGObZdc0gCkTrID5KOQtCbJ
NEQ0tFAd6aIVBGd2BBUDyK/cxGTAWMwT6rklHXGKua9iTC2Gsan+YzB8u0azaH0g
bKseAamxq1ABAZkLzL4aaPvrcY4n4TW/GQugJ9Atwz+C2s44FAmu9y9POWPStfLp
bIJ9KobW00Km/a7UyBd0cA371Ng1ZS4T22kP4fyyKbiFWr45E2mum8B/FYE2lqNs
zm6cc7rWfwM0KPVLb5z73C8VBtUlRzDrnYjgxesGzK89oNAzGdSlBKHsLa6kstZ8
aj16CoG433cxd/FP+QdXMEPfxt2EpOscQkqrVNcFacAeTQHCoy1CVX3pAPkj911B
qdSVfmSollIKTsRzFsFJGPRFhMg2EuXxo0r7HLnTmxuGHfHjRWK7SvqIfKlyNl9c
bTeKMfbm/fIi64oUi6PQ41aRAcxQRNLe8h5DIUwKF2XDSSBtGxu/5OKGXUHFYcui
fA94ykHhLNsnME8VDsgW8gBUsnsEK31CZmqUpME6jdQcdWOImjSou5fsE6qm8SUY
VNxFefm+TlCi3PFBYinVNHuomINJ/DDAzKJSWP5yTjBrDRgwY9pRlifr4DIiI9Ia
sJwVs0sq39SPxjtEjSoxcJX1vEK495QG08TdXZ5grya36XWYde/3C9eRTi4PYwM9
NGu0TMM520GBEvR8RMAcw8TlFnwXyWRTaAicyRmsR2kpeS/uV/7nK6C/30TASX27
uV2/brZ+iKiLBCFqUr2pRXbTyzT/FMkeOK0UvxqGA6f3QowuFxT/xK6525ykg/Jg
tV5ktdy0D8ExjApbHfbNLIs0nzXkMcQTS6sBVFnfP5R4CVuYZWzV8olxm7TQvHno
O607QmwC+olSqNJQSBU7d+CMXSYxTZI79AXKOhopJOPHYusLHCarPTlu4KMVtZL2
6dIGViCL/AyheuQcFMar9YOn3mg3xYkE3OhpToJ090BVsjudEjkO2Q2mFzbuG0ow
OnWXr+JtXfmyNzCjM3Q5WGpp7OMDa5gK4JfYunX3Z+T0ud2BmQ1j781mdI6lq5pX
BZoG7d6h0y+LlSHEF1R29ftF6MNtxvYSTygNme6P8B5DwT0UDVutnT2Jek11s5qh
ELq+jFEHITpyH0jpyW8fqf/OKWCWoimqkBOoVrO5pMUwNKq9Hjr26JUn8puscsCH
rfma3Sl+qWg6FdRmC3fNjti21ImOPZMppTWlN135P8g6OysLB0YZHf1namnbne25
oZXXqYPcvk1NZ3eC3Qo4/d8idNOw/6ZnCq8fQBxjMSG+bMwUEkqFXpM4xYW3IvmD
gmMeFX6lH6IJWcmFNn1YmedsCpCbsXylo49KK1SyI2/zWu5g/cZSaa+UhK7qnfrY
F1eyaR7X2I5539bhzbcDvscdStDQD7CekZNV6e5FxsDkKeWOEKYMGX6B1+jq+EKt
ysKKpKlPND6yVbWEqFuDI6CMpPlfWGGZUm3X1kNi2AhJlJ90L4VZalFFEGOV2lkF
DYUH1BeRaVK2qwCb6XmP7Qw/ne0NWKQwkJMAMByq4FHbBYqMlUpdVJzLAV18AKuY
mU9qnkx5H+IDc/Iro8AcCxQA8Qug2Qv7Ad432z9Uv7Cuey7oeWOyJnftyD7iUiBB
wiRzYxM7orblaEdddw8DUl2PGJbeTkYrrBgeCJHPZuEAkRAsTvQrVhskrNebJm/g
aMBCTISekgaZNVFmdc1vdg1xEmAz06Lf23YGbHvDwB0E1Xxy8LEAT/nieZjBmSeQ
pC02u/xSRiaCfMEj1Z+u39Y1/XinhH+HcoWNtxDz9pqWZK0g28EtmCQOCWD74h3O
FB0R/vhb/h3cT7R5wDCCue4nqqP7UhdC6EARGSEyi7U5ufpLsJl3Lgrl3crKQuRC
awX9TVC4J9gHtUs8O3IV89/bwa2X8SDdejKFAiL5ttkc2TiqzcSC4D2vgBqQyYgK
sIE/Dzx05B6YEAor2jhPa1zRCGhrANlpu8ACxJ44D7K4Hnco3Yndl4hfPIIV6wxH
TETKDNtbCijWncC41LCMk0/Wx9ghJgu2cawyDbbItQ8W02ZDd5s/GwdHEPsksmXB
5msWmqbJMlJE/Z6mLm46ujQqo77smDRSYv7zsUAzLGnL3pXhTC9T+kfRFeU4zHMQ
QhngUO8X6LTeRaMgEcVcM+ig6jZg0sDtSCafAJIOFjTAHS6lLVF8JIeSpnQj4pQ0
Yc2PLPnwq11hJIvNmJVZuuSvFchYRkqoWGYvMyecQMTBeMfY0Q+AkLL286SMgfTu
LhrZkXDWNOGhMvphLrPnnuPZXE1GSY1ldu+5sofgPin0/kF83Xh63UQsE6CZ0xFc
TFk80yLBW1eW7uSRJ6jMYxsOlULb3WnCNuffl7y+wxEfDpkvu7BH3pBjIp2m51l4
+QSy/Q90tv2uOTRHsk9TU55d2lICBWVVtLHmc0fE3OGvqpqWD9k1QyYfzdjjWaxz
SUiPPwvOa8crt15qBsczLPkUlafteRRx72dypgxLPQgOsnzdGDf4RNCKJCOt1HD+
MfziTQ5C6kxdDGY0SYlDNlYaTpZQoVgjFIz05K2Ndi7aIrG+8micGHVzpg+lYeqU
9Ao86a3iQMJ2OTljDCD6wDGxEh84V4UNR3eUnmEOW3MtymxsxPdEbZtoyz+L5SBK
rRi2kRPoTjOgBHC8gs0z1+jnBoL3zAj8aZubi7pwi8k5BZ9BFOJsiDP4Eyq5lryZ
XVEV4ZLrx6XrOX0kGPVS7UVQVJoEfODlRYuiqyl9t5RzdfGrFsW2zE230otZCu3g
AWLQCm/0MhspyFjccNwkTfTdshXiGceJKRqP6pX+y0nWy1E8/KYqOxY3laEzRwYr
gu+/bYY71th9W8lKGKa1PjLcQzE8P/kChjEtYacJq5huTN3nQ3vFYsV+O8ml16C6
lTm53gtUxE3Bi7NU+p6qGBQyGmq14jefbzkC0qiH+jgTmJ5jrxyX4/xWdu82BB6/
KZ8q8QZESCi8Ttq2jxJMkbaqwlx8ydQAi2v+LrznIz0mQXeIxD1Htofe+kAKko7j
32JwU7mwSAebHmOtzzEqJpMozMZZpYMTmjIedTQkF9ZOgfjtruGrmynUqGs25dVU
jPkrJb+et03u8Ne3k5DVVul3AbBiMODMZAHYwuoC0NoI6UCoptCnPbfFCPQypCpA
4zIdxReWl40Qb+PCEDRdKP6fAtP0tALCFPyH0u9yIZ2LvY55CQvsfDCuz0oDcSMQ
pifX1eEqddlWCFvd6pWPyMm8v1oYS4soLfdHhg5AVq9r9t1UNxWOHV2EZ7rE1Lx/
6ma8cZreEdNvgvBR1RrI4eSyugfw63qN/EzHXzR6sdJFyAzXsNv0bMeyDj0+bj6j
QT9c6Cq8HbBYhKtLrWwJRBjfj2iF1wQsDyDB/t1gWHurdG3YuwUcW29toxlXbs5D
EL62MpODM5b1DXAWtF0/z14FJGCdOLA/mBIf6RO8+clAJKYhYiycyUSUaJpX73q2
PNmTjPTWxlznBVr490ftVdOHBlvCRCJtOT5vRS2JNmXqSMTQRLD2AMLCjyTbqRz9
Q2t/Mv72v4FYyOoGPKnIe3zwBlwOXSwzMTAGSBPIu5klxTETaQB1HaskPfq1yZNt
rRM1DdxEqQxA+ehK+BW6ZwqEJZM9Bv89zerZFzOecdXO0k8SC6trqL/ab8P7ZCVc
KbfQ+IvQRL7j9G1apD22lSngkkTbVAm5VW7SR2IrDJBsa9T46ify01nUYjtuTIIL
h8XTl4a4fs/btQ3tkLSa2FgYim93I5Ci2eBTbhQG3S5hz+jMx2mWq6X+P6DNsrpn
vFMloFw9TDZ5OwMcSpZeoZAsZ56Vnisds/aXjW0xD/HhOVVMJTUaV1vmxIqN0UzI
OMFhIdfRQ4OGrKTpcuQRDuE8bPscvw7K2AO942jLt3uj9I9rTXmObnfSQ4K9VQAh
djA4ehmeIlmRHrYurwMecKIMhkuSfURyqHWVZrsLmyEUyr+thUAoTR2wFDsty6n0
Mm6pYdqjud/1cT75hOE/s/TUgYAmhq3Nr5OI59/MZpZMuAEXIPSMgvClaMOqp4Rr
xWsr8hfhrdkhJfbs5X2HpQxFm4hMNvm8ZglwEGl8Q4MF3GAuvJq/6vK9rfDpDgIM
yNepvcnAu22Gql8sASHqu7FwgRRpzFeMSKmAQxE/limIdFBphRhgvGuwj7a2RnsX
zGay1vtyr0UfyaedPrJKlvG6XwraPZW4h7RMfkWCfMyQdhFp6O2uR3H1RkAhDizf
ew/xsZ0h851UGxGW1bHU2ec+tgH1d6P4mSC1303scVVVG9yTuKpQ7AVR/9aWC+LM
RF57E7j1RkWAkA4zz4G0+E6zlMi2/BChPY4esEe791iGWaLvJRgSgKrBXdj7M34x
oDQX5oxx35K0dHNQRlD0FR46aM4E75+QgrTg4PkJ+iwCCrRtUdDa5bQ9XN6NkdrX
t4/Or9s4/EpTRwUYjBfCjzn1s7pUyP0fa0H/H9D9zWD7D9R1Sqe9apWGvpFz/U19
lKEgavNZyS6SYH6wC+/k3Qgt7sCEzlMUgMDqj3Kp2POBAzDCJfjjhXb9KmpM+NGZ
rrEyg7oB4x4n/bkSE7xq0YBnnwv8ia5C8zo3JvFuKpxRdtAA06iEexwK8AWHb8p6
cwuTd4R8UHyaqtHf48pHqNck74hCCXeicX/pNgIw+L7ceeIQNE9TUZ21NfWhC3An
e/qoesNY14IV8Q49WyJh40ItXUBnl6Rydr3F96osJSx0yVMGkFvKs6fPqpSNlmyK
4RqEpX8eUNZ/V8yjza1quxBHvRcKsdq02hetPlz4dt/je1PG5ZYxG/PzovHFVoGU
COTDDBloLWbdxVvX8bK8V1KOFQzhg2vWhJzv3aPlL9y7t2ghzZg3498W47FP9lJB
N8ldAjNxKReQGj2atfj6OYzC7R6x75t9tV2YmUM7IogqvXpnXHkPiyZ8raKrbyFZ
EPXQkB537YQ/XSHpre38jp6Zx26mhrlG47m87qM42d/DQ+8t0VulJNmld9N9aQ5L
UzucmUnxzucsos22ni3BdhIPus1nnO4y1xGUy3VMDDvt4mAiLY4TurLrupY0ETtx
WGfOhqG7lmHF/0WUYU2WvFfSm2wd+qtiXT3t7Ez7SPQ+98qTPqShpaahpjyjJdDn
sBKYfYXOYgoeoUUa74eLhWE9UHrf9loP7ghqtZd+eTzRvz4GGZ3xhlQ9Juxa9JVi
sxgxSGwVUs82Pd9ewpJguG/Tccz/swF+TGTaHsR0OpPMSJe/UwERh2fYGhJhK9/l
hlCCea7SBhOAhJneH+E1b219OazRVkzc73FCkjKakHhiPcTESS3hzepzXcHV6C0e
GPHP+LiR6WgVFbHOyjDeKpRNniY23V6+w6DmD7Q24vBy+9z2/6hgljv57s3MtKe8
srLqmdS8w5fucNUuZxnVjPMc4Q4ugObXa9AhMDaA7iIFkxw/Xly/eJnorLf6KkD2
EIg1xR03mv65b1SoVcn1gECF6U3taJEFXjMG8IBCtPBqYS2JxDMmsVT9yT9OkBQO
bv6ouErt+3da9VtcKNMIlXe0ykTkIpqwWYVB6PT/0L14eZFnbKjFW93cEdyZSTkz
sFDFhlDFeFln9c8DGun+1/6q6stb37bWoFEtS6vtSVqx0W6F9jL9cnGHB4Hd3aPb
hmp6jVDba1ux8Fm92x91LFePk0taSaBZ5d7FWbiaM0p0lFhcFzZ/N33WeR6uaiUv
bhlugIkaf3UtpL0CNGTrBtb4CMkzDWUy5vpRCYJYUePxNyvHrUVRjMw1sR2o3rge
Cf6i05/OTn+36NGiJY2TVWPAFF+3QB/dhGma/tsZtHJrBnLSDrwpaI2HKHS8L03S
RQTb9aGOVjssUxcfA4+qlAUFUSliMxLsiILyaxtPtX4aHpGPBMSOxnsTT96GVSNl
ZCyzBXeuEfrNT19DRmoH5jTWoeub4ItUwGPM+Xy4qbeJri5iutwnBpNN48D5Fwg0
XT+ynHXlV8iGFgdAXwNlpz99kM7OiJF27bPibyKRBOm6BdkpdRROLFqSVS3sghyn
mVpm/WMOLi3fRc3encv6r9ba5VK9u7azSLUM+kZ3EzoBefSq/G0r2B0Q7ZfEktPo
8TYMTlyP53bQt1U9yJlm+5WMm52SoLfdJ9Ezw+ht7tKXgAWU9dreyFKV6nZA5Jr2
kaCrnxwWp4/osR/OuQtjkgvMCvW+BqL8PlECb2jeLIfh+PofX875cEk0rVhwBGop
oZgXeIqLZx9FDV6j8SQc0Ja+GTBpwukMpD1XoPJgzgynvXTa/WDFGPJdy9s5Ki4E
/QRrnp4wWeYnIrzdrKooMuBs2OA7Yn/5DJ02CH23QNh2S+3won/d30fDDWiovrcb
iiVzjjJTpKMHY4lVjIkzDeu1h7V8/275miLlIrbLpJaLtP+9vl91z3mQTIoLNClC
yvbiCXmG+Owb1XWR1hzEcljIB1tGps8DX9bM7qVPWbYVTpyC2IvrlbLVwNrjPcM/
h5kC8knHZMtbxN3xdh1oDzr4OObU4fVxb5sHNCeoU10V3KBO/2Y8JyahEQIfT8Yo
Fq9OH6EBMbNgQeZyAbQ3dcqnIemZxKptrArdoBxVI6rB+DOBS0m8e8iLTlvExTRD
N2uKf3bN0z9Xf3IGNEt03eDWEq2RWrURSQCwk3Jy4DIwf+Qg+sLdVFTcJl7D5Xbk
+W4SCnLnxb4RWiEOHUEGwJ8DgvAAjfsRic+XExDJf7Gm0QvrhhNiav6T872MNiPx
YNxajl6L+QPpDT3nV4XXN2NyVBBGbbXVCIn7Bkdon7BRDXWUNRUklhU9lMOB+v2p
WaHnONd3v3liftN8JnhNArBmdvFpWlGQ1ZTuxx2s4WoxBsnDd5pLnl+FyrkCrPFN
zAWn4oeYKPkVXvll1yB6UrKflp7yM5bOUe21bL4tEGkAO+CCcgfAoCheVHb0lJ8D
N/3E8GUPUeBLI/TJlehTONeiQvRYe6fRFin37Xm6rIzgdbpZtHjERUnFz6QB7eIz
2pYskqK4XBfXRUt8cbIQ04TgS0WfY9cxbRis9uenHifD0ZHXx2hH1aoTY8Aksp0F
CibtYCFULhhCYXhK3sWQSelHGebCtgy3Q3Lp4GhgVsLWTXm3uZPdGd4mi/TlPKE1
PhCUMpOo3Gnx5udSIqln+Jvnv9tcwLRO3hw5OLiY+dJvlYVTO4WI8IhRdQ4Ic22H
Xs61ICLEGxjalNPQ1xDvr1PgXAxB+mVF82gks4yjWi4SIT5SHN14jLVClN8d8duE
OchxS8FoesXrNuhWS7Xu0ggEeqNsaIr53F3PJXORLzoCUCf45IHlNU4QzSx3iUFe
cqs7Skm1bEWr3GDh2vEzHgJU+sNk8B5ZvG7aeHESAcbX/rvTVrQdNi3u2fKTGPzz
Irco4vcTXnOmPE9JBS6LlGNvo5jeOXoPkrjIZxAqhRHEH37y6l5lgg8s4wSdxXEl
pKC4GY7vB2VCPLBPUlR940Tb80qs3pA8irA5nNIywFRMf58iQuybohWySUlfivWN
ox5XqCx+APxvrz7vPUWXHw5dfuRPtageuvvJgmAmOFPwH/ivvlkmJ6fgp78sQ757
bJV/r+l4x7NDvqVE63EgoXmrV1b5GNNmr0Szd0pzrb/Zqh83WKvz1Z+FCYSVQu4X
PezsqmbmiAnj4bTfE0ElnnFjAtwRjrKo/tohH64rI/LRtgTe+9m/xJhvjcDePcHT
MdR+gzv/WZnklhSmj2Y+o5U2F7GWX6fO8GpPO9TATq7Wj5TZ6bQQJ7/0rqN0Tolm
2gSC+OZM8h/yBrkB6VTm46xSEk8czNAZjYyULiyEum/rpMYsKJDmDm7wSqny/F1H
mQje4EG5PPMDAuKAq4g0aWII3pbFm9AY2hHk15sjM5GEWZKwuYyrqsLB6oXQdFl2
FlhwkP+2qeYGkC6Xnaf3AvO1Wb/OQDlO+qG1PStuWR3IK2x1pvMu+R9RjcafzC8K
4+/HsnIt1s4UrliDtXZ1MIIywnmfnPphMcD2UJ8p3lqnnLBCPJDRxr8x7PVtyXuS
PG6HPpl77X4BA91HVweyHBBe3N2+HH3w61MAysoL474uBc+0mVYmPY6j0bj9Zc9W
y8xaEmlBQUK2F8jRN/PlzRnfCNjRKXMazt/TJTPj7zgPY8WQc5rZLV+Ll9mjCGND
bC4Fs8YGcH04J6IoN+cHQZoq/+WfjxUjWw3J9Er6nCDL9xcN6go/uhL5R/yPPorV
bhx2KrsV6YKSA1iGZ30cpzIfiCvJkQ5B4N/nT506lQMeBqsIgoe2+w7qh4An5F6r
7kLqmSuQrE+bVbpL45aXSKJWrbS0Yzq3XVAFtN1pftK8Tm2otvAOItZUs3/xO26u
c6LnLVumYmHz9/ohQsVLGE8M9THFv4uJ2d3+w0upmT9psYiyi3Y05fyKnrBMyVPp
DtNiuRlWDGQGEHUTm0iESyimgF+45Z0a9nx7PYfVfBdYDtiI8hTr8UzCA3vYIrIl
KxOkO7HxEkec5VRnFNcDIXj/3M+7UKehDphbya6zksa7nJpxysoR7sKs54tgS+Fq
x3TMe+k7jp4CVG/Obl/zvoSKs7pPfzUKoawN9QtEeUmIecFMfYL+25gkjVB7rfP3
RZ9B0wZYuvzOpZRYWm7L/MeOh/0OhtIRU1kJRLcLpWuKdjpX7CDkijBKm+yuQmsF
Q+QxO+rr2hHrDrEE18SlswEYLTvRyguvoY1suZmG4YofeypomlCZsdzFhbR4YxJc
PQeDD9Vzg3pGsiBmCM7DmJASJzBqPHiVR24h/dqzZ4A67tA7yVwUZa2t3dkVWt7g
JQmXahuJ1LKO4vfAimmkEb34XdB4P5JMc4LNNVsw297tHoYxq/4Z8yzIAa9Y6Ic7
rlDJFavMU21pBM5rWG+9fqnigfahBFe1y5cRxAoyvPEFPZLihcRo3Mj8FISGh3dI
KPBtQDhnOF8akSJct8z14xUuhZZ2mH25A6Sq/D7A6X5421NttrgzGWugijZpq96v
t9ELAm32iI9rPU4ksiZKDFEbtGB6Dz+kOAOhHaV6lmJzxGZAQ70rGOnc8hld5ViM
noruCp9Q53UikQXMaWVFr+VkTxBxBfaaGPr3vvyUqAEmca4rQGCfUD6quyYjw2he
VjsD4I8ZX0eoIihV4/Q0SUFs7wN/xzKDOqsGgJ4zQdhECcgqAHYR9ozcOEL9KNE3
9FXKbt+667rf5EOUGhvJIBir2hF+s/wtQQC80jzyLJG4cXdpWSdH5Ey7JPtULB4k
5ybGMWd87Jjx+6rjrC91SG2WEnG+rj09KBQ8cnmN1w4C2aY+OLrT4DSLvZAWK9KP
hvqnSG8qDcu60vyv+g7mzX57pkm+rWJL88XP61ucMdnA0eALGtmEtly4cuie0x2c
h+R5iu31HhD/R6GUPQYL1KpQHh4Nq+SgwMLgeiccLHk7Rf7zjar8INSwihR1Tgst
TVYb7pe8xzqV5XP5weQD3/MLsFa+YzZC/OOmdRhfonKXLv4aVavsT8xC5Bc6v0mO
LsoAAc2vvy78ERor7G0/EXMElgQlWgC78VKsAyXmxG3pQ0NDulLMLYhIjAiFaD/s
A3Y2yd3ymzIHpKsl6xJK/HtwGDxMrw4YnC7comeMbKt05z9u6E02M2cD2wlN1Ogs
8RJluoa80YR1qG6orMq21Zv6pNQt7iDwxmkYfpt7vZZg1oBvWi5EbcAQtQmLA+sq
TwneJcehfcRKRqatMHOdJpBgHw9syb7oVDMwop0P+FuEpjYPnvkNyKSTgQ+ujMu+
FWIqVqjKDop0FyXJsaERH5/J2T0d+7OgvbgHzEsHdIKyk/t4HU1wUniu83TI1iBP
ZJSCnVC1HNadcO7TYz27evtEkvkh9KakCuGLX0SbTx0MOM13b+P6GcbEtkMExXoW
6ENSxMSnU6cgdh5QP/cLTQaF2xwa4c7+VQzYjJhIDLD4GB3rZUn+9TEHJrK1ztJd
orjJaBORTL0r+tI0EaiDcsBia80KfnsH1Reh9YZ/usSMLp/eUlu4kZx5mec/gwT0
HNswCKY0loxOcYzZjV0izwEYGf6LW1qup7LwIxvQy3km5T+OKe7OB4Fd4HCIe/Lx
m+JPZtYFrYBka3N9g1REYXYw4Iabt0StF40X8Hxu1nm3bnGxrnN9T9sPTFybP4O5
PA4QYqNpJc1YfTXB7ODACs6aGJRD5lPH1owEtM2LEYo1wU6Tvol4ibKkKS3Qp46X
QtrzkdSEKXgzXpEXeDYilqwh2qrYPEXomBDEPq6SdMlx97z8kXI2nT49742seUPb
qEGdYQILcwdpk4NLLtFie88hvvjnGRIet5p8xXkX4A5uz7d2XHeCvuEz7EVsmodb
o8tofzKD+3v5SZRhrFBwTuJRcRcX0fMB0TGVTb62phxBSxfvPjW2OOZdUMuS1v2h
HlNn7IFtqUIvlzZ88b6hTnawvUlXiVITbeslR5DQLFzi9sVg5zBcYWjg3QU3e6yX
EvY7qdhQBuMVcbxGvfD5D22U8grRkCccffrTg8SE7OVpZsL3W8qU38d6mRc57voz
mqkYGjNFEjKFBhovbL2ndi/dhP33NC+YYpfQNn4TfiUns+qFwL29Ce/Y2AzFO/jY
2wUv5grioOmiRY/NgeTtLjeMxgiqGIYf6ATgeGP9U6vTQPL7lqiS8qFeuKrYvI44
1kDz6s5NRRfu7ZYdmxJygSUsGg+lxfptowBJQOuv/k7AQ3jQezzGhVKCpJwtqILP
JjcarQxOzO65Gz/wQseQulRJyETbTRUjnKK39dkpB5+JP3AeCoGKwcXokbT8qff4
ywPiaiNSOaHvlJotGdLvekeHTkEirjaiQCrfvdmKm/PXg0sBk0eECojeswyrKIMJ
ypWrR9qdgQ1Kz1Ygi9Sr+W6goK9DwwZNjoKFvwJxXYe8hUpa5GapJ0BSLNXRWv/d
nEnVAFMe/RTkSFTc+PWjN0ykIukFQreksoGFyFnPaXVy8MYrcfm6d+eEPjiNsWoj
G98wbXYamTLzwHwLB+PeBA65zO4v20pE1Ypmy6FWgSpfu5iBxHVpyip5v9k4Jy7Z
K4qSCzpFntUhI9bcXXIteWBgW6nNrxHxF8eu0XRL1OL9vS+udrQ7ppETQEBnvF7j
I4jVBO8bxdZ1gYNCPidoYib6li8pl4oTIz989d+pzdAFczyKZvF7cnPDUd4D1lf9
eKhIMOcQjXwdz4lQiGh9jeXmwJwouHMgqNRHlLs5LMIhhutXoKWrP7z5xDO3n3mJ
MRkQHsPhv8wOlIFCFhjcTrO90Rs+JFIpH+4fpPjC4dSAnP8mTPYkxVpHoGLRH3Ez
QliQOGXKCR9GqrdM/xcDEa2p93W0RImfbcsyAnoo69i2gt2Td221Qp5Ue1PPE6f6
4O6e3XUkmrKUBPcPilJatF20uxsPlncXeyP+brXhAfaxXPhM8PVOFmV6AQuEsBG5
A33lICunmO/foTWm/rmLH30HcAUdluq+L1V4cbKngz9ugvneI/SDyL0vRKn/Ai+m
n3f94R2LL8ude4Bt2qRZUouoIXlSywRYNiywOcmWr3hgT2lbfOqtSIjf0ecg0yrk
5KYvFuzOubZaB8RZIU85kdwx/6L/xJlTx2WeQ+1Q/hx7w+QHrLEvpTsI5Xmqnlg8
d9gBVqEXPyUPaFYACiUZPQ+N59iD6YMbZiOw3Tnbk/n9hNRn8b/0hMrgCi2l3knI
axGWC5rF/8S7FjySbLBTme1TRJ5Uhv5sV98yi6LFLsOSH4jDu6UXP821EiyPlvlC
QtjYhiMpwJRSGuRQ/RJL3asFmv0Xk+dKU5XL1EQJDrkSMsd/3yBLAoHxNXNeChn+
yBswdU++qccShJG2JAr4WKAOy1f1h7t1TcmmKlbRlUjbdEzwv/tCMPIUQf0k+qmu
LWTcc98KmB+NtZjgjVb8FA3RqdlMjTp5Ua0kGRfrhvups5I8b9dISLg+e/KrSdZj
ywWO25RZ0OLDGyoyDd1YMih6g9S2+w0hD9COIj7tEp7RPVV0ePcvEVp/zZZCwOFs
qVW+cY28yadmFJSuarHA4XJNmtIw6R7lAq1NzTzLF4bZjfDA/LZDpVllVZEn6kzQ
kKqCurVSAhxKZHPUNUAWX7xYPexFB2cJx8ZA9QNCBXBBSMEIiCqK3NPCPwgF2Wbt
TMw0HZV6b8U/fZ+CZstU14KJ2pfjY+wGdSIupNtwJTplbx2tI0RGSoO9PbSgyXQJ
AT2umGd9IwjqnWJ6F97fiwvermz8i6CpNXJXOsXVrdcg0aluHAxGYQdf3AnFbm98
22lj2F1uA2ZsitFtSMBKBP3QSx8tn08fL+WTrVvJC+cLnOBZgPxtibJYLQLTAeD8
wFUIYwfNroyyXt2TAKnko+nu1s8iwfVcZva5FlF5IpO93xzzQwoxTAy3byVSPGjN
ItteM7QTsOy6Ni34bD7IVBH6x1ul35HoCX7H99qcGolN+WU347q/PY270NN68fXa
rjyP4//9VPcI/Td5FOyClXZL35SKD0EuDAfEyQBR1wRYY0Rql41Hk37RqBhWCCVB
G7M8l+i2lPZTSNLiCQ4jXcQIHMYoODqH7fp2mglggasVsHyHhtZ26Qrno0TWUQRz
OHus/hqkCbpmzJpR4fY8S8vDV8qmMzAJMIEVaO257gy7NbwiZUN5mE6wx4rrDs1E
w5YFg0MXHAtZHc8sTDcEvrKRsuLkT4rI15+kCWS8n2XkILadHHRWv460G3Qrvezd
ep6tghBLSdwDQdgQVzpjsa7Ys9hMiqCDeaNwzrBeYreU0xTnnG1kAqMvDdS9DCmI
lWi0R5WyyPjGAcn65jlO4mnxTyKFYkIQ+jqku5YDDTDESGcxL/bPrq4YrmHLqhZh
qWqCjaf3ikn3//wTIjWAVTd+HG9iMvEwMg7Gbh/92n3keFcsuU/+LealXV62902a
C/MeEF+nnU+Zw/USEVvrOwpFbxUYTGZdrB5u4wMh78DyGWhKFNqrGF8y30vPlLMT
FdCaRKgM62bfaeX5cipE2fv9sOQizXAgThHKdPS7pLXiCe0SFyoNDFiwkZXYQPpG
Zuh4DbpFubM84z682VKtr7dq1iL0iky51/cCBKQe2NM82roku7uQOAtP2tj5HdF3
MUlY0JGMFU0YsXaOWzEWhiAqLB+tJtVO7XfN4X2rSeC4lF8NcNB9pn/VeLooaVNu
s1sG0HXb/bfEVl4XZTFXSGx3LvGO6TsCxsSvjc/0bJDFo/m4z/jg/Xlu6unYCQJ6
2mDIY1og2vXeEA3v4K9hBt2e6mRyr2tpeK6pVoOEG50lqr8h94ShkycvU9Piw4xl
KmxFRACLsFdOkNxOXv0cAQgpliWVK7Wej6qSgEbd6KhsjtiGCJVmzXi5uNta+d7M
mt9dUk6/d6jsFlkgl1RVAsY0tnn1sSQR7ImXBcIFuCooyqinSA5KCbeiMoYqnOmX
+fW4Z+btgk+Ed3JY3RnxuYmC04WO/FxWBMA6QoqUgjvTKvpSxXSCqg+v3MZyKj/B
C1sFOtQ07v2vjnCbX4UB9htKLWT1yyrV+LxvojjRwMTF5MHSDRGaPzPEpp1yINjx
h3SHvYc8+u30saVxmJ2MN3usSMlc4mO5OKj/T8JWTwkKi/vDJJl5ST0skxLXxRNA
M3xg0zIQGzfcQW1j9Tqsyjbzg11XtEhqp4JGPLM0qgFjIUHRRjsfQ8vHt9x56Db/
GCV6lyMsVCykA8I/sZaQQ+mRvuLboOnFB52uycYO6EZCxBSSMZIRcDkjt562AdYf
8ARqe8KHRzoa/MIZsIqyxv5uuZLwDMM3J6WnnR+BH/X+SoLwNkv4qlbsjC6LJv9p
U4LJlB5h9RCLjqh9ncNuAn4FGKZ/dkAU8694SLksmj49knW85eQbJesrUlRiUiC5
wndv8PBuMwxfbqzbDDiB5K07B3uImc/MjElSM2a4XLHrbUrotVWX/qtanpJf9grr
qbCgcaphlTqXULq6YYXarFSR7ecxK1qkhIYvruUUT5oFcvaecy1hxwLLe6mpiJbq
SxClQrGHJvrkgQX/NhAv/D+4MpLdzqYOeUr4coMrk6NcSU1lEVSZiupxFRcR3pCd
bPq4tip3P5Maup4JptQtbPwsPCDxoRKxoDLYeSuHvXNVg0JR+keW8SimUrymo7yw
efMWSd7MFB/lN6P4kIs27ColHEESbrXHr5hJKcod9w4+PUjlvSVRaFQAXFWRycVx
/FvlxG05Uc77PA4mHuzHJZRpicKqJR4svml2EtJZdX1XC0vm76oTL5aw0nWa5x8/
4EeYtrqmvdOh8MzrAn+OLtlcF0UX7t7Z/UNIxIE+i8dTOvrnqNh9/z7E8ma4RZNi
lVwMz2TJcB/gN0yorQ+7L1rtfSLYfY6yAckDc0OYquF9AnEct6lLRInin4nv3O6C
PMvA85b7ZZgDBFxedGW9wgMzKRaw2bHSzhjMF6t4fMaMZ4vQdtumI3jmbO7Y2y3g
HgdchntgXaQaczBSUgHj7dwAwa6Qc2gF9CRd1Svi71Q6xn2tKVlZecK8+lv8eRua
GFQk3pUhfeSHXARmoz225N7wp6R7g+1qLP2t/sl8lalULPQJCKU7mwtNmuug4RVf
geFC5KVsxyI/Qd2JrEOIH0MjjMY6H0VmD7i/H4wEcE7gtyv7nlDrxJeuDb1+P2Tm
xb056oWIE+8i2apPI9Doo2yda8H9bj/dl71Xkd+nOlg7CmebqqXlSnYSClUHt8i4
W6MrVFQvUg3dId9A5Q6JZYrD9q7i8R5ZE/JsRKjhAdTIMtihlV6tiKsQTfTqQ0iA
SpXo20kkmsCDO+Ti4wH2jJCh9HJz0xMF2JTLHxwFblVwZ/e/1Wq3cF/PVBejvULy
x+VePAFe0DJoAwMlQ17v0HlMJD1MGVZzTSkBUP+qZNDXipZrN8pBV2T8GQ4ZCRcU
PemkrDxFKLPMFqYZt+zhUIEbCi+m9+uvhQrtlEsYgUaYyxJeF96rUBQVcTfuJoDS
rHpSE1LY1D71A0dgotVLbYlYYuRJQnyiVH64f9hrYRAEkxSH/sg5jHo323FEbRq3
65QBMpMIoOwoJjHs54/cuuEJ/+pf3832BDk8yhv9MMgvpPkfy2B49/j7WxC/d56x
vjqw1gpYpb3vfhvbKIYpSW4JqhbXbb1yedwsTI88S/7RrKltLWAX9nnRvchiiywx
CcNP7ryyoGgKX9au/G6GsZUEu3SFNZ/hyK5fZ0htEXIdv3oME7i7Y1l2Uxy5sKTv
mEkDJtUtwILJnsKh4ybAoFCxAf/JhBbOR+yOA187YHwO/wns9zbsT7YSXBB2qSsn
2KA5qU9mvziy51CQDrGHC2+iOr6V28AQkjFijZtQOWXG4Eh3GnKgxQzxegtBdgyQ
vYppBFygYa3XuVpvwDq2W7B9gvdkymSI/WPz1JbYTv/j03/lWmH4YSJpN080BNPr
RVbsyC0M4oxI5Oy5+Zt3Xjj1Rwea5GDXcC6FBvf8gagHyGRqjuCl5cOGbgcBqlHY
DE2OLpb3QE0OFhSrlyLvYb/EXw1npRGosaWHhu/I+UccMgEd419M/E2U1b94wIop
jCFjMIAf24yJDdIvFWciWR20WvuuGGU6aEeqjW4V9X3cgjFWT7DxwKrUVYZSAIHQ
ntmoZcv4LvlgItd3gQBBBMrXWIlAEp7N0DNHWX3GPHEle28bY4BMvXVGlPs6gwBZ
kuGjAIH7P3+MuBWhv8rpVqmMXlh08zWsEtYc3dLhFm3cEtpznLVRBZ6bqBOzUt20
EVSDMp7wM14ZaQWWtT6CAr4GZx7h5Rk9N9DTe8FkEVuYIRr4v8DSfFkINSV2XJhX
AI1RTWbY+ZluIg1mn/cuB9FU4gOWoYyeF2hdhWiGUFq82e9I0XUObIkKgp76JsCm
0HZ6cBAAepmh9LWI6PZUe96FPGYmNLuAv8J9T0OFJeP2ofheBSn1FtAiNVlZi43J
983vu6DIfSwYSVqAgP+d0aIBkcdOr4ohbcFpLp6QxwKDWLio45/H6DwedEWYgiRU
9ecd4/bPc3LIoB+J1ZX28dZ7Eteg2OzMNu+FFVM2ZAy8r2lNHWS3MBW5IlZQkH8/
zdiDb6nXvz8NeV5EsA+Y/EPA9cvvXgIoe/U/BZNwmSq8EbX1EpRnDDncR2HtiXjw
4UXdjhOKKoYaUHuzpx0DcM+Bq4bsWMbnUM8VlCozXkQnmSfTGL7yq78sWnWKC1xk
bNWBQSoA9b86WBYzyfkkI0cHSLLYUm06oxD33F9x4/vvNAG9YoeGuh6A6OS9w/cB
ZFMb/qrAifqJF0aFthqb0ABpY01OmQepWedlQY5ap3CEZHLD0v5FOv48zyoatJ5U
0BPrGJQXjiaTQZvQCRkroqakPIbBtKGUpscoZKf5dW/9BctDC/pCAJhrqCiluITs
6udnohIUzFjnHykL5Eva0Ta4xfDrffiYp+bGRC3A/7gOU6E2GM+OcgtiQwtbj6Nl
620zpZ4vgTNaCIa/qu10xtPljKQAWOciq1wVde6eWLXv87TrRHf5MM71Er9N+T84
/FKn7IfEL15KR9yxcbnlxgzk1HJPS0aplz6tR6NNG0h6EZyeWEbNQySYCrk1WC9p
K3RmZJKkXcljUsnQMp41+CBEKiA8LeJbhcP3XBIH1+hHcZ+dpVQZKX485IGWPVyi
4SKy7QwcJXlX/wruIXhTeOS5EhRYRLv63tLnUsRHfWgHCZX0wYbrGGQGRT4UJW8T
JzTCi9XNAEJno5ZreV5XK/0+9JhYg8h4vagiaiZHjgOYPdYxYDZ0Z7uDgQcdGJWC
fd7PycgHMhxmjo736lYlU+N+OIpqBtznohWW2ShaDVzTDQGmnWNbNEgCAL3/9XxT
TB3KlgM0i4CUoOKETGvVwn5yKLefmKExD1qwC4Zqb+PISKTA4tIP3KyNx3Ez9cFA
7k9m351NLE72gsa68Ja17kdxAvBUO3aWA6mdtKosfQx3hgfv5W7joYDBtm/f5uiC
boE6x5IbRM+534Fzv3DDcfSgCRzS/o5E9YQ597cpWpjBC0oASn879OauzFf/p0pw
QMmrej0sZmzzUXciaF9Eei4RBHlxtugJP5SNApcyvf6jqRAhmXg2cXM4wDka6Lrw
qgNPrF7t9RrsPnxL04XVTcVaBli7XR+O5sGmduaT583rDIKLitXA1uNLgOTVkuZn
Bf7/a8zpCwUW9ICvsDmdkub7gW5WTqANUJnlyQkZj2e/rzEf2b8FVVilDwxoTZvq
PIiEiTOckstxcW32qFYFCdyzfYcoP8D3OCYpDmZTqyysp6b5yNNk5qdsf/6bU0cz
Qc6xlc9xWMWYlMxyHmLht+43j2Nj85+V/C8w8QmWPRQuPZEZ3zKYjCxDQPB/FCPm
oKM28McdOOWsQnx+eCTSLOg8DkEaKbAdf3THcSXrs1dFy1+blpj0zkq7Ewz3JHEi
zEKH3Y6wKGaRf9LXDcb+Es1srV/hOjnCe1Mt+mnp5s0Laxy7M1cLC7ianroZ2zKt
o0vCPzmpu+pyq9N/iAwObOXLjx7FC5AZs+bVl+WMFmxE0iNFRSjRIJhSTsXITQal
A30JNaQSH61UfLyER/ZXEC5wUNqNtAjMM7c6wUwYiajBCUv6fwatfONz44GB3AIM
TE0IH9x5VXHfvUIJYKC790UTelj3ggvQbRGkjX4X3gU+bjLtUazehrCgEksyMNZP
IQZKDCt43uC1/VzWjkWBFGqUF5VB/1EAQTw+sZs1iXOrH+tBI/6aaqUjVBdz/UGd
yqHoB3+/BhmCOjYXuXJdlQK8OIBQiAO/0i65iUpJlF5GlmUvyUbBB7QrULYbwYVY
E1aVLIk/GwxUmSIRhZIn1Auto/6VoBQ0A5mwleIILkvau+NJAfj6AT0s19QicUt9
pLxn3peHBqRqyJjwt0MBhlcFhF0lFArb95XypdVTXSOZ1ZuBW55yoIRmWLqKo9IY
KsRQ6Gl11hiOg8EaDNQz5haEcWT+N2YgzsxN+8mQA+vEIHq27q8KscmK+tZN6yde
tcSwMy1QM0Kpa95CjQUziFofA7PzkGUtwaEkslLYm5IITDArOHhnfZo+DpQgjszG
EMymDfUWx+hQEuuL5qeo/HQRutTgUIDI1eKrYQzVo5YfI+gRT5UukkVq0ca3Xgb/
u53mfNJCPPxIpVIwrOzc2amLp9LNX9PkV0qNObv7Hf7411oXz1FlbOuBUPrMfGWH
ZomDkSGK2BOVj+rdeQxpszyU+6S8aAQ4Dv19RPtkDZtj7Bb5HGtUoRjLBuSgnJt1
uQ28zIdTl2438M/v93r8HhzYBU0VPVcCXTEOy3GzAMDBBJIiURp5Si3aQb078Bsw
Wp3YbKPxenIlzlG3tkt/7dzjFr/MDpNTXiIRy6hnfF5ikE/c+7LRh+Qf1DDyT5lC
G8TsRkUeFE0Tm2ozunjIDtRa3ur5gMe8WuCFU3o79KiE6wO1kbdujDvVKusO0vho
gNmuqV+W/KGNIrUfl8HblRqoCrxrxSg7Mzhe2Jug+XQrDtl3yItPA3r3CFNTkSSb
s37qRmTUg64PJD1IMEabvG005iyjKp4xJ5msropvheP5RSl0KN7IpNbz/kZMoTY7
Q8ydAs5HzTtzCHjfhtpBgdFb3y9aOmYqM2JEczT9WJ7pLCVWB0P5zqfGeUckG4iJ
HklHPl0ENwtqCZDglP0B0IWBvOIbJoBqMoNp4O3XWBqNH9zfJuD3LWYCympSZTNZ
XJuhNDl04fdPUsoj2FhGi4SAXbN75r4rA+jzesO/bAxvj6cfq8E0zfGPZuDczEqX
AkLFQkacnMxMauGXp33UsTCsiRIE3eyJj7YMWhz2+7pXL2A1pwuCM87JPyxNaCS1
gAjbakwbKFEGgsJoKMvjaeuv6GyXlL5umei41UhNcXDuMEQL+OKlbviXDt6gg79s
JmUFq6odVomZP0Te6DXCRSWPjOY6a68dothutxT+KPS5FeOBGy4uN7pLodgP6w+f
6WFk5bMRjgKC6AodMIucStZHmkOA7bfdwyTdbKkHsnAj8r4p4LeWm3DKNxba4sn+
SE9oI2VRmf+cLUyrVk/xsAwYchki/HLOglyvz0EwGGKLXo/VGIL2dpnLwbrU/phh
tqVhK4XYJbwdKH7hBDJ8Zbqtnr0l1PII4uHdUE0WwmZZAPg/vHf+1xJ3Tqk7aAUt
kLXSuTXbyQjkawPdiy4kyocgXyo8cpeUJrsRBrpQbNBmb97VmeI0OhfEvfpaq2Dw
bBVE/FGRO357AGDOzft23vTgmfYrSZoFz6zDKMLrEFLkZ56n9ZlaRZEApTwXyK4l
Y0xBgCraNxPOm/m6rtDINOTXhQWE2E6MmO4Y4ZydGvpQ5WcgCZb7W7wAylU1x3Kz
B2swLpnUFyn96seSu8MtNb5tJw0c6NAtoTni4KGrhu/PxfHgZz0RswDmAS1Mpdja
efoKieldHz7I9d8HWn/b2YUVF0LOr5jG8cXlQInu14lT7aFeQM0CvDXcKKuyEp/l
EAQwDprGniOn7xUf5XgMsRXxIzX4tbm7YUuCRAvFxksGXFZVD74v1zsYDKn3fO1D
RXFEpzFAuYF1CmR9zM3AMKLw6vTXAI3Uww+nW0YAyqes1++eqXhYgHYlf4z/iX/R
jK/MyZ22VDHgsugexen8AqrMleFqEnB2kbIg3Hhk+DjSur4MzUb/hojZhVNVb5k4
uUpvGh1PXGtKFfh8gY2IXdYgCRncJvqJs1dRBFGleoINw68cbt0qAPL8TJWlUl+w
aZ9murFvycUZ9m/8KVW3yabDyCmdiOqXAU2ZNVDDKIeWnQBHfAVG9e/MJjYqQR6H
Cby9r+wflpAj21JfVufjM48GIG7aM6+gSqKk9InkD9Oe7DAuMDxaspkZusxsWXbP
7oj8wF84GWHQJGxMZmpdOt/RngiG+MJ1V6wsTDy3HW8I3PfdMy3M81yHI7uCN0G+
8SmvP3vbvegWxe+q8lV4pQwpPusXL5noEWSv6JzoOqEgKzs3jP8sLs0vJHJVTYhB
ny5JiJmCyGcONXwzY2OyLWpgFOfoDY206R/3Zh/JSebsQXSMA5IeulVDsqFJBAk0
Hyqxi3BT34ib+xSpUYxalSlPuZd0ISWZNurSGDMG2q5RgHMm49JIs5oCtLvs3+fv
vDbSODXKB7BwxT9XROzLNWTM4O3G+njJT+v0ifrN4NWGE6ZpaGjBNLqfQ6+gi7hg
VHv4a3dnGmjJOjTfq6F7tXWWEDmb2trpkZCgNg9CJ10oViLZdl9+6yvHcWKtHyso
xwCUmbXT0zRSAEL3/lMwZTmvDTs5La4tDf/UwmmGWUtPC+b+Efa2eBAy3C/7gDeu
bh/96TP3XUYu7J3FQnTRSXPLOjYYWOPGblIlIRdixn7XLX5pnTM08L8+k/UyasIl
u/123RfsZp0RjhE/JinLaB12bOdfC+vGzyyqW9JFUAO9fIQTjSHG7rMyzJxfa604
ndwp+XTncmTKDoYlIsb+l1WGmvEqbKyPDCTqLyTJCbXzq3ABLRgcqNyWHE7KwX6M
Bu7Yb7OLsDZqX9yrrC0nyg+rvO897QbsrOHxxAi+uBLguYu2wslWppAnLY5L4GYt
jM06DDoKLuS21RWIPL7EEs1zsRuBvUx2vCrT1wMEP66Iw+zJyJ0RlOkEhl2mkleE
DKYobG3UATAaMH6Ii75MONdt8kyiwK9J1M3iyrkshgMcFOCv616KsGK+wZ3dOmYW
imTwsguBCSZb5NA/4pIak2XRX74hXgtKy/rx5g0e0VpsH/MshcefQ9FgctcWocG9
DwkRsmdSOa0E/YomkbXEmM1rm5yXkMnxnOvAupaddSziHHFN7oGZ/DyEbkakCB/c
IwwMrIwP9s8Q51EUvWdg8zy7nd+NYvCp8P27O8fUr5pi41THZcmmsCDWmICB4FZG
DjS7Z13tKRosA5lG6khvAT9XKiXd1fv2Kt8LOE0xlcauErytuSFHy8uBmpUDpcTu
/x7bNyVL/svVpq7yanozwiQLv37XkmhC2+CNGT10PymsYqQ8ztftDzZAlqf9A0R+
8ACUs6lUEmIUoYJimlUoZZt9QeIv/ihySDXOqatVFKhGtfGAUZnpnnPxdJcK7OqM
0aU362jNk8I9icvSKrZuV1sAdOU4YyLx9Sia/BY3+dj3y0wonseveR7yjDGofbyn
3XVn1E3C0LgEYjGfQKgzB+PBO3/owpqZ7+0dmenohy/gjBZ0iKeFF5vxZ7SbmN0o
uZ1U843PeLNClSX6eNM8p1sV57Cj6KuEJxIX2bX93hdoPx2XSmPgiftEjdrm8zOx
z8FKJoGR9a8LRy3D0YBXWURmB6c4npbf0ub2EEYZqm4SDVpPm9miQrZabndvJI4x
0YBUEtnIYOVBHRjTam5zVJptgbqbf/AUwhs6PXdgoScOxEEwsTNzzcPzG+Kg3pgr
6cphG0UfUlBKo8PGrjwj1ZBF/HwoY9hjGdLR95IDWmNn6q4lzlXuxVfnZtQBsq/H
oQZ1QUOaLRf/SRlHSOjOkMHO9jXnc7sMz/m/aa78oIfTQM2YVeQWVXQJqvD9TXXZ
6ckh0b/ROc+900aK6semfA2btG3PYnczPxdX1v46EQ+lH9fgSoiaTpQ4hlb3d1Pd
ovXFJFhoKC48nkDrdXVIpT86wE+0QPFFUHmLJ7Imrpmk942PEzI/so/7egyOcNBg
HfyUry7iD19c9rTQ02ld61vIriOiW7d61fiFfSxph6bgZ5Ua6KfCmtld0f9xmMOp
mPHgBAwo51QREZsSsFzvfK4tUUXGFaKph4vEvwKrrj3wZbylOiTKBAheOJ6s3LLi
t/t11kirPf5Npj7GGTM2W3O0ks5aVy0wMA7sMRNZKDWTB97TjwfB/JU4RzhCh1Y0
8dpKgHlHa77hadQMW2rav5eNxWRt868EIfnYubMrxEa69QR5P2uYzWsouHg5fxUN
vuPFkXjFOyGgia9a4Vc7s1Gb3HB3s6ttZKixBT30mashHWQcuamHewwSPgckQo2U
0FCeoGW22FCGzuKIHCfqqH+y50OZP4j3RHcaKWekEbkUXIIeF3GGPzzYqXQlbxWD
6MBEf++COCgTWCL2NLUy96F9FA9GevMLFRlFQaVWUJCiN4bObB1iGxDcx1kI+HEf
2sJw9ABl83u40OjQlmN1L3xY1hPs+dPjaSwl2ZaT3+V7T8zjTu3vg90GNUeXnEQr
SRzp80A+AQz42DM7nBnh5rANIq1haeuJz7evWUsEuJvp0mTpkFqhG1kdCCwxeL8N
A9I5rVywS8L0hZU2J36B6ddFjHxgJ1pNQgeARdvhFbBEAwLWduRHT6WjYoJm16U4
uOlOPteGEB1iuUosyjw0RMyIMw+QfAx2qJitS0XfoMBsozalhH2mSWSowLVnCjQx
pGIWAzU6+oXmPW46rAEWJYjGl/DKz/hcaBlYNV/eAtmRm15xAzuS7/D2aR4JZdGz
1tLKotqbRPXPtntn44H1BsElWgFE0g/hiwrNOC78ohUgs87Nq+JrlFd2SyG5fX5T
Syqpsdrz1fn/xDEI8U/HKvLVfkd3VxyrY9wpFZ2y5/9m9rvoBsqPQO06yIbw8CnF
ra/uhx5J4EAk8LX9rZi1oMVQ/9rZf/uzIGGpdPcQdkwfns4UE5/I9MpjS1lXBBZu
thfJiDUfhcJpOCXSXK4FZvRiqc18KCA8u6eh/FxX/StlRoa7HJF9Z8rryk8lAmJH
v0w6JR6Kv3wb7fa0TplL2TlY/BifsJ/K54G/nclMr7FgcqasW7Mv0177lHgfpNuO
vap+WgUQniv7vUciSupOJmvm77wLTMcAQ0dWGUxpewjqrpVTSIjRr8cY7phkHkzI
a6RhTyfo6ZnY7yxRE3E6mbo49rWLkfnENyqcYQ2f9nMMDytAUDhcCpegcWVIZ4Pw
K4urLJlKLrGq7LGHk/ppdxc8JZHFeHzmAfNBjKNbZL8d5IvQF/spdwtcDBTsaRAL
HfWtdg5+CH1ag2XWKOTPCfnIisek4c8mQE5FYcX1qX3NzdnFx9N5cMHbDmJk0WWD
zLcnngCsmrGFQQRlD0Nz7NYLxBN9hQHOsFzg4qQWojAt0VSzbmSsWHmEVzpQjyby
AYqJNJTfVkHXtLLOyu+dqHOR5BmyeAHYKc7wHsnBRcbfnAxq0qn/k2XjMXiZgs8x
4XDXMjcfcadETsPa5fZy6PpdjCnHrwXr+E0j/SPopeCIyy7evZO5RhabkkaIhX6W
y2eMwM/4z3pv2Li+3sq3etMKuGCAZrE8Q5UJOFqjUZ1KRkmykOBeJQiidGZqq/jS
C7+QO3hzKH7jSiIRLwv1ARET36xeWN7vMJy1Md8qvuxqS/cwbQ68ddUnJ96Y5Sq7
wVGqf3Evgb9whD35r6NmJEtKRW7MODVQidQGxYSJ/zVvbYo0vO/bfTXgLXZYDrKO
weNmWZCGT+Bki7xh4R+2MXACwDIdrTgxSSXHoVsoMCxI19ZUzgIjnKj4YMcOz59o
tSMUdj++D80TZPM2JZXS2V8WxMHsPs/lnSHktooq0gDVQXk/3Mi3gSHc1HtXsBu9
MhD5plYjugnHR4H88/l7Eoa+z/HrbQxWS54cIjHkqJPXC893V9OJrUoDfGfh0w77
On7tCsDVDuks5rqRt9MwIcZ/p9bjHUAG1fhwMoqYXlTEB0hyc/T5q70D/cZVo6Yc
3yq/ASzpFvPF8RiWa2DC91UAD98f2x1rM9x7nxMF9CdCVHVkoK8bT5FlCWHZNQOT
pVnnfYGx1ysKIEadXb2fqL9+GpMygKWy81c6g7Z4MJ+ymwmvTsACxFErCLj9IrQz
UDZ7bmllKEO0c0paRumSJG0l/E43bTDSdcMVGAA6oq8ZFEywROdlYn/6vW/Wqjw5
S2adhGpH7JPGTZdGnmJ8ey/VcoAwsT+bESGUCNnqBDCSds8tBiqCyikpKzosLjqH
cHqqUyk9T07takw+jzs3V1M0vdPqCUJHciBIfVKkTUCwPvOl/saL/rmxwUWrAJTS
/SKjVXPrdm8HTzfB3snpivrw/UuEYsvsuqqVFttIpT/zcyEdnej+2TNlUs7cFZwn
e0gjzr/zkRVah50u/HR8tG6jWjyhNMx2HXzsDdu+vOCgZ6DVr8voi7JRV+Lnlmb5
0WkFC2hv02iY4w5CKwMi/qBhSwQv6Up3jo68NfQXG1SqsuNRflboHCXsY8GOe6Ya
MyF6f+vLtuvsKQByziQzcdaG5Yom+nxz0BwLFk3vObkrTWH3+1i2AV0dP0feFV9d
DzQSdKMvxERdHXfWcFblrhBKdglyM3nD2arPEWqI56isZvAwHSaukZA4fgE5vb9F
94x5WwL7+rmZVVjbZXDGKOtU+gFT2W7XFhpPJyOG9vLOyg8XAN19w8naPmtQ5zoj
UuZmGSgE/Hmq6J7R0UyQSeCGKXd+ReZJnkZeyimQE6Dp/Xtw4Nsx/9fQhUQbpPbP
Ptg8EFP7Cu+cBjYV+0leY+JDIv/GaCKUPNes2QeAm17KWfrQso4hx+hn99T8nV0s
14OdgoEl8+/9bQnzk3bQ7x2yTfe8PwjNzTLjgKL9f896mS/pf2COXg+sVzty2Z+P
TbCyR0QVIY9DZCOLpPDpL46qg+Ai8NWleT3TUjBGWxCBT03Z4AgY+Do4J6KCipyk
9JqFpERsYXZ+yIE2T/nOVbJ3ctedQhx6zE4+MjqVerjhIa7Rc+B2SZ03t2/k+Smd
JfRCaSKqSdlgKHKOd+3Co6ozZFPs/MMruh+yYjY+igtef6Q4V1OvSfXIC1q8JMEx
XkguINmtjARi3RR5tdz2mBBsmCDNBFC/jG9v3hvHN/Y55Hbie56zv3SxOX/60Pt5
oWFH34GKc4h2o257cx3/uXyU2Hm3ndJ9kG88sq76A4d68S+pYs22kn7olSO4Fpd5
4i42OESHagR5jBDQ7569YzqhddiywHOCE/Op9qOjrfkwcNF3MHMbghD3FY9n2up6
CuC9Z8IIZ04N01ZWgmA1TrB4AJSAMbjhYN2Y69vm0jWBaMnrnaOsA2XtGXQdE+/h
91ujGCuI4osb0Mvo6DYJ9pOtgi5YrC7rQRcBnSjPtSxgU8vYiCgZJxfEmD1FXSlV
a/dodT9VwE9iLu6s0Yyec25s1PpNN6IeAc8FvaT1G+snYZLnBOxhfqcAGbsf5REf
arfFeEdWpAeehS01z15FNBSdmsd8XqLKiAY0voSrnwOUWZ+F4A1NETTgq2zaUfDK
/iPxDBMYWih9dGIq6enKaBW88hEmg48kQCGCs9XXMTELnYiLPCrmaBv972+zUQbM
P3qRXJwjMlRfWKgdTiyWwQXVT/QI7cBwA8mPHseE8roB2XyCSlGi8ouheaJLzPm7
m4aFT7L8iHVjB+Kcs8b3gzoJUMqsBUJUmQ91bQgFgWLpy2TQIjy4zxl6keKU0RrL
I3B/PfN/xBiRfcLXaPHbCjEuQI8XmopC5rjToZXBp/p0wcyy+nOy+pGL5CMdBfFO
9dupkrsi5hbMyeEOD5AzKtAMh+vn6hZdrm26JE53Cb16LRsqAMUDBHOwIaaZJ0CN
ihOI7p7aY4+7A+4qCA8ERvyi7TE+eLY2mZJGCgY57YnfhIuy9qTcXeZqkT0Ted1b
cqxmTQrEWZCj1xw4ybwknGMBsUppVRvVkxnVD2OIb0XTjSUlgdT+mvUQSd/Wpolu
IHjxTGQJ1hkuh3s00VSCgUCQlJlBoHJJHDQfLt0c7dNuwrXc+x5W1C2/fDhh714y
BxiF8fiL4crtcNfrbr/m2mXVCEF8F13yETOv/r1z4PdHwv4e1fXcRODIW9aRMd0u
30ItgpdEDerPNlpgO7xNUkRdgyyVvYOt1oheseX/+b4O0FPbpf1TAJPLJcwNj0k2
ljqyg7+ySFLdDg8uTGHrp4YAPfku+hIC1Mbwzj/hCXYiH3dH81xD1e7H1drhBR5+
dz6DGivB22O66Ycswy3ZDmb0Iv3WJNSKn/UgS4oaD7WFXxqI7Rh3XzvGui59tkFv
/TibcInerbZNhAicLdOgS0mUZDXWM0a5jyFuSo1ThUICvIHaUsJYMMtW5n2LlHZM
pUOH3s4ueI09eWn9S57Rw3DhxZsF4HcdEbUMPT8+QLPS2/aIvPtoFuEZy6uhMO/C
8UtJjEoZQR9yFhvcdoIm0oz6eCMBxp67KD7a8hoqWdZK6eChV//17mdW6/69Ov8/
/T659J1ZzFNOoR0d30IPt4cK27VZiYj83zoUKOJa59mqXZtkjZGcJeUwRSQCv6Oc
wnSXjfmNJTjzSYxj5ApQFHIcoHnaCtmywYiuLhQqMmY5Z4gZ9tb1nMtWBxUF9Dcb
3JRcGWd24weJBpLBQ7Vot5ZGqZPekB+CNKdebkxfTRKctJ10NlzIgJ4nf+tmfcuF
maPZEkSW7ojRT66Ejl1xPO4mOox5tvKdBqE8iNdxPpgL69nZZUA6SLc1XjfSyAwX
ub0mN1VgoOwVoblt7hRPnIV8XLN/f4tqDoJ7vT0D1L2kyZYR/CsXrppbSukceDUs
9qFyWhrCeuPno8tqHEQDJus0MZspxgmmLByNtgwqyY4wWhuUPe4MLDrVZ5qRz4c8
B4JYiXqZo8iKYYQkH9rg1AdiXBe8qsqLNWokyDX0kZueWJbJURnfVdla1MXYQ317
kAxUs/IMcGtSwCrygVk/zTgOUOpr/J3JHmTmF/s7q92ST+4mRYpI2JmWn7UnHB8a
Yc+yi+W9Shh0xh4+srnBRHs11X8FZ/kwTj4ugy69W8hirjdnvcZzLkTeatvuci4/
ArSlrsUYOyf/WtOnNsAE1zi97gmAu9KU8jEBWprnpcfJf/J0gixxXPVvXgzFwrDr
BfZtxXuvQVVqFYHCEf68EoNA1duX2LLp609VDswvx/uCDSEZSWeeXdpR5+SBS5qJ
7cFXTr1Hkz1bTNyUt26LTZjG4MYob/oUatavOv2eXLN7Qc0kLJS21i30PkKdfV9z
TnRpTLQcre2OWzUpxSWMZ4cVnEV9Fz3062GF6tMsXL58h9PFjZIUdWqGWb06MIdY
8No6meN50QOGc5/qoQ1LsiVrMr21v2l+eLkJhIWNBCKQJ3K7c7Y8+wwyElvZTRz/
g0aNjCY2JrBn+y8Y75CKY5GzDa0GTVcaiPN3tkX7LpwfPrtI9kddCQ4bgIOuQ2qP
Cgp6xYYkJNVy87LxNUjuZFCrfZk4znO6xEuRRwQgB+F8EcYE+Qyg6CCc/ed2sN0E
g/nZFReR3z5LB4IodnzMNTATQhe0Dvw5MWfpxXzmmMgwPAv797caCTIoxhSNzn1h
ehfKrlVIsqUk/+nC7DAZSjM/hBoTQaCxGPJaa8KiirufUX/QCwu71IfycehrN61y
h1ColnuQTGq0DBdt0r8DWeOaEU9n2onyJlU6LeiIkjVB32rCgKIBypWOMcaXgDqq
RLFXozSGtlj4PImWK4eXrXS41WXuTY/X+4kkLMJtUnI6MkOvTy/DA+5/ozn4WYW8
+BlHzGwwAtX/mVuNDGnL8BS9wnOZhKzhmA/wwb1lZOEua3CxF5TyJQb8vwAiqHkV
8zv9B+bIdgU92VtjZ0BlZ7Lf+C5lUtOGZmCz8BJmd+ZQKTkPVgIa4vUYQ7uyjwyE
rPmy8pTxp0dK0+TNfh0YlcfS1IbZutNZ7Ry9U46OpTmHi1uhyf034vebme+xF8n4
HO4LUFITlz7RrKu8f4xvhQnYOXO3UwlFnxSkxPFQeAcfnRAClznXOHLgTYk+VJo3
S+wl7eXep/S8gPJcJyM4hkSQjJT2T1Lb9iY+2V/Ac0BbxOw+wAdt8ylIoxAemccj
Quq/5M7YwO5z4woX7oKH+FH7Yg2ZZ9H2JVDK58NmeHJOibvrU4fxTSuBhfiv6TZk
aFyYhQQiOHW9CFQt4RaUyOMKWTmkt9XmCo0vhynZiZFkzKyR5dopO9XxyCvQF39X
8N2KFKvwiEMzlsM0Z0GWB05Gm3HRoNTHyCJgF9btas+ojse6I8yt/htls635vHhy
uxzmI9uNJ/XixtqW7pcflTFho4yNaHCYZoiXwF7w6z7UygLFfPr11YoxqF2e1bmT
joJEadHK8xLKt2zJKUtL95tjQSVZTWYCeKQqSRV2YsoBLjDOJLLvu86woL+m9mRn
IhmaowCrvikD3eqEwBsjMXlvumnaCL6Ho2J3I5mXI/GPm+w00d+yEfmky/IoZ2lq
aH8bqsIp/roySLREgE8abqbfqqjkWFvlK3JTzrc7yhWgW42PpAKVmgUmbBg5DYLd
c/S/1yf1N7RzqzH2UzLJoWejJtbbGppv+BxPngENQ21FNFmRGQDoy+5c/TJ01KCo
rlX5vya7ca1R107IXNwuJXo8tfeGGBXxLht1IyrmjDrwYGyfpxMNyXaED/TnEmET
dJep/fxiitN1r+76k8AhprhPtEuMY0lLgRd+rRNt+vvcDZKqXXLbJFvW0YtLZqcZ
zNwMgE5Q+cjre82xUJ6Qlq0QqUWZM7mf4rJenDoRP1Xb08otQsfPWDEMWCOX8M9b
wcEOqdhAnzOfPJQ5cEHi6VrEg3ZgpiS2DmOrhJ53S7WFnlxe9amcJYksQv8vJhKR
jwH5EG2KRTuupyrlwVlCwnmdbJ1iMvAy3Mauec3ibr7XZz9dNdUPt4rkd2dUzYfp
MkebM8m1u9CuT18lIk81HwEhZzUel8F5aog7DSFFS4qiqFsO0wgA2oXCjAjo+66f
2W9FfGTYS8NCKOP+0b5xLs2zX7I3C0XJjbTFyi6+p0Vzrh3O9Bqdm+mMSlnm1rmN
u0M63YAt8Mr+XeFkEEz7M1T9RP19NzsSPTQk5m3XK7KPZ8l+qj+VG3ZIKI6kYkdy
JjLxQqN5GO1jFWvnIVWzn93XuFAdqsbaIQyaT2Z2tkKMiWieDUXqXkwzVeWMiVNu
SzsKq8WbxREWrrT0CTPz/enF6EI/CJgw2RQSSCpJ5zQsbi/PXYxX6hOlCLqJDBwK
XZ09Az+XjLND2hfCe8mQzoIOJ86GdgmRMfNzLOOsfJDczFG8hvXQv08+zultKYi5
k2HZD59HzPsaktY+iEJGccUGwOEW0+DMBg/Ls4/hHuasunv0CzylMTe1sLzDSJoO
HO5zTWgT+cBPk4PQa+xNwcQD8zoY8vVzZuop2lrk1mronoi+gVbRjvIVMhxCnU/t
EFa+9T32rvSJEsheAmOg74FJR57pwPd0XasDEP7shg/3ApGP67hRcXjbEzQpxZ1O
XFo16RUrhxnl6kXFKdy0XR4odZ8QmLmWhFnWhNbPJcvs46WeZ7NfOn4jTb/ohIGj
VT0Sqis4vOcugjMyqDecQPywU6nWSHeKIdXSw7ZUipDdMZkdGuk/EK46WGteHNYt
pj/nSFyT7nlNSXhFqW0pxVQAmTRHq6pH5MhQ3706ZWk+GIPawAexYiMJdOtcdMJX
rucBU2b8sJBrfhQXk+TNiDhEpCdSUlKNa9M3p8uVlP5bDtA9ni7eqMYC4wVH2wRC
o+Yroe1IWQBCEX9g8toAudWg5GDgBaav28KAgq3Cru5BtLsnILl7/yaTE00ncink
0sddz6uPVGwsZl5OWKBZk17HBK6pLqi9YcIcnW11CLqA8aH+WpNKiTk6MobcTc4K
IQgu3ATZD0vloz9+V/Cujjq/S/eRhkcsaouYrxp7WvGMdUW9fd/18UWNv8+Wuy6P
qkggyRcjxqBBWMSYBtwH1dnJBZqSNFN94ZefZWUr2x7Bo7a2hUccYQYsmG3r2AiB
+XLr3vLC/REBB2uvSnx6ROKo/k0m/fFua4u1F6gtGitAiJP0+wfcHWUT9xq+K5md
9CdNHe5K37vCPgzkW3ttgih+Qi50IkDyPbJH7yGCcmmorFb5vcB7syhiUYt/1cjw
6xiCwJiGXj5rkxUF3GNizx/zW83doqXTXOFKAVQNMcl6OxVPec/gf/cMFK5iaIvG
HZyhFRxGF39qQ9AT7fo+jFlG+onekkp4f9yIiRPatJrF9W8Aqw84LC6Py38byoC8
uY/sX0nvM7szL2ExHyQZPbiwDQLXyjN70Mzn8weXug5jeaAzWfnkWmzfCHUSHNF7
SP9GtHl0Cdbiu1fGrgEw/MUWMb5i1+TD3LrHbetyt5rYQ7L9Q5P37ddzQJIvnpWy
Cjd6kDbyt9+gswg2mhwhO6HYSySuyfOSx4Ldx/fheRfr7jElSRgBzsJN8Ql9RfQw
WNXVcDWoFthe8EKQzHbnmFrAUW7i8weNgVp45wDA58G+fLhwPlP4NcyJtDbKW+1C
Erii6zxfHc6BIoaQm5WxSOaGGpLB78RMM4fIv5nRcCn/I3EPCi3bx6FYsXm1LKQj
kfkJuQ3MbZCliZGbiuZ8pCyqO0XcXve20pIFo1RjIgJgjOFli9Y9hfcbxsjrxyXM
nl4C3tV+KPdOLOjXTFxXQDwanO8EepJm/QcdwYXlHeIi1WWHx3wma/zHafabiN/7
7uY8+YB7AmqnTv4D97IKylo+65Gt4GQRHpiFlWoLirCSoEBP6s7mJkCgx1SA3FI8
E0oYSp7VZMTfd/liWwrkA7Zqfu6lZfYa0f+3LgTJY24MOl0EnE3ybFJ3PZBXPd/R
bFSkayB4Bw2n1vHZZVoefANuzAlARIFXwBxeCadYFliPfpbmtalrOkopSsyCmBPu
UmCFj8J1hOdyhWG+4FFoQuQDwro/JVhO1zjihVto9f7N2ZZjiBNSy/KZkj+G/UDm
sP1WfhnfEPtmFY0J5BxlJqZDfXh20aCPKGkeaYIbISCldVXiQLkSzOy+n+eVAP+l
wpblugc3N6c9ReU+gkTKqH0KcjwibvThXaKGSTP7CMRtRney0uf65QqPdXOOLgpO
2xPpVVvabGXjCHlq5a/yidwCWqEENqhythBm80RoAB0uqGhBQkfEBWX62Bt+SXQt
gRdE2dZ7h3icNuobOHcdz5F7/8KN0jnZC4pgzDny+kqig1QHADtpFfF8yFRhDzZX
XtarJFM/AdamlTtaT8wgMEKdCN92ua+Wbgjc3LS+22yRX6uxo3CK9QJDMBG58qwZ
7fiODU9XGm5giPpUhQQ+Z18OOwcCUlVcn5qSn9NPzvbn6negvZiWbfqLYrO3wEuY
7nJVKMWQVtqLC3tjGdH4YAjoz9G9InPjpf277Qey5RBdYeQvgFKiHLH11pHr2a0O
ssCZu4tjl9J3yfUt9o+0xxWO12kWh9kbJVi6/4MgElv2xLBCq6UPlCZmwLFa7SSX
AK+kt+ygQU+9zkfwIEwvtPNIdzyQ4FxDpW0n41Ls8+TSUErTzMQT3FbgX9Njiuzs
9tg2/pIT4JQTnoC58DolrM5y59wVzzlplW1A5b+yml/tEnNKkZ3GZJM/sYhfNWBY
RZJFbH2BKsVqZ8FcJ5fIsyUf/pM0Ua+L6k8KKYzpz6FolMw+BAkVR98+anC8gxVG
OHAEKGDYhF7IKcF3YRIw83jv0QoyVILei8xvOmCZkXHvDdtWyMT0ORIRwuPBc4uJ
VOtpOQSueF1txWd26E3lNSe/tl4j53K9GVUmr8IBunJEzZm4nlcR4ru2HrKidOVT
5CRQTVgFCMoXoDysLcSf2OsxBd7UmQu5rGPklLILp9F4O7+MisYjzZqRYmEf2Yjn
G556sM00XkaVE1ON5zdYsdoADBr5WV9LfGQyTCwLM17ljb2TNjfOt/ZVdMaDXcQf
tUzHFrGPw/0WxL3CHJok54ERAzTgbjETNKEQa8Ufm7ajysMzZRe+5Cwau5tn98bl
D4NZW8Qw+ejqNPsUGqRdbZywdh1BdwqWdkItnPDfJs/5vErmxrdn2iJB4pUVUirr
QCuEEjl6lVtt0nAIg9G0GDURZEDQeI95YcYgXvZtUAAWki5n6rLdj75TlCGtxLTV
GNoI0xjgX0YpDJorMsFD37RRJd8QFogH6y0en/0a4wuuKPlykWOego0Tfuw0FaYI
GSTRF1uRpzT/rx6pGOUXFVodlGhxSgphhMRt78vu5G1Rx0tooyEQVi2Xhlbcy7gx
GpqYXwIdDkAod/iJrktKrh6Ccg/DkAiKAEJbtOlenDmFHk6PzrrSNzJ70TLpQU1G
57NN+8m2fIXAg03PmTvQsP7K7Sr4lsYPVCXYzzvHY/fKDa2y+IR0v1ALIFkHxNNs
oMgMpdizSphh7HdRfnvXEa9TeuM5ANfDW3RwSqQQMlMLLgcZHDcOdWP6wcOKNquL
xxEuepONKzq5E5h/oYfdFTUv7IdySebry98xUbEgM3tiO+u93cK1quu5u+QtENVW
mEfG1O6yR6OuDyojSVF+32491FW649KZsxvRCnv7Z28JQjEpNbnT/Oxyg1ZJDNuq
cg50z0XpJBrRk/ATpm6Avx92gddiKkuY25j54rpnt6ENJqJbRgPREfPJ5KKQ4lkU
8S48So81Jq0qPmDlzoTgocpFZSltV7itiqV12XG95kW7zPRplrmPWjDvyRbYK3M4
oHKcb5QeZ7Ox+lfPKKJRk6UsJkBNyuKSfu3D13ybT419a8ZPeKbA7ayeJ5sgSXk3
mUyOW+ZlRCog+I0iFYloRwMLkxunBxMvEE2NEQXHRwClDURBgHUY/0TrHo13YiU3
bwNQtdJMvuVxaUhwR8s2dBwmWALCylNdOcitgxIgbJNyWL0sQ1YCzA32iUKmnQYW
c6GZoQ1xx8lrsGHnk2oZMPvnrcvXNI+u7iJ6EtMHAJLBJpdHGj2AYTvd1JpNyhxB
99FSQhB77ea84ks4cdeCg7FMJqt0v+yGrTnvS3YoWtj1NKiu0HvHQyrtEnlVUbsh
NXQCsDHLZ7F2GFjmDi56AFU0cEhufy9oM5HUkjN9gshvmqfncittTbjC2s3/fMIj
BwmmHZg0AjybBRYl6PCnuaKTG08H8JURqd2byrL2k5gUolPKpE5A+gIKky+vGYJo
J1S42S26MczA7wtl44X3iCQiOqkh8DVtBrK3P+tkCQ2bL1WUzdFIL5OsGzSM0CY6
ukMC0Z43Jj9qOBMNm87hHFna/I8NHF+qInKNclDQGRsG+qqsf7WrFq7EKRtMwCbv
VCkVyCVv31bgWsdsDtDasR0T4S/3NYwF51MJohsSHbfSucJNRh3OiCK3IKMwQVfa
1prcs8YE4g05OIYj423f0RtCpeimE6kLjI3aiC0UEopHISsWpLTFXfEYzGOZv620
0DdI0eRGDwnT8ybJF4TTsxk6Cr+vjfs6DZPMfZTd1SdeCaO7mI659Q8RuQcelEb8
v52UDe/8pnGagZOBSG8xC8U5/lQB7s4iwibSjH2UwXQilL6lhvb5G/SWsZaLviAj
bLMAFbPCCS2aVDChNPowuZICPJDy5Cq9ECeWNLAe0ZwTHn6jqpSJPW9yj1ZDRRbB
DbZDFyQso0A2Y1P9ZO0JciB4obyV4cLgghaDIU0Z1weeDXmR2Yvgt/xhanXLloKj
Djh0baEYFTZMnsPm7Pi6GPFf1IaGQVQQlxHBa/JfHEkWP2o6oN+hUDAJtL+nPGgu
cpNMY821c6uOVqpsoPsqLGxAXUM62VbXwdI8yI+nX8a/IUIN0hGrA8Ve2hFzMMr2
tBKeROa7cZoV7fCkp2oqYzopJZB8S7heZHU2kHH5meekYaqKrK4TYkWPTAoOSlQm
3EZ0qCthOD8i2OEmVUMO0YODCVE184KqR4oUq7LhZo6BHUI1OHWmuT2GxTZelOG6
M64uGxWUnyctTtghGpek97SQMCy/1l4+jcUg6oUKCDaDR7JeSekx+dRql0EyhchH
Ufc3gGYPsNZWUQizM4S/Qy8ssH+auOJ1U6n1OPCXuZ1qe0NeB/kNqjHdg7wR3HpW
2JgOwYmhmU/3wtX8Io0PVCsKqk32B3LsGN7YS1ghED05d54TaWo8FzqU1MpFg1vC
KYiE7fWTwEHaOQP/UU4HMzgOU884+5uqbvLqG5Ry9Wynm5GA/D/uwzwsQRz6dN9q
AzWd3CIyNWrdlxU5h/7/s7Fw2czY9OvI7fw+NsxSv4fc/OmHboa19kMjO6hCteFX
k65BWQJ3sW6TrWmZPImiwdEgjYqyyqKGmDCIe+miH6bKXzBXQFKcF5tHD6Xt+lNb
hPKpHZ/N8NSqslnBX0JoZ6rGYdu6QGXYbViDfDRdHRjmArehb24x/mwwrRmMHHj8
0elza3+Z8zV8ONZvfEY8cKn+QotKmOSLxCfiN21MiNlIH3A+CuDMCo6YRtZPR6qV
R+CIYUqry7o5zQBgWaaNIR8jvAsJnXc3b3nL2MbgIQ1X8AbftmN+RKx69LwzTmRV
s6b+gr8LlVCpzmDDFmUG11omuwvridXFYokZHA2Mg3jFU5sM8gcdGgj1fidH0FT1
7oCdsYGKFxLy5t3RmQ7t6ohoujr+uXyASbZwp9c/sdcsH8rBqLExA/h6tJWdD/QZ
nQlp5IUvaZcPtm0WVG6lyu6rR78bh7Hv6DkDC813LCY0//6xQwJdPPJqoV8/PGe8
ckJYA4Ru/cWb9RqUZLf/QKveoh+IcFbfqiZMb7REDux6k0xTh4htcM3kcsxe0d0k
l+ieRT1GDRluGhK9HEFmcXPcPDeZT98XE1j0DepwYUwFQB+eNzJjp/2ZAYA3Qhv9
0mhp4A1mgmUfibqbGsa2Ysj7IWUbhEsA7VEXvWtk5cx5SsUvPMBOcpIcTzj8tzfx
fuNrcwhRPZIYx5X55YjC0qYzFKcfQPC3GCOFGcOpAHfEUMpQjBrSY52ob3g2GSCc
xjtxzqFHxKil30YQ2MuBaAJIy9x11DiXE0YAQ1eiOrHnQZDUvLBoe7FbyR8bWhSc
3RCYnBZPH2SE6QaMFJmJ/uSUuPQDZw3Vb458Zk6BMGLXM9GccgaRcRSrf1uAeSA7
42bnjZ6Vnbjf+IY5cnj2IoUqXO1KV6CdvYfBEEYOrfqsSJ0+4SPJD+P+C75Dlwwx
HvqgdoR2ReJhBpMVsG3rbbrJkB6nPlqwx0TSvk90x2aTDNEoag1cn3Y4c254xt3l
2nx8dwA/0NC1spdTs/NJ1V0r7HS4gH9bVQ1XsOEXLdBGLdw5GGEIXth4+1wUbhzJ
ppCS+0q8eEWNWrlQvhIEkOZGDU0CpxmQACOAKJrzUICR/viTZILwRSulf9jYooO+
PRYk82Y1bxf5rH+ZtXuetafBkn+KkSdgxbYtcC9qQoG232AYDcwWxuYOvp04VyPe
Icl/cee9vBim8z/PM7Ancrx9BsWTPpvJOba9f2NwG/oPF9EYfDSWiVqm2CsN9OF1
K6f1x6LVASFVyIVn4z6AS8YgA8AUhasp2HrWhfQGZWPdDB8U7CY8RTiXtvB10mGt
JvDhHIvgiPj6GgHovlV1mqRStZ83030YCcRB1PFzupiwlKA0QTCdES+6bSW6/LA1
id89Kik0E+dI4HJhZUFmcrskN6tw6Ywxv05XaNcYrjQF9OSAR3TEXC+oH/euKRdT
yvRjJFNSbO0MeVmpBzjimOtHCdJILlBPCcUCrrLzoAD3G7UNPLn26KGJia/BWFAS
CqJ4J7p8T4mjh0rnAGrfx4fM28ZDio0rwoqoSC+/DwS/sGmfC6iIHJ+AQlOazr6U
1oLvppdC3CcNl93l4m+fy1VHCiJwV9LtPE+EK4ZvAmXVoxKpEWpBWn9NVCB2sjx3
+D8vWbwdp7iJOPQQb7fb22NdI86SkwfQSTKeSkehqquEQZReaLj01StJH5q0yHg1
9+xHWrVwmzVx9JHMfT0wJPrzD4DgnMHh99USC5F1neDKYnQEeFd52GeyyWHL+rPm
SXcQMGoi3rlrsCzF538NJsRJwKCXMQBDqky2NaoGzN+sbz7jv1nh3e7JfjxHvRHa
U2M80OMsMRr+1QXlqn5HJQIjg2A3INN01knsO2pwLhxhzokOvoQyev8uNi2u/JcM
igeVfI8ZHvfNrx3PZQLitsMQQRtYji/favOKIdFOPNOLnLkYWDP7qF7lfXWkklQI
uzNZeJD/NHcuduNt3NdY7WBwc9YAwjNmRWcPZqIwDSHi/gckZZgvDu7N4jtUWNDl
YM950dIzGQelR/hCJZMtxZFeYPMyOO+FBThkhskVlXOqoNAzxN8U3c3XsS90EDaG
02Npg6foqVuzUzYrLTrfS8CrTC9hd8Pfe2IWmDmJQxYhVJcuZc50SS+rti3govKE
wKzhYKCDfGn03jw05K6o5dvyLBN4TiG/oww98oKv2JlqIBWN8SEtooJjmDvj48Sc
dENNeQvDM+EIx3V1cKO0gDVvVvlfBkWJAhkG8iquR9F5M7pyyo5pi+uCPOjY5xLy
t2L2PAPdSLaNhPYkWOqtWbfv2q2cwtCWQJ5RIzfABtLmzacn+qgLRBr9GY/KX4Em
MbSOn3SeZyECaQK+p4acGxPOT0cKCaYB3KF/zVpkBxFy7T0jpf8KM2VRzrwy7ef+
pCO8ukG3ITskj0Ka5eA4HgdAhFh+ZrYDeT+N6bxGcDS2KVNDPOMVMfJtQb/DyFJX
0nKoCr8O6lvrYUrqvOXLVHGUUDun965Ifg7I9m6Pwsr3vTS7VdImtF3EUrFbUNlC
7AoARdHFl0q2tHz/jnOSHJrnIkP5qBEGYE+mG+LDmIVNE70C6eE4sCfdGMCV3S24
8qSs9GBJKchSX60DLfRrBMFwtA8F0KCp1XffgUC1Fmj+dPTde/1QTnyynf28Ad7c
3vvAZ4ODARO0C6aw+B+W7HKRIs6zgJXmYoW+5YbQHFmGSfXCNd8e9TbCgirSseTV
fuH4XtoccmPCH/SVUkxrTnbJk/xQdJufXW/4LlvRSB/tzrE518j24YKz8xBAPbGh
JL3tdAsMNIzgn612neAAnB8zCDWIMI57mo5wnGk5zJvQlcGAiJnxCzi8WEvxlIno
MfwZARuzYEsenY41hB7NbFBWlLYnNTXbaqnLkRgNKRmvP2IIl4pkFzR0TczAUCpk
055Tgi/03SoR41RPb0HOb1Zc5i7nKMWBrVpQ87w/9WMNtINlLj0is7WFXXi1OmXM
J1PM//zEKotuBCwwRJar1pWhG1b/k8K/A9YuhQP1s/mBHnWWcUnXAw9mkz8fojQE
fxw2Gud/jrSnFBKlXCS0/VYL6Jq645LrD9e1PUQyXgjCRryMLdbpZS+UKT+vobl4
LRLB5u/8vtM05hWZSKujDQ7PxNbvuFqOIns4z8cYEpmWrVeeY3QQ+HB6IKcKg3gp
2QDL+WHPheeCO9zNFCzO2gvrFgW20j+nmRklVLkjmxQpwfE59/vhm3SXyklVNBIv
kbxSxjgwWXlN1e1vB61DOKi6xu/ElJ/p1OcU11SmSiochhaFWh3McjhhhBAOIPP5
CbPQStz+iIhzlryRDz4/ThAXO8XkLyDGO/Om3TOC4Akw1xhWk1cUCXwSb8+xW5u8
FNmHMSxTj120KpLun2ZuleMC1XTw1XhklrBWKSmUdDyO2p7aApbhJebrUl2Ky4bc
wIeWSq1gW0MKOCBK+7sGIm3Z5UMwSb2FFGN/7Y97NJnCq6xEUdVR+gC/KqUN7ZTO
saxk9ydsmF0dD64lqyr6hFe5Uf4Gy5zTJz65nVdBzSBAD1WS8TVFLODOrsQqc5IB
EHWKMBSU9nIef4KNgeRwgrfeqH2pcFnqVmVI/9eVK8w5spsUOC2QoTHClYCtwVbw
dPk8KbFoiSYuy9hYFB0U+3Fyt2ZPuzL5DSVCOKDaclF7kDVD6aIaeZ0V9ujNoLX4
189qB6vjptGm0rJgCR0epIfAFfH1whRhfwvmIHWkwyUwcwdojJoaVYWbmdtgStfW
Jzt/ZeajtEXBHglnqpuw6U1OSvunKG+hzH14KonE0wjL1P/bwQrhzOkZ3eFHSt+a
212EDLfeCJK68f586D7MIoAJ+ocw9Jfmj8FbcNymPNZI6lO+Ww6chGXIjek1JuQb
Z7RmsDaCvCvogklDARNchd8HmCilB8ZP0RV2+qIe2rvQXewUpOamuxbJhiHjU9Yq
MTX4sFKanJxH86uyLdiKxwOnTmZYqdMeKiLJsJV9OjVtIXcAEybkrSsJ+mujmFoB
+bs8v++J8I1KsObuwBaVgyFHlrpARngyXKp03MA2SIoVofKcVAHY9EQ3a40ejKTt
y34JWubmKMqiFLB1jHupT+vOGHWvWd7aWeeDd4Swqqmb9He72KLq4PmcMfN3015n
GkWC0XKtTniHqDRFzybwp0oO+yctKtA9NYVijL39Zc4K0Oc7yI4fZxzkMOn4Anda
3tsl/Q8+gCusHAvyi83gBLl0Fj0jEyGHhKN0v4nrWanELHda3a5/fJr2jds0nKIl
mQV0aaN7OmdBd4G5oFcHNIt0wsAUbaw2cwHBMhkydOe/uCTFy9nBTJfVqtn8Gi5B
chnlC3fou0vSjjtgUtR1z1F+QYXi0ZoWWZSRu/H9hT6MAQ1wedAYkLKLdeLQPCyc
C7iDErexD/dHULhS/qXLBgJXAV6fxAPeRPiSLXga+IeLQwG7UJ3gaK1t+KiizVzG
D4YH1S3G8nIhq5a37LqfWp1s1ir1zGGvlXbjen4mdBvnLOx7+AiyrNGkXbAI9WfL
Cn8PRWbIc835JaIO3slwbs01Q03xT/gsFud0on14SqrYTep1NcmYQQrw2Y3MqXx1
68VQ8lYrovE1muA4m7YuzGBiyvpqG2MI4S9gKhsZW2vkDYXw+Cj6chRQyDng70J9
Pq53jlIZTrCZX9gZRXkFaBMg6CtxErIa9T3TdIaijRNQJmTF3N+/hx2PfH3bMhCK
XD9AGoaTqX96652kBNFXhNdKDYraOsfaa/Adn5fltmVAvEdX3EIxM8hjIr53EVy0
0baEFA3g5F4METDm8vjKzYdi5p4Go2aUC8V9X1j5PV9YoC3FFc0lILw20+xuvnf/
G5RPAbgtjaagQdnUbMB1PBkpcEg0KVe65fDVIoyUJ10GMoMkxEnn6J0YmLe/TUBK
W6TLlss+uOBTrjvNIVvChVNElVEZX9sMSer33eeA/C3JtlmFNQASBMorp0KMrWMB
xzPV/9GdyKT36EHj3Pmc830jsveJ6geS0OgBFDIDcfYEq6ACTaYFfWcIHKdKaRi0
aYYit54oIzCVVtDWlc7XsN0ysgzfGiVPq7Citk6JfqYLXSJ0xNDSP93xiDSKb1rg
TO9ikb9VycH1pgXOrpbEOpgc5E5VzBT04Dn05kkXjFTdKEn70MFg5gqT+9TLZB8y
9Xzqts9WLTEiRw2WGcER4IGjfD3MjXNnS3n9Iz2IIBF0GWsPt8E5wZEM8bv6Elj+
s5RHvgo5w8cqlWcatNkc4MBuvWcYRqkhLyDZ7NCa+ByDyoLwH5HtmVo2N2cTcUzp
EU2M/9r24vcFUNca0P2T3S6qP9OFYwtMKzyZFdlXiXE9mlQyPBmHTFAERIR2ys1v
bydzjJiE/ddrxi1uZQ1bLwa1QuKIP/7RiQcVMhqOTHBaYYo8FgnHO7fl5FIXPr76
zffry7Ar0ROPnyPKjMdvWCCUE7BDWwcgskURQnq3YzRHNMfUEv/SpxmHsEabgiGQ
PACXHqWcAy6qpYOSA8IDI+vutLMEGMCuKwfcI+htey+UzjDrHFqUObxuNre9K8Ck
lJk7hWh4tVIEIe5KPAXzQ2ObvqA+Qls2L2a20E/gazXTB3Dk6wn8oAdsjKt5jW+G
QiSVK8jOPB0AqkG3F+DlSKPwVIxdMNx/HbB22feCz4Jwj8W3N0tcZgg2o9W4KXcd
eJHOV4SuO4aZY6PneUUbaUQKWDuyNwmNJN2XUPLnEZDBVaZwnZ7DC7OFm7szzpxy
+2YPp2UdVCI3oNOplt/hV6HnR38Xowc45HP1UHpub9sywtCjcF4Wc9z3LklRkeBI
uu8jDb5a/CEo8teGJPEc2ibGYhvqNInHLH9jsbJm7ilqNg2Yf3u4Qwj2YCW6R0oS
C14n3Lk8b3mszvB4xw2kdlsvchSIcFD6kfeakEoxgiGIyWU8xq9qNQh9rlbv4tH6
mQ5STaeWVghZudN5pRFZ/feMyOLDmo61B3FaXGq3YDAR7T8ahYiXP1XnGtBfMnnx
+bQbQ6I1PYgUEl5FfHr/De/yO8HO74zJNMmkv2uFfa3zYqsm1qj8AkInizN1D3DY
ZaZEGaC5KRRRYO8qnMyuAwY7XYh+l37RhceB6HTufwErE/wAygoTzwe2N4PPWzIm
/Lz+V8FjYkMjPT8rN58x5GHHlgcVCkpQw7k3CGMI/dJQiRZ2SnZ98f3k8HKN82PX
+CCK7fwUBNwVjCaKLcE1O6Jyf/SDDNFElOKQMH0hYNptf/cY8g5WQCIPi3/5U2XQ
xEFbmPkAPYoBKU2zRSJ73yT6ZDP9wNlop4CcZa8ikuyPHD+9LWFSOzLeHWcNtlBf
dnP4jJyIzh83HyGg1JBmigssXI6+/dUslBZhnrxP2WUPZBlKjymfCZJImCmngSH/
YWlhlWo16vEs1kHryH9v4w/5NFr96XkrfBmq62sm2SVenPGG0Iz8T+qjpR7Mgs0p
nLeXoo5uidJEAnpm4/via6eUpC0qEx7iXXLQy2xVVaedNuDlGmez7TQee+TfR73o
VLwgE6fEI2Q3rVi4GjuDvfMZRfAcToaMhtTHMuJ/TVOIfKDUQ7daJvTrlnA1naam
ewF3EjCNwVgDhIDephe1Nvbl8RaBz0o5N5H5e70WuFnDG4fFiJ0N3SeOPm8vFlpR
luXz/ZZ7n4Tq7ruvYsoI8teieqKj2dI8STsx4i/WWtoYguRweme1cEwXZbXbKHfb
0AxGvntPd8klVfkEmOgyJVZUYqIls7XMZxB6rV3lkk0AwdnbPXu378Yd+EsYeAeg
dUB7DnkCRaPxX1e8t6U/6MutF5F54D8IqV5ZSI/e0JB7sQESKiVVYRu3bQDJCv6N
78/0nVLEyls489MkR3OWorXpJjIc4Yt8hWl8YT4rBDih3wVCISdP8P4h7hCh33uj
eh4o6wXKSnL4Ts7SKhjF/af585m21AuM6xpt6mug560YR1C9sJygc6dxzzc7bNFN
lUQVQ5VYSVuFCdu5dnaZgj4Qk+lmzOImNDfOe5EG0pE1FZ5d2YwZD6m0bwAt8pcu
THuzUNpd47StkQhgH9GPXFJdnoDXGP2QJd6VX+3ory0h/HnLR0TW4i46Xmb6kfLM
Cc0A97TpFh7VkSSmo+ZiuT1dd8agHgEG7bBvRtQnNPJ4UgXwLt+qhEk3DN2TEChf
i+iNDG5NVHt2+uQkCZ0J2IrZZs41hmtWFkiMClPj1okqXOHV/lW2WN0x0Jg+7WiH
Ka6X+1ij311dZ5RRLk3278lIN5xZmTEo8a9MMEDvkkMQ1tWNvZ0PNMu4ZjaKp2Eq
fpJuL3JeG0B3+fh864Fmc9Mspne+8Bola5zzK6ZarKFUHzbwJAWTxEgfC5j/hl/2
YNXPFLd1/UujqZF8uGHtTP0h6Vgb+u05fq1ogrrkom32fnsGdUvva2KWvPzlK1Vf
r1NsrGyfAhJotS4kuQ3x/Ck3FbGAuvk9mPwLx63hcVenucwiT/S38MHvktBDMzPv
XeLjYt+jF6FI52k0wfPYKzS2rGTzfhYXvp/rBW4QRy6HIki/o+KDsKABMDEwuOHK
e6utftRiZoHfmLo+y0Nkl5VMGI2duAnBzP9Hy0CDIyoKTAQ/KPm62dIWylVImE9H
ZXbxT2oYMOdOkRUqUCtPDciPu2HYvD3XGyx/+9aetCgEDA0Dl1kdt3nUASDhA2UI
morI4BhSEmWj/uTlSrwUY38x5oCXm4fHoObgmO46jhdPGrWB+S+0zqiKfYWK0c8x
rbDwqW8MduXull2LaszOP8PZ3YH3VoUDzDFX4+pa3bH6pG4y/JDKCu34yW90RnwE
X8Cl6NQrYzPwjTjMVxGwRrRB4bMLbprQYb2wmnlJykGyvfaGAtLxWRs19VTwA43n
v1CwcGkj9edxizUbRatxdw01LaDrT5D00nFjJ6fscHLebsmOuMMzsTN0VFFof1P3
TLS2o7WssqLen3eqB015Q9pMsR/mbv0wjxKfVVRkrR56oCqM4XKwLeU5m6PSQRSR
3OcEfRMVhG2JU+hIJaJGiTJGGbqK0ixPjVZgg/SEHhLm6xGp1Elc5xMjlT7BAh10
fqzaNvLTHhgSnKePPS7FC2+mpLZMKw5VS4Bxvk4RhYFSTYF/BIHCdhWPcZJxeNoE
nh+NGQmIhNwDV9h5O8B6U3c741LBkVOyplYdEw6odxs58ZmJd3VYGVt0R/N5xYk2
ohRUO6uBguvIhg0va8+R4P4/KOudhpTHcQr93aG1OE8x34s+uMzjJjnVSVFl0whU
/90kdjMNiCqACxBm49EA8kmRuGHiHWXHktda+H3zEZ1BpovQ/FGoqPRzICTml54p
ZsAhOpNGiWeAxmWLQnXNr4oqNVTFsI/niJ+ZXYlp885gEZUmJTyVs/MRBX/wEBWy
+YnqKKls2HOzv9QCYMUrLxSCa1XGKXcATw4MXCFNrfBVcB5AiDAWJd4Jyh1LAU04
DKOE3Ljcw1MGjJLzVCF2GgtnjlKfdi2jTN0ShhEPNr/yZjyVBM0JYwOwzyqC8b36
xOOpqFtjAJCns0szraPi+doyuSGr0J2sWpMxZ5eQBa86SN5sfoXAAhJFvvyGKI+u
bxe6U3yOAWRCRDSU5PlFsZ+Gn5nNlFMBLQ/G1DwOrC5L46lRe/AVlLzPcGFdDXpm
QRWXGQ1gUWfFLYZck6ECkeJa3Rt8YiWTITq82P4bLjHk4wSYtqZKX8TRRFsKknDZ
f3g2R50f7aD4TI/E/fBKhhHGjrOsLwC7lWsMEavsn3iR58xXYd+aB7RFpYyHVcxu
bRNP1E5OGXGodsWquB6GhpmAnIV73DQHg5yvR0y3A7+I72/mpeaXXOun+bRv8rrT
YfnWH4+MIUiX2AB5u6KzL/wvY/bB8PFnfwRcPBothfQA53FjqGi5b3yeizQ2KfDZ
5l0ywZQkN5X1vA47lKT63zXuScgt+xKvToLZoTyrcOtmBvw/yTC+LIGO3lGqcyP/
7mfpPCGK5z/folcsNUi4Ov9+Y5fd0sZlGad0rwpEReRI4jAKTrSJPAyziCQUs/lB
d8nTXhU8WDJ2w/CcsCwFA6nIiU/juhN9IrnGXl0y0KWgpuJJXU11Yb0ws9dIO0PQ
h2prfKElXMEUJx9HSbOq4/8l5Ql2jBrxk+0ZhlwhlavVYEzpFYVJpxMEV1Z2xuYo
0RxcvZSm9PW/EaMZ1BX7mhfJ15/4H1e4rkKx9DBI0wXmYGAuqGEQ9dILnd37vtJH
bp1rQ6c6D3rwoPRDWU/X/0eT2pfyqoUxEA52PDqcJEuLh+V8IlwwJmsSbRXXSr7h
b1LkbSMc3T1RWw9+VDnoHWpFKsWNrEcFdNnF+S9TccZ3lIc9M+ncsWum5Sr9Ik55
qChcgvq0ZRlF6cNEvNUz6fU/oDbTwUmgH7Lt8MwhcJ6sm7pqllYFmeDYmTIR9btV
z6niAQfWbssmnTHpsM7r46714D+NwQs0/ovx85n627yT2JwiSGhpZ/JXkd8AuBx2
ISs9bmpn2Eu2hFgZfR3EMPk60fz1ouqeyb6yaGmtMycYXJHJLSBnjLOkBLQ6QejB
TJa5mjjpDV19AHkEjZ40a1AlB3LiPaZXKqMV37fBALAZeS/DI0dzuEig0KRMLS4/
8HGqNLMk11xlkM4HI8jrpwP/Y5D5BgiRwy0GhSLv6KtLjkmY8KzBYNgjsVqLC3oT
J8YuGlGRSgMmhHg5Z+ht9rgY1YJGn0Ecg9Ely733Ck2J7aOgCFZZ1bwFoHy66AhO
iNMa+Q4h7EHx01IYOEN/4RNb8EdXEXGP/9E8Iqo7ON5DkUKwY7ZD+QSBYrdQLfva
xDgEN2xLTmE9vaVd/POI8zVfQ/drK6lMR0q/LIK3MnHtDW0BbOHH7HZtkiCNtdI9
hECTHAdmkv/UYlYDNiPgTsTpP4rCwU6wPQ68FbQgUfykY3z/cCnKNvdUXoxNozut
iTZYawTBw9zYTEjMnxiOnlHiHJJ4uVk3caYc71T96dwwQ0SA3Imx5L7OMXkvG9qK
jkgRu09RcK0XZ8DHpYKVdnihvHPcRP1gDZ1xHC48hvxp+F/WwqvFf306XIK6MERS
GALttVzAUH2bG9t1ydzTdhMK+VHPlSSXk1eY+HYNhv71uo6BEKNW96Gt0cpTPYSq
NUpt8e4D0ddhXMQLLpmNwgnmbTqZOje8UQWviRYuID+8A3ddYtGxJeX3zYEVn38/
WZ6ruh9iMcWrlked9bL2LZpDjPDUTuY1Spt/BAAu2PL/+AnzWxDYmPB2pR3hKdJT
TkOTn621Wnp7K507R+vnRdy5vOtaIudpSd60m6jWYr/UuvPhaegVJ34Sa2r6MtBQ
fw5MCD70qUHhbEqD/fnEGEllE9nKEa26yexiWQenPQZhHy0jX0IzwrwOZ4coj8iK
z9HxM9bvFkqHa3NR7CrT/83K52blkGtvi8o6/lQK+CAN0y6KrJSGfixoTW6yW1mx
Tkb9CJDdcnO+0PsjLPUZDWEF2NPzXGcz0WQdqkKupR0wiu6n5FsHg0jZK7FGOZ3w
XKy5A6WsOONLZU4WneIAWVJSPYuXWSQ5Qa074ZxyGHrR/HqSifXs+C2L7rScahdB
9rfoS/l1LZKDtH/uMMW3zojVmHozXXNVS7K1pGVTaNuAJLGYxDoP/9YVIv3gbghh
TPxB1VKLv6sObSdrylEWs5dsL1b5hqRwJ6IjKVaElxVwXKjcH57NLo3rin/qK95X
r5iYmTjgpWkXYG9rq6WGRtoPQmVL74LC5OuYSXW9BSXdvfvTrDvtV6X0z497EBCo
jZbTnslSL+Nki1VqkS6a0WN8DppAyzjNkVNVrEgTxlW3JaF6DVO5LuA6RjDOSSWe
DJ/vPCrrwdJcNZ7xcm2k8qGK9+U6N4prKgS2H4AY8zzYZ8kWUilsSKsPInIfenqd
+Byg6UjaGKG9Atw+Y0k2+fnglKw3yO0qbaoeL7LHrlVD8VW5I7rD7SZc1GlkPl+a
//vHGn6pEvwXEVwXlVc7sAkBx3cFWbA74jOOS0Vo21zlzYhS/If9gXGd5/PDNF71
5afobgZyfFJW8kGU82UJtcGa1eAnWJwRj1UIMaWY7433nVEuGWCRKT/0aNdP4sNJ
NWymsK39h9R8kEWv+9sRg1Ef5jcB8m/uF/0o75GsD8sA7DZD3FE8xywN7LIGXxPY
CJvh092Hw8/7VVSbEzIxgOX7txOiCnvTvZ/vweLm6qbWdu5WBpDq8YCd4DRoe5Uf
cPd/rdR/IoiSYuHTckYMrqGgvEiVqEPcedKbX8E5nEmUQCoQktGLpJWdUkhqBnWX
MagyB24H1zq24P5fClgkzFVBOI+D1ZIk6pTbnaJV3CNWUIM1PgFRbsBuYmCsVayY
axu2OzgVYetcqiLV8Y3bPNz58MecTE8XIfvlJ9kvrqpRoZE8ufIUyqhMv0uWUigL
4+/xtUR2cDgpru1kwknPEu89hwv9vpEA93oNk8LqdGzzlGGj7FB4/GH/s36tEYb+
pcvC0VNSP3zL7UR8mM4ee1dtrn1BH6Q+ukNf6+ZVsczA/MaWiRpW0NMGBSdQymrR
zhoN/tdFnl8Zl8gRAmyifgq1EyBhBtacYdlnl1wGSJoKMuwtR0ubLmToBTJEGOmo
Vd/558EJ/1SzzNDoo9wSCtNt/at8hom6gqugplC94i3UVjNjo81FFWmFFsw6QgDp
lG2neKoZ08WuVNgFp0QbNBD2/or2AOH4azShlfRvejaeYCAL5zvBujqX30KdQdVP
zzaDiZmDzCv9uA7UvHXDuGq27K1BshaY/qPv+ByumloICs8Ucr6k4/C08CsTqXRU
bDHRCF2Y8T66d2NhqxCvODTyaE1hvrVZpiP80mV6hpWyopPaIGbIaowiLue2DfIZ
4bXstmTRU4AmfmWGdEVCvkSdB+CRGDglLIZkttASMtmlicmOz/jJ5PA0A3/19QNT
5r+vJjAX2JGIQH+V6dY3MkDQ8k7DAIVphdbGokW22ptW62JRZDFCOuht6LB6kHwC
yCgBhWkldf7UtLCczocl1sTJHpr2KI5w4xj2aJwym5seGlJRmgOnZGzHe6aP3YjE
LW3pUiPxiGrpBVsATzzSmPWpwDYWgtGdHjSeSlgTsgzLq3Q675T3mU1clCHXa0Ys
9def/Y/QPy/3ZohcXptBJc/RSNCAguj9qAx/5pQ8rA6emEKzn5x9w8omAD0E8HlU
A5Ej1N+otdPKE9w/yWf6INPaHDPrrniGR3OIHn3X9jmFACtyBcI4cqFHiJBh6AdC
CGywgqAXyTHHplA8/nnuGsuhfT1WC/Vm8GT5ED42lJah+duV++MPyGIjmetUSUx0
d6wf4jwHSEyTANbd/e+BIxYYbp4Axnn//0PY7Jb1G5MAAuHi9DDvNOP+s1eObSfJ
aEl3QtkjHS9zSyqu8OegYutP06yEyrVx83A68VRW0+n7hqm6XlkT+vC5rlPStNJ+
kp4Fax6iB/RwpQ2QQNS3hBtuRdGz6UwPCEv/X8ThLSqj9bAH9AgS16Jnr3JGmUr0
Ucac39o6t80R25VBvfvrhGrGSg3+/OeiGQ5TLZ74Gzlm8DW8v78l3OD5QeSR4qqP
CyHQOv5EDOZ3QuVagri6m/RAGPe02w/gD7bTvNxBWzS6i0apn5j7AlF9P7Eb8dQV
DaXkXHmh9zKEDaTciKzanpeVZfu4G1t6gWHmEAS3QbotFoLM59/OWE/QKezeOXVa
4KEMluN4BnCKrWPWs1vZV8sx4r5B7bAurn+ilWMj/TXOxbJltK1KXYzTDCZAi97A
Ce9gfv0u9kXzxgWYSo+NGB+kwR981kN2P/rEvpAqTepAYrxIhnToa19U8KUZGHR4
qYqK8Ckh0XiGPMJVxsCRppFrmr1mRCareup0ZiHMp5hRAPdNQm70rEsd74TrMwLg
6DbxF0v9wP3s29mj5pB37IJS7DtnQ10/P9+BRT+jUWPohHXDUX8/Td/+xSVjQF0W
a4Lm4GAA3X0ZRkYcyKBJg04W1UckGAfTWikcFcgP1+lAnFzz4oWN8+ckY1ygqv4S
LJ6Jr81BtRi9dtj/pQul9crTGKoGrnPDBrRzvjOdgJdDKZHnI5VSz6kLq0edBkBA
ZFO1MHE2cDIOrwi/sLi6tp8GHoD7TxFGKmEMUxIYmtGFXBp58/r299AWZstTWdV1
7J9RNgRFqLxCwCFX1Q+zghuOSU+6wOvakmaoYwfO94eg5g/PKEERTXgSgV7b/hAl
oWDWo3FgOfWTj3XXy+daSpmDj5DCSbscVHm9sDyQvVLrwo3qYLjWH4qC1N1C6IEi
q0az7HdLGm6ZCMxvTBFwDQ1TowBqShypZkul/nITm/+6gmqbJZU4vxftGHzQYvHb
FN7tuU05afDyKJa8e9ggjssZO+Yz1B6LRir14KGmOgPvGJBKgda7GwnIQI1F40RM
O80AJjepwr3f0h+m4mHO9owGHEzXibgr33Y+0Pu21WEdIz4Bhd/8AALm2RKMptnm
VN9RdV/EtiK4mn3EonVaCkNJs/fBAtw8SuIq+b3+9KGeXlWTQccdMJZsiiqXjpMB
SajNF5nXxGiIMz/cdByLC4ul84V8LGi3SUJk6/e5g0qbSD9U3T1YtrZpzUiMjfkm
yPtjBa+qfEjb2oZXClWWqY+8ns6QxdgUmrpcrTCOL9h5iJkpyyrwAc8Wv+QrSn7/
DGlvrPo7B53U5Y5pjKAGDLOFmKvt1iwVNLHX1lNGf7kPgAShs6z/jbu1mCZ6FVln
vGToL59jwQ8b3oXGfK7I0qDAWoNWZz6XhtOKOBcZoMGPLmur09fVliG+0G5qxoe2
XChKchlgpm84yfdG8GnEXoHFg4czzEw20ZZl1wgrJXeWev3ZR02NbWVctDTYdisl
9LNNTdulzNtMyYoOg2ZGj7IBFfThJz6PrzVTuKkIvdkzkkqgtwbnicwjsEE9c6r7
Ec+wQ3zakpYURzIkrMaWXHA9ztE6k+Mcpa6MxSGUkwbsmJusujalmT/y5/w5g2iD
LB9cSE7vSJh/x39nsDrGL1gfqw2AZMAVo8slYlJTLou5GWiNvkJWyLSzrBm3ikFx
/y8gPoQYkY8bMOkr8Dm7wrd1ZJ7EUHFP6JRw7AEFCQ+SUXUN90EXg1qh6VXt/Ks4
2Qcl9y0TWvhVS2cCgq4fe77Rt7chMp3BGomPcEg74JvYzQhzMaMUaRDpQXQR9ejX
PAfpZvXsVlSLZioyrdcTIVhQdOiJDO3fYLpwtelbaStQ8o+WfY31ZsZCZEcauWpr
d7Is1JhKbtiuoPIVd5Y2GgLd+rXdA8lg5IWXorK1YakOc9MkS5HGvNByzoeUF4CM
c5znpW4D6Ry996xbHVyh0UDd9EDKJ0Bmj5XZ+9LlG/Y2dcvW+YIyyp8A9YHprrbn
1FcP4/W2G1+q2mMSblnNUeZ1kMKnsEJdadoxTavmMG9r+tIF53EWgXy8LKzbo8Tz
Y+ikWbfsDymgmSzkK/xFmnJhZPWjEceZ8eQSoQZJXJ5DruWl5YXC3lSp9D39hvXk
ImgJtvZBcBG4Adrx1zE57+aaby4wf2nmQ5/w/S1vKB6EqTCiFa8wpjNPsByx2W7f
YV9g0W8rQOmZhTwuT5nuBkL18mRxrha938igBmBzvWwnLmOed1I9hZctrKv30/03
GY6P19FWjhW7GdQhSkXufAkd7PUdYxApj3aJuCZRi+oCKOzmpfa/xsGWYA3s3gwN
ql4HsukFN6k9ojKkhhTLvyvvHEI11ZMJjIM2R67vYwyc3TOxIQ1j5n7i/HW8KeMw
DG2VhG4oJKC56DxqLF1/UkbltIDqcoOB8N9paNDvyV3IdRgapQJG88n215EaWqB/
MCmdmdyhd4siNpDo3BtAhJpYdmFsHAblZskm9clU6INAt2D+Lp/7pP4ZePwmcqN2
62xhg++saXtU0ZHnBE0ZcS1zyk2KX4JeJHpdoZYX9N2ApT6bf60rWtNCpAL+mhER
kp7+DUXiOQLYJTgrsykltR7fQ1wMCeLkcLr2YtUIY3QP/G+AMP3Yipv+btjM1lsr
6QekWVygrdSDjAJrKvWLowrHwGEVrYgoxh+loFJFbm0kvZUt5CzSQXWgY6ZpzGpK
FsvAROIgUB4HwHqRJcDt3P6x0PWGnSMWPpRdSvK5T1eQUYBlST7rS8vvunmA01NG
nfNT/KygX32vFTZkwdFqt5dY/RqDS4IEcYN6OMbPM85jp2pM2od219bMuaRwZs3w
fBjnKv1fkZX0DU6jzyysmQypYwzxoa7nE/V7hn+r83D1q1bufamZPu+b6+Abiw9J
kkkcNX+YQhyn3+PyoNsR3xnBp3QRJbK/MT558nsHGaDXbH82YU3GneiNhrEerNfi
8kWty3ruFoKoOta1Y7fSHwnjN4fYVagn23J4tdWtKXOHlJEXMRFGr/qpoy6u7iaw
F9cWG1kGIR9zO9YP1AtBF5jFOYZ6scC3Uin+BOfFqhRNE1LMd18J+dQPF03E5WS/
htC29qXDoPEwLey1KKQ/qnDid5bYwr8aFgTHFJv31SFE7vj9qgTlDDMm/3Yad4H6
LmTawwBfZT5kof3b2kFbUszOjUo/x5PTGkKNf7MMzi57NN4gfVjzWHaZzlFIxzXP
sWpDlsbCpQGOj+nZtai5OvJILEjN1LQxZZd99FM2XOhuCcrGlPeivKBoEEkXWZrc
lAF27KVWmmwp4MrIA4vqa/bWYtrboPjnu7UqV67afP2YscoZowcQMf8ROEVn+bJK
BtiP8/hPF2aBiIRyM7ssW3jJJ3CLfmxQa/eYMJQnNYeGC9tTIYjqGBwVMdcI/mFO
7hHTXrhY4hiBJpGjFilYRYPfe0xoxqxZQxWXyJVUW0O5NXlusWRkJYbh0Gq9PEbB
E1V5ymi5zJydcVXl1LvF/gS3uwk4OELX1fiU6QPJrftTNZI7j1P03x8fEd8mI1SH
YqIIM29RbLYKpIMTuAceiwjLax1LuPhF0uYiuM5Ef9m2gnbGAc7ojb0aQcGbbHkB
59yX2IUiW11uuVdyaebEQftf/1ZROGhUAeQ+SyQBC+Tt6jIkwTOGN6ds9M3WPpi/
BNFFMigiAPlP5IKbOXbOBX9CZ9ogIM7+pdqJUbKJauAp2d3QChrZknmJ66vMTSo7
/2OE68qLE0rA4MSrk1bVzYoio0kGwDUlw/igMsarU8POkzyqDLPzVmp4yrB0gtBm
JJJ4cMalvcWK8JzgiGp8LF4nV6QBqgTbcPRA6j7zD29tUgbQiMYKPSJyuJQEOt1z
Yh9wWh7dGAHwuzhJE7JnQNJUO9ihuq9uhaOBS5UL1C5sY42a15ARkKBAaUaz5tQ1
+6kP/oq1h+x1CPP95vskSKYhDqcELpEitFjG+gfvyp6B6jmbN1RbAL9ZApft25hF
hO9L1MEEAZmUxW5oAbQF4kmv61WouTfZPE45k+2PLe5ui+zy5h1Qi/fhTb0O7qVg
v+FlR3FH7tFbul7Fk3O11CRb6rhladUXYY2NSaq5wNPQaFOYuON1+l3QmDt9jLva
oNXsTzWKeHJ1CmJcM/Pfig/pQjY1kgPbu2948uIRgjwVr5Eg46jO43bYKHwyr0Df
Ggdocf5DB6GaY8s0+G9EwBBQTkIMcaeNTnmllNtTfXyBtUIaXx0XpIESUtc50UB3
Li1ma9ogbxzNourP1RPYxqT5wrKgRE7F50pns1jYaEq2SSrR+tII3DA4KXCFk7mL
TM7mavQ1MhVjw8UEuXQn7B0AWRX22GX05oikoCA2AFbdlZSWfkNpPYF0e+rudeoz
H2hp+k6/h6bQ8q4T5MmONrcheSRhAu5jbp4nLXijyu0j5insrJDN0vmbl/Gn8Wat
YoKdJdeMPDcYzy5hLOHTwwGfxiNYso5LqtDhFgBsfmpgTIKHODJGb3BNXsY4nMyH
R/eQDOyOa7Hj+PMigL63TyEmYelcC3MwA89eivmifZFI/NxF92N0OhkCBVglJDjZ
DNtw5DkdQr2jmbsd+RMDq6ksW5Ft6gtuSM7d70Ql7XJKu394LXZ/LcW4++NjQ9+t
eEUz481jkGoLkbBZ6p/TYoySHRTCDAs9pfP2CR6Eo6G9EuoX7RGAoMKeOJnMofxK
1GhJec3VCKh6vYbzUzOF0jeVNp2thmW1uYSP4R/zX3qs8ZMs2WwBfwBm7Y/35q3a
LcU8k7Re3mcUnvoyMCaW8Yt3byMN8rFm6D3lg5FI457JqwZA4xZdDdiAw4cYbqzP
DIdl5ed7KQjTfyM0j2WtoWjgseQnIunl7rOvv9ZugM+bhx5mpTS818cUp6FBx4/I
2bpJOHjbV4uCu1+EyK3HClgNSxTvToucFoOMcwU1x/s/0qipm3evlw4kF+ZtTXEE
XnrhPjdvEB7juu4GGICvRAqXhrSK0fz1oUKBRPst9zGvRgf8wHTSeoBtxga3gwdH
yl8YlePMQ4Q9bx+RHoqVBdXGNUKp3+wKrkhOZuOd6GC1vxosyQ/8IJqVwvr3MXQ8
tcEXj+tc6y540+zEJpfPFZ0bqqTyGZ11BSTAPSyhPSLhGSmhuxH3EDZtA1PQQRDN
hnG5Pzwohtzz5ddvJ8vh0nqQmkJsdZE3XTL5Vy24pWBDifmFqopOKKN4xz8EV8c3
dlAyAW8uSYocAcobRUZIAymLs66sfhLapNwUEo4Yp8zPKqaJhQObr1m8CPaI7kkT
44bG7SwN5F4iT63IGYqCzt8EdkJose2FdGBNLyCdnHYL4zSiVKtrIzQ0lff8m6b0
6JFIa/N9inLyZIe36ABGP+oV9HIHus0XJjfP3QXSZXnwXZh9vLSSoG2pjZiswbSe
YHQAnaB21fiJ+FO0/AHRQbKXlhYyVS+UUIgGyV5R8hBpftfyHPgST0Iun3mtVufX
jdHhQ96SAs9Z2O1bVxK+/FQXhEdDJXviFmvr3ifRCWaBSJl/KBXso1ApfCsIDzOh
jB5MKwTMXRwqw2iCLwBU2mIuJFX4sjXjZcO4B8MtpDlWKOp67uR5jfJUYQyrBpiO
/GC45VJbuIsgrgNLulnqJK0gZfrHJEmhE734Jew7bWRyOqKdvlSZKfc62TtHGD8Z
iuS0SuBk+hTWTI/IipkHZ6rmJqu5mQ/DuDwK8xzf2d4MVFiQ/7ZIDUuMyOm+CBan
eBHbTCtxi4l1NEkqNeDY++MW0O0sm1mC0YxyExsYVD8Uyqm16z/uFI2YwBi2B+uM
WnsRBTyHrwdyaF4aB1fiLFV6MvNK3m8y/IYx1A9mKwjkOg6K9u5L9531y40ME85n
5HaLj2JKazc7+ZCK1N/JEFh40lYPVH3VKfEI+AmdvXiDqwOz9ArTdu6kCPYZXAvf
fCeqWQkaAK/KUk82wQtSFkBTkA+pasIxM5Lhsi38ktSmaMxjG97n8V7U8KF7Ya84
b2+zaYV39wJ+YWo/RjWvk6hDsPOajbEdZnI0obMCBfncv6HnmDDQPlzD4fQ98neC
vqL9xshTgIEcAXV5X4v+M4eqATrG5oUof/rqLzF1eQRDyN6szkREUPNA8vzUaGsk
tZSxiZf/Oa3+alNmBo5Wu+rb2gGDnMLhLECl+u4T6aV0EAJZO//ujMGpSzl+18j4
zSxx7Z/7NGHqw00N1i+O4o6CBQmUGOI1jFd5yb9YiY0k5A1L/RdP5xUeeXlp4TXF
FB0xJjJWzti1XeNXrv0CwFlaJTrUdzDWceUNYCvQDPcZVIx+Fl8Bjt7BjVcU1s5b
4UdTb87TSoMchbtYK6mHLCYLA7Wvg6QffDxMAUTyoDNA9Ppy9R4oKB+efmw1vPsZ
vOP+jV0ShW+j1X04xLrlTRmnmPI8Jg8aUA729TZrT7slPbvY6jEHVhawPXf0i34z
lSqPheCGPF74TwuCgBps6AxzM6ro2+zsIw/+S5mOddAHGR0mR2wEg6I85/FTVs0u
+qP5hzG8cJzLjAdnA+Eyl4AYtp9fx8Fbr4n2+7/A7NFizMBlzjNat8BYANeOE8Ea
kt0x3x0xIcg6idvsbRleBDAD+ZhCaoRlPukHp04/M4xQY/9PW3Yxby++gFYWWLJX
PMxch3GTcwdXl6r2q2458BH0WsCBGacZ9/vVto6yVTqC4JdsWpW6sS+AD5zgzjzU
SqMREfpQT15/5kOt44PI317XKvniQSup3Gg9dhdFMU5VcLNknkeersAScB1uvttp
FKEeRzk1ouri/p0tskZyyV0sn9k4j2rqKY8+kOqjIJcrGOxWk1zUvPP6FqXrmsxM
R3P9NqIB75vrZjA0QmvAZvCccNi43seVblWNUFJfqeWidhjuRoh5r4R3f5GUZUFS
r93O9J7Lc6i4VQQM53A/cyzkLZ2egv3MOp1e3wxdE58oxPxAWpJILzCZrZbUc0mU
vx24U5SF9nKU4FhbuihsZUwrHZ6ScbekK3IlmnUMy2pWwjg87yfFgWvL/i1PVoNj
NVsNfoqo87HL4S8f8H1hVxW6c5R+FBQQyIvdGKtcL2JyURAnfQvfhpkpxeYA5VKr
zi/QFnU4N02YUGe24M29aIyEuGteBziAjb3nO0nXYFpsuiTSBkZPe2FtWowgZJmd
BmBpi9Np2wzHDmiB52jMTRN/mE/oXFXjJhCIPj3KX3SDet/An6EgeF8t/TWZ3QgZ
R62Wn70Adyafx6YjyUVk1jOXuO4lrlxmR34tbTq5Piuac6YN0egM+h47nrQiVUbq
NdJSgU8gheucfXmJpZvmS/20bogDsc2IzPLJxwAaJR8fs5AKS/jcibPEFjTOJ/jf
klQC3ZGxFVFhlQybMFmFv41Lr617hiOum3+VXVAZL3VxZFP6ub50EtkyNn8Mi1da
TFLBTX094jiC1G8gYDWRwlMkZSzfL9fxQY+bVUExt6ptAo1Wt9+hH9jFWa/RB+cT
0Y3lHpFS4ZTg1EzfcJzTndfY6kjpvZyZtxpTOQbT5ebXHnU2P3+qTOg2QS2kPn7H
uJ/zr/zcEpjJ5VZ7iD8vzro2jb0QwCA6N3J6emzvCyKdFNlGhr05qat/PzyCgA74
XosSWx7zdSznmppYndJjyyHwnb1DE4In5bDOcFEGViu3Fs1MeWfPJu0IoVssE9kw
0gMRi/alfefh3mD5+xSbPqkbaC8TDoXH4/aczvZvPoXGZLLhQTCtQfCP7Fk3m0Ei
AC2HJ6xxNqgFAahcvzueLxelYeZak//UIOxeS4JSl5FrcN+HEzlP0r5DQsxqliSv
fGmKJkNlW3Z5BcQn7jPg9wGu3kNLf+8pmNCnseovpO4IMeoF9TgRtyBkT6txHO5t
GORHHsMLhgjUmtAUgYbYpGNMNzsXCyRo2kqNWCPcs2uK8RrhEtCbGR9Tqha1hPin
zo916wsagpWfQuNcJD45pDdSRkoIdsukro3bYXpz4bO3GalzC6uftMf9SRVAcRVZ
nkdLYzAFa0q8A6tOjCGls3IiD55HqBM/zvdPOjeKaYTLBI81nBBwaSNApoNDxNqq
kOTTqN9RWyvq4hd4fqRhclZcyNkYUU/+nIkcam4itZEXQ/+iogBQjp9I4xM61pLa
M4JB6ftMQYMi5SVt1O++X7Rwv6V+dd+vP5O5llhtQy2K2py0x/MoJOel9JhC7LLx
DkMbtYCyCHGeALmV4UFRTqxV/YeUOjItmFbVrQMjKrq9llQndVp9WW4meAuIuSu1
yFZRHoE3UVvMyt2RzFJgkZAWlVkL6noVpIkWh1J5QZWKIo/zWxiyS97TRSu2C7hk
8t9EWDTqBWMSL2s6XMdSC3u4JTdK5R4yI3shCeitz0dZkIfWEQgPjl95OGpKMkkq
SmcsbjT680Am9Q+YOVSy0SVv+f0F7qJB3NYPb4Zz+gE7QAuoMekXXi/m08xlfdd9
qtH01Pax7a/8asWZiqlgoVZ/+nihYw/zaN+FdwqNAz+R25AfM84aPTXEEP5Mv/Yc
RM1VXd+LmFoEC3PWuc73pyQIsN4vabC64eDO0P8JZRq/6FmlSQoAZFpS8rQ9K5eW
YaVfElEuSfM3tZbz+9IMe6NhSziSFE07u8fmHmYXXRBIoaZcLws9Ua3IwD+f0B1O
IzDGuUdY67jbE4TpSB4Qp+VTJeWecIEBktugmBg3udidCG9mAecxBDAHaFMI+y0g
jb1ry/0yNDtMP9FkUJSAkj7Xi5TwEOdQlBzjfSAzpHqcD6YYg+rUA9UWaxMrqCrX
osPtfmisgSnu8421KyQDFyP5kP7fpe340zPjVBs71hQlHzFQXrOQSb91Qv4NVBAt
Pw9HI+kXDrgEQw1Nl31FbkjZyESDKBtULbGhov6kOQIlkRtOStj6ftUYFrW1YkRm
HRCg/DjmOvh8zH5XNN0mA5kHVILN1y0+gcRhbwQI9APmB/26bdQdFTs2YIqPItGe
HNJHVeH8hx5eDK2gUJSkztz+rCY26Ghto/YKuYBFWEmsPmcJchkJzktUF6FMqrcS
uH3Rc/p2m3NWOSw6PalF5UYAEg7XdU9OvFA70ARQ9p16xGlkYt3Ie27ouD8Bj/Xc
4NoKARaAd+B3U5IDXb0uzZc6wy793E13HAH63HipaVy9RMHfGtKiCkcnhSQShguU
RiyNOWKkc8ZCdwnYFMNsITae4eS6cfLSe8YuRMMsQVfTEMBHfNEPkxTvCKxCobqm
ZhZ4f6NW+OeNqdz2xp0R9yNfyOik8Q05bmipiySW9mY1AYlx2mfQvQ2ywUzSnL+E
jWNPqEQU+eRIX7HPEqVLplu1gacbxCwI/DfYqHuqrayFqhFScEwLbnE5PCWfur+u
DBM4CH23K862gUWF7qLmeuLjwd+UBSeVaWXB1Cj1aYbIZh1TG0vkOiPFgtt8WXBk
uTTSvRkMo1ugyVWHbldUXsJxfqVLUmVn1B1bFAt8LPz5uCS3ouKWDkMi1xmc8IqG
4SznV4kjM6NsLQpAxk/oMiGJAg7CLegYkuaHwqCCVbEWj6Ry7zGoeaGF7fz+xa1/
SUFvK47d1jCFOmeJsIuBbnOgV0Fy2FBn46tjWR8JvlJrGOnkfUCu8g9qrsfPhtBE
zAjepI8/vFqDsKmYil14K+WguteFayD4afedijKf3FEPUyoR6cUwHRl1BoqLHuph
Q/Y82H+Mhkr/NJ1ea+kTHD7C9JClhHwVQ3RUWKyorR1+1cgXaSxKNENINqUUXLMo
vX/PwkvDfMBSWFEjv0nd5udHqL3j2VbThuSujAWOhLxFyaKS0nJGLnOMjqSkLSdt
QYUl9RwrQOKqczzXkrdXJobZNvRr5wGOc+WdjQBXKvhzYxOwwpW/bDVHI2yDBt62
X3qPEaaSwFh9Z9aMmQMZwxPnx5kTKvABe2qCVxU95u5meukq3WnSjijjYtfNcqdI
+urXzuBK9ulPLAw/r0g0/XPODbmGA4D72M9mXNGxG5ua6Rnv8ffI+TzTgYatZSwS
4SLsxBv5xnoHTpqNRiDf4WWMU8jSOsu+0+7/yf9NKKaxDZYT+R2nkKpKqlq6aP4Z
b2mWTCmqzLj9h11tDbyT/86i4/Vl9kNQo2gtWcBdL53n2foDCKp5oCAG6rNb9co1
KGbga6FgfZgqnx1+FPm+5QB39SO+ZmOey9AVpWoFi/fkcx1nfzIuh0yRdRrghZ4x
sj9iNd564dMEXRZC7tpcWuFXYDzFyneR7kBsBRH1wgCdiMmUlCJCcntBdBC4k2HA
jm2rz+9J7BRGLdXdqU5CutG+hP3dxi+mh08iPN6/d3qsacRwx0ivNbI4kx33cqmW
hE0zYcE64IhmWuAXDlC7Xpa+vUH8XvEGExjRvt4ySTf5cHPKEl1yx8Mcy7gIb2NR
FHalnF+A2/11fZCsOZ8jydCOwq+/QADV+qqqbU/nZlPa5ycxnAEgDjhjwKn1vJW+
be7dFCRnQ1coOoTIbBO5cFISKFyJ7A36hNxeAuYcaRPhMY7O1cWViXQz0ywdmRb7
hwZk36ukWM/gvxIDKWX3kFIY80kpdr/Km6uAw3xf+kkknmpDB7mWnhstkRZI25bC
bjR8rix1tfTBq1Dw5vtRw+TyqfHJ2NS6xOjgUMOVOjtrbH/NKhz+26pEymodEf/J
x17PcdxLF+pMMYymo4T5pHy+OhWsrfEV+rcf1NIYxqx3L1COXswFQEX3NcRbM1sK
kMe+8tcLKyWrAZ8RZgaF+yZPlEzhPNtAlw1pbwO4t4OXSOXAXWJ2nYjH2c++WPzn
/vWjTpfJ5k9w3288z9pO38pHzwQ2EgAzQgArYq0Ojx+sAirNyYq8VAHZfjTY4ZUr
MpQcy0W3NAo4hSORFNylOyO+Eq6rSmrzLpA7I5re/wOTFn0phAFyTRO0rsB7HiGA
WhKNuloGXYR56hihCKC0mrTQ+u2G01khCkaX3mvz9/Dxre6E3CkKjBCB/6NoaZjO
8YnQ7ZH1vrBWDkCzb3g4q8jFQOmpRHvuuCE3wiOs0whgKzHXqPuZ1Le9YZXt8wyo
0DGz8/za/ojqN/0m3o/C5VxmfX7qSeUm01lr6QnrtSwdOKSQkKFxDRnWRUjwVvOJ
fxgo+kWbmTs2KThrYqeCGntaxXYD6V8MjJbYMQV2ZEcX61ERnn6QaXrsqjt7i9mt
CQznG2SdhDxy0/koOeiTabFSl6BzOr8o01x9MjzM932eJ8EFmWZKaRoatgjEPU24
lbTUAYHb8+oDLc9E6kC42jTrjHyO9HblZG+UqdzzBCQ19KaIW0Bs82hpxtfK5Xmb
KmMjbHf+jneMrGVXtDL9lCKdfWdgA7aT//Oa4EbUJnXhK4upIKwYKT/3ukY+e+PV
mCkhLikYAoB1LO8S30/C5BEIyg85r4kdkAPetcCquiFiDZwrGRyI0KePBCeK6G9o
7ayHdw/wxHWofg3t2jm4neh5v/AoWYVg0nJ4qG2yJbwpBxLTbDhE2sMR9+W++YvJ
6xs+CTkasSO40I/wNy4Pj8kp+65DKSroG7HB4q/WKBIwhyXUCYhZAdei93PBJuQR
t8pFKhN0lR6VOiX6Qel6B7+qPQMgtxw9K3WVj8oJuafi8cWykduecr5wuVyHJYyt
+xkNkdw7BgbROH6hXwiNQtZ2kzyMyGrbvkJy8iRR//QFJ/JzylulkF2QlQHe5Wiu
LhofQFv/tmR+J2E8uRJmIu3awqdb2kaO4CpSMjmghFxiVTa/KBXxj+D11ySfPLai
Pun8p/uIUBbx81aTur+8/028A9sbMC1KldKsyjAcnu0mJubXxeh3Lqq9x20OEE/i
2d53LX8dET2z8aQWpW9w8BIUKfB3JnluB8JIIQhZckZ46ZqazWXopQ6l40CG4g1D
KqIXXMf4fONpwnFOdMM4zkXLFOZNPsK/1MKLqKjKb+VhHOAir2wcnmt6/LzbtC42
GEDFNqN01O64d5x7O7grtfCYns65jqOs5NiBW9zLYzCWjM1D3SineBPOu5/mGbLG
D55AqzDKDgzOdTGNNV3trN+PaZztBIMJ8AaDszDWdQFojte/4vSR7NTj38rWcxZQ
Qbbxz/xlhvqejnYUGPz0nVB1HfFxuA1IM/DdX3dJGSqeyeiPki8hzmkMDAP2JW5p
Piu3qifoKcZ1oBfjd1wo+Grk2BiX7I0Jf6pf3d3PI5tEyvNSJlsc8lj8nkwcBRyc
hav2BBFjczia9FuKIanCePMn4ZiMTdOmwcA6tbJQrkZ3WofZhAt5o/6W14ZzVE5r
BwLVbrBVDMQes7ihNIYI1G/DgugP0Yie7YpsA4NcSk1KpC+gCEv4at5Zqy5CoQZk
6FJW6BzLTd7GfRiwS8u/Yk4yjpWx32eoCCcQ1dzDeqZxEr9tx/7d1PFgf9hWIa3G
6MpEXr6xA2A7MJoMK6LBwue97ilerhFM1ucJ0LD9S5tJQ6iXPv9dj9+LRBw9edsS
BomLjBaloGFX7gWynB1a467PmsUioszRhuJ8X4dJfJ+XXcOa/1TUFDOlO78fyK98
ap6TkbV5RG63iCKF400UWVLrHmARMinUzOfqXCZcFcQK+tjtPKDLXMSicdhUqYwl
zuNzcfRcsseBWyloLtpYPQpDeB4DyfXNnAxcq5CS4yBklO7HusREHtKZ8TSO9Bki
Qht+/L5x4Ije0suou60pGYtH8ds4OZZmsqx4XD4W7txZ2SdgZ3KCAfDLy0nu4knJ
rmUHksBw7t0AAqMpPwLg8Lhwmz72m0nEZ3z881apUS2ViCkpmQtxQ9uHjNC5CO8G
DPynldlQBBg+z990yD3eR2lJu+IulajLkkgJxx/Kk77lJif6F4/wxpn1U3zEL8S7
vUl/90hTppPLHSJDmrH8+yGhbY/MR4JfeGTMfVXRZ/a+z0Itp8EuYz4wHtfucsJv
18FQavItUlnM0tFYFSnfb9SGDoYlQ1qkmzcKPd5vQp8aBo+CtxJuJ6ToBSjOUmfq
w/ysuBGuSqqkDfY07RpYrV1vyj5luI0TiiTqCi4aoJ10X2kzUVSRGj1AdHRq7E+C
yQlcyTf9Cj5Cgh87ILWRucVkvBZpndy0GZcoFkFrm9oDX+LDVZ93/u5lmakfa8yI
xXRp5pkJvj5et+1l9xKTqoyxb2FdNOY26vAH4k+1soIP6r2Qn6ooSWEVHDV8hnKs
GyXwhFQV/E9t2Zji4KHUfgDbMFAvcMOe8ZgANvDXgiOX87owiu1BwEfzb8kSago4
iw5iPCmgq317ld6Q+PmL2L8PCASNF7fCFzo1mjofcMhjeqx66H1sXem1XFYAMFmt
IUNZ1f4PWjH9sJUMTL2yayMbM3LI3IRgHUVBb5r9t1PZZpvG+3xkiIJ+IoIGsOjy
eo8cq9SHlS61FFNjLXW14Eq5xhc8rD+EHN5cERiY0PJeXa9i/67ufJANYRm5H919
EfowtDeXsq9wL3N4wwGx7kASpKeKesP2F7k/kUsdXOxPWfYgeDRNo0sCGqQnbDMJ
jQbo0KRjXgRAiMjJEanZ4qGuEd7PZZK7+cj8jpQIu0MN9QMC9yGecvBlH2IRAWdr
AgZrTa7WysS8RlFWyphrNXCe72lCOlwN+85im5WeZxqaO84d0/qBqPptGCuoMlgD
dUs2ASci1KIRM5KjHMk7dEcKJcb33IhaupHJqgKTcMFT02XWoFH9nLlahTxUBHoh
JdIsN1tB8iQ9rDPpl3bCsECmbK1bInG7pZ9XFSfyH5/3aFiq2klxEzBF87EA/PEB
cxHOXasR/8/pIFXQz5ZMPO3+vJfxH7Emxr6cfzviwh9/eDHUQ34jnJEC775fbTff
8B3aWYuD6uP0bYMq1Nx3uX3zJEVNQ7PbdqRJD5ScxuoHPO/MDb9TXsZ9SEPHd1st
DXv9w9/MchoqkSEZZ59xheF2DqjvAQ47T5Ru3m/KZIPn5dE+RlRfA4K1g86UNOQT
Qqz9n84tyogfBbmB9M9rBesta3cB/O6r/dphMiCCA6L3pntqJs1KsHYwjBcBZnjD
/0aPBlC728NzqQAchAKQJyxCL6E3yU2Ln9sE4VbWOl2J6U35imh5Se5Z6MPFZ8hc
7zyuR3htHms7R+p5uu0dm3gkloFjgAHMm7Cd9OTSZUHw1o57OAGE9L3IzXXJcRFj
XbNpRalrdnTSWxZvmBZ5Z0dec769Kl8Y6dqrjt9EEfwHDRmTZHlMUBhWPNrMICTR
g7hBR/2lVHjfamG42dq3l+LCk7ZOtUGn2iKtITa4C20pkCY3Wdt1RmVttVi161k8
2BwLjGQNZQCJcNxzRdvOAKvzTblkpLsZlUZMCF2L+tg0Szriz80DOenbbJTur0cK
eMLMpu45g4sIPJlyImQ4ssS7HN1zwzS0uEMgmKbmB1uJ99BsWWorUy+bNm35KO8x
Y+HV1wN1214GeKgvdskbz8Mqc/hxq7cN+S8oxgE7gixxCCd7Y0L6uYLzDtM1f2It
dB+X3BldEr6bAJGf4f1WBpEtjhEUOrnUIlCnkoi5GkFEBGKFh6NWSG9ClKX1g/pn
fTV/s8WS++DbknWWMqLYt31gGHFDA6AG7ftkx7nr5vOGfvFsUlsvfPo3ogIz3SUT
MjHDGTLuJI9smnAx16bCrjnUUFbWwGPweBNxlC6havBWlKon7ZS8dqXI539EmVa6
gtlYtcgAX9rgQCoXO/abJtEzWAEuci6YL7qSv8z6R+uwU4h9fb8zY18sk0aQNbhL
c8znAz5jI2VZktDr3fdGo+x+xYi0DLHFm5A8ZtYIpsVNT3G7SdMC1vavoa9oi3Mv
vpsDns45EUZMwiZCTUMF3HmkZE9uECZ+SRUIhPLBVK5DvO8R32cCG0EiloEV+M7B
W30fQS7wHZQgJ3PieUv0V8HDYs72laL2SVhCvGAlmaO5POpAY96Uhftm7ZsIPUHp
u0tZtEIkqRdEGUCxjmqr7mXrzlHQ4y+WBySui8GPHj04xEyt1GUPAadw3RC9ijjw
bXR3pHL/6droKknKoJyJjcZy7eH6jr8YvYxM2DP6KZZm+cJrp6hIoafn8EPlqiUY
ZpYhgVe28tgpsQff812VF29axP7Dw7H91AqqldriA290qOx/4x5VWD2D2ZP+6apk
dcJ/vcLS54qEDt3PNx2VLce2ombV2Jn5bxfSMq2LPrcTxcMhkoV18LTxjtzttqDT
a5ZRTT8GDSC+nXR0qtsvhlLe98GrlVdn0Hn4TJXt4KDGiGeWuacBqIZK7WSYbs78
tCdYqL/OIrjNXjbnyZEleWTDu3JlKo0AQT8+jcfTvGI2up2eQ/zoCz2HEWOwpkB2
pNxRfmfqEcCjwKGVFZzInrB116gbPB6cJlcI5RflDBe1PMA0d1maoMeOyLd2bpie
oPzZdi4lF3kAHru3frsuVKnKbnvACdB2H0m4XoSsy++sq5jLHVEGhTKSj7ZxrCQM
V86FaPnPSnsDY0d3SkM7pi8JBIzdYtXQxjVltWto51NZwfzB2dXLtman/3wyjA+A
Wv4XKKLuAt/+L/ZNZX6Sl1tNcIMpHSVo3/9+vjQ+Ac+9XqjVUIWsKca0S0FQq+t5
a69zMfzCcRkVoMGdxgbdBortyiZXqcGAGgtpW9YDFB/axkNFkYqYxE+5koO5NbHE
Fxha4sGM60AigdU8f/s1iHl/BjbAmv0M6it5DcCuPgXjwepW7uHNvBhzR9zaesd8
e9JGr8pePgsWmJ9rulehpnQFx+nBRNG5AFNbAtw1MI5Kjh3Sjed+rvYxsv/BG3kj
yqwDaMZqfyqnDs3PN1IB7pA+czMphTQARkHxUnLPyW9Oo7KeX6cNkVQbNc9LH1uX
h9wXv3k+pH+pnozufGwVGTeygktckBqOgt7PVlsV+HoqQkS54KpOgE58Xzf47cqC
ME6Y3jzSiV+7pgmxSnezb3pGDPdg96SPdh/ST9vbxKY49HPVIoPnXZiFQKmW48E8
3y0OKTyATnOCwUxFFfIzl84j3t5PkzVC7o+oxCReieUGV9p5GPA/uWsydkV38H3r
zpm3ra6EBr6R9HG7Wv4gEM4JB+oGQYS2aAlnLQeniBBAWTc+0VfJXa589yt9EGJq
D1g22aSPNbPvEKKQJ889Mug7nfzuqrM42YV7fAmps4LMHfAeMYlUPXMyoGIhR5xl
pV9KZbWmmHa+HIf37DDs4gH5haggwHd+QqKM2XkYeGtDe3Jxl1HTSpf+K3lnrX/f
gct1iT2qzb4grTOox4mfnWLeVlNfcVk7K78ZdTDhwZhmGf2va12fa/YUZkCgIhl7
v1OxwU2GreEoAZUpJPCSjTIDiHFn2ogxnZn89fH5cSZD8Rh1L4InW/X64ZeIiL38
aRSgsrx+Un7h/J4tq9Aa28Cq6MZ7C+FvNZ+caKtS2ZA2jMHouIpfGlL55M8X8scE
rZy4LgTYATWZCsaVABM/S8r922FFatH6dtWK85vz7bs2cOCipmwASKrl4jCe1HZD
UBNr9cmyYgI6f9OOEfbERIxMmG/Pc6MdEwgJ25VyWZZ3FsjuldWRqcwjJUw/TKMn
V+362vvGn+SwVzZQUAw66ASivmHvESBx5YyBlFYihwaXWN98HKzCPi+H9MMHAUtM
r2ySuhMBfthQiila83JYnftakOLQJL4vRqJMghFaUCnk2iwkaSClpLPXoXMdpS+R
FQJm90vBPRYHjV9MW826JHXpY0BQQnfhG1uJFklBZewo3c6b2f58PwfycJ/mSiFF
tv4NYXKSL42ffQP5cmGN2EjMwO091TOz3co/Ri4JIUmA/7m5a2EueI6YLnJurPyW
qx0e/qjwVs3agNUxoj8KR+dgIcKNA/CuD7a8kay6c1Byta49AnfyRU7/KKvgqLap
52rnRpabIphf44G/5EQ5tpFQRGE2Rm7wDbADaUe74yoMf1zl8t4I3xtovlMB3ORX
GvNXAt/5SwDAfRdlXz9Jrgzow7Dm5dktU1X1okSQTEuNl+K0M/bib+DqvWuS+L8N
lwp4FN54F8LwOXnPM0zm8E9gorU3AYnUTNBmtMgoubALQeCus5mA6Xb9ZL8bfh/V
5yS5SZsIQ1z7H7ntDv3TAIXr031Vrs8hXwgs08wS7DZv+O8XeS3DieST2lxuCHdd
sizXPExu4qPhFZBfK8gm1JlaWbKRrGFrGZEpbyua3sQtx3EOuGkekP2661tr8yqY
LGbVRs7iQDEFprKeGq6bA1oJO0qvymXoly0joe6QkaejPruqnBd+OXYo5LV2EUdf
3ur0fS8dnpzj8RQcNubbN6z1by6XhPJXmDK7QwMgZnlZFbCog8gnA2qDgrXfUaJv
N4kjFE+/1qB8uMPJ/kfggAelQ66I3I7K9XyyJc2VZSwG7rGlWPSTpYO3pDTVgS5F
2ebRRiZDjlmi5VLm91uxoi4flZwNPEXcoYyLdC+PhFVXgSvm6lh7YvpISZ2YLLEc
ISJOfarzhCEvdkU9JNA15VtZC8Sm1eWWqDHmfX1hxyDxgDkuZfL7cC1ArFQNNr90
gnlPoaVf/DHww6r0TVHrkFTW722dKxqVOMrZtPxsVGnNvRzbWZ4GNqukePa+RYKV
tCeuIVimY0bM0LcANAefB2NnSRbdtfHUkJqVb5VXoROvHMHaN5jHOI8evhcdc+me
CM7rRdMPoLISFqIpLh3lZyH6FSzR/ONp5esE2KUeS8GRFJE3HBf9YWdNC0oZWDBj
HPjmlsv0rTACcsSDzD/Tmcv31YgL2uU4BRDstMh73hPNv4dBf22Yq4y/yNfHLgfe
Ilngz/8TRHBXcxOE4owLLf/KUYYRvM6N60SZiWHBGnySMD1Y0Bgp2oLK/Uj684y+
fawox2Ppf2hyp+V2ybNoLovv1E0n8svo76dgzUX3vIMNv0F2ECBV85WwCV3MNfcp
dZJIojBhi0zqBDdfvJWgJXXu0cnt+dSKSj0nYLmNMcipsyppgid3IGYv0VIaVFTM
iVaG6ZmLPsK92rlxjjqMA8WfZszt6Oq/fNiGnf3ASo0pt71G4Pr0ZPn8knCWEZJS
nfrZDgol7dcihpXmL04y6WUphVekqHWoOeJE5WUjhqqsyzvsw4Vka70XsTdnb+R3
5laDc75h9KCAVAmyBNxFFOJ8S1aMObmGVhB605oxFEbcAGqXMF3q7Xrek8eRgcqw
T2kmizWvSVo4k6+bIulUZnNbOZpWfqTArOcPrmttdQqpd8MJyl8VE4s1VlzlpmV6
88lAaWoMwJe28h3x+cXryK46kjVyoyTejZNWDcWT9ntXkJ9XUEZgyIiZqsWHJoJq
sFBr/eW1iSkTLj3w3lRcXIFCi2af+Swy1eC82dIbU5zYtLW8eCB94ll/mw80zbJ+
ym7/s4ya3zoNF4q6owDzOGDMkhB1M29uOODdIRfhG6atRS6ww7nd+VXCJVSsERlq
+TB/0vEb9LQnI0b/yqfvgZAPN6qCTOqAbh76RQCYAiKv9ISkXMyin1HyiQB05IR+
Qqgv3PbSgc4nwX2sXMePJziqjX693Juhov0Vt12SGA+73C3U2JFirE5+0qMVvH3Y
rESZ/OtA8zhjvKMCK1JJ6Pp1Xb1lyn2VRzqWJGqe4ixO45PkSZQ3q5wdLOezT5Cj
5ZUD6OnolegOhx5bOXsKVMfvu3dyvH+KwdEegheo3lbPVDmoQRkHxv/oFkvGOUUZ
gWy+PkZL35BH74gKPhYYNRKgmJZvpH+VC9s8a+MX2PYEX7pwuMrIsFmmtpIpjHAs
HrRjK/C/SCgKbDSwTnH9qGl8dAoYWUroYmVHsqAmQvZ6MLVM/YxsuKwRGzenVEO8
LWRmxkkzFZjvNbyqvJAWszeGPuzQN29jBKUvHVrtKGE5ZbyUj06UwB+mxr2SYR+K
iLGJz/ai5I89g6TqGkfrMoq+xMSmw0B6UiSyr0jsHUIDnOJuIgcbDClK9whl5Yuh
zXUINZr5pyIaSAJqHRoDkAi3xMBjCZyrxACkINXj+aiRReg61/jPMbMOa/GbppJS
G7EswGFnzKQm5Ku/Gcae55dzflbSXvqODOSl7RhlZHNvInZnss/2YVUCOq2v1Xae
Ckjr+H+5iU/OIc0trmOsYozcOFYpgWsqNeLGbkIQMYXgc4ZbJ84eyOtDjmdearWy
/XfqzdslM8Gk45l50tsd2wc3RUFiRohRpwAm42wuuG2YsaKYvG6xQfXjiHvHNuOE
vc1np9KN4XAokJpLdIxeVVPiymOWyzOiGfXspMk0l5xg2YDaCjtU5AMaApoiBKEL
7vr/Yib8KyMREPA6eAqg149qauTgwmvOSTjfuf+4oRlxif4DXt5hkAJKWQfKKMKt
fPRszxuGvBPrb3MJaQnZArFGHoO5frPtpEyUXGWCE0Wgodh+AGwg2QIJnfENrHW4
BKA58j5TGkTMywAchFGNgDb5SGgzREsK43lM43kW4kibrlQZ745yesuZAu+OnQOD
XTwGN1cEfKyatchbgej0vLvTl3epK1ms6Sbr63M7OH01ZjITdYI0uk8rad32TcyO
V26DJXgkpt0L3Gm0i8waupsRRH7ewaKEFbCDis5t9w4HFe2Lj0tUmq+BUp2lBHFP
VSSEukWQ7tBK9c5CuXfRp3pTwkJVYm9/MdiiicMRWYyn4gcz5o0OrATp5Ud1dTn3
YrcEcxFVssFHGXF+HBkzDnIxPgztIT3Qs85/XOI1t1M4xz8AsFETFmRoDMucgIh3
4mk057C0F5i5k40yp9ix/TGwTxUFJi2jZuUYOV04crZSN9WhH1nMxdPMSx4Jr32K
zf8ntXNVHkqup8coGi/OchQWJbQHbfh91IHqDcVuvcs6X1bESXRprjAR1CJYqycz
mdNGW+X4LKSgURlxURdG8dfJXxRYdmcF+uwUzWY/DK6tCOsvNQW2wOjthN2sVNJE
5kcnhjxJBPuJOU5A5Zx/4sGW6XQGYaaJ0eClYDKr4JOenIehKWmEce2q3ZkyeEXA
OVI5oMcQV9jhDPeMWPTxb/iBzQeBgzRkmezUKtC/gyx9emFFqTGzjCQ++FzhnlwL
NSFSLKFb8JhCcc9dzsWH6DiIq2RkhR5b7rcpjekxnyHgfzM9+Mk596mP2vR+VqHD
/Q5QNDWOmfM/cfXnUB96z4WwuyWItv2wN9PGoRFtbO+c3FQ2TmJAs6RgM95b13OF
c7uuo+/SeZfRJaii2OmEh3NvDbaw6L+aN+SXCkHNYgg2u20m4cCcsuTlcy5WGIqU
VSCKKjXKgOmZf8ywAa60iRv5kAR3iL5b0wBSaVNpUoROvD6gaZBZQFHyq0532xo+
lQaqh56V0csoK2oQ46nlNASuuOmF/4SoIaA2pseGosGhPNgoarWqyLTUDyBxV4DC
JPdAdRHxiNs/i/TWmJ7Gbr+8HLI/nYd8pJBGt0dEJQUsE12ZYOd79luOH0IGZo2e
t2R0nmOGoSJoRc1WSsijVpwtV9bZETMwpOxjcZ2BCgFNep1YuSCwzn2oQ9FCIOVA
4QcigO3erTIxfFx6mWBEsoT3VRQhOFOOWELr4ChnuR1ar+FOwjfi9DYtFVaJJmLZ
k1M6uUfiGtvy9XhTmjWyMjFCT//cQInndUoIg6XVCGD1NWZ6oFlXNleXTuzfLUh0
AGt8KtDK6gcbsC1rFXtKiiQRnOMeFGKQHL10kadliYQqAUqmR4RGgqD5/bNddxYd
dwQQImgx7rDDeyYGfvhCPDIUAnqaDTQhLKhImbKk4bq5ngcjkTbB/gi4/WLD7Lj3
bH5jCetD+LnCMnUKEsS2jeyd5pTzhXSoMB2+s9V8uLFOK4JqRKo7iwCZEV+IakEJ
x/WiGEI2z1KFaIoZdHBiXStRM9Q+ZV81uyySTQ5tE+T1r99H6VO8DgiDAHoUoRb2
vHqE6xLKDMU0PXvMH0f+Rr/zVa39h0lk3FnYVDTiph0hT4Ix/HT1zztc/SBADtgY
8z1Ui6KPbCpH8ni4C611K+D6k/spj9i7Mfbz1zIrBrBSLw4RUnDmIXI3rU9KlmzI
CU2Npb1oj0uMT8gAtBDRlAOS6BzvuGgP4bVqswQTfeuXjxWbFQlJcY8fMvB7GPws
NqAXKGCSACyfWATqUqMXsvdPd5zyrJKtipT6tSA/X1zhKukAA8uyTr2qzaltzeq0
afRXaMR8pYw7e6ZdwaiMx/mKB2/rhB66d13Hc2P9EJiGtlB2QrFByu0RGq31xW3o
GB2Uiy7OdJhNTwArYPKw+Eal5jDqOYsCtguMZWyClN96XvNoxOC2sQ0TpgNw+Yck
7HubMW0qgOWfPTMyKRYOZZVtcqHTKQ0ooKxHDyVBlyakLGseRRjw1M1pvqj9Vav/
O9Mno2ugqugGWuXO8k/wIICJqUXzx4Y7ApEV0yvqFlxBvFIHFpbpRoL9YlclXr+6
8CysdsJx2DKG1HITyUkNhRKc30UpIVFbXaupWYMsl7MChLSKPWcwiEMgV8jpCHxF
IAWynVA8DZD9DsZTTUIImpEdkAe/rBmllJUdhWWG6Rs3IgxAn6I1r8w7pmCXapJF
nFdVE4+JGcKN7RfJOIhjGK2JGOlpLwlw7TKpP8ekJb/NoieQBhLghVwVZ6ehaaua
4UFPuB90B0y0DSrHGIkkyDRlzjXdEjDXUTay5YMUnPz4AMHW7umnpfw69sMiRXeA
8pDKv8bO/P4DyDGzmmWNZW4FvuhfdiFf1HWE/hI1OCmLUotRcXebAFAdhoxFrsib
o7mqe4E9SLFB8xpK0dLRXRfmG7USMaKfAVCLi1fD7NnPVTZf0T9oWFdoVwY1EJZJ
Ifm4gyr8FLFxa/MavN6ulJs2PymtWSrKfgaK0/i0ETqMsvyR0cwewHbsTGAxX69O
oI6bdQ8uQSrOhBytMa5H/22cg5vomS195bLkVa8gMnYb7e/boUHXeDXtzbqPNx90
4WgMWqcFgZjKVh+56Ei+zdAlzNNKuAbr6BCRsugfq0JgMdzNEqX/aADEXpOiDXPT
n3KIg/k7wwkoKBU6BSSd8qnQ2cyuxaTvFF8Jxb2Mev7bgM7vJ7pCbV7ewIOGdPNb
L1EnQBCBSmMo0K6GARNCwdZj4D65FiDaj/IO7UD4zBLYK2Nh+umqFSn91G2VBAQb
rHWMB1vpwW2Ew3V+Pv3mWCI+6xL+Jw7qrkTEnWffMFPcF76tDM2MKZ4uSd4REWlU
X38KkRskxZKM+4gnZ4Ooq6jOEwH2+SJf4Dg2k4tNwV9keCQ4V0EdNIIFn/eEvGUs
0GiiI2f8qCB8Bcyr84Xm8gBZ+pSCauFCPwm9O87DzanhxCUh7sPsBug0oKWhEx4g
QeOrGep9BH9w+JTgA9nkvkqqL/BG+5ChcfCCZ0Qcp8UE/w1pc8gPnDWhj94hRypU
Dt4FN9FrgHe85sMT9UWoBxMWJmF4/HrA2qEw8gTCBByFkxFzIiNMtHbXCJfzbo+s
eT/7uF1S0a6k8HQcItG8CfNRyNC57jN9eVyhBUDIxdqKeGQ4MjWloa7j1JFWYypP
TZCNWmdWe0ZcX5hLcObiovAya2zcQqFTRCRz8CbtLpfE1vZ9uIw+hyBUJvYqXcoU
BnG8+mha9gTW1j2mJofR7mkKbiaVyb0mlnQ6qEAytfFSwuaR0qWWdb2crnJNGnaU
aTkBdx4Q+m2UJCsc1SSqqltV3wS/RnqY8WqpxO3SrKF/5AOKf6Q3/wmJ50g0UGKb
9DftGd0fYRRfwkQMEtpAfz5gQIl5vKtwqHL/nHbYbuffj/2QiPPdo7T68yuy3qdb
K5yDiIX1XTDIrx1Sa+YjjzvgRHvHFuPsDqycXiVAXn0FV6p+dBGIzK+ejIMVmSII
WJ1u6AAX/fsXMkReO59O/zTT6yoxBOi3vvcUzxT6rI1wvnMUC44s1FUNu+vZqxVY
w+eYd7vm04uK4UvS7h6d7zwySHhC1zemR6c81VeGmDQM3YD9rFpxXHFZDLiqoDWf
Viizivq/GyJ4+ZgFCZsIr0+M/ViBglsZWUzMsGCyJajKPqprmThAs9yrp1VXRahm
/KZxUbQpkTM8HsAM44i1XEDy2CXn2trJ3uDWzF1EuGas1ZAppAJFdrwy/XTcI3jr
8qZhP5BZ2p+M2wPyELJNa2N3+F/NzX+aG76WlfO+3WE3SdWpeSe5ghV53Q55wlgf
lAR50TL2ZqbsPOz4zGgCJrHu0Pze+Zt8EMrF5hDM7KykVaoAlShk++1ObH1NqFDH
TeMJi9R7Rgaz3UjI6Ku7Gg==
`pragma protect end_protected

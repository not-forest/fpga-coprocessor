// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
GzYtkvUYPQ4nAL87BaiwqLY1dYGFuJ11ZfaH9xq0S0p4iyTfTPl6Q4l5VCbL1cyKCt2MkFePtkPu
SybPKipgliZPnSlsYXk1PDBrLVMaQdmY4BcbtWBGPzhLKW86OHeH/DuFOY23npKCvA8z/fyK+Cwg
oNzQR15oiLU6XTaaZagZpe2TGgsXX+tnpCGDNkqF2w/HbGrxtdfUDhjVxY3u3eOU2QtG+ESLvHKW
B2SJ6ox/I6C18TcbIovyJEF5RB88oVWYLVgVO2tPbJqlSuTmEvQ9rsL2CMZkncHL9yNANucFwVzn
ACZxn/agqAvNB++ZylYx3tlA9Oq2lWaTZI3lJg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 4976)
p1qJ8ybn9nKU0aYPj91GmoXx1q3GZOQjzqgDcrD3J+ZQPDg0Kqm/wQ8yHVdRE5guhwiY1kwSeaEI
F+fwzmbCphojRnblARYkjJA9IxpuZq7A17nL2TCqNXBIE0GXZme1hf3YT/Gff6eEnXDVbBZ/krLC
wjluasUYpBfyRRRKGPxbbUo/d/B6GbFWfMvRcyKiyPz9gBHX3oTrJ2HkiJ2/+1oQsBSYJLral+jO
h6cmYTHv6rHYLakeNWWCxoaSodNhhxYFSzhMfiox2WrNVGhQ/3AFTSsA7Wc40Qe/UjekvaDjAC2i
T4hbLJl6vl7zRJFl0M3LW2k1hO4NL2rangQfOkSJOw7InWTu7RZ90yL2GvG32NXJlW4ucxoNoAGE
xlzF/3zkJ1cBWxsF1tJf89rpbB2wN3h1nWC3DAVuHJ7g5QFVjJtazthWVrPx+JgH10MR1/m/LmoL
NNfpEjkxUIbG4kEnqiO6UerCn2SbueIzarNlwutj2WOBfd7KJ1SS1Zqs5TwDcuHGXJNjuY2QR4ky
XaH8uIrSEdqCrHuhtCgTl/5d0PFwBeWf9Hgp9AzxI4PjLDrCGELY2huwO4BM1zFNRtAnmXDBEzhZ
wU56m9WYtHLLcVRhjH7VVmWNrB3aQV4wlCoa3qQKs2sozy1aNs+rz2WNKWjl26YOH0mCxUXCSutf
8Lhy8RxKDfm6GAjouVqTiPL01v3yWUeeoFkZUk7YQoXOnkN9y6dN6u9xmoxChtp7dx4F1M0Fe97l
mSB/5ThcPAaJL3vHzR8Yqg/VVfO8tY5TCVMFj/nUy0OhkqOgsp0wdk2TPDgrI/tOZso0q3QIjoSU
nCq7MO3UJQvmTxPKh/YFF3Utuo3PYduqe928JENZNfJEPYScyMhNbFE1Mif1IrU3DFKdmoE+pFQm
4xKwW41h8HuuhKO2yIBmSLdffex60asz+1WTEo/JMmSE703zwCyG3O/NBU87BnA/UtDqJX2BrQkG
iiLbZLqxvbRZ9arvMKEzdu0iaCBc4bd/y7xdLakEDT9VLCoNNeBjlE1sfDE9eoNZy7n6XaGgbWmD
0JCGzs4vIFyDFtr8FklCSpWcGpOF17swgZpba0RLUw6sb1kai8m3C2mbzLCq2Tyos1ej0IFvd4S4
8MnuUvdgs3hcgNwzHFRTTk3N8+14io+nI2cd8bUBQx0D2/72EbnpbJ6s/i63kKSg+VagmJgFTlbX
wRyTmiiDOvN0Dnxnz6PPPpcOXODbSuxmpxEWmd9uwG6VIMeYiuTvh4JJRlbOK8ELJZnHOiS+ALsr
rRMC7voJ/pO1y1QELqgY5wp6Tb6guWGGJJOEsDnaybFeKsocpGKrSQsK2zcKKkVRUhoAImdQNAyt
cNX68wlK4q6WLj4V3eKg5FEVuCvbLk6dFRtejJ6RjRC3DxJ/FlG2BaRR3AYtDX2PisyTkw0jN8WX
g6DNf+eUr0f+FxJCXx5q9LZGe9dt4OwHu0nExjkpDf08wi/D2JQUyi48D3uhgbn9N25OlWDvBUyU
RgZcrsmE/M9VqJWJr3qXo3TOPSf0AYDMJnElO9S5DFlVjBiUOUYEXahA/V1VUkcdmH6pzFyZqmg0
msLIRPbW4PhGSWUgpGq9QyUbnrI/C++9j3SUCYz9WNW/8nPvMxgYrYV6WqAuNukXPRAYRY4z8nuM
RMQN7oH6/J+EI946S0icKJFO0QQZWqPVtEOAEpoo8AV7Lz1TcvJOuvg6350+xSLBdtjcpbgDGID9
nHP79MjcLScUuHZqHKkI5eg1bjh97m0Yl/0K4tSUKgquQfkG4wTzhxcMV3yH7pupKN8bLvgvyemM
R+tmIcataLs9hJQcmOOzrQJnm8tpp9EUqbQClNvebBVx5TjUcIeLwWedDxXUs6COazmu/csNWT28
mgTcnUMbDmLAlhX0UjGNYiPJXOqDdoHB1xOYpTEiA42yZo9ZRjZjvZi8ozUBVkluKhxg0GAVgJ9D
01Bs1+4nSfX9dpR1GmoMB0fBePpEDVyKlcWr4IycVAAj24Dr6mMDjRcCYvcWeL/jwr0dOJKOnO8a
kiQjmDE95lHYplKky0dP0qv2VXiADJu7FNM2LhiMq8P98ybIQJvGbl3K+jdxFvXG6RAmmaSEobRm
1Mzd4G765nu9i7bgraXYLRAwK2/MU3KsPvWpKrIEw0qed5SWZttucPPlhz42fzfzOu96aeA4BKpF
9ksQQnQ0OQ61Jd16W6jXdg/l5uM68+XsagcBJfkJlKfq7WWwf47BXzaniBzGhayVQLm+NuwPq0cw
UhWLm11A7EgWOEMw3Z8sYdD06Kgk6l9pcRyQPWe7ktv6+G91HvjDiL9OQDIIT+HSGUd7hxHrMAV9
Cf/3Vl3Aq9aYUhzgaQUYzLDKXh5EL8Poduy0ryV6T++Y+AjXGZyrNYyDIi9Z4wtDjS1HX5DCUstl
qMijWLfC+hD04PQv0LhIrfBkPLuXDtJcw3czAdOBsxUfcHSvIR/gBv63X0IY0ttlnA9Bb5W4aXas
3Si4zTCvnlh7BdEJsaJw4JPTKbujwRwtO4A6PozuyaEyTW95RcZ1IzVkX1prWS2dHVX/OKVSdJRn
XfGW11rWKnKsINhwMMySMdG14RgOmP33jWiZ83ay7k3HThtyTaKFd02xlMKzAmgi4wR9QSoRuDBK
8Szp9p1rVUn1AzvpSDVBlC6cVPyO5f/Tyh8et0o22HWAuxQxBb6MKIJdTN0HZPI7AVtfgqvxSc4X
ls1qSmkKAT6mfQ434TwDD+PWQaey3Anabi680uD67QB6Zpn1bLNsVqodHtIprQDUkMcYKrg0NaAc
X14RgShzaAXWZdQ3AIW7amhCcyjA5LGLVqjA8MsDn+P3l6W/KsOUvCul/QG8kM73p+/QB1tfdKd1
7e41EjteVKju7xRXRadjLJdXFai0K9Z1duWN86KJNcj354MiJn0sNLtrzCMv/sf8zMYT5LfvvPRN
JWmH+6RKiPcylOd62EU1zNivOX2MI/c+Ix/+htQtibiAWI/wPAe087s4qClZ4vlm92kljAjByMX5
ss4BdQDKF2vo1XB4Er7IqtNr1Jf/6dxYDUSuStGP2XC4GKuh34n7S9UFFQPZYpEZaGVOLTEsr4hk
DN6anTheYRAbqSTUlafWsLi27Siz4IB6ah4k0H6n7zjlQJ0RKSw1DZQFoILou86fsm0AwF2CwNst
m75AJnUct/HQ3BCKfnxVnsElSNPPEUNwwrVCDCZSmxkjO5GCLd1Koi27M3gkLIVeVTzEKFOTdj17
2drmOGLZCbcCKOWTO3+HgmHDm8lRoMVG/AFk/4HLxegBj3MIqwG01L6NaYp1aFaZqh8d0lFb/Co+
rqm3XBHEX1FdR8I94bhzLG3ioBpgqPaGLW6+TjYWq3+9rO+Z6FTM4+UfcKtmn3GvIzII861ItoWX
QBbw3v/4/m2mzqN9z1ChXD90Qzm/cECVyMUR6bZe2bSPwd43rpLZwlqSNB6/0ntK2KlF9aGShUBE
z02TD3aVDNd8pJnX2t2RVuzHiDNYMu8xQnX1Olodcfc+qGHtfUKL8wIzauyx9t1dJvAugqRPdRXz
H2J2fE8biE3an9pgyeHLeiSBXZKwbNE2c8t04v0ZOpSIR48MibWM0N68hghhI+OLBM8nEcJHTDY0
YktXo+n+acypZyaY4se3epxLdNCXOZDuVG0OyNp43HG7x4UprogyJK9CqkEAm4AAYw68qxJMk1/q
mw6GyYQRZ4dAVl6yalZzHja+SSv6Ej7RvQazXwwxxPBOCdxEGQHWD7e0ZyCM8PYA9KeQCdmxZ3L9
rEZTThHqOOb3dC7iMYYpH6KWPqj1kyq8eznsAxadrF0O006vSRdKkPTB6pjgpuIHcaK/Ce/Y0I8f
lQJGS5IxAjWoFkTLQBWdrp3Nd0Zz3qDdlGMd5ho3B4sRyXebjqbiXFyDlrCBXwmsRs56Zabm8Boi
ZMbtNrn6UxK3fy2Sff3EY9NXPn17jrcThagzscWso+6TAl54YtyLJ9lIekj/Jr8ZdIQP0duxHCbA
i51952S6qRNg6/G9oFNOBLjmtbCodRxy4KNpy/LC/YBDeB4XtvqFcfbpxNlS4WbH79Y1oor0fXDy
avyIaWTVVBToNx6oc55We0NKtA/fO4xcomFu5EHp2FKJpfIAW/PhvdExvT9dos9JHDSwUEdmblUY
RUI0v1zKu0/HV+MWlmjqqI2JW5KRxPks+Pnd207iYHggVBWkTgPrdD2IwWitRvIrJxRmFsEG5zso
TobgRHeEVyz6Go6kyhFpD6JPCx8DslS74Jx5DS60SYjA7PK0uzMLy3SnUZw6BcA/LaZPxnbYqkgO
/0H0H/bUGh547nNkoBpUb6fKATU/dfAuBaPpm7mKf9BYZ8UCI2KqvX077KnXhaVmD17ZUq32qtrA
HDn5MdISN8CUe2yYIomA+bwxD3y00NqviijYxyyAj803b/l0C2NDTsuoL/0DALP/YGaiUkI/lt69
LB5C6amMniNEweesqb0pf0Nl4ZFt1z2ZxuyQPIPxm7jAGTBnK3gPi/OrkB5XHuYi8Nk4P+eyx7dY
PzooYaHl8giWkuCwu9NVp5o3tYrAvb9eZVTjDBTSQq7AUBn8zFO1MkrGPnPEqgVqSF+t5+9et+TC
X39g1HwOlYKsG2SGL+kTIhxBIwxPpujdZqn1UH3TPRJFMzEzl9Ml3WvV96TSSUCIaJWdiUkQxvsi
GPyLXRZulwMsrb8UDIVJilWqVho+aeiT10uIP5Z4Wm+urlXK1BjI3NY7lwCbtDLxbqYI6E0Gp+e4
QxdTD4qG7HvJcPH7rA1Uy9M1HGGTvenSJ3y+k3w1jA4n1jrarx1/R6tka8Bn3BraBI6ZFXfZmSo8
LN/L/SAj12lBT4c/XQy8sctyEK7nojuVlQEHyrjTkToZ2QGbqCDyNE21ISpVmpVLtX0Jzagw9DX0
1Vb1DiZ1d4OCEbpOHGbVooqbnc3SxpMCNBMKWjJlDtBmxlyEsl5BJ5z39/+tteMw8wDt5jDY3UQN
b5Jqv215ru69ryD2kKXWtCID2AqKP4/tV+8lQP50+ugMkIzPPuRv4T8Zbs2uZwqYHbJERhEcMd2k
cy4gEXfswVkgvBVvxi+vnLOaHwNbc1buWu6ZQPNaX6ENhzmvedGE29m3kZ/EbaBoiq3q+ULEYpNI
ObJYOLFsBDcPs5+cMO4mcYmJES2pkSFTZvYh7LDahKwK0v/egPJPP/MisWTE93BBIbrcB2nRSncX
k1wvsdITtzHTN2fbHfPUR7towzCywb1AhjcQCwBIyLNpjnZwMlMz/fEqwK+fNrTZ/4N6goyISo0M
7+R2yHfgmuCbZEPupqEegVNCz1vroXabBH/oKweg6/ZlTKDzblyjF2Pn8TapsElJPSbKm09ttb+3
vQ9lnJDgg9fsmA1Ff7O/6EY38JvFcsxDKeC+GVZD3cRK3S88BU2kvNbsnqNp//sd5mj1T7fEQvZJ
dSbAxlFkmNfFjJXGw4i17Sm1Yc5HperV7jfMGE/psh2MqtPWE1xLflMnTIRv4r7XIg3xChCGC/Pf
YQjbg7iX3Zt2GtR8xH0BElyexwxuG8LV41rVZJcoTwavpFEO8aiHb//AkdkYWruJuhbNGRbdzPPN
rrkO0+Pu6h/rqQGy5pYj63YvmUxdT/V2L93YsSCHiL5bnOizWY3YBtpZB1kPxKkM0mwewvHPneUl
G9fPFvFeOa7Jtzx3cmy8DxCbpcnSMp/GiDMrnWVlhuB5MDyqKw8NEhDslYL+vFc2uPdrRq1UBml0
npFdKCK/a8KbWyRBObRv1V+wlIzga+6Sd01RUmDjPuW1TaY0+vUS6PVMl5739xAqfOvHuYBIhb2O
I0mro+tktY/IW8MJh1R/20qrKHBtCu6Ye3aMa6CkjJPQ1B2jkv9lZ8o9boVwwmHxjPNyRMOZUh9t
JlozRcGadkHdBk9Oavs9PDD3Sbpa5skzlLwViy+gfVFyl535puz1GtgsnM6ndMgiljyDUrnyelSF
61nyB0wgrnXSPfS5ZbesNGRP/Ia4pgQRKmTi1zFvDYg4s0YFLHEyDSs5zZa6y5nYwQdX5N5SU2vn
PeKOViEI8ASEKj0ClDLcPM7HIi7LAsLugZQ2pC/GH9+OCEBwcgNloSalBDFGBGtXaktHPzpn1wdP
3p2pxigSd97WF6N31li48Yl7vrvrvkghU6s9o0rYG2hzndZsyXrvHP/HGX1n7mRs0X+vwiUfAmG+
UNs0+iEbH7bNj4ikGDItNmdWJXArxverTNBw/xDzyDrkHMm+IEHjmo3UM+m9itgyUqu8w5+TjtJs
uPO6clH7NPVyB7e/iVLXYY71CtNVUPhIIwrLgF5+EpLn8S8KQ6jIVkYda3PfshYLB7xFWXeL2yJH
s3VzFocoltumfhmPS8iwF27KBZDhMnf7Io9NOce/VdV+NqxXuxHjYwDltOnwBEA0qtmZIB7+l/8H
wIpGucz3rIpf01CdEVdU2CX3mYGoLFxWswNX0zS2h6yQ0ZNzlvSv5F/1RgZJnmOrM1eb2hKjWUG/
g8jikGTl6McQbvDdghXZ0iyaX9BGbr0nGRkkWVwSSDoN2AKZzDzpwzFN6LB28tgdWds3rvV9PzB8
uN9PID3X0dW8EQAs/NyOdUU=
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
hSYr2QqRUzojIFzqFTHBOEOAD1FM06b9+Xq3jr1fQI6QTrS0Zppq2vwbzXgNwBJZ
cViEQzZEUEB8cNpNyVjVDvmujnDu7juWsaJVsc2M3cmneoBTyRLewxGX4vubxqx6
lA+aiFf7SpHvnq8Ak9yyNR+x5TiFGf/mpa/8r3zNPle3VHhaRdDBdNaCH6kIourQ
qZOEM3U27cpEUM8U9OPAUw/o3yW5r7pbhUicrWDfvtrJXlqu74AAF/hXGzTa2Ii1
C0t84reqxK84L5aBH/j98/45QPRB3XSojZgUNo8l3n1KZHDBgODOznxz1ZvlyzYh
rXisLBpqMAavqYJtgAgEoQ==
//pragma protect end_key_block
//pragma protect digest_block
rAcrDkyr/iThjiUBki7jYGU40Ek=
//pragma protect end_digest_block
//pragma protect data_block
4fJdXElXFlgDWxSQ4f9UDpvHIO/3N62eHtWbu7xilNg07IKbFLPDNtGoFhqMpMkb
S+VD3qJzVqfMqRxUTVxwpuCt+ZyvUui09rXtIoO7bD2OLRkMOaadTNtL6QxJQ7kE
4poYHt1tOILC5GgU7ZuWR+ZitvqyYjgx1qRX92fleYckkrWcgKuSEukmGNtSxLkl
IbG/ztzebEIVeTa2iRAoTsEiGOjztQP67gYKvXu97CrZQc1cB0gKkmaFpyyFea0T
D7kLiPHCE8WBXHcyKQ3ErYurZAyMxsTakean1fkVal+qg9zPIkUxG/WvneCkUI6S
tDBTaVXrlub1Bbq4p3tavN1XOfNtYuwJYqkBR40HcP4dWXv3NbIjNx5rZC11mBRR
sGLdEpgMZfNc5q8vThlJWlGM36oS0CARBEu8BBiNhZo9jdqGwf94dk+vodCyksAZ
enGXli6LWvjSrNYudgbZOxrX6AFu5m6HfHGc8rvH9W6qwz30sRE4epGAT+OTBRKj
onYcYLyD73eBs5rS9gbKPFF6fe7kSE+YQWxJJjtX+SfZRsD47TU8rpFhdu1zIbjl
lmYwG83HvBwRoP8JKX1+C4UAQvnLwXLeTlAyQ7EhoX/ZMleL/EoVmZUd0RciPxZ0
NW8Ys4mUgslxKnreD7BL3xJXXKe7vcYo/AIt44bUzVmfv3w13OYPKBO0OAnZ+xTv
ktxf9Lqhw/mowKnFYFTqSv2ZL0MkgXv/UpYYH8rAoP88z+uImXld2xY6GS7YYyz5
Nm/DjR5SlsSLQGCzmS5WZm5iKItDOXuyV3Hbb1ghsVgE1g8eEBnLRLhxpay8+0V4
9G2ZxEagXZr6rJIerbuKeyBZB+X7m/JtFPwmIzg1Qj1Xf5stA183DYRWtv0GVgjf
u4shb7rGReuiqp3zDNkKCTNSAmf69dvOaOH8VR01e1RQ5C+r7hVpes43YBilhOZy
t76Q+ySLdZN1W4uzl0FGMEtXaCiquUup3c0DMV30oFEEkviEcjOOn7VUKkyf7qyp
bX0HkIBpTVb6eC+eKR4fdXLcugqZtmBkamLnzl+KVpq3024tdKAUKI84dhu7rbYg
8EarhniOp4tYroizT12NutpRk2n9KSRNKghWjYC/k2ma0Bucetq9BfRiqOK6hxBt
7/vzBFeOIY0bTy+VZj4cI3h3aYfKmDrLqwoOQHwTvr8Cxp5zHSahtq3hSGBDZT+i
bK6e0KV8xZev6+klD5/axEw2vL8mWFYnYlSGyAYmSMWlQr4tnBi+od4FbxfVXVVi
uhCZEvqSCQKIKdUJS2SGA1Y4yiopK7l+Vx+kb/34jgwBcN6tLpHqn0RrVd7Pe7CF
d9BoS3pKXhFjraDNCsyKaqnPNQN88vXcYQl1Mzkq4kuK8+pfjoUCbPLAto/gy7dB
y1QDZU3miflHKxD1rDEZ2pxfp8m47w9ncuESukQ3cD88HC2+r2WFIz4x4Xps6pSs
+hfdFDJgI8TrBrIXNlNvKIf7v4ZoscPlK7rpc7GCQOu9WsV1BliKqI6hBocMSPrP
5qy6DoXZo/n2hgpYSZE9gDJR+3j1LtuF5lWVDJ38jOoDZnwm2s6vRHJ0m0bi0E73
5qT5ALVhtIjyH5Z5139+6diz8mmgAPjlpcKr+EaQSO6MV71YXr/b9rcs1k8csKEe
FiF4m6WaKDkuc0yET6OaYuRRomYCIiMZPClt2kVC5ixSAYbjgf77fnr0ptEwRtW5
xprGL6KfRJq2HlWCm/bsbPnxs/d1EoNXFlPdCixYNAjwa7+dYZcTX/PItbwTR1St
hZDt5YglZxQgWq1G4JaZ6r72K+h+ZSSwBGY90iYEmsc0TYIbf5NpCgUqVGZK5l3j
cJBwt/RqQeg2eoLADdq4NIzducxTyEi2ccPZBN2LXCoiSdGpknJy8EKp9gBGiVda
KsUzr+1y9v9wOC0iXwqm7FGOxwpd+v5A2v0yaKRCNQNt9f49wCHb9DTiTjDzx2pI
KqqiNJurdOyhR7sYbqPIwkonoXuRXN/de+axGQFBwbATqkQ/DPo80oBxO4BSdvjs
AYSHpqp7KykbpILzRlwHUYa1yvtm0rqMkRXxGNtZCjb5c2U9mZbWmYz/ttjsjls0
F7mAY4am64kmPondySYRhgvTZ5nvHICIaWFh9DQzrsPCkjQFrzdqpuKlMhKwyvuF
238huWF6RRGzkoGWchVxN78qLzp8HVxIjfM5joW03LMHsgMDOPaGoH89cTfPjn4R
6lbQOgMakdxE+I04twRJ5otrSzwmsCU+yCW3InijeNqrXroTk6tvzTvviSrJtCQi
VktbJ8H+pTOlkSnO1hqHPoxh/3VE/79Tut11mFUXE1FbY9qWEknYEKzfqENFbf7c
vLTZpt9QELgEAPN3yi1jiEzESjQtAuMVmVWa2630EY2/lpaojN/nCbnCHxkTmods
mX0xPgmp1vRXmP/w8XKQMTzuAisce1ZGUFJ67TjZ+VjQk9bbt0RqLgBmPNrPetTV
tB5nTdin6VI4NuIi60vHjjZpGYyiS8JeK8w+MFzpt4ZzlleZg5ByK6WZ0KGxymB5
bW1Rqar9r2l+KQkhHN+U8M9q7pd/d/JTIEp6AqCgcUFozQOCFx1yYzwOXyKh4pHz
4gmoddX2PW7x/FJzTOIJXrLNxWTA6sT23XpFzpMuVpgwRJzI1hKIhuPD9/g7gkaf
IBdEpxGSURLCVDziURMUnwzX2z5uo8QahLZg691MK7z42p2QTtTt34g0PC9VTDkC
R5ZLCvq6YhD7l6kSM/FO7AdKy/LBV2aqxqDVzJzeWKuolDJ1wToJfIf+EZgqFpdt
7e7ggKaZ3H8ElNfp9Y6wRGXpmdVMNJCSuOHe3l0x6ljHseigRHn0I3PPkzAvnv2o
0vwRmCF4oCVnU671p/z9gp9vk7EB07NXCmPCKcvmLSBGWwL4ADuiTGsHbkP0Z/vS
UxWDclO6DXmSqt5Se7kG7slMJorBo7ORgq9eqOWsCNwyZS5MEFsDX7A0k/picteG
4GhJXBJOtZhVTSEWmbTidAbo613Tf5bXY+GcR+cN0bFGkcAgzijIiJtTKIw0fD9K
VixAreZyG8PnV9owxaWGzwXj+RJLU21rEmASoHdeVGrNqfslq/n/0EGma1uaRP2+
cw2t3vonptJgo+iGcIRlw1jd0yncjJ/GFLOO5bXj/GDyMik/A2PmvF4ogQFtKs1w
5Ut9X7Qg3XIVMyuvEgUFD6wgyeEZJo6XhcQn2saBMaF/Lgm9VFljydPZVwS1+S0o
UWQY7vJHOctbitTlFbEZ+/L0Us0Bqj4YslvlTIriIiVytGQg2l4kZE11bQeU+9kR
dgdqpAweLFRl693pSSIYzqYI6ECJRcPfe3Pz3lDwoYHWriakiSUmS3DSmnCLSfol
vno3/gF/Zk6CaVrb1pnXw7VHvhq8mGZ4+YV59QhpAQf0ASzQ7BVQHDg91DFwdqMd
Dvth1WLWhHmhuSXUgAsWDeBpKrBBy+t8LZZJSNB9xgL4geM9cdrj0F4BKhT4ajqY
TSyESEWcxuITpYdlmJLUfSKRfzmV/qrvSQl1D+zppMdTGuaeCEl9PvdmZjvF2uWM
puc0QKz4BFMLGvfoxPqPZ+289te2Nq8KGCJKwg09xCuLDJv8uz3/JJqF0c7YGxSg
JhrRLqfBNttITMlH1hgKjJmxAxYyagiLQVGqILpv5BEZWXL/85CEstmS68kCsSWj
PcufZfTdnQ31LRWGl305NKhm/8ogsdIbdAr3fEgaxk7oAyYhdfFwOsNbUg0BIYWL
HJc2A8dLaPLMlf44qUXhJ/UJgbi7dVYxP3TMZ1lrK2TzZ0C/7K9k7SAjPbhpf31s
7Yzr9aGLzr4ypD3da72rtq674A+BjpxTd0f7jhFkDD8Q1h2QWyWG7jMQzGl2w78a
hHm/v69plvOkjo7e80OLVQ9qXreA8iN7/CSjCcxTx1g+Ycx2AncQzkmymcmGH1g8
xKve6LhnDAySWnjspS0PE3baDKmOwyF6hhl22c13GXLQ7JZP1FkbestdCU1DDUa6
TqBvXn0+J3JkTTwD5WmULD1QsKNaXkaQ5TEXsYrASz2ZrK3ltB+RYI5qCzNB1vgh
b378BZsHgth0t67REQQsVNfFpxLmb/AuY8WsfxWH3x9jc/MNU4WSQaWr+yyK6Fcl
TDuOOUfO50B3Xgi0CS7pojXH/9VCwY4xpc8xcodFLzXKQB5YyyP2PKn4O0mJ9nzF
X3GDg0xvt7Z7hp5AevfDwFRwBXiObRb73gFc7RBfvxIGvTk6WnsPtzExXdfIxqfZ
iVuASgkxCNLJvDt5geDo4jjC6mCXlkiCpY7igrySKSUb5/r7Nch2Z3yI29QA6FrP
XWjiwpGPWsH7C7u5FG2fN8xpDdCLPyLiAGGcXaaK1TRqymFl4ijpFaMah8ND63vY
HimhVylSxFnFnQiuKkoC/6aQcAg8a2hNg7FGqc8fXxj6djvai2jUT4shGP+4WsYN
OWQl3n9u7l3VOi5Mz52ZnN207xzK4D14zzm2bDKSwMw4ncBLVhwe1S675BJcKn6G
OKA9xgTKkZ5BAUtAGglBoVZZgkwIiGyAvOybTm7GdR3PYOYCfqt1rWbGEhbrRgS5
n+kArLE0LwKwtJOWLPrEhnJgLtca5SaJ1bWrz1Gw9/kCRHJV2PMdDApbdQwBO7LH
NwYdzHkWcU6/ACMn1ihfWkPchMGSzGqsW54VauvMn/8KJTwSiKUYaXxwa1AGpmby
U/g3cUIXr6CYazZP21buGuWABhciIIpAHxLjGOnvL8OMiZ8CUp0bwMauI2l9gO+z
ZZCTVGI2lIJMQLJlCNxoX++Z7EV7NbMwvqczSutvNdprq6xYk0vbCQ09pL9rm0bb
XJ2ThDL7H/Pg030RwO04CjCgLh6UXFY9BRJVKesrrlsvKQqvaQ37V9iut3cNYREU
1udoOvDMIYfC+ecd1AV4gaiI742wxkQdeugh7o2uEhMNNLTY5IyIrY3n1Z5yIwvw
YpqkrqtzJvhVeefVtpT7QTBUK8IS3mHXRt/DaQt7KnQdUM3NjndHc3eZvRFdHmCM
Iu0rCi0r+M3HmkYbTyqenyXB8qbP2EgeYXXjJf2d55TsPY3ofJQ5yHritSbiYxFC
LDjKeFtA7vlzSK4Jn35sCqHVEM5y7rWKpb+kWQFPvm+HB+tYYtwoK3N3q/Uei18K
a7+i0sEnqZh8R33o6Ymdr3JYq/8BeB1JNYM83j33TwQ0Gjwxm0u8U2jCyogcD+Px
IwWyK0/PLdzmaxpvOyBHRNrnhKUuSPLxhiark2Siw8xr9/ykjP6G2FcBKQzjcNvv
WPCH26YZ85shYD76lyRVfZRQBKk4dmOa+T+OyiNy+w3x03u7iCxNrinhyP3+R9/f
0dr8pTRLHJhxjZVJQwKuNxfk2On2rWrpB/+FOepX2kzb1ToagXXQ6FPxi4wBCxUn
TS9Wva0syKlf0p5WHsf3Fd197JZz/rVv8BGcgo5bc4Ia0pllArGA5YQlOAVjyhrt
p47e2c/UdEpl9AtK6+y1gKGILWHd2QyI0tAOLtaxukGiaxxDXl7BPd4ZHGeK2e5X
eub4aGuiUcz0ynPBYeb9GX0UYXV/sFd1ntJzZD/PKozO7cU7gssfmpMmlMCieGyy
6nkTB8UuskHqYNUt+0HA0/fGAoC1M4pDqRFSriyjf31osYamOk1v/wyAMronDjTS
hQcWe6j2uKWi3HpI1q8MpQqLZ4osO57DNOJ4vHK6g3JT3HYFBde4lkpRmzdTGyaI
sBqhBj2ST4XINTDO/5POUFzFmwMbQuF0FwyyssufLSdUQNPjb26tsDsNhdxAlzPW
3Id9zrV46p5QkOpJ2zcMBBnvaRmHYI9t7bqJxTrvQXOffX49bDacLRJTCPzExqmJ
NIsbP//J25OtAKQChi9FYNObaPJ7TBMHLwHowvotDL6lpHzouB6xKRWDhlBK0+/x
HDvrANEBEpaaesk94oMo4HYKtpFF4r0iIZtBef1WWqKV3Mji20QGWFX0XGLN1YeT
+mgo1copJNYQjLQfbjqicwmYrPR3U6V8e3zZn5Jg9A76EAodbIr26MylR2AGsKcn
kAB/TIpqH5E3i7OdW7qB58TPOmclcclKYIuScokHndUDcuFX4nz5Z8HE6RZUJXLd
OWwGduVdP9VgiL8ULr8LXxVINbXLTMBZhP8KBHfX3UnNrW42hlENh3PWI8zZFuiI
v9JGNhRDVbyxyK1kk+oZbzEdfED/jAIOzf7g1opUFdpZ4x6ewEccNSw+74lRsIO+
/D/i1ScbE7nKqyVAkq3v8XbFbpuYK1SqQO6evFgL1nmzAUbodNZE/XRFC+YTPik2
I9aCRxM0wrCflVTC740JokC+FEBgtkDDIH7Bbtblsgq4XutVsa0u+lDf3vZRPObb
8ObRurELZX2OrhBYaXiRcVAL48rkKWU2I4HKo1ARVTW2ghLvWyqgdv87HEot/J3u
Csfgoi+hYqq3ttR+9FUGnhCyi+9ExZJ389y7k+OmhWLB9/o+OXBeGs2LwYb+n1Uq
MUihI4R9aSdM92vbV90ECA/XzphAmwIadNa401nT0bkT1Y6VcRWSHFXJZbh5od6q
CMYAI4OwgdTBZra2tNFJvez6l3GI022cjRzCe9y7MY6zdz6fRU4CmJgSLd6jOB2V
9euEcWd8MPzDxE31tkKNRGHlKncuGkEursue/lwZPM4luM07LYMKGuw+EcaCbITV
IzZSbiwFMKl53yCDi4dnCimoeMVMIcv/nMOXknmiYdHvGjsx3fHrq7P4oa5M5yIl
A/Nl6089qRYIaqFPcTXgr6Y2WncgEvs+ujELMPOXuoEPgQUD13RtFx5bARnwYp0a
WpzEZsoCqGfPEMVU6FfZOPjfu3JBeL4Ou9ZIKMvhWhEqdu0EznYgN9Zv0sXW284c
B3UZYLZ32RRO2L031RPMRwQ3i7Zw625hkCibxHywANMLmXwTb61MxsfO72X550/3
UiChB/Be7wfk7Q4XC6Wj0bfEqB2ErH4QiN4NyN2zkDSdwhdl1bUIW8KjpzhYMjpd
UW6bfakMUHbKrWLRcXsKNR5PR9QFntQ/5FoqDE0Vlih6sKGWF5v/Lx3JnH6WdlcU
u1Ne/U1xXXDO33ZOR/K/ZNlkJOYpJtt7Db/Mf+vCDCnL5ePCMc53UBsKiULawYpw
Is056tQdsVeH2VmeRSMyWxrz/2kOINtdHeT6aAB+vJEOG7ccaXxpFxenY1BrK6X3
1i+hln0KK25f5iX7vDrwYMk8Er+ElfdoLHjF+nuQPwE0iuPJuPCrv3rm0nzbddqB
y8OsECnWFKsYSO9Uo5Fv/rvLPMVW55QnrLwE2Ru2tgMd2ZBe6ZcZeH+8cgm5zMXQ
AS5fGZ4TUBKnUvMcgwJUZKU5s+5Auawx8KM3y1iNiBC0eVMQHuLDH/GSWgBCGFv9
lO8qEXXtq4RwO1suYapJpwnjlmzjiV9px0DQl0KshAVHaC475EToSCaedobkl6wU
rjtYlebaZ8wWSOIOJ5EkWJ9dif9CDoQYca+sGl/3QhJUyLwHDg8SE4n/5yblARWS
otXyq3rKMNz7AklSwfxIldwyrG87UT5jP266p+DpK4AUnRcZ+Nb8RaXE7Z9gkWn2
zgICdTSOn+7pNguznVn0FA9nBeACGRlw6GcsnGEzvxEUlZWzT4s/slhd3+dI8MLr
GAcIVU6AAW+8LHHNBFyuUR/plBf0P7uHP5O5IZEtiN7ZYlSwud5nEq6j9UBnbl8l
MawfPfh8ixA1XMRlnn5QIs8Jt5jmwkDm4VHgGXm1URHw9dE4Xe6ZqATHT0RIqaUw
B2KZXi6uakOjB2MXe3ZVDP4NCvS3qw21UBGu6NXC8HGn7hgmeZfmRyCg86Bj9f/b
62DAvMYfUhNWKt20rTZ9Kpj7StMUg1Q+OV1JeKosHuBtW9vLAmdH3uFpn2Q+6TLO
JDPmSCbveqFvwhx5gH6OYLXwi+jxwZhBBCohGad/wsWJGbq3sGSVKyQ8+PRVPX8D
z6bZz7B/5T+ssDStY95nfwXtWPiITwAiNcrO1p6Ol5fOCerd0Cp49lytxNiYURG8
waUsyFezLWqxiPzQVvZtgFSeQ3gb/Tf76QbnDXgkYVFKHWW6MgorKspTl1snxtkC
rwDVVaQrrbICSpNZQzz5cH34cCIiCifOu3dL7vzx4u0IPCCp7DbzZN4qkr8YEJvG
8yMNr4c0K/oXvuyihG5W8iq7BKVRG3jHtVjvO+64wQRfPPq4udpm/uiC9xPseErr
IXYdmSlVm4Z20IB8Z0b8tVa1Q4Q3S6dq2OU9CKK/2g78NlKI1YhWkQbLFdW+SF58
R4E/GKNjGc47Os7HSTApg3tVPHXxuIVCGlWFWcmxCFsIkXarVcbldRoOGi1NcZaF
XPm5kDdyMhc/jNz/EHhweOUoUuHKGxxXSNdyx3D+1tpvYeePDhqE4ipJ6G8wO3z6
tdZJG0FtOy4tPbuj73JRN21cNQ/D1ZlF3kjsV+SIE5n7C15jZ9cM9BgwSz+DVNRA
lk21DWlzfxeya6WhNchFCBhMuFHZr6nkG0lSYISIhDpawgK+9hxaUGg5Zqm0OBIj
hP67iLcRlc+puc7Y13s0dm7TfYDrzCn1T9oq6+IKiHWzt3wyZZ0Jn/FtdObmhqJ9
Sz3tpxgKWTBmnmPGaHBOYXp0lamAgEFF3VZNpTt8zXfy9/acDb/F9S/Qar3Bs4Go
ErdxsChuBoeK5Mg9TEPbod1mzJB4QOuyJGl8hyESrJPOIs/oSepoBzbqQ60gF8Oo
xtIPrjrKV5KZ8j+ShLkvEaengynu23DDJ0x0uR3+U50hwMC33+yuT5RuSgUU7Gf5
H3zjUqyHiXyDR1qo3SrerA==
//pragma protect end_data_block
//pragma protect digest_block
GNrKuPIC1VnJDyP7c8+eKJUFPL8=
//pragma protect end_digest_block
//pragma protect end_protected

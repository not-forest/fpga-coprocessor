��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���X��f;��on�# ���5"0 �T�PL7T�0����Ǿ*�Յ�'x���!�����*��w���0`>���M�I��M���M�At�YY?��w�/��
��D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F���r c�Y�mI�1M�Adb�t,�i���ʂps"����1�BEp�e��mN�Iq)iv�������K�W�Z��ö�?�柋N�5�Y�!%����A�"��m�I��U��>M����ѿnj�D�z*=b	f��+���Y��P�T>�����&t����p���n�7��%�8{ȞU�����X��4m�b�ד5�H��L&F��B�8��zI��XU#�d���P��
Y�q#�+N�C8�����M�~��ۢ����)�^��I�4 k�ս�+�[�Nt=�nr���7��<YQ�v�X�r�ʙ�����$iu����6Bֽ��T�o�bl�Xy��~��,Ll��R\]�3��ww]�z���Y�"p��2����C�jP�MWu��0��;����̩pA�!q��u��l��)�S��VVYVԣ�\�p�=���h��h���,R�d�$~��ٖnU$`.K��Ȋ��k����݀2��I,��oc�-��l�-�<ʷh��l�/VVH��#�ie�ig�b����V+�����Pho�����vD��N�H������s�ӁJl���9G�c8�/AQ>.�M���zSj�~�.�]AF�m����ȖR.�}���q���Ja᭩�:�r0��W0��V$1����忁;�4I��YX��~]J�\o���]�S��L��"w:ʍ��@c��&�T�,����TZ��'�eHQM�jHX\�J�F�6.�'�QRR`E�� ���21Ea� ��넄AZ�<�U�?�.�íL�����8����w��V�E0霒�e���BGr�%j/](�}M-���C�'pr�W
��"F�L�	LF[��	��)�:3��rt�B�'�$�)A{�u\	D\圪N4�}�oV�K�6�ҫ���K��X�hs�O	�ý�⫸C��d���Ug��9�?���)�J�Ǉ�!����$�!$  ���a�؜\���{�/R|�W�I���/�g���C�`�������@��|=�i�N㔾����#o��Џ�2p+��k7�|~إn7�^kU{n�Ŏ����7�&��T����/��[���ż'�+�:[�
�X�Q��ܿ�|9 ���3{N��@���.�nU���f�47�&�a�"1J���YcYq���`�'�9�Ck2�J1c�*?��Ҥ��JN!\i�)�m��,;Zj��@�l5�<^�r�d�,�������SD�|nVZ������#5����]�Z(|דDăn���z�VG#Dn�V�6z߿0������xK_�<�����ȧp��JI�h�k�xvH�K3�s��z�3e�Ϧ�k>|�V{����
fNޠ��D�`�����a�WQi���sF��`��3q�~)g:m[��:.x�)�@�N^�	�祗��݁G�u^���:&3v.�|$x�J�BJM�X>c�w�
Y�Wr�,X6�G��W�`!���K�	ٮc�F�\�����|�7>\w�[:�&v�0����͔jJ�kfO
�,凢���նu	��CI�����2�:� ��@��-G7�2�:��=W!Y�=rbo#w��W��f/�o$2֊���5k���l!߲T��^H�ق
�,�K=�l�b����:;<e���0Ka��TM���`�_�k��d���Gg�	Y�'�I��;�7V�k�D��m\2em�T�a�Pٙ��d˄ů6z�E^�c����U�����8"���d��L>��I���̫V G7T�N D}NmHy��y�g�(4ɡ��3�"0�\��MĦu��{���̽��Ũ`��K�v1* ����������n� ����*�x*�
��,��P�3hw莗�5�b�C$��]?��j����e��շv�� �S�R�b��*V]��v�Ph��SԒ@=�´n���es��1��O���z�)`J���r-pp=��}ne�N��z�0w�vt��� ;/X�$*͝��h8-~����tAkߍ�G�1��,N-Fq.���o,Cqp�^GEe��P��!W2���M�����oCx#���Zs�bK�
)`(����"�����ߥCw�A�����8��D����4ىQ��2$�[f��<��Hb4=�욧���ē��)()�$�|QPtm������v�@��!���d�<���`��i�O@��	����x+��x4+���٩�(T�ϳm �2MŤz��������F��]���)�c[_C�e8ߴ���(�	�e���ǌ~����G�ՁJ�֥?�@�#ʮ�?e&���d˩�I�Y�e!CP����Upx�4h�s�z��4_�A�� ��ӎ�0U2�B�.�9vQ�3BK�S�~`Y$�&��oH�X�vP��{/'��Lɡ,�f�Z�{�&(����K�)�w�� �Y���6�-;���G��L�+}m�[w��%�Z8�RUjb���XcC
5'�88񥶬�W,
�����^3oYR��!���0VT��"�>��>Вu���r�G4����ί
����;��
Ɣ.6�S�{�j����{@V�\�n���h��W�c��b�rѫyO���bk�(�w7�Ӿ��; ̀��Ͼ�*�w�]թG�B��[o.�݃� ��<&��E{�l���:�����x�r���;L�Y�U�y�̧���S��ZW���{Č�@I7��+ ܡ6�nBc�l�o���u� �0����86�n]��D�ږ��x��\�Z�	$ﺞ�0a��$���AHmo&H#2�Z��,ǟ�P�b�"��@i)����eF-�7���C�/z? Yw��P�f���m�xXr�ԙ�=��g������C�@��B́�(�HC�}*��mR��n�l�l� Ǎ�M��BǜJ ��.x�"�����׾��Ж1��-���}㤂sO,l�?��5�J�C��@��<J ��m��*�Η�1�(z�/�0\6�ޯ>[[0_o�\�fz���*��Z�
��nM�m,�,ӲԜL� ^?÷��z�{��{\����K�a֪�(x�B��#�FIk�/�7̫c�S5F��"<���d,q��~$�7g}B�A����[u�ï@�;�v
��"��s��eɐ�� �e�gъ��A6~�]1��-d����{�z��B�lZ#m6�/ɵ����ߠ���F��3�B8[F2#4)=�	-��8a�C��	�&aO��m�\�	�z//b��r�L��n��	������!��~1��ښV#�穨�@�2I�< _���0�J��p]�J��+%^����2X����g+���j�.��^
�Ǔc��w� r��>J������E2�_��x��2���w����hko��JU p߄��D�8>��7�ۈA����-r�͈�w����1�8�r%k�����s�F�,�Lț�ը�0���ۈ��˼~諸Y�Y@F{�1�6��������h�Gd?��G�5�F�-���V��߂R-u��d���ͤ�e�0n�`5u��|�WP�������®ŭi��s�ƴ��T�g�X�=�v�S��V(�	�܅VXؕ��&aѠE��0<yF���
��I��3D\����J�B�lwr3��S}u��O>C���|�v�:aW��/
�Qg�ܘ�i��1�;M'֫?���2�i�8C��I�UlmY�R1�&K"��(ŕ�(Zv�����jڅg���_v<��,�zq/2��]��셠v����K!�Nkv����ĺ����I�w��*|�1z�b�ѭh��"��3J��e<�^IO�� ��B��o�g?d���ƿ�m��nP�����֌����fq�:��% �V��E}�:P��?�I�4s���d�T�4�!�	E��:i�`�u ^�L������P�����}�!g4�i��5�fס:�&�����M��;�	��v���S�ސ����}Nl�%0(@+4;��D��2Ԋ\��j��HI!�eIΘN�!�I2/M e�������
�")�x�?j\/ȁ6�7����="tϰ�e� B�1�w�@/�Hɞ;�H���):�m��k�'�zs����}5T�)Ӓ7����Op���(
s*^�'4yt�%���i���ʒ��[�9헰�k!�;ʱ�{]��-t$U� ������vu ��p=�q6��w)
dF�����v�x(y����吴tH�lBZ��a3��3��Ϫ`��������28&�60	l��ܻK�.�a� ���
O۠Z��?>����r52�[ȧ��#�c�+��|����W}��c�����⸡�o7����v7��������J���U��d�2��>�!�-,�����\���)~htQj�a��ҬYl#|�%y�L.�gf��a��Q�A=��I��ٓ���#�Ay�Xy��05m��Z'�j� #��� 8&�a手�j��޷=����Ъ�ǎU0��J㪝.�OY<B�l��՜��
i���zgS]�;�?E8�=�#�����	&vGO����fS�Y4�/R�xl#I��4�W�nUѕ.|�����*�i�<P�" ��%��̤}=�SjD���ȑ���C�`(G_b�����!i�* y*��v�%��tW/c�Hc�������d�TVJ-�o��!��<hh���(�yz�⯻�F��0%���y��ɷ�'�~۷r�����)(諪�(��>:�P�� V�h��(�J��h ��}��\�c�\��޼M�d6oگ�[�]ǨC�ɉ�\��mY�H'�F�]���b��g-���,�� hUOx����P9�����Sg������ #�߈O����E+.����F7m���2[=��'K�F6e�����2X#3d�9��|�Q��y�cpP��x�D	=Bx�D������YC�(~���]	�>��ӊ
�%�q�-OE�p�]8g}Js�^pz1t|�����7���$T�D�]�nc�6cǻ��9f��[��^����xW·A?U�I<oͳJ�S=~���>���s3Ұ%U"3����oğŤ��+���Z�X�"�5LUs���j�GD�/6�F[��|[�����bhϩ5���$�}Ou��w� ����VXr,n+H�^p�X�t1�ϟ&�0o�$���u>ܛ��������� z�O�G��=��@�:Ԝm��{���	-����Y\�dB��撾b��x5�r wF����@���~I�Ϥ��,s��+�ĉTjN�����b�W�7H(`K}DyW����w\&x��Z_��<�G��_нSu��{�ەz��-�,t�#�ǫ���������}�Cw��W���e�$√47C�x�m�yDs��7	�'��k�/��Y^���D���$�t��.��whQ&�Ac ��E��lߪԛ�L���6��m�P��ϯ�ȌJ{�|����3����P�}��T�uX�3�M8?�8zoڲ��7��s�Z�U���$R��Z|S���c5V�^)
T�T��j��1��&��2���&�-g��a~\"�G6�}&h=�Q�˷ ]�͎Q/���-� ��#IΝ��WȰ��(%UP�R8
�	�w�1�A����A��1���BE}�Q5힩~2�/�݋��b-辤Y�l�����{#C�FPָ�D]�g�.��`� !�Q�@��2C~����w�o�Ypw�K¥�䑽BjT�i�e��"y�l�>D�R���`D����5�2�ņ��V�lpr����zZ�t��m3#�Az��� &Ȧ�a/����}�+H0�҃_h��\�V�$��lG�VqPA��ȡ;��ܻ�� !m�L��{��{�uꗭ����l*��נE�hL�y���*�V�
I0�ûq����A��F�ꅰ��ϖ�������Z�)w_y���;��[��!�Ji5M�F����3E@;㽛�dj���[�,���-�[�eo=���d��a�2�JXڢ�G`9�z��{�Tqo�R�3Q@�6����C�z�A������� �/�k��/cM�"	�A��NqO�e[�����G��<�{���k
�O�%�W��!nd�s��E�H<�v�3,́X����5LZ�R�:��Μpr�%G�_Ǩ��|ɋ��/�o4�N)��5��?�$P�`��|ឌ��AFئ��BfZ�C>�\���2��˲�_/>�t�UK ��տP��^hw�[�V7��g��rgaKOYG�m����GF���_�bO*���S,X��o[t`�N�� �Y;�k)th�쌍�������f=����=��m���B!�0��q��m8�u�D��<r�Ģ��ˣ �}i����vH��}ĽK�r�5`|��9���\��M��(�E�͟;��]?��h�ҋ�I��q��^��;`Eԅd��c9m�M2�n4Ԭa��*u��Li�����N�֦��#��V
���*\%˴�X�D���]O[_I����3�޻?h|���j ���e��8���SF���~"����&k��V�D����H�z�
?�&T�xȪ��lo̭H���<&q���;Y���&�5"�"״E�0_l���OZ|�f�l�9�������1W�X����#k"
��N�hF	8x���'ɞ�d�<&��?�Ue<@P��V�փ�_��R�V���s)�B�R��Vm\�F�@|a+'"��=*�J��)�	���XN��L8/��[�|�G��[�y�;��m��{D7j�!޿�)oCH��4e��H������ڊ����J�XxȱJ�l����n�KX�C�O�/�U R�Y[N>�{�z�`�t�IvoF�"u�Xa|��W�ߧ�Q5�B�}� G�gi�����G����� ���ȭ�+�h�9�ٮSF�*��뢘:/<�mi�zɞE _[�'YÛi6��r�uCqP3��6��F�&�lQ�Sڂ�?�h}T���u$�+�F@+?�.���g��R��Y�G�r���^��r�5H��]t�m�j�$ծ!�z\��a"�i$���'�zQx���_�ńx�u7e��W�2��J�o�(��D��Jj���ʊIԇ�|ְv}>ȫ�։{�gk$Z����"������y��/0�ħh5�n,����c�]�\��}�k��]��+%��sw���T3�j��lA|�� Ƶ�F1�]�h���g�Ֆ�:8K�ɋFO5ZƔ�5�����]�仜�I1B��[�I���[k8��K�� �~!�UÒ?���4�"���w�.���M
�,h��~�LN�T�DEd>�h��#BC�ݖ�����i�q�^-Xk�I��
Nq(�_=��3.I�Pt[�PQ���1a��	4���ܺ�Wnj󻾬epx����#ʋ��9�SFӊm�9�/�D�E�O7EUv0��K����Ѽ�wTi��!2ױ�v�I�G)���~��t��6A�iz�H�.��2�:��N&;�y��%�l<z�h2���Qm	�m+����K��� ��B�F�^3|E��T47.6�,�\�"�FXu�w�5��76��ey��f���oJS(2?u���1>ֽ�'��&�@v�����lAv�CB�g�@ƣ���m�ڹ|Ͱ�sw����6X�L|0E;x?�Z���n�C�׻�����o� ����⹀_���A��7�*I�֐�.c
�����~�:2���v�pU���^�b�K���p�rO����j��𡊬�TxF>�vy@����@!�z��X[P	p�dp��N������X�,w��x���Q Mb�r9�W��>Ml�BE:耺;W�8�(WS���U�؊�g�G?-�Fc���4k��9��/��Mɂ �xZ��I�ɰrjD�^���91��/;��_�0��2�v#���C�)�
r�d^��6�i��4�a�m�C�j<!��<�a����.��
Fm%����A,�R�x��ق5"���&�u5k!oY7}�C��ӁҟQ��$v+U4�Oz�2�A�"ҋF�7v9��n�%��H��k��{�m��Er��Q�������"�TƜ�y���R����ۙ��^�F��+^�>nne� *N ���h`���-���#���U�v,J�2D��{)��5g�/��7V���ǟXef<5M��X�J/���y-:6���݅'�3dno�&����-����Z��! C�1WJ0�OC��ԍL�]s�aώ`����/hP=!��ye�0�?���~���-��������x
'.�kP�~Oh�	����Ƣ�p��_�C��
��&��Y�%A�<L�D�&.�Ѡ�n �&����G�.��/V#8Т�nqY�v}����i�k�>s}3�M�����Z2�"�`єF�ǀ��F4n/�B�<[E���~�q�.n�4g�f
ߥ��lX+1���#��"��{L^m,�	A.Q�ze^P�Ձ�{�3�����ZP��,���C"�`a��^E�|Zڵ0�����Bkj�Q��XCM����#��	j3Dk]I�OjX�w��'��D���RJ�j^�jI##�*k?�!/�ͅ�~ �i�%��W���|~pk�����;!�_��mн��mpW~��E��F���ڭ$Ls�W�a��LXP@u�k�u�Ht90��<���k��8���l�A�΂V�m��Ehpͦ{��Lr���v�f։jy=�o
�6R�O��!B�b4� FE6J�Y���F_�?brd��RmKN��{i6�u�CZ�8,�6��O:�rKЦ��q�ü�������N7�&���w1^���O��_��h��ʌ�����,!H2��|�Ý��;��G�Lz���XW�s�L���6����0����RF+��{�>)�1MQ�����I�LI�ڮ��X�؅�:��+�I��/.�|~��h�H �Tn<��X�����p���"洴T,>�{�!�z�m��a�4�a�b&�=��)|�c��ä|�8in��&�0Tx�����<c�������NL�8��ӱ՞.�fp͑��Bh�����bτ���P��_��j��kζz+lc15;{N�M��7hP��t�Xgqf.�P*�4S4Ć)�:e�朱"/:q�jw@�����=6��kU� 6p�A��ԍn���u]C�aDh�Ů�^&��ߦ�`��X�0�\�.Ȯ8n�e�B��o%�+v�'��]g��]+���6-�I(��L�x>-T)o��j������a#x��YҀ<���X�y���7v#����M��1�3���'B�r�p'�����ʙCp7�?��F��y��>���v��B&���_�H���<Jy_u ��uۤ�E>�&��߭^ٴ��e�A�,h,jfkY��_X�����#�o���-@�y��z�贫�=kc�W����Ǧ���Mvu@�J�Jҕea���N��n�:nW���X��f�ߍ��IAK�٦�'��k���CI��t07w�ba�.'�=����cA��R����$L��4`]�p����ދ s�ŕJ�3�xMF��b
rZoK& ���~+�#8��Xe|�����bt���aV���լ��O5j��}ӝq��w��"{5��E�«�vE)1#C��j��q����
�Zc�)c@vʚ����n#�ץ,Q�'1�?��;e�[� �����p�b*���0&���I��ae�����E����1��*�B�M����{h\�ՈL8l'�x�g��
C���,0TL`�{�2�-�_��axT��
�Dƚ�K�Kլ[��Wk����/��߀��R<F�	U��`#��f���X��g�oK9W�x�\�"�Nw2^#L�w ;.T?8�OR�4��S�ҽ��xJ����-�<��a��Ɏ��/$��E2��'=G?N�;܀�Q�S�o:.�Nl�S�gScB���M1-�èH���a�]�+�þ߱`�%`��:�����k�/� ғLz`�or�6��ǫ��9&yqJ'\5!�Rw'�w�p���޽=V	���ٟ����m�϶���[��e9�Λ��h�ZW�q�`�/��:�����x�TWi��2�W}�ň��̂���]2��L^�����jv�ϵ����Km�]���;+QG����y;�Qr�W�.�=E����47(� ��5�l��@�Q>;��-������/T�.�+L�3��xΠ��	�cY�\�{ؽ�ۮ��I�x��W�_8j���ˣ:��2<�['l=XP�}	�8�B��0m�!k��v������:�*#8Oo��&=l_Sn�B��sM_�[2c�W�&</��ٞ2Ͱ%�Jf]��Ί�W?���l�a�<*\Y�3�7�O��{��z8nj64�5�'��Du����r��}z�SF
���KŻ�dh?<(;�D}��x���a�\p��L�;�^�J�fk���ʅR�7��p��N�&���Jt���ʺmO�ά��R���Fj���%kRj��0����~*ߒza�-���DGS��B�3����v���W��>���Ʋڮ� �<����R���A��Q�3��	�ϡe��x�w�i ����>�|{��.(�/��/ڍH���9�����W����⼪��WO�L(*=)��\1�d�,��0��¥-��ޣH9i��%��óM"7�(�f���4������<�ʫ�1F��7�c�4��N��"h�;zp��#j�O^�i�Wmw�����]��������#��!��W���0_M��BS������T������
0���$�3ܺw����B�ȟ<�����v���y��_�d�Z��3�FZ7��an��z��B���` tl�I�g�b������:�w'��aV�JI��X�d�_�Խ��̀v(��,w4���/"P>�H�h2+��_/��օl�fW�(L�Ȳ����n�y�%T���G�=7���h��S�B��Һ�M�I�`䂮��5���9;��"����꯴ڜ��l���x�t�!9�� �S��H�O�ٴ=�p�A���_'�
�T(&�k�l��f-�뮹�7�mߤ馼V���J�o:~qSݍ�)/�
����X����7̺s����o:���/�lbi ��*U��h"x��0��c��Kn1]_;����X�&�H"�+k�8�����H��Q��a�!��.���+?�M�J��T	��*�6\���/"_�`��2����#p����?���Sh)�C�]�6��@4>�qX�˝M�g~b�O���R�G+�7�jw�Ġ���^�����q���=��IS��P��l18�K��l���1�c���yz��W�"�)���������)�G��D�Z�c�p�wF3*:���S;H��Sǝ��B�3&px[/����R �vjM��K-v!j�n�&��qb� ��:}�i�:���&��,�`��T��Xϖ{�O��,�V�s`U)$3����9�UX<P��X.���.?���]+������`\Axt�| �q��}�s�݅���ޒ�;ʸ�5;�����-�批�v�����/Ώ&��[�}5��Θ��� ɋ'�lJg�^�H�|A�ʻ�|Rzt���[�\��iXS�o��R�F{�U����ƝV6�Y�Dj�V#�.B�I7sS}$~���;J�K+�!iߧ��5�/�k��'�M�K:�^$G�P�	�?=��ۢ'Zi@��ZQ��@�˄o��!�|��{�QOf��p4H��C� ����8zL�7'�2�{��!��T;��򪞇vmI���&!��(L�	��?<G| �y�^���8/����Id	�'��)>(�d���-AΛz�,Z���f/�x�){Z;U0��#��,s�؜�O7�;0�
�c�>�v� l2-��V?_�����#�\y��uy��lϽ"&�Y+ �y�/�l��Ixo�~�J�矒v%(�S��kM{˸ �$�m��46&#	>�O�A�S�N;���v�� L��~��(�mC%��!!B�RR��{�*C Q����qWw�gq2Muǆ���^($GQ�
�1}н�S�aF@_#�g�l{����K���?E*���"��G�[����n�!��)��q���h/_5���Te+paE�+�H�Z���N}yro�GHOÿ,���OR�����Ɇ/��r�
���qw!D����ϟ(5mRFQ��_F�ˬ��+m���7�*s1���X}ס$�_�{q��M�k�/��4���.�X��j>���G��X/r]վ1<ׂ�p�_��u����Y���Ǳ�\�
��>�<9įe���رBS{G�G���mT
9(|^н��_�?Lwr�*I��o���/yUN4���Nr�m��%�(�Y�I��f��s�$4������j:����$OJ[���_0S2�"&;�>�B��[�^�NI%BX�7�A�3�*�[�u������ע�+zTn,��D���+
�㕲�AByT�Y�����Թ�ҩ�z�q㦳.��PқJ��Z�G�{>�ꊆ�'��5;�Y�o w��#\����U�w��Fg�n^������*W�����y'M��/J���βN��I}�MR�Q����1b�4��s�Vz"��KU�}��b�H�k�g�vo�UO�l���ǭ�	��̀t͚}��~Be�|�6|3)������e#�%�V�^���	��`�lXn��w���~v��	� �xw�.)��)Ӟ����<h.�2=�/����#�'e
�w]d�np�F
��sv0 S���@M�NǨ�/��l a�0��~���� M�f�:	5�@��ix	��`���@-��$[$�3Z����*�<Y%��#ԭil� ͈!h*���)�_a���f�I���g�@e��	�v���B�dX��$|հ�/<�1�okuۤ���'
yZ+]��>��^G~��mcY!���ר�_~8W ���4P4�u�ci-s�)�]�IJD��:J�j�Y86��ݬ�fE^eF��A�D}1�����PU���Sg�c$�T}�>�/ܸUxy�m%T�o7��h�v�iq�����Fܸ�0_+K�ʞ��j�E��ͯ^@�c�b�Z�[��E"��Hp]���x�⹷A��f�L�ݫ�P��k!�[L�t��sB�d�썍���%��������Q��KQ�}r�\_���W5U6n,(���
:	�!I�A��\Ÿ�<�o��������) cr��ݚ9���h�q�P$�u��XG���������S��4��L!OcX�ꑩ]����V�X� �b���k9�b��_�mk��@����d��g&`k�8��� �&�HǓ��}U��P `��3�3�/a�:��097�5��zba���}g��&.�3
��Z7z,<�,��:�K4>t1��'t�m�v|�3������.�qc۾ylMmU�R����D3��f:�N�s����!:�=;�M@�z(`eE�F��X:�6"��k@�akJ�:7����A`�.��d!����a*A(R�~��3�D�M���O ��R�.9.@0�����eE\��?�9����Md�מ�v񔭩��dB�}D��l8c���#�p1t5P�Ds����!}Ф���0d�	��L!����_\��R�r�驭���H8�9&l����W�G=�*9�ڍ����*��1�O�e�I�j>O
�g�t���1�nς�c�Zc�qq*�B@�x��ؾ���i�f3��	��S��BΔ�˱�5��&��3��@m�_-D������5�646���.������&B���{�@�'?�~�z�8�^�3��o�~F�&�����=��&l�<�k���v�ڥk��G1Q?-����~p_�bE~�%�M9�!Ƣ
~�_��@�Ĩ"��G�� �-�+P���" �zs�����b	,N�G\|��N3:Sq�e�a��W�p�d���y?y�g�*_3坏'hQ&��\�~�%�B�w�=������L�,�=Ĳ�{�Q�Vg��@��%�>qF�'���a�of��1I�'�E����b���7��9�%Q���_S��p�����TE��$Z	=���� R��a�3����y0���J�R��C�W�`�^X��1��	�� k�k�<ϒ� �P=���=E{�?���0q`��]iT��Utv
�er��Q�r8���i$�&1��Ğ�D�E�)Ę*n��?�S�d̙4Ҭi�I��a/�K��K
־�5`\�Y�W��P���)C�'ř�c*�&	,u����/!ΐ�^w[�[��*��NOϺM3�x������ �K�НV��"��=Ӭ�8�G��m6�Ey��5J�U�[G���Kq����$i-S�-�-�x�ɵ�#�g #����D��,�LOɧ��+��n�k�Tάh	p�.NZ�d-n��y�>vڀe->�N�c��f�$91�P����zpbF��{�������^��F��(f�m��`i�T��<̜6"_�
y#��W�7�>� �Kenvv�9���:�,0v���̒�4���������i1�<�g�4�p���C��Ǡ��aK@�>#�/�h����i����05���r�L��1V<(I �+<M�/|ikR����.W���͊ɓ��n���cӧ���a}'�.�THo�v��K�K%�����U���]S�_/sr��� /�Q�O�ωK86�~xt�TdK�p!ڝ�Q��#�O�d؝�j���r�X�/bBz�f/�" H��;{>9�6�/R-��*ߍ���J�%���;x"@d�.�[��ս�	k���f΁V˄�~��Ȼ��Ab���Z� �=�3��H� `W���^�\�C契��7 q��l�/��TU^�e�+�F��Oj��t]�&>a�ٚ~'#P\|`�ٙ�aJB��4)~7��Dָ���`i0�q��o��Qrʛ����$;@��:1�Ԕ`u�l�B��b]�:܆�[x8�'L���x�$�4�Y:s���B����x=2�ic _���@�f!����*��~n�u�K8(܃@s�������5ϾE���>�B�K�3�2߽�=��A���������iI��[m�E��|Y	Tc$E�p*+��&[��1[��^ہ�=�6/L��O������,��i��pR�_�xR� B�x�YM�$G��]w�g*$�o&ق���ׅ�U�j��ܖ5�Y��}�7�����4�m�cS�D�)!��}�^��F&��4�Q�H1EWy���J�C�[�ȸCx@6[{c�:���t���͜*�X}YO��� �p5�B(Wm�5���s<�?H/o�{x��'�XW��^��������h+$�J�TMi��ws+�$/J ؾ-�ŵn_�3�y�a[	^d���T1�.
V��X��nR}�1M�����tcU7#R�����,ML�ua�K�s@C�mm0e��d�Ȫ�����R`���a��z����mx��X^4�~��z�BWV��"��,�<�xG����G!��)/!�)�f��s���H2Z�>���@�/Kec����o��^	�q�-}֐5.��N����V����g�WKB��p(��U���ó�ICHc��5����v:�-���8'�>�0Oc�w���?��E��K�R!l+�߆�R����G�~k����Ү�0O�h_ND��(�K]2��E#0���vm���G��ЪV�+���3�gZͻ�͏%1ӨZ�z�َ4�G��c���|�@�o�s2��v�|�t�K0��J0^e��o��*�]�a���B��X��D8K�g+�+�dЁ(�p�x�����i�iK���d1���&(����qt޶�QonXE�6��q<e��s���k]-E7��kҘ��Xٓ�.p�dH%,�ϕ�\&@��u]���Ma�2F�0
�w�Y�Jg���`�0�]"{�w��N���cq���{�PN�2"�=.˽�&�Ӓ�k�? _�]P5Xjۻ ��K��d���0���j���ߢ�~�*�{����S����J�Y���!̯��>�_wu�� ���	/#�	b��>��=�M_8�=C���p�߉��6А�	xk�jD���0E��� ��qO̦�/Q�9��aA��*�L4�F �uÙFa߁z���8�4R:vC����4({�e�f=iq�`�K�M*DZQ���_t�V��"�A�$�>I�oX�E��yOD2a�;CЭ��L\w��Ѽ��VF�5J�$�[ì�[�ﵰq�X.�D���3Xݘ����;�������,�k�`�fm���A��.�O�?q3�%u���2?H�"�Sӥ/ �g��a-,Q�AX*�~R��B�xN����x�{6������?���ӛ�b8ܠئ�K�ԕթ��1�K����r���HfY��t��.�y�n����eş;��gf��#�\��ڣ5L�Y>g:(*P�.�kt�F�+�{e�M�qo-"�x���	c�
��ڜ�������!|1���w�e�V� �i���te�Þ�+�6�����S.\��"��zs�M��t��O�x�(�ܘ6��b^�s�ct�����|정{3��eX�g�I��S����n��Ưg�Ǡ�8�M��$�m2v+���Iȋ3��){\  .��Dt��`��-D�%XWY�wy�h�9Xce��?lf޼��;�%½�<޷���YT:m��Va���_㒍��%������/)V��{qɖ�K���)1,�c�l�xM�a�[p��G����u�7�5]�+Z+#ˇ���N�ϴ@j�,�hT\J�����LV)���A�ȯ���|:*��֋.�|���j�e!^I������Q��B����={Ճ�:��Ԕ��6˼P��t�6��o����@�_ ��*
�/���Z.>\�%--Zꢎ@˞��؋Xf'(�\�U>C;�:�q=iK�H�H��X�/$ ��r��A�L:ʏ�Q@IQx
��p�i B+��UD��nq�Un�ǅ9�P@�lK����x�����|�Y���he�#=�4hO�����*~�pT�+�kc�����#X����� �q@̬�������'�$�ذ���^^�X��b��=Z5q��R8Z�l�P��U�����?�`vE�9{;k�$vqe�[�|A��g�A����?�� z��"6�5:�y	j�)�V�²��������e0rs�O�)n0��|R��BT�[9�x$vQ`R�����S��	�h�����AoH�!Y��*Z�6p,�ެ5�"@0������v�޾��!�bφ(�=�y;<\K�H����_zL<�݃���o���@ @-��vD@�(���E�7|����2jR�tw���j��<1�1���M>�z��������F"���+ph�@Ko5f�Зn�@�,� ~������ ��nb��w��Ū�����K�s�,����jh��E�*�6kr�:�2�|X����\h��N*ae��la]E&��7d3C�?�s�ж��\A1�������Z��r�I�J���&�Tg����	2�f���.z)���(�do�a�*��дl
�T��ˀK�ǔa�	ݐ�$"�o��`������GV�����:����
��C@�S1�ǷB)2�� j�Y����C�e�mM���۾^!���V�qS��K�w�7{�mY�?+<@�,h�Z�ؔ�w��C��V�FTu�Wԇ�����-}|��t�|�2�����A!���������cG5i��6Ȅ_q��І�b�d��V<��F}ᫎU���fTq����"�X՝:�`[�+ؠƕ;\/���>4�����mW�00�`���6ܐ�|���!ш����]��5����`��й�~w`�y_Y?+�U�� *8 �?�*Ϥ�+����׭���3�5��+U��X�m���\E���<�bwn?׎� 4��l�Ce�O8��S�i}P�H�%���)�Q�%�Au0���*0 *�k�)`������#s���z�� �S
1�;�5����;b�"�D8|[3S�I��gR#�5i������r���1�k����	���q�Gٷ�j#`1>��a�$�	�;η>��"zZ��G����fӺ�L^k�\����N�%��� ��B?�h�9|<�����a�
�#�w:�FJ䜾L����i@��B�" �U�����0;�T-Ŀ/'l F������`�#g�b>i|���K9Y�</@5�ܞ�����Ab�	G�۽Ǖf9:y�,$Jf_U��M�j���3B���0��<R�Kw 87�"�̋&�J�LOR.�ŧ(�.�.�4�&_G��x�m��=�������J����J-���x2��Wf;�;3$��3���\/+���lM��L��D�Q�(d�_��ND���4�>I�ad&:��I���.,��>v��b૨��~�d���T�v'�D"h��,c��T%��4	E���ՙ�r�ެs�@�����C�%_)��p錧+;�cj�K���D�؃�ĭ9��m� ��-�m��B�䯇2*�:�گ�z��Vd7!��
�\gʧ��zX!�����I�g����s�B���!ɛl��^��m4_	(�(�o��E�h�j���'�༔9rM�ל�n*Z�����_ϴj�������i�=��-�烄듿� ������̠�G5�0�H���-�x��0,���PZ�Cm�GnjޓbvM��]���(uz��M�4JIN�1��qc,U�4h�����m
�g����w
�����F���2#e��"ܸ9�`a�|�y㵍�ݎpH�f�]A�9)s���Q��.nT/�o�/I7Y�h��?�Hڙ��SHϪ��v?�x�wN�_�鷑��D%���'<x7 �U>�,�ӽ���{��؏U���_Y�@I�P���G�o��|_����0�'�,�$�،�h�9�p�A��ԤB	Y��put��6�2�Y��Zx�l�?��i�s�z/�c�#�!����zk\��7b�������7bə�Tu�#y��B��z��6@�-���X����gx6`7�L����4֗#�+j88��[���on}�vȶ��R%*�K�7���~Uk�Ã6I �>�
��y��YP��@y��ȋ}�JN��y������n��>~��^�em�0+�zP���� ��O�@m[z���78�|6Z8٫HYpS���+e�
�y�Ոt�FN/F爹�Ih����1�O�P!�cm���LϜ�+ &�F)�)�}�y��C���w�#�c��"�4�؝��8�J�� ��=F�q��k�2��x�,��]m��Y�(��|:������Z�G��z�ӭKO��t6g���}�g�m�yէ��c�vre<,q����
D�Zz'��\B2�ޓ"��2��*�:�1�N����1l4F.�dW�/���_ձ ���:�V��ڊk�ԵP�̅m�#��������G�kF(@���V��
�<c����?D9.�4~�.�\�+���OX��m�[1n� �h����>H̥�����2v���-;�rD���5�_cwn�
l��vd���&����a���L܍�����"��(����:pk�"���S��6Т�cMe�*��"����eu�S�ӽ(Ȍ����,*�K�����(c�5�S����"5Y�@��2G �C��	V�����fg�G�y��/N3�]+���(�1.�tm�:����F�ͬ=(�:lu>�Ɂ�Y���饚%�%��#äM���ҳ��q'�XA��譳
���Au)_?0q�[V~��������]�����2�~�J��v{r��uJ$�gG�d��Y�*/����A�E�}������]���ϽS���{��ak8.�@��b�Gx���������[)k�F� hDG�d�)�AJ�����>wu��,�Y'����+X	�mp2��_�U~��eTQr��t&~Ѿ����@'�&!gui#��
�yG�/��=���:��`P������E��QhG�I���31��>�W��SS��4I�{���Ŝ�G�?����*V�ª^~��Rx4��O+ؾ῕�~/W��cv�Y�P�s,/ic���f��9�v@���!�
pE�����
��/0*Yv��Q��P���V"5�.q�t[2U8�3�!��iFc�&-L�{w��D@}v�2W�cLܐ�\�	�]����st�[$T��|��R�u�㽹 �i����F�>q�mY}��@���Jim�>o�p��s�˿l��e�O�n׫BĶ&6��J~��"���i/���=5R��ojy���Pz_P��(I뚪pbkX��_�+��5}W�hZ%]/���*hT�$<�9/@�%�/�i�0Afm�C��J��[��cWT��B���E$�R�1����"59Gԣ�r�}�^�+���S#�>ӯ�##J����aZm��zG����R�'�g�?�ӓ��b��n_�.�;�9�tg0�3�K���k%$����"�Z�����;aVK��vW�<��R-�mi�5���X��6ےk6�2(6'���U;C� �d��:��gu��6 F���z.f*e�_���w������: ��l0_�T�S���m"Ƥ�Z*'\�r���K��ɭ�@�a��+���*��Tov�i�"��ϛ:���-e�P�2��	d�~��c� 3���a�IvĞ4jr���U��7��������~��8�j&>��AJ2��έ��î��9u)r���M�3�\@���Y5���]`��H�#��r���^]"*���h)$��w���I8��VѰ��瀣+��1���nE��SR6�U-'�yn��t8��ҋIP�m_�8p4(��]�����n{���j��+��.p: �q}�����:1+��LI����Hj�LU�Ň
// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
wcu4So49QV2Izfxj1VHZAzj4Crkkm6kspJ0JUGiThAC6+zabbSz+Q1kCEVeO9WlE
tNMIhPm4l2uLgR0Bpj25AQO+0PRP44Qe8RSz0N6EXpYDDMQjcDJONnXOXHOgzZZn
Mdbdny1i7Dre1h+fyXFIZF+rEDPEksYC90UKzB6xUzY=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 36736 )
`pragma protect data_block
XmGUs97nS3pC7HALE9AF8D+m8VyNNhmIZs8NZBK1lNvskyMMSFF5lNtmAwnR7FQa
xbjU9UrfLtDl+21YyzZdN9wI2U8DawFj73hYnO5SlbI1NFG8ZMZXbjduB6oWb+F9
Yhna9T/yEETMJorch1v44Z5QecTzpJNk66la7cGxP3d0Ibhr26dPnGXVOqqJgiZu
4DGknByu8KSe0R7orVcszRnnCGeyzxUTuhz9aHTsCU20L36rI9QOD6YQzT2HBCBg
kP5qFEYPUtqRFHLkGq0MnFCP22Dy5CrH8fd+XLjwwABHt3zopCisdTgO6vi0uMRn
zT8MV9hab8//PpqPa4KyyAYPgX40yopydSZxbeykRMpF4uYuD+UDeaak8Qg2EF6X
/2lUgKTzJZdS9DZmrodnfD299Opy+K2Tf9SQPtIpr0m4rfnkndi75cZ51QtObGxU
gY0S3g9D6yQt3zLQUOrfLQaRESzfIMWppJRkLItACoQo87NPM3p2+uh+e7o6Mw+F
cgUgG4u3cvloUPVQLnIOpQ1TJzqBFFUghLWIVTCj2KqPupe1oiK0lZfUBcgqcutW
+zIle/mA9Q56q52qKaCqL6CfqR2dXLBZ59OKW2fDP3pEF9uydDnBTDQOavVO7OwG
8oaZlQpHqdCnv6nS4fZpx0gkOozJ0jXQitA3Ck/qCdvvxF29+njK33h1NfHWwUbZ
0eeyb9+JR/lJMGaf5TR+3vQw+sxPJf0aECwieqe2ER+HW7M1ua0OknRfgP62fHa+
5y+DqRCmnyUA4Q+GidkbV1qcef/B6mSalfH1VQzUIuf2CFwzMdt2Kt1fRP5NtDSX
mXnfesBCZ4zrX9JWkqJLbZUJBLq+wneUisTSkYoNn2QjzAOH/5JdQsT1LTAX73bw
jzF5813VZFyCyoU4Z56ooQ+skwEw1gyo0YqzWIL4y7tp5mvCoYnne2wdjRVfLLGD
4LjG7Wcf9bgkvj6C0bW02xhXVX4g9bG9hvc/m5J4itJB1RHC5B7DXAjbc78oOn63
zqK78cLFxGUiG/6AKOuIwoslaJedaEi4D/5tOESKsCUHXAtfBwzn+iVu1qk3I3HG
K/lsJ8IMKoTpruJpuxZcHn3xv6GdU6la/lLl2bhCx4dy1pIhyNtsvhqsyhPI2QCd
M5d5xBWeOK1qvBIIzb+kXBct2ViD3kWTSd1PXlghzgEDsRyUhH5lbE5pijL3104i
y19V/eV1nspZ1HCyNDZzQd/fWN0nWUYUvut28DU3rA3m5LJMxy7c1GzVwC/az61t
ETzqcgy0OA+aw5YVWiHIxh9vIuef5gH7ve/eODe6Yk0mlIGQ+ekOf5D5PonBvKNR
Cv4AVy+OHh7vnlcU5JSOJk0BJpV4RVJlks4iT3V8AIwSM6RSfmGc3Zp6hLOMdULC
GvEqGZjwcYzS4kEmtiW5J2wUlDaII1V3r+Ne+AjVuAxDeyG1v7nMup+M0K2eoqvr
zPOdE7yg+B/0i88t5bAB2sj3T67gfiDfddo8bnNg+oQDQWUhZOi1Z+2BIMLsDyiU
X5M7zMWDka911SSvCtC2QdeKLc1W1K43J1ZgbxD9Du2gx7fYRanc9uL57wgbnqP8
vj01/ItMf+F295YsETFWpr3sJxLva0NQJVQGPey1uLaBgUlSYTSnavA0LpZTOHDZ
fbJ0emDspX4FiaMYEGkT78L152E8D3HfD5i0yvkFpBs8cncWDCKWqpyWTQ+ZTgyH
cE4wKtGtaE9k66Fas1GlsSv9RkHSWCdsKBqd3AummttFFBiW1mIkQcVZ5b2yzeUs
6eMYbFSS3/yq0SgWrU3KMwDl6qF66VUsy4iWLbI2o1+WO8mQ8q6CTVoR0ZOmLg0D
yDBX2WaJOQ7XHJuLmknHse+UYz10YP+4wx+ezebg/tFyubzSAAY5wxN4BLjzFlsR
MYv/i13F2ytd+FkPgnKA2Ay7r3b2eS0vjMgRYxDTzZC3cxBCh/1N9Tsn5ydvqOsT
xki9SKp+JaGZtkOAE88eMZrWaH8sVqa76fxTitlRB5NR1ERcKpwYo2LnTc5muKiQ
+Q4FGDybjXmtLfifpzXVM1Tw1f5CGUjL9st029loqYztktpx8s4TryjFNFOmIQi8
tsIgmKtMO5W9NgsWTezjj0sMQeq/sIi05+D/hW0ni3XmckJUky7k04WYFGK9cDlS
dj8d0taklEzEUm5tDfo1fwkrS8ZsAmJjmnpvpnChFO6vzSFhAH8eDYFSeK773Okc
YuWZdwOhjFErBABn4P1wDyfdIubb4Nz1PiwmlNTd/eerq/wE3Uda5gP6napKP5sN
/ms5qrGjnhqix+h4UuvJJGsdDj0t6CemOuR/qLByUZyGfcqmfFFmQJHC48DD8639
QeGOMk19u/DtjYOtCDeIQ73XiIOP/rAsUL53goD/Fr6U6FFF/ppFeoB9QSycpLUQ
MMZQFjN7IRvwGSB+3OGS3Q4hgLZod6TnVEy1P41VueXUrKH4t1sNT4L8xHdxYCQg
kGv0MPzudPeKRQSlys1e+l9TgxVSXIClnzgkVjBpUMvSQpuCKBsf0yHs/+CyobEK
WMl8eSyk//+z9SH/sRzT5ed7gHazPOqEBsYjk3MINrbgJsIG/Cw2uroSX4vI2VoD
5c794XeojqwfF6ZxmsGviU1riCipDRyqAZD1MupI/HEDuaLvsOrcDv6sItyg2u55
KvOZ6W/E6C7JQYFUwYHuJQYS0KmXm/PuFuyUOiFntMqcygzKZPhoro1kLCulDPmQ
TUbNndjOJKQ2ElBNYZx+YNY+Tt7OibSaZMIMh1DMRJiC0N03AoR36h611qhaZh4Z
3PeFD2kZ48svwlW+QPMM3Hk7azfHT34j8lThhbqLjPMZoDK3mEpXZxmoVzSzt+xy
ml83VwZBBQY2H/BxFq83cvyM9L1UuPzJpuGSClASVvwnGjBx7AGs9Ibmvjf7Sy36
B5VrpXXsJf18HAQ5pjNcg4X+GQ/bEpCGScdIRMte5cjiv338NzKGpQ13WtMrWwhW
peO3Ht/LIl4c8M7QAqHjOvu90G3LsqIreru+McajPuvUKG8RxRo4tZC8NcNiG/T+
ATT/kAj5pHs0SJd7conQRUr64Q7O3x4aXitkkocJP4+hde6Qq8RpgbLDiNBYZHwk
sU/QckrGyItmkpS60ny5T0gLpQu5e9GKLixhnR9PShH7WpK3mZWdXSKozvFrQ6kQ
hva9TzjiELvOcMz52DDQTqjd204RZ+nne5mwuvjAvALsI4uPQosA46UnF29nkvzi
vniq23dsX6CSHl1udC4fUyhPBxlayZ8NvTLhE+I39mSA5HrSpZYj094Q/t0i1vzQ
WTTQR/KWw97D0jQUQr2ZmXP2yTxi8GNaPCMUSLiVx6LkZmu18U6r8TsMPb4DDDXI
z2c7YXtZNWtFA20EYfmb0ZdvSbRyasTXC+NW7iz+Xbva/d3+NUwtL03MYlq5gT8o
++dsDp0R/wJu/o4IZ5D860LbmGDqd26/9N5FahuIkwaEicZOq5c1Us9OgMUnTnZ7
iAYQrUnc+3h/i9dJCdB82x/M3DwekmFFCLfo2qxzq1mjkBWNpOsyl9ZkralUi3T6
AWtZHW9Ur/jve7BnAbdgKrYUkiCq5MyePaJrre+ClqoVkWAt/looAk8m9h2BEmE5
KKtACzoRw4pXe6Jrro5RIi8T0X5q7FDxVyKh/Isf4duiBPCz93G2a6XN3dGL+gfJ
UfNDOiO/m3wekvqnXcm2t3GOoURpKERn44sXarvGfMg0Yay0nDJopY8n0HUm3pNv
iU/PZ1kPImta5fvw+BeOgby6vqEI1biIMZdZiIRl1YrZOXblH23V1dExT2QQJr4E
YyZfwz66kW0mp3zLTi46dWN07NiY+wzc4ZVSm8GRi3BpnlwW2T6Jtoz+Q72CroFa
aMtK55DcObN9ZNDP9CvcSxaOoywXoViJegDDnhXV756d90WPBD9SZgQXDaET3CQ4
Zwj+dnN3HzXA6u62CHNHjRj8r2uu1wDNnHGtJNMJojPsxpU2wn6Ws06Qoigq7KpZ
gbb+d89dZtzs3c7fgk6UQREJRO6s9Jikgv9LazISdNIfE4hlzCulhDA6HtHNZdvY
m3Zd2zOGu9eOd+260U57rTnKONAVcWBznanE+tE0hqIAnGEsH4iNg/fevM4K5Lro
hqxug8NdF/my4mEslY5BzYkW/lxzf7X9V3BfGAF3BEG6woK+MFLpu/9aTvpMrDyv
HTw9rSZWZMZ2hx0ZkedK0y5wdfjdqgcyDboltno8vPrORGBNKuy8AOk9ElevNYcZ
3aXIsI4NjA8Y6kGze7+xfIs7AaJ/Ktzwsc/i+ooFXwAG1o8K8p/npPMHbJFPgnMc
i+YLiQiWtcRRBvK/FXkCYnDU4TOtGNXc0SV3WJPLy0bkU5yJhhlNjNZaSkqxW5ti
m2IswG0ttKimaWg5ktUdoxsOzLvuB1z2yYQRivVAQmoj9rst93KVtWaR+e5Q+PeK
tnk4p84ZUVb9WTF1L1cDXoziIHdpk/w1KCb8qO0a4MJb16ixxqDXmsaJYeirTMEp
12+m055ljip/XF3XmMzoHBHJiPwUB6pHSyLsrZJGG1V0AGLClZk5QTra33OFTDTM
TvOa6RRgIm7tyEY2D+9ysH9wli8o0zD4UNyllbHStj9eE2XNi0BjKI9FysrAjTCC
rACy2nvqWFwzC726llQxmAT6I5yCUIbrI+yz7WV8y3Bw8nKXDVhdePJ5UfE2lY3A
ceW8qb+gmDz49hdj/Jtcv1juyyX8+ZORIpjto8ySbBxvSH4WbhJuaJp2lclUp83C
1k4u9EHTk0Wathu5C+wosIDi/g1jvKMR1XYbAQsZ8ltBvBR0IaJI/Xkk76AFy4hm
+El0Jo2/fpjLear8JmNxmkIEhHTnc5J2NaMp8DBApuHaisYdUysme5Dk2kU+NBpd
YEnj35s0ZI9EIAYd2lrimo2Z5hOm8VtkCdR8Q9x+pkwIpQwfKAA6R9Cu3haVGU2Y
JUq7g6cdAScguOxEJ2hehI9vttd0Ro5+lG4KVht355+NdlX4HZcptNGY6aP6/33+
C6kGfrNh6/tD+mjl3YQpbpQB91Gy9YVduBODMXLtn/nnP8pCyR3lN4tBh0qCSLOP
RL0WEx8AVWFeNx+euQeVLktVlRil5rzQb2QmAnk33VpZYkLUQsv6rjmeqBEaX1Fj
fDQ0fJ7zYfKiNUzSpk9KNJh0aOOsP56LTkZXhb8WnMsk2+X99v0I6PY68WQPFpLu
inhLMOXiuxLIh8CidCIYvGiP26oc34kMlIoGIAwKrKKw3v9tXbGAihtDE8bbOmst
UYKWjZBIpxGK8BErVyNclfu1T/TEai3LTvw1/YoqMWemPHhsBDxT2sWYLFbDBpZj
OPkJ7EqJCdtH+1EOMCDthmQgv6xk+Z7sPXBlUU4fue/k1J6eyOR8+e6bptjrplI4
zBE7jtahOiDwlSgE59dewzg/ijAfbM9Bk0mSbbJGrgu3JYjXiLflaC/LvvUPfJAK
oXavFTuYPEwOdRQgfqdsN+xFwm2yzgGhdQyCauJ1qDb1cMkpCTeKPTQIuwBd7nQo
zDm31xH1SoyWfRXg8okGr7FvoJu6a4jnRhjtQWe0yPdAJ8SxRVSKgcbWc5TdYLzT
M7VhyIvc1t6Eur6oebLgxm5SfTxglOcEgWaQe+HqI4Z/AtuyQQrVTz7PxcxtXjtB
Xz2sI0VHJB0pGRD6K5g4WUNXmFsaLJTmxthOKXKVi0JnuMletgoxpQ8aBT7vfy5X
1RqQueLZuS0wSnVNDkDvr/Np2BfgP4ZTZrmFICKvbQ8gV7oL0c8gBTuKFFFi9ZTq
0O9Zz2FMCy4Xg/cTcl2jXaLSi9GvmoGEKIU5oCsR917+b9v1830M7sWo0h1Zri/i
Hpg5L0JXsUpeVMdmUm0tko4x+Uw9tYbioOPKazfrD0jVi1fvASOV+Ucr7Zc9PH2n
A1dAqvYobU5thJgAYcQnDiYiECDYLHKhMs4YJl4d8jPPVD1QUGIQw+dyCXr1/erA
6MW6LxloviTA9YzfV1ou9ggYEH2G6A0YCmFjF3uob+tn1f6lJE/aVU7IvfdRL8O4
HsfrmNGGCWdwXqfF+NU48Ntf57Dti2GiaXEvNvBXtxK3QnoxZ8FP190G5PdHXtnI
OLIImGDED2y9ZFFhYMgLiBRfp8clUGjFRGCCve3j21ZWopfN0b6I1ys3xb+wGtJ9
pKtCQ4x43KOhv2pOQaciyJi/6tJs7Cd6NDP0gP99FLYv4E/ylIZoIHMBHB+gDnBu
i9c+FEnpobtYhe10IAijilSIvDC0XgwzLX00KyjHaePwAqSBYVSvPsn0RG7KVVrg
wS7Q6hGlq+xT/kUnGKYEfv6wczpFmGFLzXxorMIc9s5e9M76ZeCnspbeYYIvF052
7WW9wMxHB6/kaVG24clW2kDiTqTIRXfvDgrsszoSLL2CXkVIdYG39cNVu4Q7RNo/
Gx7xmU8J7sQ6LwmyKtNWju8i5yOiUvn402MBlCy4/2v4JWVbpSCKdpgcqg4HMGW0
+Ps2BM2/nBfsUszGh7ezcGCM4Y65JRk8gg/rPr7d/AZppj1Ei0z/vXCNlhTcFem7
pTUzGBz0sTRzVGLl61YFrXPT3vBcwGU8eeRMzRdfahT6PGc20YAy0uHlTcgyDpT6
+DFiK7O1sjuVxkmNSdwZNSwGB4PAoU0ImrS4GjosDPLV/gfOasburWaeZAQglIUA
aPrhglXZIGS/j1IQoOFyoxC/vQXBHWYRK9RozPqCcEkxQiD28z43IwlGsok6mn/l
sfiXcRoha0WkdCoy81nUrAdYA3DEPqiBP5RcH6W789fg+On3E2s2SlxIGYgSPFFp
rsgd4PSzV+7TsFFYeaCDmVpE0FWGml9+v3GhKdF3/IaWG3dVY7L0CQXRTqAZOh0y
0pb27IPaBlq0piphREJzBT4i5SI2QmtbcAlpp48gaYyP5z86HeAgiIvk7AmhDpCB
joKbt4Bv0Qb+0KtY5I0VjDMfMGXC/6kY93vG5iYb2GXkxQYixEE/trmNiwO/4KZp
VWrx8pdd4nRbY+zyiPLFkoH+xjJZvrWoq+Ao7P4xf/HJBGLEQrXGF7Mk/MCr9DK/
xKCH0wp0JoCBodWQRFGhGDhxQ5kIEwBQDnMflZ37gwUcPbckvK55GJP5MPx30gpw
7nt8oTl3b63YIExTLQApKoUuUT5RwGsnc1MCzn+9Axp4lsQUsi9rE2/JnoLN0ABI
qCQFXqSFEXodvxvATFiKdScKXLmSdW8GLcoLJ5zltD+J6zj0ebIIzvAPqcaCK/je
Y308yZHYOwAT0yjXRvLw/YH3LIBHvRsWgK9DbLEEthWHnoAdszOa+3rl7DF//Tnf
Tijws9bQwmdwtz2Bz/A6ZkFskklmNj3jSLg5KSKc7+fbebOv0s9ZUl77yTSdUPab
AouKbfUOEPvcPZwm0mgla8odevgBQOUj0YP3M8g0kDlLuVjN3BNgXbOHpamnTEti
Fa7cIHcrorCXlTbPAglng+/IT+QR0SsmQ93Sseyq0Ww+ZVfcU5GkkO7ZuXTuieuj
cWoSHtjne/fNApvncGaExnPNtuxvUcE3i05hIilIsLvIekymZHBq8Azn5qWkggyI
UVmEaxGblrh2vxqrTXefoxpLshRHaf8NoyVNdVj2DXltK9BkqIfm2Kfy3ihAXuVz
he4RZVgjIcDMQuHHWloXv0RjmobTXllNdeEqhnP1tLWkeC0YyNeT1R5r9460XMT3
iTXysHh79rS+Te+STIr1o8YcfOAJht1waQGoCNPRmuECxoA20LKXcONvdizvBFsY
rqBGAKDqqJUlcz2QmLyVnpnG4tBuSrnPKyu05gbmhLYFNrEm9UXkOKEoy3fPXvfS
wHk4/gmKN4xaemak1X+KWZ7A5tRZt1akGjID5LMD05jl++ZQZOBD293ZoV2P5vkv
IhZYRvbkFBMomsSMvmZnAQGrWvNpayF2lqi0pkPYyk9mCX0t5clq7PWYjy6haT2V
n7E5KX6rldr2wJPw9c71TVZV+IfvoSTTOTZ2zOO2k7fDd28ajI3ywNvT7GSopLz8
hg0owF+hlxj++NCXAe1+EHgQ2Tk4UTBoNAMrjHlLbgvHnXQclMr+agAX3HQJN6G5
kqB8nolmPTNtA31AufmCtZpOoSrEkbb3zT1mvs1M/PTylr7ETUC1xOH/ZIp3vEdP
alcD1u4UvvroPr3oou7MLnt94TC/aQGrV89GsTa9ZRUgg6AJFVLoRXT7OyF62UMf
mKDnagtjGpC6zicSvIPEdJyE1+5zSPhfsDeyYwVCkpNwocbQ8Jc7ZV12B1Bnqn5m
o1ZwC1El443lyjr0z3wDOfsLT1Vh+wX3Ea/BIJOb/0vqCHKl6q/ZW9VvObkOvZms
H0pUz5dew5B1v3urfi+aIc6CVDOsYYdJvUCjoiD4/6aleyKH8srcc9OBc4/qyHDF
+9JwXDaiO7ckNXy84gn20rCTb1PkDkk7dAGogumNal22qTHH+W9XjEkbhi70ww2U
2aEB3+RjQrLUba094ZRNluMtTtZo00kVvfkWSUHNDvMVhmam0NrtyEG503ZUXTq7
NyMAfVENNYuvikhHha88j4PbHW/dXyJYdMcOn74R4ry+ltDsPq7316q4ZMNxFqrB
I1AhxTV9DkBKKbw5PaVCeQuBBjTxBNsl5bgquYm2vKmf9AMPCQn4fLiNuuI1tTot
4DBlknKybexssGc0n8NdFoaTcrxqwtcCEdtKUfSNZMpPUgXY5PA85OiTmvjActzk
bZWvg9S6iniQXRqX/lEooZ9e0XMExjhdh7YXFaR+hixi7MLfAOz7L07Vzr7+oGtv
MiU2CrRSUV6ngC+OzXP35ptNZ4jxGTvxW6+1OOQ+kScp7xElKrMA146UoqpoOrlV
dLDSCKPF4PSmNDuy3tZ2Q09mk+3dr7HBDgP3PPHjSsWTRSwS0Lost8Gn7ae4z7+D
9NUXV+oMKehHJg19pJPa5wopG+rvMkhmBcWz39isntgaYyeFtAtsgEpl1JZKzwB+
hn4g07avkGOTi7dCft3HXc6OjUDs7auUuaZK82D/RxDbPi4csCpA2QxAsArBX7zy
w9adcUBud4SQinTRteJ1IT+S95HjkMkJXkARQRpPgNlYb7V4jqZjcpf4DbzLmMJ/
Xk0fyTH4BvtknwdJOS+eI92A1vHUu7gEiLr6dHyLn/V68vRnWCPft2M5ifDB+YIC
KxWbrksDoU+tMepGm+eVXAPY4XM3jpndWk5vawmDAwzf4O0H8dFITAu6JYDJxJ9q
L9yk9TtQxQwdrNOCVu/qlSkpyiPk3D8zULXGA+qgnKcz12dpgmyhHV2+x6qytQ3P
qGJaLfMzcyEPUuc+i8ENSnswNmRxt+BzutwiN1HIPHhaA8UgLbrPbD0NAWZWWa2z
DOwXaNWUed4HX8x6F9dBMi7Yi0XbXMJPG9eerK9eMBt84hoPlMGH6Nq5nJzWj/BX
DXE2a3in/C2tUnjM0sowJ68ahGKDjbZO0+CkIdkp7uQ2YJzinUs9UyaCHXrNdEDW
BQCVRw3eSaSHXAJXYeQ/YjamKCTCd2XzWP5e73mXagZBWykWwwEadXuefStCb+/M
8NTJuDkDDsCJd3l2E2ID5LJEwTayVZmu/7iPhQT0uDWuzOxky2o+xvkpYIlpSjq+
sl3fnoXwe5C1lOriUt/2NPvO43E4SSN/S5QiaE0fZxwOFwSSKGEG78PNahfM5brz
Z1mkAlys3W4QaVmyTlL2YM6LHH/T5RKhfLLOOoevxEzdnl3gQYJouv+GsNq7vS7I
pOHGpuNArv8Tynid3ixlfbu9Gkvzkuz9UYz9MOxCe1zVzdk1rwf7DcFWC6PQCfeJ
819avNFcuGhoZMSG1nfNfM9gTfu43V86D0PeoXLYf3l1f7tBL+pxRtrGlT0V6QRh
eaVTVtktRcppltt3dXZv2BNPxpn56XrnrUi4f0FW3c0KVVGjvV7tsg8dhcxaKQTt
Uq1oaeEtdivntB2JFHvvwWgME+WFvG04Qjusxa4EfjBZgb/UINAVO0vH1ddiO+KW
VDasofKQ4ChiAchx559OkR3uPSupo+Tq2z0+mHrc8jFzDds1AqOlZxdXs+4W7o4A
bEptSKgE5DaFlYKQuFGH4Xk+PoD69cUUqycR0WV9bOt3zkWg96zxAI2CTjIXHx5X
mW2iiKQ2xO8AGsfZFO+u3/ufdW2HR/QGewH3XmZ3jSiszha2MFi6RiwAGoOpJgiP
Js87XREYt0mXoaTIN/5Y1TdepWrS+f78oX2MIci/Gqi8Va4xwB3s2iBb4UuOndwC
NVilaZn8PZffW6d6dwNBQH3TVh5RTdugzUNx6vGvm/yztbxhAxrpjT5fOBNll5QM
By7aOL00rTfzHFHb/TblIA+QGihyWSY+uTG218f70dV9V1hqjAUNKi9Q1wXpXuy2
jDkS5JXSaVU+cDdMeHBRsMr2S3Uw7N2DvzOECwgBLV+Uzt89FCg8E59RVzdBZCBn
pU6A2xI6are4VEQYqNltuE9HS0GC9KW5UEuwO8iDdJqf7camn+a7yk+3MeDJcLoK
Kn7cL/jq+mm+AXYnZaGL9PzhZx41EACCDnQ/KRaGOFNRDGNIkwpuEX9R5T+ott07
+mkve+r9pIabkVjN1Ard6IzKm9WpRMorZDQAeVr66ovORsxFVSrJfp1MHwC10mtM
DC2JulBhHEi6E89HVhv/f0sMyUOT6TKx1yN4h7l774KQ8LVWAAvYExBOS3eTDdty
XtuqAozmI57SYxJN+zg5p9Yi9IVcbaJvCGRapNbExmxjEBwQbUkZ4dhgupGbmkRq
DWbbKigojsDbNT2e7AeTVz3BL68DlRRh10DsMVmdQz+KlGCN0v9eji1ZVKQXVuP0
e0Whyn+RqWHQtMIQrbyCKjTO4gEwlmJcyUvsYF55d/RMJ4x3mnDCzZz/W9aVA89i
lxI0bfx6LebtLebTvN4qsmrS3dkthhre818FrJ2Ht0v1Se5AsTWvYvtAJXCcQ1mg
6IrvpJiLoYXwBD/aeRjdHAkrcZUpj/XdnMMIlntMkYSUn7TYIFXSrwkpQ4PdRe3L
0/ne2qokaj7ZcYhVrFsrujEgMcJH6V/7sVZHqGjhTlIMTP2d6gzJZbExJ+yFaf7g
HaNtbaaV8eiCgg1DTxTZFGyo+jmDPCIhvqRdwCKcqTiN2qP/FEqzi3Ii5eOdV5tt
bGPKL0/guGoWQixFlW/HIJdn2r39Rqo+DyIR3msUCHhsilIcFw6s8WY25huz5Q3E
uwhZ9erJjeVkbb7/P32zNXQobNyBXNjOEVSoqRZ2fTwXilEdrHBSe9cSYUlXFaFp
fP3XSP5XDzKrqOtTyGeHcE9raoOogPKlbaEafcNzFiTYxkx3kXMrHqE9XvpCLKFP
OB3+VaATORV1/IN70tH26MmbyCijxiwW4ac5AXW9fGa4dYHRb+d8G+ulaM+AF93P
i9qY9S1Mo+R3PsRgWcLHJiF0JVRd+E6SCAtMRmRzK7apQBmMqGyj+jtCXt+Pf7CX
Zb/exiHblujhOUkO7XRAF43f4KoxBPhAIPkPUWQAPwtkhzzT07kt70FsV6QQmhwX
VaUXDSN2weriPzjyV4Nq0JcoJYEZq4EnlcMjoNXY/sB+ygGhsLBUWGTrokviml2n
vu8UkCPZN+2xi8oM3A6pE1Z3rO7aLsuma7dNxRxm5oFqNCtqfh6jTvD9iRw5f0aK
xPZpUqEzLR1s3QDMWNnW6mMoc6Y3YQWo9K1PstJStdpFN1P24pnAI3VfOiPsCGk7
ahZDEpX5j5y9pAuFquh2Gj4VQPai5guJ8+7LycoAvadgZ+XHJLyKdG8Xxk6PT3Z2
0crlnNZGHFQNert3fARLPe8NkWVq2v8Qukfza3q16YF/241KB8iDl23KoLpcNRpq
ileus2gV8R8Tv3Jwymcj1PohcDNmVe1M734JbKBYX5gHEnLFcKJ/IW34brDgpgAB
PVk14ExiJT8njaRz/x1dzEJ/Iu3kIAHGXODm1z9A9aGT75q7E7AO0WitWMstU+1q
sZxHvO8YA7Ir9Bgt35llWtsiNU4vMcHkAofkHlvIifPQX2KwdyKUJsN0l/XIkStB
h9DWFTnf0mUoCD2k+s3zEFgqdhbJSUhSqxarpEpFslbqRhWt5hDA+bxaQWii7Egj
mErlSq/H49qmU3YtWH1ffVLy2ll1t1Kc05NrwOsjjdp1WeC5UD0wfKUsVDO/3q9B
W/unP1ej17PspAPYaLbIBSSH/M84w5EO7wdL5qQlMUDf2XDX+ClHhLkG24RDqr5j
fji1Z7NCe0MwM1xOWEDmdXN61m/rLDxe/LreRWQ/Qv/hdq5HNqHdKTbbQ8+yCPca
vfP0STlaVeo0fBVbCLsjb9K8q864MeVYQ/Zh2nEfoMibAUSUtpqkwTIVmAEEuzYA
/sF2I4jlOcdWrRs/gefCLR/fgCKdPBkq8cQqtzuk/wJzx7vmMOQme0LlMXVODdMQ
omRJX5HsnZIxkqvCYOarujbxz/F9+zFLpzRCVFCvRfyB6iqRoUWqEQtotqU+vy6a
Bnp6PQmhDyvGe3MMsplhzWr5qq9O7gy1vQQChR6CKhDgRu0no0gTyYmcNbZqyz0I
xAkGP5OA4OQik8vv/tfCh5Yw3aBTSoqtk9CvXgYjvxAqW9reM7VE5hdvPQL73QNf
tZGuvwGytDPdmrSodyuvcuo+VgQ5tf/RmfWtUidIhGsRkJ2xApp5evqOc08qIoOC
iebwkgYQAmodejY/pWKJ62po0ozz6WR3zTmbvfzM+QE1LeVthzFofozLHsFzeUu6
zB1FLhYTuJSO5P8L97dQLPQlb5ruBRaBrQNvQIuleAUja92AJpMMxqUVc5VZxPmh
GLTohIP2lklaI2R3DcGYQa+Y9GaPn8VmEYMh9qsL+P7MwiD6LXSk8/OUueef4ry9
W4dypODuj/4mhmd8DlhxKXoHDtu0KAs8LNbBvb94MxItXS/rjMpQl4c6KQFrmEnD
hfK1oWQgXg5N3d+ZLeZSOmDOMasknQVCjdpQhj7zC08aH8RGAD3l/ygViqEaJpqh
+p4TAtTRIoWrbac0GwSK1OSQKjTXu5QEzZwvI3gxuK3IYTJzJhuhhho0/z+MNojE
Y4NWj7YoGVedvENF73J8/9ita/Vv4ysUBSVno1u2aP4EqyLxFp8UKK68ljJOZdFA
5pVk8rZvJPMcNWgyDpeNy+A+Xi1b76J3FKcAE/yV26NO/kPSCRJopCSGIAypiA38
jgrJXUHBSqiQd3Uf2yg2y34M/87vXauGWWym120Ap4RUAvbDm2+ufxgfC+dPX6jK
HUKDEX2vfg4vUq8bVckZ9IAaf8qkc2/g1a+F4xMvEt1rmkYepWZL0G+D1V3ZID0J
VbUBzR5Zdz3lhZkUVqxPsIrzXO/F6wjnnY4VLu/73yiIl3CTe5ZEgAflCn5nCG1D
r8e54+gU8hgpbzYvUlzT4WDS83duJx1aWRHXwXWk9o2R1uF70khgAV6qup83Vqeb
ihDF3stSv3jJQBaw3N1uiYNgEdeWDgsYDlB6G6V3hh71VMkefBtk2XUgUnF+f00c
Qg4i0Zba49mlM3x3ebSTZWl2Ae7ZtfQZM5z4RKQPrG1phZMPTcqMkYJdKIPAzdNH
O2v+LenqL+H2gbZwi+By5b/CD5uy+OueS/lrxse+IAJLDXRNM+zFzOnt8a7N24io
UpZK8OA2C+8LexaZOV0f23wy2UYgc8FES8uaUZVMdPE81mWG3zj+43gD70BbjRpC
43Hey9iGt4EykFw4sd/xhwG8+Uf8QnXhU6h0RfXLE3ULgOmaSb7cwRiUURVWlFKZ
fMO4MLAin4sHGML3DEZLOYJZqHfdwvnAq+tTTAI3HB9edVqS8ocQi67wa4G+JgZe
Ub7e8YibtHA4Ur76hyF0Lkxe+0Ql5A1aKofqOzpFBljhyp3qfOuhdpYn0E2u4AY2
et8jObFbelxMOjHJ8JYSTB7U7sBgkkg+vsW/Cxag3lv6b89v1afYovbyW1iztgc3
u45/7zyjfbtVe36ac1SuHQp4bUfLrL3iYiaf5kYxCLEsyk5Wj1ItiHWOcrrxiIo+
p6N9G5zRe1qOHRS8llusPi/JkHj2SU1h8dlG7FgmBX/2QWVTcOAtwkGY+CYAdXcG
TA/yyq/Yccny8Q8vO5j/sgxzNDHybREQzgsoBpHLUZbdNwXtwIVdLFtgJAAHSPv3
PDcUr5uURvGrclNDH0rHHUGe20rZRP54ARplfy/vPB/4F+vfDwdD5545zU2YDrNr
7Oh+UfVngbL7NXa6hYBNxo5/HR1fl9+KX/qhBgoMOkVcf+nfq29rY8QGovzDGImN
aZWALhxCJXBDJsx47siREztt3rjLvQ1ixLOCim4km5xey/X28ef36+5UP8YaSPZ4
17csUiGLdq0Kuvs+Js7pl5u2mYZyq2m1h3w2Qz38xIK7Cq1ONO1sMNNg8DZYGMw0
I5RWNRPX+mlXq6QXu4hyQ1WO/+9QLYjnA+mVDrHo3V8nEH73zVzOc6jc2G2pA7DB
v4HlwKqOc8Nh68zhtArK1KPj7jTF9o14ODj+v7kESqkfBZWeW5LcOty7kibOJT3I
2YgXbz870xErE7N+AiHbGJeFc99PzD2dNR0fGztx7HIiA2hbYjaA1ACqn1Jl/Ak2
IGadk8gq65i/TKvO5WQax1SzZP+xMA/nlfsgKTMlrtRmnxdPuyYFODZeNjo54vml
tl6De/UQp5gI6lzAtLyJ45SjaJcgy4WBZ6P7ovD8+q4U0LuvoZNaAJGEhcDluDVZ
EgGtFVrPFcupirfblGEOxyZnYUZ2uAlOk63ZEQPcnmTi+9Wa0Jz7q6MqEGb0R3XN
Yq0WLMBfUmNr+BJb+iRyfAxklNZc3wa/hpINhNBsSx/L9gkygRztvocgl08Oh6FL
3M/XA1l1ryxutUuyl/jvGTdmQpVvjM/OCm7XwniQ+Ou1hVnYBoL1I5QDckttKBoG
Kt+e/YeMqqCzJj0e2K5gOKdzAMer4J6MgyhvpLV0+m70BvUhoR5sRR0q04qFXZWp
ymqsjrosn6A3PBZadaP3ACzSrG0HFKjDuCQD+qL/K1wuEGGf/97WPV8OhPYeFG+n
QCetdgXWZE9Hgt2TjzqekRt70RjFhLCWUZD8lbUPo9vGkvIBtrZCyWQiaGlnu31c
LOlCHwmgR9QT1wsURugxTRsy1QEu6OiUhr6910frf66T4lj3ToYw+StOG317EUoE
jm/MTcurC9lcda/jpMb1hSizJWH+PDdRlsbEUI0SvYMvZN5SloI5QJE5nDNHNnbN
0PNEyOI7oE5EcWqT2O516R7CJ2ZOmlKauKQtRXzAlHW0DNA9Slq+lDt8GnmIpxFe
AmxfqajFWd8NvWgfFnxISN3vM3BhIrl4jBD75xT67E8yg919E6eHSyxKsgfV3odu
bcSpKTxgAiL/xBcAEJ97NqAn2va3QhcPOjr1raIjhtrVd3Bbo7FuUcXldV8XXzYJ
cvyHjREliqJ58HGy+1TyW1SSsqMNoE8kkvcWTMWs2O7cLvd/+hufRlln9yYYJuz4
nRXuxSLXg5vaQ0ZBSRYWHVdWSpSaDFTRWD+IX6OC79/pgKBHrsZ9CPXAtlbEtKce
5JVolRNkpQlbKXPSfVoHq9GQSd1yLSGrGR9ue6vggeKfLIOXVTHoIa+mxPAYzafG
Di8k5IpZN0cQTeKRmThMgMdTklYKDFe3sTIaTSun3n3yt9h8Qa2wwomL3gxraWyw
Pfzj6cfx0kyRJn3zR+U9B/SevJh9vdsdAUqSwhtwypjT1d0WNiSZUEJDbtbY+OrI
vO+rkLUd7jzz9yNIgUXc59fx/hiiNXj/gb25aFkj1OTMjjJOdFR7RgkrgWt4VXwn
aLuvJFiEQVGnQKJbR++EnPffpzdYVDUNaIC6ho7CyhhowH0RSzjUj/LgjJlkSwD3
FZt9UIsneBq/VzAqDZssZqFoRcSHPfz2C5b4oogJSfrnDPq7BrzxG4DrXXp7d+NG
Dw439+UVsKXtl6gEezff/NWXjjPiGGNaiNer/cRv3vB0nop/tGVIqt2HQ3+MLD45
UNIlaYDegE6iLNZPk+zgenfclkzKkVOz0OutW/lRl4EJXrxpzKZ4aMhyoXBtBTD3
CZ+qRN0yeDJ0jMzs7lJbkLEyiGztVXS/Cu7OdU9SxJ1DFrVPNhuIQEjv+SgiRUCU
NgsWBHDDsigtBL72Az+6SHUe85nlf8zN86PEQ0yGqI9f+PSDX9MQFXZ05zH9By7t
MRQ30cA6Q6KwLrgrHhEcm9v8pLpugkJWAQs3RH/fnhmNSWhTbzTi5RoICgh3S39O
i7RkkGyzc+IIvUpITR/7H6zeipGkztrvJ0Tzx9QcOHfbcbm5mkEkOzfNhV4TcIRW
DpcN8g6rJoRZZn2CpGb9kaDulBCG1T0IY3LjSBH0z8VYrvIQ6bk52L3zyuNaKdDK
hQ4RYNaOUY+Q+Oq5Z/17oCjRyHUibjINeDjWkyawCNBcVamFgAqmt2gpVkwP5Kw/
vMZ+UBXM69h/XIYTl47bzt8/Jx37Wj97AG512+YgSCLUfly6xbkA1mIhiNykDwHM
TyM3WRTtKVlUq0eBDdnaU85EhYmGsp43QmJMl1vaTGtTgw1Lz9oaxf0/aPuIYOTr
wNru5jXDlHN9nKVivhuyZ4k8bOQ6475PdRjtd+zHCkmxZxpaH11ykEQKmPSkZ9B1
si581i6uizc4Qt34WzIJKZ6gb4u8GfVHxsbKutt0SthGUkLTwXFKHRDaXtpxa1VB
jDeilSpAJNbpyXsNCkSKbdazw4ZrNSHoSA6dPBvcbZFt53V+9fF9noBfsJHD/ww8
pnyT5QfakIbqyqIC1onuX+Rk9jW7Lp7KQtQwmY/SF3Xj8QbOuQd+8M5X1141QbVZ
m8ULExysTKn6XKVTrZIMCk8aRvLlI/WxXofo8ZSX0stlsNEtI//Fv4KyXirsbjeL
xUdlCbMtnW/hHVdhiXWlWvRfJL6zpCGk2vxzBtunHjK4PchTKhgVqNrYdeNeN/Va
2mBEBCSfE8tN0GaKGgLGP//EteYf4i7wv33h6AB/NwPqmkCO+ufZHJ1beywFWHVr
rHFObjb2s93ZFBlZB77alkQEZ+tIo9Al14pfRhJUnAPh6DHtUpInjZlpyWVLf8R5
F4ABYlSUwOyQPyLNfG765L3VkjhluNQVVLGg2TGcC1QUnA62Dz7WkXT5K6qi2qtj
9BEgyaqBltXAfMFMsKDcbTJuHdxuUTUE/PElvnwf9qHq07A+U0rLKycRy0WfUp01
aCrajvohzjHzVknUw51UyjOAMaT5gME2HUYGMwvLSq/LhBx2zKnMTX0cys6zs+Ns
+9lGqWkmF2sbKY3RWtI6+kSwxraSyzAAGjsTiL98PgT6UyvgJGIuMp/3FAKxXBh6
9erNtCv1QCDZgqQXvdR5yVvNXfuNN2nD/8UPpG7lm57EozdargI4RQi8pacmVKrn
aynGL6Pg2LbGTKNsUovUBoYkHDLQZWwyWcT0Ghjyjqa7zTZZcLpxn4vkaYKcF0Og
MUw8yGj3m8DYenqzEk1v5OdAyy4NL4TvctssJNBq8DfIE3PqAaDtXuUbsMdBfQpT
LgugK4rKwf19yB6g3NnUy5ZSzTukGlKzGKJK5GJPNnCvlRwvw5LFIlIZKACLbXjx
kaQMOvofSzu2tjJgbx21C+n1/QOxQ2sOdGFquCvXFZ2hmjJ89XxYPmJPJVFkz32t
eJtcc9UTNk2qJYWdm8xf9K4GeIMceWcwKcI0sjZW6cczMJHKDgtLSMt99oKlyBNT
+CWI8NYSCabtrnbQelbsDCVAoFxTsvexP5f7soRDz3k+MMQnPIBbUrF6t+GL46Fp
xHKWKSC0SOouR6pI99bXcqxTxVFBnFJiuVcycPcaWYTvUrFKGqd8vY443hrH7y5D
+JOEvc7GDeNkev1QO7kavV9gzdVYGecH0qJAURWoxSzuiGrHTRUrCCY8sowdwu4P
klJ4j58RLWej38/kByBrUzpOvRu7HUo0P+aHIAvjf5E96zMrnuKVjGzCZ+62R6f9
H8lUpgv2dqmMncWyV234KOE2t/k5ehIf104PHp5cWR9UduDYLR3bZtPaSjzL935d
ttOtewTDLpJtgKH85E2sp6erT5G2TJEjDsPRMn3ZtOr7lejhyLmvd+LidcBRZnOK
nAFHDZgp117aVHbC4Z/4RRn+ALBhv/Z97gZO/otDaWNyrjNWvhUb5BwPa5osmN8M
eC9RSAuYQwjobZCvYmrVV1Qf5yQIUmvNSkTPXDBDyh834NT+3VpcD32XMjAp9aqE
DwZjpEyMufumyaovofxKH4gFZwClsNMqnFCWGwjRu9Dr//mS81yOtslYJa5vGhZ/
/NkO7ZOPU5XSGf3nX/G8CFPOLIVEwV9l7qw67epYhSjtA8wYbUmHwAtLVccnQIMS
hfy4PAKXsZWIN4iVV2cdp5YcvwrGer1Vj4s5kMVLrFFHSUY0OHRHmboCAPxPgii0
wkSdlL3lhpMiPkz8OjypIq0QHvxsI7NOwmhTzabyI+J3QfNJzesmBPGWXW2CbXUL
PvK84IO0tvpe7OHvM/OtI194kFTji4gMjM8M1UFzq8O50hcsI2uBcIXhRKJefBPO
1p0q6gqcOz+tlfkLD+2tifafne7W/Xzj6g4lHIY5rQiCkOinW3vG5VXW7T15QVjP
T7AFaF97Jm6wDIUV2B+QtL21RjyTKJf+ac7kbyewwubz+xc34TbUQ+6Cgkcv78pB
+j3IRxRISEaSe0C6jprSe0xv364d7rMLl4nPISAPYPFgJf/IRYtiIMQmleij14kY
VYWOcqwPuaBzdAbVuxRBDZjL+ZHkewkrmSbFqACb7UZ/QGkrbu4xCFimO363lkby
TQrReT8k2PpcXV/LMFszcfdud1NKOL4cXZKmuzVmmwTc8O6cXJKEJGQtf2wAmPwF
VdYO+It1Zw0VSd83F+Pl5vWBemaaf6bJUpRpPF+2UCfAtLJVmFHo35NHx4qkLyyg
L02OsZ6I1BF0lGCkLDeZEi/W5LxbWFFmXebcBJ3y43XsI3cMt3OIGDAaSmKCydFT
F5xNFD3WIU8so3UjhaxIJG4Kq3DzGYK/Fhu/cqpWKylkFootdtxHBpo9ygKstTgp
pGg36qoQGpqd8x/cdPvfFVvJD9uncAu0MVx/Qyb9dcjLGNkoFVhpcCSJqMa366hg
NmVmO3+/wnEUgay7WmSelcPTrqfjLriBb+vTcFESrjsX+wZrIhOk1fm3ZeKVZ8dU
EZLK2n14jgTVm0WQNa9OiXTuilJCByv8RFOHSKdpInoLwiR88mMgkcssxYIpPeHN
/T0Axk8G89ssDQH0shjvtX5u+66NBQPXBHn0K/hszSLATmYV617lv7I8VfQ+tBIm
9wnrsCqvJVWo0EBxQs/IDNxXJ1LYIjfPOFtd0mlbkH5mzLEzTYRLw2vLmYJCb6Hb
6Tji9Tf8iSTkrfojbR2wRbJBhW3gjRa6f2bK9xKQ89BmAbrcMTJgCWA4SZ0h1ONM
bh0a0MIpMQreJk3MUMZiA+R238gk19HU+DUqmVjcXhrm35EScw1hQzK+jP2Wd4ED
vj2c8MdjuTJoik8/6w1HCrJEFC3fGzAV0h4HbauQrtdS8/ydjonhrJH5R+UNSHdu
4OCznQjg2vRPAI/0J3TSopKwoVLfFYNH7Ttgw2C/tK7GSddbuhq2oc1ufQy5ouM0
UsJEjzqnZOtMHfaR3IKlxvL1AXOqiRHdlXPQIed/+ykCeHaHwNcq6fQfw8nV3aVt
rNIBpndG6ePCzBOVHO6rzcE1bZKyeLspPDAoUuLWVlQRyqi+k3CbtLQQ56pmgS7n
FJqYT+z9DpmBM8a0E1AD2GvzCBihAiuT9psv/3DloVNPHABjL0v5XIrY0PdDMqiL
WXhtUJ2QeQHcNdTrCX38t2jpkyisNSpauaKD7h6k0AEoGl20helpizSjH3pxr+WK
ng4SJTI7YiVJPNGsoyeXvff2PReft4vcq51TfZGBBTPC5A3Fbg/bgL32mnKN/Zgr
2JNevUPgiIEMWEWfU2kI3wMGNqLUKrmUbm4xoPEm3x4iB6o/GvTQYPfE7gL+SQcx
FvYAw5HUOxMcTb4TEADU5eH2/AgshA2kXxVGaE+qkJsCn8dKVY3qhtW8BjoH2+vX
bhBiSX/n9iYukSlmX4A/H+shrjyq8h/+jRz7sGTovVd+rZLd0+ZO17aI1BdKfhQ3
rYzNk1c/+ioOSfUNgIKiwv4ZUQgiNZb3UFdrm08bnJdjHSoCkjY8/t8lcw5wapoo
VRgf8XmyHnx5GXtl5MhYM6FJylhyl7rg4H76nsbbrlFUa6J4uDMFaJYtUM4PcYRV
Tc9e7yCC8EnUrFmJShR8zDh4QgzB2Axe9PZDryR0W0thTNmf5DS24g7X36fDqDC+
JbAujAAvx0a+dXRPgQW+uJ08cRGOVyIsUILEoBdsrSeON2wEV0cAvCYTv5NMLpWn
kKUGUhALnlKIVPmfITLeeCEms7MsEUso0idx/xkfTHdLnOYQF3q4RmmbMPx1qsrV
WzQxaE8kzw7SWJuviALcxrUZ4Mz+JOt5MwkbRGvzzmJlafXEuAf1OF/tNZaGi0B7
x3bmS43p2/HGxcmXLXWRTBCABPKQUgZVf4oMQegbhOUGupLiWFim6BjlnXnYXWym
qBUf/NBYD+lBmsYw1gV4Isq11qLiSCKvc/R5d/IPJ0OiemK/AY2TpGmxnx4WQjkx
h8kaSjc+XGljsNMBgbv598PbzuRZt8Sbk9IQ6UpLVt2IOJ/lSrtlbruqkZCdqDGW
+RMwkE/kbBcNBYCkUEDdHuRWV6DClqd6S9jJ9Gkj7Ykm6vZzICbi56h3nWsRzzjY
2W5ypB1LZQBSZ6P0K4PpiZkzX8ZrEKe5BPT6iZnzDzGwK386PEIIth7qyGpVxSel
/qunfwSEvyQ/TAFZE4+tB7Q4nB3SLeIdGli5rHnmAMhhqDgRN0+yhkP7t8r6QQ9i
sltZiCUMlw3UuWcLpRKX6HAgS/accUF5iL2GmmU3BydfeKYWUj4Mfp88ir8oLp8Z
v5akeh/sVgR+v7gtK0Q7agKqETjJ/e8Jrh+c0KgbVtE0flTDbgkoMJKOjg4OI9eq
7q4iCK9USJ/yBO8YtZM9VlqUFqSHQfC77E4nM+wfHvg8Xchg53P0Fn+39xnz8JkO
XehZVxJJQcPUee6oxLjsHiVlTUoJVJVEaT+DkGRsN1AGYztuwXhLeuoFbkKRtJzo
BwXkbVVRGwrabTdhq0C2Lb7VH5s89Zb1qXxAh4xrAvVF1CoX/+G1/hmE6W4vWIRO
FhkE2qdWKxeipPaR7iUvFl0/i0MSkKjoc3ePlE8Nj8MUh5pynhgpYQXzORIA8n5T
MdtF0hq/fwJf1hQB7h+pmfC3l6m1ZwpRwXo49MlhuSfzbLKDS9af7S73dRhfuHti
SQq1T7BFjpQn1bjeB/Qr3AfSkXWZO5kCOCSW4cC3gL/qdJPay4JmBslMUWvKJYfd
YOvjNXj7vgRRVj08s4fZzU9BWrRWjoBe2/OUh4sRQGgK7EgtyKiEgOCtnsp4jdN9
RXVqcMnF7O78OcVf+xk5XTERVk6RpgtUss8xZqFH/+Ar+YSHdufdG59VMotq0SYQ
/crggt0z1TE4DiMYbA5TKzTehzHcO5KOEdMuN8xLCHl1oNQknyRQRvyPC/RnU6K+
LAdh5aa5e+LhuAiGyobqiTjpE/0silFht75WW73n7BZ7/eUbfkk625k8wmkIGMTE
AHVRELcbaAOXyOOrSzJHpVn+77bPqaSqAcv8wgHwQVJpQbx0wKfdd/EO0RRfiWUK
YxeL3g2E2I/1gv0nIGaVDMLSba3Dd1ManwUzOBdYQyz1cLGcBIa6X4z/dq8uZH59
rLlAi4lklrehxV81yDTkflW+TC2XfM5zNOy/DJE48oGgI73OMPinjkf9pXC7lCVk
I1HV3gIAONKEuqDnvjtqetznFcV5DIwLuhgGlNQWPaAC1fkbvsL5Dd5+4qt2bF6H
4KY8GNwDLGdcC7btZlpDCzsuBd8DsWpA84pm1XnDriDOcAvFOosn3Xqe7YldyEYy
FOZZueVEXb3xHNu0B2qdeIt18FgQnRcBhQP6EMxpjEoQNZklUNjE56P5ym5uNrcQ
nxNHQZGSbKz1A2qsEhqL2YmqDLb8Cc8bLgYiz33Pj0Kv4N+wvPm2kbYFiHT+YWwE
PBRxrdh4eWiD38TsF5KjaMp4VevzQOXjIcTusc9FyRI/CqdCe4Ge1E/7jhwoStWb
OEOnN2yGvWbz3MVDVzWS7euqg8mwxxq7JVV5/n3F5WnS1GrxtmkzTWvWjqdHlb4s
Hao8IjZEqv3LfNbGQUtqvoGjQzpCkvMUnIvlBZpXUMlubfRsvnvcshto74WiCcgM
VXOFnVsXo2EpSlGLEeLpyF6sclPeaUAMLtdtaHCAtgsNCU2+SM+J+k7B6yTdlLzY
ovSQkKzvsUY1AGqTuhPylGVXaF4ZuKQat6FBSIsnjkkeMVxRFBN56cJgrQqOBe8Y
YfdzOFbg/9q9iNBND3GSN68QiZC+WtA+CO3C8hOUINrcmMolKIjDxni+FjyJWtcJ
j6eMT04a3UL4s/qbZnhCMNsN6ExDv2J67qZgFK6WFGCTXitmSL7nbJ2qDPkODMNU
k3VwTkadf18dxxbgwkWoFDFdBKbkzP86HmXWp2f9g2ckx5Y0PnORTnpUbita3PXB
1GLfTH3UjQ+Eu02CE6x5gVaPzuLlUvMLyKV2MUoxLqgTDVtK988F5yxlO9n1VcaV
OE9ocW8nsmCNyB9H3uB8Kr0QKccRvboZzbLapBxl0+dT2NvWp5sP//OGwR4mljPL
HDpgLa7/1lB1MSKr/nQPiVfrJTw4fGjTV5bFmQcVRPknIXsDWO0YOgwa4cVsEohr
+v7PUpR9TD91WO0Yt2nFOJDPxc8/rRnaegbcQR72fplav4Mq5BPwDYY3VFcoVmjG
MxpnfTTVu5QZKn/44qA+mXKiitQc0wbWs9LzgZNlBnd8vk8qRw5HjfCa2IRduKzP
Xq48k0eA+8qa8oT9H8yqrBSltOVhHNWx0yOlU4iL4vyRMfpEwuQ1k85/6+ARvq54
IXDzNgBrXutmfGQfmOrHwOIZMp4cxUNA2UCB9lyGdErlPs6SxzrYjMyldlg8dcQE
JiSDkqj9edrzKslzwgrzXe3CPUEYvfhUB76OQwuM83+Q1mhZVcXYLN2rbj+TL6Su
3cnW3AT+wydE35YJSCoTHL2x1DM4CV+P4MCQGEVCxUIHwy3EsqUY1+txvEfrdLc7
jIjw2Pd6SjwRtfBzSq1mKJOQrmlnjY1uxmCzhEqtUdVucwmOfOz0Hzblx1JDKXCs
r8nZz1IW4fm6kdqiwUHwZtKwLKL/jscpg6zA4dW3TQbg14ksogGEBWfg6gl8SmDR
6V6rFUVygnAKvnHM0kH8ycFyfUNHcc7FNo/yKgYEQ2hnh7uoDh2H+SQnojfl6CRt
fZfF170sddLoHdJs1oc5GIKD+wJtW2pW+PWjVsDodDdyRSRZvrLN7/C6+TSCvhuW
bt9xc9sfl5520EUXS/g6ocdgOb/4p4nIsal1Hbx6q7X6Nj7VcN1NpeFS2480gs46
KpKKRRVXkIy+owTj9CXkx5moMDehHGNHkqHWIZNzLBHPVoTJam3yulIVbaO8T3bo
HhPtocJRcLvvCrosMLo+DahkvuBEqc5SsiC95GQFfNaIut72zL/Y+gUoX4uPa+jK
MmEa15JPFHP/DRPKDmJjHgOxF5D8vX1bq6i9ae+RoFAxoI6+0AenKu65IuIOjutK
0PKH2JgAL2xrqq7YLU3dPYjC77l6IFL4VPQ2cKAyxXDF4qprsyUEcq4MY37hoMU3
vkliT68oNBJLA8b+OOsXSvapCRbNmPsLJIPUrPHYoxi9Fi02qerpLNaNHErDqTT9
w5QQcI4iEHrXkxh0Da2wtUjYBeHcQ4P3Hc3rBq0ozZVCcx1XiOju5mjrowIj97TW
vXa5cRVNXsOT8mByvbi8w4iB6FJtdwEllRjZxT6sGuDHYxbN7FmQrbe1iioZJHGP
wSIx++qbp8q+XY4dUExYzuOD5P+hFN+caG9tuRKR3o5kV+Kd1o8dugF5pXObTEo5
Zu60BEzJ9rO1cwcVicopGt6yzjvpsgfru6WIKsXOPDcxTbpr/6KPGzw4HjASAmeX
kNmcPiSE9zX/teQR1GyjpcdI2DDenrGW2kHxtVVfLGhg799LWOaVEZRfEWOWHxyu
PpX2XjTvK5bwIPxGHq7VhP1q429cQgLidOlNjmpkNAPKyYfxynES2buAH/ZgPN3a
LXEmcYF2qYjPBd5i8WpR4/smiy2K8UWu7nMpgIfpRYuRmrdp5XkLEf6a6x7XX9VR
yHCgedPClYKonGPxALDD17AhVNN9lu6nHSP4lxy5KM2dWGhXE0clsrlLMk5N6HKN
7ivWEzDnyNnciKDKcaKShOkfQ0sz06MOqzYYTppunIctDdENU/IpmsiTXAY4GPWA
yZlx+evdScsmKArJacxgOY2dww+IaWBEMbWbaNwiWRUf4cyb82T62VTkeWrM3oo/
EPpJErMBwNlnirX+lTHNyn9w4tADa5tLm3xVdFf/icngWHBWjGBIr6U4So5ZoxCv
CkeBkFTiYqHZZ3S83TSThIcJOKjZINqf/o9JMcZbsjVr+ZLEy6M/OCtZzUm9VZsx
014LJsELST192/VXTVALXTRZsXYXIAOQ24wRDwIz4pu/o54MqXEDwMUGUYGIOh45
ORaiuxog1KUztbEX8cLx5GOx5Aza9mFSDrYCcpDzcdM3+pPHyDxwkcnVQUyWWyTM
7w1fbLRirgUoxDQC3CnuNk0VzjboRh9OsXD1ZZe95IqRi1TZugt1+YIWxt1MFyKX
TrMazmszhvxC6M/X6CJsWT61v+HmpRzloPIVfAAS/DR2GxXPsTgP+iPmteQWgeTV
T320kB/5zJOcOR6bUXnEGoGF99kfvx3RA3LL2kCBU7tYKhKIlpqRnxVE89RgMyYZ
07VeTbDB9whmZwhVrrVw54ps2ZGfUFIrRdJqg48cAWRFkQUdSTFFvDA2bfjiH/de
nPcbpGnHn5l1LYRXkstCYBnuLRBe5g8MTJ9p/lt4knYBfHuYl5mt2TmWwTDHUlH4
yvkExmMGeF71EwsYN9nNndR+3YXzJSJKFue7w6rbAs600CkW6gI4fgjkRLF3eBYi
ekTdy0SwIT8aIqqGmbAf8mv6GHN9tZ2ZyAEKQGk6VRCWfcIRFNH7BxhOmRdkHF2z
I5Kw9SGetWpGmTJ68qLa+Pyaaea+E42uXwq6ZtBsMXHjcu1st9d3OXFcXoR/jt1k
94AUqIC8WHfowOHMXdxqc7ceLg1kuxEp6j+dSp9s3ss+soY6SgVCdAKADfXjtX6g
Nr1X1/M2xNiVXTgFnZU8CbNQbjtTcnFO0V6rACYdIrHnbISnHtyR15LCUyYw96na
g8g4krNrracemlaAvtdzru06UEqByk7ebZAthge9lyIviiqABC0CNNRvCla1Tahb
qvy5Qnp8LnRqKo1uQ3NYgUEHfnZeimjJO/piq0TVHWAuhvx7704HzAWpGMFfTzQw
+sK98f+cyEDhMXnMzyEt+6DTS/vfebSQlBgcvzA/IJ353zh073BigrrhZxlfKWuC
st+TAxDpLl5izpg5V3ZxNR614VFYGEzYZ3GjtyoFaUmNDLsjDtp/RHgUlV72NnQH
ur1PSKq3u4m38E6v4xDSZ6POZbbqzwa6036+/vulIDYDB9PmwDla8G8EcuaQinB6
qpiCwfvEAiK9yzbObmNJyTXVd48Uu6Vj6FW06m895LJKDptmjp5xGW5oiP7wN0r8
w6kjhFAt8CmQh6f4in+JLvHxW3OYS7BoelfuIThadNY32oo0JZcyneudsscMKnY6
tF5APJ6ezB27NQcfG77u2BLa40RNI0fYh+kl4hlO1z7n7Y8DByC8dySOHzHXpJIN
BFhq/hLpytTeUmNC+C1rj/iGVQJLcZ0yaokyKu2PbYfkzUOhilRWeMknkYjsWNf4
RVpFCxHteTYKVUUrUDdNdgKS+f/mcY+DWq6GAhAyZzt/32bldvZNrOKq9hZmgZ1a
/nwpEzUV4HI4rvYdA65B9ta3q1GOzZtGRmLHRowaq7JNFwfo4dIZKWkQbDrNl/zj
a57VrvSUbE5L5bsSMKaMaby55Rrh05b96Z0SvtH2JQwF9S7UtiabCoAF7xsFhRvq
hz9YOlNRTVQaGvWkyxrm/byZMhPRf6IPkhbDAD1qk1MuZMbO0gusmbDwfLw1LAHc
qoz6qdbDJcc/3bwDlchrFR/bXPPaM0vGF4kUr1XeykAH9uzDNzZp3xETUkhJh3HT
Mi2wEsjxoD5JG5/E9RXaVbuu4FSLnlek0OCt4LiGuJECrkE5ITvPPi0gGyDTb0Qp
c1r14I6HTgqoxRZNgBYbDfCZioLAPY/ISZCa/tVtKh3eZfarbyXdyEy0x6nUgJL4
ZwjDppslOskDoiTtdi8obqpyfAgDstH6c5c6iZp6L0cE0sPhplkYkXGk0OF/TqHK
RZBMDIH8dyR4z0un1fBOSiSP4upKY0RPvcT77jfuSBV7AS1id2XpFeBCd5vpqgeV
OkcoMZG1cp3UGYNd+3K+lS2RfnTWKySiTYuLly82QmFP26KN9I1w7WAWsggbvRZy
UkCxpYTRUNCON99qsFnXHUGHS73flEcQukr3JG2ZCUewuV8ixSh/BfWNxvKdOQ6D
LsEXjC+pLez5SeDAH4NxffHVR/q1bab8/77AfsRGkaVlVpLE7DduLYRRr5Z+Ta0G
GowxZ5ktnrDuewVdlvAYj5fS+mxU8jmv+RZKkoTKW7L1YjYANt08pR4oAZh1LRTJ
xBNr0sHAxFi0yG1Ch47vq7GTpQ3MEcgZraHUKrxLIidR+oce6276MJ+9Qpt2b8Hi
4Kf6biqe8uow4Y4ycRn360tFJ7j4r3XUU0ImJ/Uduj/kDEyES17+wbhh1YbLSBkE
4IZ6n1JFIJLAg/L2U7vwAF2dbu3n7nf0vutSrpeLJt/xc1NyEnC0WMQtDDBy5Ui9
wP5ZcBsvJ5k6wWdD2isjluhMkSK4Xs677EZ8fEWAWiFekIUJf8NFkKfjJcDSczAj
CtlznKKvRjtoovUDkoIycNUSYlLsRaEOR9RPORwbwLzD3eMeNgXjJDG/xMmS1p9Y
/VrRuHGtLvgDX5Z0eykcNrjMLyqp7S13zsw3xMx/xPDcerPSA1LVDoW8qOiGsck4
fh8KQGEgVe7Y0tQWEgAg0C1Pw9i4ESIIH/CmgwlP73rCY/uAd3R1sLuySUWAHSCq
2a8lpg/xBdrZgBSb9ecR47bw2HwEFTe4rKhInTX8hmSB0KOsQfeiZ05v3KZYxmyo
4phkYQP44zRlrqU8XeuVqF3qX101W8lDUbZdbOzDVuv4j1nLVYg5YeOvmsjTwCBj
LzzhttK+XtfRVLvAGCxLe1u7WEMFcjP8mVWYGv7qczkWugh4v4TMwXSjeaqLHx1z
fA1YjwQp48LodnS7rz/JqX///oYfz8yiKwiWE9BC5UTIRuahlpIKa8mncw41+Yuf
NV0My8bkYXPzpLHvBFt0sXMjKg2SuO++EuThByRzPxAac1hDrC5ScKMsJw+7YE/I
rzELJWaCdCBhJXwK9dF1xLsDNXHrtmB9DwLCNgFjS/TQnCZHl3yq3m+LwABfmJnC
hRJemNtZIA7rcT6GXu6jZ63Qna1H7u1esH1rsglplMVXvz0wZKwKOokwD4LF/lI8
PJR7BfKSO6sWr6rwkMM17zKE3RxzNzbTrTWfsleYTjxxrbVjEa1lsMCdM00F4qpA
IzbKX8jcZjpMEEl8rHnA8wDpibmG7ojscKQrT+zkzje4hS/3vud/h/mlpgyDfr4g
DllpDKhioBHvxXrHztoCMsU1VdK+poqtaCL2YUefdFKlBqX+Z1OFjzthYnOCkQH4
djlYi3OEgixSp9P8Cx2593msd18T56c54FHlnFv/4zebhjfXcRKWoSglBFMxgmga
fXT2lgm4MHMiToy9WH9gN/blMsCnplprHMj1ZA0AY+8/PzPVAF/kq0bLlN1iy+E1
iwmhcyJJlcaoS2K9TTDLAot2f7ljI9uk2pmT1Tnv5Nz+lRlAi5/+RMnXm2vd19h9
JmZGv0CLwJK+H7R+WD8GMzHy0RvtUR4XH8idjoQGS3/LFXPOIahaHdTjrrdthTF7
FamIQNuMzpdnDX84g4d2PG49iddvLcHP6ltJssGZMIX+IoXJBqROFL2mhyD4CJl6
/9wlQskQxTdaNw5LYT8PXtAEvdnfcgzpRcywhPnmegyheLEXoMs37g+MTXaRVK8s
jdxEKldzGrhLQ4MEdVvoW08oinQdRo3DXkE38ehxplINf9XC/F6CTifQ1t9jb5de
moq4SvRTh0xrPuFdWiwqNkItD3O0ZK37mwLAwjFYc1AuKYFoMG4pcEaQbhcO4UH6
06GooQjDj6CaRYZTlbjIZ5jOOGfDd3P29CKJsdl40cNdiy2QQgPzx6JkHRn4pvob
sKjZQAXKDh+7SmYi6aoN0lVhku0pirZiT07QkGiMbUShVWy+YQzL+nZ5swKH+SP5
NGBPOC+dsgUgeE9649O8/XwC3MBknFP44fdV1g5y0NktqRJlRIbxVWjEz1NPksnT
FeEFkQYPo3xHzpvrvAFE9B1yZyX1Rxm9inZ9/qWxaV5zdI1qAYr/IZgRt/utuBdY
nOk0n81S6NBOoF1wgDF4+gsKVRLH6+8pQzfeoWBT5F6fgNcgsXhJRDpJJZ1uagqq
GWJvoeqOJjMQn2MGdhUxER7+OckpjzM8lpMBA6CiPQdTSuxeYqd1yb7GFTH3FkuJ
nkSTJyexO8nD1kj4Bna+H5tTVcDYRJm9qc9algTmrsCKJrH620MalGTfbgWAdrzT
PPAx646rCfic/dGAKN/e+Br+7N5kloGiibItrI6UXGxMdeJzq99Hy1e2piBmwEal
3Ez0KQvW++il757lxGUP731LyvUbN9pY3Ml43HLgEkWCwNbqKliM6xfVF7Zw3BLn
5GMYILv2MeOSukS9wYvTGmT2dYeYE5QYH8tCfh+38ucGdLwdmJ2KDpwq19oeYKwD
JwD6Qk8KRb4LBAawukl06dpC6l0vWrfmAA04S27FDuMAor07ZzQ8k+79BR2xez5k
LSQ9MTNcF+aqEAFP87JmF1D2Nd0fKbJ+bBZFccOmg65VfZoVbyC7FRYG9K5Q+ATu
/L+izCEScS9NTcAsDlerbmTpNtiKcqW7dA27BwDYTCiDQRMKqBw61VdDmOya7z6x
CuIwdGLdkPBuiFuDZSAVeQDpNcHwRA15oHXRj0dErqOD6QyAg97gBAVDWtfYWUb9
zgCXi9QKgky7pnmatn54R9BBzSqHSXDkKA8fxvQF5/jy+V+Is7p1WpXTGVbEHuhR
mDFuDDPEsgKYAaaJk2SC77zSD+DTucmF2fsd9+dki0BBxN6EZLNQ92rszem4vBpr
GpbLQx8AgD5cWXsy6V4gWtqaDx4TN6ehNAE1ENGxcmEHLf8yqNxCKvH00nTHRSri
GY95xAx0IlV3p0j6A7eaDuwI+SsR1W0h5fbEQQFxT9XOQPmwet4qXZmMyy2SVQiE
/tjJ41SfH/LiEcPc9ylo+jX0CbaaCR8edJ8bX4nGjdPS/AxVjnYUjMBx37oyIs2g
FFEM1g9aakBkhqg1K1ehqH36bAQ8WntqPemZI9y+jp4XQ98hZMj+PavvyXg+g8kf
3OnJONLXJwt5A04xM3YblmlZFxekm9LhIHOW3Hk7sb8DSXAlrI9pkt8gXQcLJ3xp
86ll2Kyyk1Pa3oUhP/kRatn9H6KDNqUk8YRsfgJo0QBvOZnkn/+E8ZZS1PM14VaY
TIkF9zppuEi0HuQjhuWiq3hsLjUj0qyNKHCYDxkZ0wXb9xWnOUV99E2rtBMr85pQ
4tm8BV6bfoVtgZT2ZMrHfhWwJc3xOpBLnkJIh2FIe49KwLCmYfjt1Ho4DdvGE5oH
koH+9eFE1uP8bdvKAQtBg3JNRcQVng1YCLxBfOlt3WZGrkJdQjQynekXa3x/4KkH
/kIk1MmBzQM77ja3BoCR0dmeNyGBX5Kuv7YO833a+4RZyUZEPwcrHMn+Msj1ZQQO
/8abjjfZm+pPC+f8P4Zya5vgOjZjOFegDfvfKuu/RE/RqBfGQHzPu8+tv0UyLEQk
g9K4gcigHf5ByYQvhS0Z6wPN3rLDXwLDrJZNysmFGl+36ngQf/PRhJt5ySkrZjww
t+qMfqOzEzZPIk9F6pAqi+FiEDLJ1xP8J3bcB5jlueqtciMDGdG/yofZtyG27zvt
5ZyNTIF65ERY/9OPi5yLko9FdtHnjXA4g+JBhjA8wxJtabxdwH4Y1o9o171lh5r9
lqm4syg2Q55QG1u4gViCr0eltgtCDseII1Vg1lnxseIsJ3Mhud73iLH0YiBpMpGJ
hCbbCxj3l8m2zMsakLsrDZjtqviBoLaxyQ5xwOKSGGcEoIqeZwmZIuc2wicnV3dE
prWfLbiDq+jlrcAAdTGWkQRJLrvhi5LoK4jXir1ap1xOasSG8aufBJ89mFZukEcO
oJ/I+OFa+xDl2fvsx44Y5d3NLGg1eOmeksNkCIfuwbosk8BgH04hPuXtd65CeoIF
Hyr1Uk3W2Orh+ZjyyTKrfgsBWmD5MPCvLZOAlGhom4Tr0g1PfFhlUF1pmG+NRhak
m2fCspGtNHcblqyA6WMjlgb3hye20LTmOeKNiU6IBzvbYLYUFOOkTvhrN4Xuvoc2
Y83G0YIS+PQGZYwLJZl9mUipHDc8IvhCIk8pbxx1r9HezldsLD/Q/yGzeGQ3Pof8
WzsboHNESyD9TWZn2RHP4OTqiUVF/Xw2YgInx9f7yCWByMOPQJdVU/pwUX8woGcf
kbNZH211RTlGmke4TDau10GPEft+VMU9+4rCzzhrc136v6WHgtwhAPRJCOWz8n2x
RRFXRmhBId9wcGlkUi/za27+p11h8l1RbyM8CDAKgJ+CHftxl6ONLZruKKEevNNr
3SVTblDuj8swhlHNegW1kaj8bLyb1px0esV51cbChyNJahHOI2S8NhqtNBtX3/MV
kAICUGradlW++wESJ9RUKNtA1A3V4iKF6DJ6+gF3cRQoqYBry460vvccEUeWkEBK
21cEL/DrE+nYBbCABEw4P4qX6nYiouhUihYw3rScfWmx8uKV+DSzBoe7ojYRlgl+
/xXbRo83MTSxgPThMWV2iYjltO0M968Pw+iu/Dp60mYq5Y2FTAcdVtV+KAYZOe+v
DjREktujujr9ENMa5kP7mP3yuJH22xanN1N+DULf9aHrjlrWBai/SfDgHNiMsNXF
yQoDXc1hul8FbUkGRWdXPgPjqZp34RVc6JT4PvjynE2rCwjo15nP2BYKx/bM0I7t
vQ2qggiVVVXnh4hLHmfbw8wLb6DHrHQHBvX5bpeqbhDbl50fp59hk10upXs1oagK
uO+eoxtC4+QTChOf67yjhpWN8rgJqlfEgNqV5hCrPmtetHtHMXbNS7chMoifQAre
+3Pvw0mTg/Km7MKib+uCXYy6+v6muYNRvTjZ/h7DeBLWrIFecOWvScfblt4/PQ95
HQZZsA4ty/e8JHqtZmVeEf1ysjpzUVmq58AUFBFX1FT/WbbsZsYpaAwRaZfGphaB
DhYdvz8oA2rsmbGPjz/b3PeHqXHDsHaaFpp1YHjZokhQ3SAUo2kvG921Xg/lzWY8
vSvIyyElz8eFadqVJubBrAje3BwqlpIXugpEUzj/PSlj2K5/+1Qea4PoLNal1qlP
cNGBC4xEj5VhNnDx2BTD/FuXPWNTTXAMbxloPw93OK0R0TBRyKoMNr09HKlJte9K
3SrHMKhSqPl+l2ogpZ6vkR4f4JTXlpqHNi7NPFKqdxWR2fHHRUNWEYXbQzn+Yb/+
ZjO6DkWAZsMWol3WqUFGPifS+kLzQcmuZafqCLk+GP50FYZqyi54MES/hVH7ZhTt
iu4NtVJTFIoIT5PUpqowTQzgpBQXvdRgLlYjfEFM9Wqk0MStGrQnWdB3NNShEJYh
bWecdJszkyknmdR2Y7bVDauaY1N72aAtklrYUsDajx6JJIWaHKxUfha5qcSNmQ1M
C6tIxGpbUXmf7joxD+s/cCAwbkEt7zJA2YtoHvymf2OzhKMGe3fN4Viq0+WSsRlY
40jDUGkqKszp6ijUiUDbd57Q1b5+vtk1iT3AUKb80ExPSHxYQ2ZpdHB7iHMRGEvJ
whj8GemZqKkfOP6oW/nsnu73Ujl6RICRQWktk9xNDWqbCcwxfLIxPumU3isxVYI8
doMgMVLsblckBMU2EyUwgImdlCF97mSfZguwY7pTqaXRV9XgvnJiwuYi2wdtl59J
wgcvI/VftCHlSqDsQZs9n07hdh2whwt9oEi8b+rxfo5HdIVSGuI2xU1QS+4vO7TZ
xjbcqQxnjhqcMvG0Hki8gRwXQY1/KKEHknP/sdnUvYMuSTK7Pir4WQRjd93KrlTy
oCi+0utHqZjiCU2i02SP+4yz197YXbIUemGSgMqtU//GjtBC7EqeWG14Rvz3e0Ks
bw3yae7aoZrEZiDgSRTt3Zdu/nl/Xb3oo6d7FtPuq/xfwtl0NqCNJKb4chGR1EJ3
wZJu/jeCBsJQfxMF6f7DJj+Hq0CLI4u7Oxnz9tHvgcrDTolvk8VE7LN0KZh7HWEU
6CXbqCo0cZEVax7D2deahAfaiLbDauSyWFxFL/DFIk/GJti43tgWPllbudtVBcpJ
1s/S9cnZc1cvAMT5Z9MComQgr8FT2A/4ERI590ANDzyTy9R0QJYR9Bv9LE5iO/Sy
8m87vUkykhtmK2DFI1akbWpteQvwlCbc90Lm4VNArohHM1D26WOAHm/8ybk9mjsM
fP5LEc9CnoibWenSGulJHzVamS7dcPM8/V3hb8NTBe6TU2JohG58IoWKvljAXhMU
ZBGfEdurgsUYg3T/GJurd+v6LmlPHj8IHcpdjhtiry63mUllyGApWdEy7rGCHxP9
TR5s7TRKjE9AoKp14BDTuzEb1WT3rVhdgbH7kljDSaChrcFtfOxNKL4v1EprWQbO
3CH71r+xz+rT31lrlU0U7q7AaKfZmoPG7bCEkm9Tzh3r3hvwjEy+4CrqiOJjYClA
eLrHSd6z3VyHyi8WUPYbew0VMbBLmMujQJtB6WnN+i6umyBaU6eoB+DC6mzpxiKh
jfFvbfpe7NDM2a4ohhTWQDY0kKqFm+GmLWJA0hWiobe3kcgixK+vk8taS5V9PofI
MVPKsb0DiQpfaf2eEYrt9vsbFETRr5fhhTVPjBAoEqoVF8TFEP1ugT8vXwCf6XT4
p2wJNpUFag75zd82BsLQqRrsU/9SFEpAmYvH72i1mkVETuOF6yaul1NN5Ab8FVKn
uD2+oMO4f1vugygl48ITuTzBBe5G01JiTgZ5gn4zoavHdv1XHg/1UMGju4oXItF2
n8NKPLsFHHXUbORXWOZa8PvCYWc8Ebcm6bcmVFgmiNsjsnPc0Malbaso3gJopiBd
9UXt/BJDt4OEDtvRBlkBqLxyN5G0/ae7CGZycjIyvIdOpthdXaHGBVAPrEq/MaC2
ngICdGCE2HUbzn2brzAXff/4NPZ1kQ2a4uE66Ggr06aR9UOlukp+pvyrv3rCH0I/
x2A0RTKr86cDxhSfrxEjyoF65mIauCC5CH0D0F8zc4lNaKmATnyodOcAc3CND4+p
R9p1vIPPezd7mna/sUtPowyQ08CEVufpvNJhk53JnmX8ghoZsLAf76LTiYkSELjm
osZ1NBNoktRnOl9LWMIAsfWL+vhCU/9Pwh2xPrhD4Vo/3fFmveUfX5TGnkRTVEev
9Jo3bYpQBQ/7xfNjnTVnBa22kUduySBQijrsAwZ8706OAzkrjJdBO3Nx6rQ6QBL/
VQNQKwv9iHEo8usnWkiPvFTbdpA6eWHOmj23gok4ZN5xysyl/MwrtpaEoUyeVnzT
s3ZmmocbaOIGWTBZIqVXhrLMQnDLgfG+UHuUq0KFsb9/Qg5x7/m5KhKwsFmZ9zrP
iYqbIqvnsXYt6hA3Ssw/AZFdqb6om7q6eL7dbogVrjTXWVnupNuo6CyhXNfD0g12
GEsSsH5k1tPIx74GvSvUO6Yb0M4rph7poTWrVNmpOpFKhd+2q/KlyHCTGo7vitC2
FKTV92mdzR/SLcsMnR5V6fec5oH9kSyep25tBdvLuGqN2/Ote3SPOUxAe4yoqbwY
Hgk6hCm+MsJ59KKMOP/S7rso5C1uYilUIPX+RiRKHeildiSzn1Sz7tkYoQjU4mzk
nOBFyW7E6qSmp48zO2mN0gNh+3urOyEQWP7olqkLvSJHtkNNh3e/BcdKpOY/bAKC
xlmBPf/E5WxC432E+/GHlW1TUFQv1suafppo/lDmUDg21C0KpsTTsI2clI2wI8pG
dn0TEiSu7RGewqYkelvN2x7ohY5Uu5a+49Y5zbEnTFWiCETi3jb3ydjwRGtEbRbu
2dhMNuLnum0/VhfSNgP8siHsUfJLerpdILatF/oq1Ts/zJ3rtLswJgZO6KKAXgfy
9exg2ZCLxNEkYCgL3sgK0nGFapUTayqyVmtGWSnDbkFZvTLM09KCFdXtgmfe2gUd
i1FOhEWbxKhfj70eNMmNrjQjFBDSlmUaUk3g8nPsisTiqaN0nh0Zv0tOBkl8TE7o
X65AGQw/jZWog5QhTSOhKhf6JjqwUG2x150zsyG1Ph0tqDWKp5FEJHCFV9YlGu6I
v4CJgIX/kzFI/ezamJK2vH3Fp4orEkj6MiNQPWjRT6BG6xHF9QQnU/RC9tT/vRV2
uq53uzpdLyoMTTKL2wgIAZFGMKSGuermnLKT3DtNdrWBeTVRhwRT87rR/A6eu11H
hk7AwNUKghzOJwiKwWRGvPPkRJ27/CDoXp0bhxd4uymMR5QZ1gWfJVSG5DCvxKL4
m3uOomkjEZHvmQyPB5oTaW+/UDoO5/f21cQh+254swK3z/zlJI+rEY42hVW2/3uR
V0pqmHTTYMX/5607NIuMb7MciURYD7oI1Qa8qlSdIHv1FM7dzxUqx8QfCB0wPRMV
EQ3Mkees/i8y1+i1AHsLxI5QtDjQzdUWbu0GnMQRA2D3La/yth2EKNBrhg9ddBT4
c3+LwB5F1DC16kh/IBR4tkdh6eyKlwqK7B7FOuSbS5rbBPJro0u8JYQpXIufGp6G
Hhhutol2aXw0nzwnzGyROAtHzSFWHophvdU8QtvxfKRTgkFFT1+Q3LJWkNdJ5byb
R48UdoRUcGiwCcU2NQShEmTNWjgvDZRxMTAVKXS2meI1WKhNvZN3ZhMk3jgY990p
HIz6JvGRsh+f35larcbdNwAmEkpeulIcM7qqO68BQxFcUukc3xUcL7PQacO3deO1
Udb7J0qf/SZnNWoKG4I/04KNyunWZ95jKCBZyoUihmKWw014z5xFcf5EX7mFdrvT
Cbp/jz6nSMBBe386x7/DLl2NmLMizansL9wyHnFEd5qhmyz2aKWncshx3yFww6de
Sr2aukEovCZn0zFfnao6qSEgv1g2cH6GShbruT99QFdyvs7bAkpl76Zy8eYETUIW
9QdDMxjSe+1nHrOXSPqQsO2HkO5oNKNNKgmPu1gCA/WEf6nB6SJLwe5tfUtAgEc1
GU6ixsbP5ApONi70kv4iz1f7Ue45hKq9I7hMAFowFSYjbYupfhkunlMN6b971jmr
WhxncW9qGi0PUDhcdWA3Eko3/VbIqfcVpyst955mu8ckG+bKyt/m/2V4oW7iAj75
pALskOkZa7etObnClnfKGtein/dynvkGTk/MEOrmJDTJCjxEKBfpt7SMns0moq19
BgoQqSHUyRKkotfwgsiVuiqD8YFBLFIYfPpgg907YIFPP2wwH21HLeh/TK7Iyssz
xhGqDpxk8FjCAEGquhat6wnFhvz2XEgjKB82gI0h5jd79b07O5RMNJCmoH9dAO1V
Lg+wQNEvoyWUvN+UXN5JsR3J2lcXWvSiKbkKb9am0H22d+8VhSmINhJw7Huhx5LX
h4jB+mTihvaJRbHq7ibAbfoFJ1oqN+MChnNN4hFCe86QuFYWcUwVExGMT8/rfZy5
mWtdRUQ67T96mtGE0mlvRQzcU0c2TSLVaf98CiK5LZ8a/0fQzP9jANxYsLN9OD5T
N2UTPsujvPtXqPK0GZ8AIxSbrmdEz54pTuu7GVR0B/HIiv+KSua/itiB949oxXiK
qMNj+gdRIzdEehqKQgV6mhsW0Jf0MhlPlvzFeS5AaMWW62oaKmEz6LJ9jNnhhWg2
bYcRknzVCpcY2Zj5w8YtPbnyZybsEoobKsY5PutiGcwYirq0n2/h7jE0zaodEAjs
GuQsaZuqL/+9VG+f1+r8SWHAtXFUCA0a+L52XdVLoowG4F2rByCRPVGEgUrVrNbc
8kSku+R07QBblcRjRzXRQ52JW2e2AfHvvwP60IhixxNKrdi6fqOt90UaG33icXN6
FvOEKUleOlTZi0fDNniZJBJMZOttZvoSpsblkZisaN/43FxaDpDNbwhiCR/oc1rC
yQJATnJlHr3pjEggUMsS6a7jj2oclMcO6WL3lpBwNgd0mWK+zdbUQeWP83bIC5pA
LfrqWPDmFrmHTnkJ15S+T8n2vi/ejr+nSqiKfJty1JeUzx8GCg7PAqMoLWBKF4N/
uW5wCGOH6+uQBqKe9g9xiNjlvlyZQx5t6ZdsHeEN7E9DNX6xXWnJ0+LjSsHNgJT7
9YHdDYtaBNUDvIL0vPVhJNB/CwdbEH9LVS+mXSBk7FTSz9j1O853+weWpvWiHPm2
6HchhRvMOJ/ov3Mzj7PJ8tp2hrEP5G2xkfbNQ153E6oQRZUdjsyI8M0bIhBrsHWj
w256Fnb698elhNIa5Mij09dffmNVOfm9nFsOLmCdQXOTBEbaYuEpC92atmojeqCB
HdOEuMDpT6goI4koYYC69o1q7Pq8BjW2kdmCMIcQth/IPcyYo5Vve/dw9Hl3Mu58
e2t0zAEl1Y4dGcX8BB2qSY+sEP4eB3m+pWW4LXmWDDSAPTmw67LR6W8+RjTV5e/l
V9VsNlQER/uuuqvMqx+0fpYX9vctCU2MlZycSyFe8VydGmRgPvvOMyB1721vMmYu
9VzxqZZxnzgoWbo0iNgW6s9kFO4i+zToQd7ULV/SmIZ/4/CUs2lEM85HATFrvwVX
Tr0GMViwdctgL6I0PBLCphVjyZQTmsV58ZidRvkchQiaOhAAHuhjPwhDDfLVRQ8g
Ro1RTbInPwEkTBDkH+PpzRrUHRzKSH7KBScMklWWoLGDqu4j7Raa12d7YOR6Rm3w
rEYT6qnBgA0JOXbaCQ5kotSz+vseHH0UeXPxBklvQuuzpNFIAQoHYNccnbegsvbQ
4Uqan19peHhC+zD8KpJHAbG2K1QjQz1ABAZ8L+RNdabawMxgZu2RuqcvAvGuIEDx
FvnWLUjvvN4jBc9+s8bV6DbvBnfMRHOFQhIKdwEDM4flBySONix/P8sl8k33a5q2
eAWzkBmUEaQpC463z7h5ayUhCFr+6rrMCzvSNlY0gVAhJ0qh+7bmv+ylHDmwu33e
qLnoOXw/PiiMMlxTeKfcGEinLCLGfdWgUMNxHgPLr99MtdTplIbL90k5l8T5WsR0
2DxA3XjRxdypWTeFGFsyeBarM/mrFoz7lJ6c25p7MyO5Sra/P+uot0SSSJYV0Rsd
Q5l8aGTEDOm5PMBE5YL7Qn4zH/XZCcIz3BRjq20FT8VmVB/P0Xrm0aReQN/1MHRm
B5kMPESbXr6xbdAUA0t+LFq3gatbzMzAtxv2s0A6XEUb+dO8SkOnSGCYRed0FzwC
V/JJkOoBUsbQuJj4Wy5HA3qZOK4SHYLnjxGhPvOHk2mijs62QtaPV+GrLuXF+Hdg
BHgMlgGCPYMlhvhrJ+Vq79slpisc+7YXvAObvCx7ahuDup/V+PomlfZe3fI0e9RJ
fQb3oVcz57SskFg6O5FoH/JfyIt4PYJxPlajZpiVBRpuTkoVMx1hzfRXfB0NhMU+
Sf/wMkDUOeN9Lr4yrTlWOPB5Is4AHiv2TZ8XS7EG4xr0TkIM/8FBhjBmLV2Mykj6
B2PPZkWMflgAO0wX7KC1Xc8XQzdhD9uBE0EcZHyFMdLwufnNMurWHU07V1ZX/7fX
8H5+KR0tm9g7XbHeTTtW28j7CJFf6SG8cSYV8eNNV4NVnjTap96ON/kjw0clDsCJ
8oJUUlla2QDoHYzCc9TIL+Rt3YliEMZhi+dtEGBUVmFQIp9XO+HB7fd8nZuUX1xd
Xp0BGzCpJWlWBw+YUyFpZlzsnTebQmtp6sA8cFjQ1zOagX0SfZeu8X6cyEZWyKM5
0h5b8iMVn28MJsyBm5DikHMIccpb714IzxFOyNE756lTG4wf5rVMHVu0iyFNUlzx
aMi2jlCFHARdIwtAgMS0VDRzmdoGbykTaUJ/UbYb+5RQmwQBwXH7hCM7b6tCe9j+
nmVv/PCGp1FXeFEvPGIaHBVctt+73YGAk/EGkh8W6Aq+YlLh0SjL8lsmQF6EuGbQ
8ZYHBKWD/ky9eHBLEzaBB2BzIbw6JLaWpwDnANuZ1mQTzRXg0HEUsHIwYL6NSnCd
Kb1Ebr3T9KhrZIzOERF5EthRSYc3BSjekzl5XqLi2D2fVXOsIqlVoRqC+2KFDWyY
TT/gYFh7LEstBslzUbfygHd7gBeAFplDvf/YsI63cqNlxjA6jcC3AlILedQm7Hzs
Fmu78Fs+jo9V117LQ5UQSFTtxYBYWJI83m67WKPo+lf/BJyLkUDK0dQYRLXOYAIz
mpaMRYHRb/wP1grf1t8f2E1vkmRBVmoMXhhNYYt1FLe4RU68dDoJqwTgVl6lnSb+
lqtlGEGe7YwSXKrBl66XtZpQJqS9K8dzHb6Ip94aelbJ83vPKMi4x7U44BSrH0Zk
PvABfy9k3Jq82G5oNYDA/YRfx9tBJpRuz+nr5d4ul2LSlY/xxwoTixX7mF+2aI4c
MgI7uP66TIxm+2wJpv0aM4gTkqPKpgTgbY66Endp6wTvM6Sehz8SHeSw9wKF1N4X
s1H3LkEF19GWBt547jw5yYAqzJol4+Eh3Gfu2gfC69tkqPFK8fEk8jkPDyAYXnbJ
zCvo1zibj9BqoMgVidldikdf/0O6FXUw+IrxB55qbYZpu/RoelZ+zUtxfDn6FIFJ
30/3FlRg5a//ilAtjM3VqvWChOJJJly09UlGTIsCWa0vE7sX2ZZysJ8DL/BUDLI9
DFGswXdhwUklFhD8usBPwR9WPfcUuxc101Rxvp2G2qvuYY8DirTK6sbBHwhlZZTI
/l4SvHNnU8I7Gh+G90c6C+14YfdXyq/XhpIMZlZuYdqcK/y9ejRMz12SQti5B1Kk
/4IDWGlwj/DZUnLR0dtXO8AC7S4bjF17FtDxW/5Y8oIiK0Py5GvSf6PG3454YVIP
h2ur17g00nuUEs1j7xOTdeiWSXFwBbgDX9DMhy/UY1Rfqb2yCKiV+Of8GqEnEi7v
rz5Mur8T368nVr/x4WSgInRk5VaJ9zJbidT6oF1yEjymYVSoN3lLPKt+60UKHd7x
m8HEyCcdZqr5Q+hA8hw6KG5Y2p6+nFX+TeJqNOi/NnWVuUvpfc+fiIdK2I+3rQpP
y2mcB1MygT4yqhWO04P1H8/Y/BUOEFWkLjdnyva/m5vJgKshdm9SKPfDXslTaqQk
f1NV/+hH2FScz3uGi2OoweJIrupfai6s/LH9Xc1EQZ06WMhuvAKkS9ToAWyMLkCF
Tam1BRTEqpaxjUXEpF87B69Uuu/D5EdUR/nVEZp1eXsLJe5xFx2nnhZMPwpC/lfH
vUE5vsBcUa/mozIeyBNAdD8rMorgITVc3NbzZVqkVME3hCxfVDWnqXw2HNg0F/B8
HiEWNNlkKfWoRZlKPDKFOFGHIft2f4LoILy6pRUGxazvyaRE95c4ZWXqthOpMgWd
FL4tjrwmWTxu6k68KRBSPMXrbeC2gQkhL9VcKPX+ClZ2grocU/fXzmHVyMG222Gx
dW9mNsOKKekZncrxHsbXV7PmHabn+aj1nDZAAnGkhUZhIZ+cFJm0GmQ3cDpnY46h
2s2gUFUZRcaEkAD0CdNufnE66MHyYtxzaZautfjWseBvsdnaCxXwLhxJXhDj/XjS
u1/QpsMQt+gpwH6bamxaQvh7ebDgqF8mUquSiRnNKP+8wgh0uK0XnjFWeCA9TUfW
PpNSEHhK1/OPI313tnU3vO92ZpfFXimjEkMfQnAoNF0TL2vgarGm7mWUxhrQYr2M
GKIZTl9rGjsLLokjxo4VbV/ugOGukWrXCs7Ou830JRWAjuPQ7AWTHcRuEeUwyQQQ
arRg2qAPOVyTquCDt2yKLZYyVqwprJ7qgRlXzes5JL+SczheMVXSJCrDb3WiRCJ+
UMdqKUk37V0hb4nOc3+HNNsScRFK5SSKJxMvXOsGdwMOyxZme2fe3NCOqVyne8rg
TyXMlZQZOw7NKsH2aIMV+TlbVdkWHCvqKl2+mcBGCXmI5faFph65wnVWpMUfK+92
4tSpUAU9JAvB9u3NMRaseE5N74Bx+1jLPmv6MAvamqZhOQ31UBtvPC6R4M28Qiga
knscCHoGzuxW80hb8pFUgPV38tly2WBLdaJWtwvham2+ruuaWsy3gMR++MkUPZ7x
B8D2GUFVFGIHkQLyrcc7AFh7e82r4S6XMzhe1qs/5pbGIKZt+2PMAKCG615N636b
IuCX9xNHrztnliNhtz8dcu2Gw/lzl7FBJh9SVyrGbohxWfkMRkHojqvz2+euFhVA
hCem5DttL1mJ94bTfJBtpMATi4s1gNsrlTmTFIlMmkmtA7nrL56ZZCZ999yKjWkA
9dnRX0Mac5Sl+BInEIrGkND8uoRdfl739SToosg1xZcZTv0jNiHwcn5UqVka3ugL
c9svBWDgviUkBQKTd7SfQziqB2IeQ4dxkV85hp0BLw6lGFVaRXVZ8Nmz7o8DJOMo
2HPPy3nU++j29o6JBTzIlQyqkailYjS0u010PDohw+8IDcTpFiUK5My8o6FdTFuO
pU5DJ9VHoLG0lJniC4eCV60jNwJPEiqoi4MtfKltrtNOR/wiGWafZYxKdiZW3MCz
CSDE6nqY18sAmlj3dT217PuCBCJ7sNApz8duDbg9MO74B+RcpqbOgqaV2OqA+3ZI
FORIW3CoB+4nf0jfjc8+eyQDHYBMgqWOQSszfPg36oEPb4P/MpRQYOJBU3ibbnkl
HqEZrFdWJd8v8mPfZW8yICYh+HYNgxuOsZIIv7TqXMnxZiYDsO2SHJ0C1yBS93tn
HfsPpQHEGx9gNrtpZ55hN3dlWGQV+py/nkf7Il9AbOAI7em1b1bYLGV9zkYJj/i6
NS91xN2S88wunoDxizrpeuFPdsuBZyAhs5is8gxhGhhtndoEdgUyCUCsP+DY5dWb
nqveVF2ZoYl052dPPTmR9YzOTmdO/rnC6a6E1QlCY0x3aZaht7VdwrncN5cnkCs0
xKCwZzMrLUkEc7rZxQsnJpQqAyEO//gpX+6SiZ2eCBgmUnA+jTOQZK5QQcf5PxJ4
SLp6WacW62FAp/pPWmOnjdEvK90Ch0bP4aIwXMEH7IOxbZVk08NFQKpjaSOume6F
L70NnHVzo6FxHXbiScbVg/4euv1hzyN9vbufjCjZg3E/awz89T+PDYsiIzexKPOX
hPslFthXIYZ+hsJlD8ML6PXlQGWVvPFijkWRMPc9tKWQT55I8300J1OzUb29/wQo
Eo0MGJiQH7aZCPfLHSKnL8ydO8zc1Cm++mJCo72aAm/lD/laW7j64g4sDZLnroc3
tR+U0Fiw9aPGBChbVxxiHMju+b77bcShZ+rbN5JSa6doWEkL8cXSyvo0neYNyPtq
mvgFShTpzejWci7GuHwj6aUXIQ19Jfa+ckj/QbMwWTlPs3/6fbMFUsrsxbOYNhes
zdI212lGHJAFRJtOIee6SOOwIzdkZoMVmZFUDjqjG0FiBM1/P4+Ubp9DkLRwkRWR
tSmxjtkFdFr8j9sb7ez200L8GJLuplCUcZ3QkKAoS/QP44kQcwbFwNXorFHuhbKh
92wQlk4a6z2wJnlRP0JPPTkW4HnVvOwLDNJN5w4k0or6pA4+cH2M7Snv7x2I850I
ZbN90BidY3DEMml1f3aQKv2oBolaOplbd7Y1y9kLBHTt39+B/bwUL6rc/oV5QZjQ
1wenTVEEDREc6ajEo/zEgFdlUJFFpTPWAgrGb4wBuXIOq+nulwOHe1EK+5vrLW3I
gsdzqC3h3nk7gQBdod181tSMfIiPRcQ7CL24/g+sRBkHHhiVHuRzGJXyTVwE2D8v
1i3fnoFZnge7Yc4478lVhmsI3sXxlbqFWR2bfxUEn3QaMr7ngJm10CbLojPvfXIM
oqdo45OQ0J0vyR0Ky76fRxd5SPzoIyDtfz9Mujt9hYha3BMyCo5AvNyFV50HPpSx
85W8TrLNQIMXLDIXV/tK+HdsxFcZZo8F60NJ5vwafOn34CsjKv6ZzcyadCcKE+W+
/5dpA/dysES7orK+uN26gRMFvORufdh5kmzPpYtbK68wL7vyW+BxIymPNrQ+BDYg
pzWHhK+VFtm2ZqBDycHO7V0mwEvNUhuWloGdiyGbf+VsJS4eSSe3LpvTbOJ9gTDC
7DLs6gC//sbbxO1U4ip+7sAspPAQxZtNKMIdhZ0cEyxlLYnGNCqEvdzEbnX8zDl+
DCpLi9TkiqKJqAQPPh3HbDIaCj0as7WbrURIhTj4ApMsP+38ELMjparWCl/p4enq
CVQgx5ucR3u3BTJjzXFMDwKjJXM07TMVbhMBW7IVNc4S4YxVxM9fe0Mh6wvG0PwL
g5KIg5l4JDmBH295XHCnbbf8IMmx2HIHHvI+p5K3e4wlXX43tp0z1j4XvuGen7J3
kEQitfvD3vQCQBv7hsZcrkwiK1f5k+iwvm2q79ZigdAkKC1GB70DKV+W8wOPzokK
dULEBIp7qE5cam2GGXBgZcZo0lf9l0v2KVz98lz+zdFGdmHfuBkzfYME+dp+ROx+
7DekT0LLkEL/oY+wL+TRploaAdZgmDfwxWZrCv3mC6cyomLV71SFTzSeX1SMienc
gIHqdwryGK7aLyMSsB5SGkelm6l2gtgdOXtYdw4LsCLvISf0fO4npGfsiPdmCEsj
y5KyK4vHVNScaK3CwMymyCYGd35dURINvR4f4A6cyG7T1tD9sbp/nDvCQ7hz5ViU
7ltS5FxKAlHEfXustvXSh7NWJQHKz4mTB2LOQo30vYsGPulDe429uVIFBeIpg3f+
yb8ALy8pnv9ulp+RZd6EIHACiXtWgFsf+irApZcEX8HnUh0CFhEGy1THbEUuOaNj
ULUGyoEuXfnyiRkaFOrEhxTzzCAJoOD7zkNt8lhhwslVVRzny5Lh4Hmj8I1JjnKC
bG6E0/gxKtvpSuTYV8Zp/82XAXo2JpnVoQZ42DsBq+N91sd031WIBBJXjGdVQcxb
PZRZZhxLLTeP+0+JhvoBwQtbq1SBYnlVTIW5coKRTxyjTjEkHXzJn+hazktpgjon
W7Hwx98N1eh5DuDBvRGmnPjekXJ7zwkQt/8ApGDormu7vkSdn5+PXFICa4uAdqIj
iE4ylnQV+uWQf+oy5lk+9luf2vQ24DaFRygPit/muz7sQZSLFjYCMmXSHu/M2Yjb
BgeD/dwvZhYbS9o3dl5pQIxXgvPVk3c+kH75/Agfd3F3rTP3LIt2FJqzYXMeIqky
OOgxJz9QLWBzDBSQYw189odlVlOTjh0S+Pdckj42glA+YUzwoOstUjYtVUprlspN
NVOxB5WIcl0iGADeWFiGeIumIRj3Hj5Ia/AIYhGiRMsGYU3TNe+sKP6Vrn1QccPI
w1mVgPUMo3CluOhKq4fpvjFQ94Qf1XMFx9zqxb+gOOhqk4b2PDXMwXD9P1U8K3OK
h2w9rd1358cxYXszMj8/18Fz6RLKyYkk4i350sNmJL1gJR/PPGOFNWW7zSy5DhzD
K7jvdLZPiGM45Rw4naGLgMO0m1oLUbQO72Jwwb41Fjk3/d998sfzIRLgVkGx+dm/
o25QvoncBtgglu4Z085uHE9BmmS0fQUTicacBzNGueGhqOi75/P1v4sImZzpS53x
p+RfV3evSNZ6ns4gDOCW8XOdRzeZb50FKcc4icEXMQiYuKWMcIQnpLBvyWyeemBA
sNZDkD4xmbJzdLPchGK2C4d4ojzgTWPh0BEgyC/4g4qT0c+waW7CKaekfOOpvwUR
EGjMxlGX132EWBTfvxnD+Z2OEKmOUTuIOzUFrHnZNm/BRG+eGBDKYw/fFmV9eVGu
FURB96VKN69ypWwNAuMuiZcFft3uv7MS9ujuqd4nSq/vVDHiYBBS8QEKYyCw2iZy
Ez4NGrkuL/Sp53elgF9uhgs3yK2xhZOtiL4jsY+oKdFT20OieXiTqmAqWWqK/+pL
eWxb9m4OpEomUqEdmPNKy+o6XEmlONO05DAyzVQm4a8u3IX3kU/XwXjsKE4ZOm7f
q4DH9fpjKztIfmvp/StKsEDi4iAtAs2ihkFzPvkl3crJvPDqbpBnXTL+0N1l4bQA
VH2C9HvKIJpDjzpvGTLQkIFK43X/PS4iX482Wkqh6OngSRAHjTvysUTkYupSTl9w
gSOg7qKmV27c1WEUY8kDPDRwDUyukH4uFsG+p2uRqETM3KN/6npKP/DG/SrQytts
pVnZMZ1wNKhwQ3GfV2qEJd0MsEHL52F/LaY1EAacSCnuIZXddW/WQBQdUPeBcqiD
xsw+dCyc5C4OmphHG+3ZmJBDDGULtOKu7feDVARgoE/W14M/+q2aadL8FOnJwXNF
6nCi+uL1ddm6ORZyZ//czazdV1cOyXelbAIK/va1aJtGt/+TiQuNYZG0YRqci2BI
H1k4gKA1yDjOwQbcT3Dz3dpL3v7p2so1MZ4BlEEWmgxnmmQlpCdMinkFwThMCyPP
G5tysK3ymynuLtI+XH8nbeYc/V2f2LgqWv+hyRAI/dOXmErhKegagTyGBHyXi88H
Nd8mNl9tBxvzZKT7NH391pe5PZqHUsasHG+2lIQr38B50de0mTCLVQDPkOoTl5uh
vKRCfuMfeoRRMJ80MrCiut62cqsAH/IFQLC3+E15ZVK2Ik5GIDO3Pc10VUXRx1ld
W0I6IyheiXIcGFRIiFXvc5YUwr11OIUiKGVgn1Lqb8YkjBB3uWR28AZtQkjRIMU6
H7UN38Nzxbikcb7renI408guf/zLoSsVvz0amh02CB8dLmCdo8cnADtMUL8qREMC
WihfC2b0ZWSG5x74z1jXnm0Y6H3/kea0wVVtF4mrIXs8/kNCvFVyESZmYCf0B5eV
9BdhQCgt/ivPzh5Qez8S4XkJILH0t0nLdqae4eSCwpajX+Ejd7G8XGlXRM0tJ4j8
69acE//oqQ5mYMARfpdk387RtX9c1akzhtakQOmRpxhq9jSCF/UACxQHmOWydCAX
LJkY1c0X56l//HDTGXieFslmYr4P2hBMFqC/89+GcNGV1dyhBoS03YdRWnUw/Vkn
Ew4eTE0hFpaGd6INzyP7ngE5zG1F9Qaz5USF7+JbbzUfwnLzz6I93WU2DApRKryy
TVi36GnDCfe6lEDQ4zOouwyUWQ4pViuxjX+XtT792fQIQHm0gnk5uVKJeon+2HgI
5mg8awJYltwEualDAPm+4OhsIkT3qBILn7KKDvx7Xy9Xs30Yz3VN9CpexO8UyP4O
I+LJuOWkpdq7hEqpBwrRkEn94/d+jHKXbrg6x1YgvoBeK88mlNRO6bGUl0f7Lkrw
i6R/rh+/nVjs+AGjj2DOBlfJbzRSo7/FTZfqJdBsDFdHCbJjuBO/eF2b68Zrz5Cs
hRqPNwU74qV23Q5iMQPNA8Aa6xRkrFgBRJN/rBo1QnlaRtdBDHXPgOR5Dv9952Nf
QWmm5fhSyHcXlGtDpFR3hVMm3S73EPXweuoJnBXsEBu+UzIzMrkVAydUmgG3OSNQ
U2fAStDFDh+3atru5pXAU7lcKU9qmIaA3Rw/KQRGDx1RHmFcPn6Qolng7NOLDecy
ccjWhs2ElAZezqjSs3aFqXX4aswVuo+06VrCxLOFkgNkxPtK3aL/7FMxI8CaA2U+
Uqa92l0ZuqG67+n/2CpRdAUS1Heh1oII+7BMe/bNOld8N3sIMUk0g3ctjaVacdCm
Wk6HczwcL1l5xbLtgZtITpMtDY7Gm/EiBpeu6G0d9KQjH+xse9w31+NTWuO1YVP+
JXzkLvRPW+TRh1rHhHz8DtpCRo50PUT5b4qvKV8a/rYeN2BUsvJXVIKL0gS32i5k
eVa5Ioy0fSVTgsC1rPRZtOSa48hLVTRW5dt/3ICFN4PiZu00/pz4F0yWXfKMcENO
7Hha87831SiNLG2IwCqSnNzBcIjrlIrLyQnHJdrJeXaZsazKJIihONKFUEvVz1QS
WfyJc2jL4mv+56atkqnO8wgvTpIzPkJ22jGadUlZkRMAnVs9y1c4wRTfUYlp7H90
EC79vipOrKVwaQPAUQw/fTBYLKm4nxtYskDufPTRfLE/+Q6NTxAwZvGaiGY3M2m3
vTTe8gBVroTl2w1dqzIDsN62p4hILLCRhqE4C24HXljNGxoSnoWw7Qqm3EbGeCvs
5rdtM8jrhQbHUqaWeXqEzqo5xyoejwJHaVmjHRCUrczxbZyAFnvSSvla9htOspws
NfmDhh7WfCppK81WVk1wwviBNCTTH8mxalvWb0Z6xH7DCdCJRTfOQqyGYVTeWK4D
ybd3HNGpSBpg0j7WC7pWsHRS81J+lnWxQs3f79+/ZPea2iC6JgitMH0iFpDwDAwz
v8iLR/x+s9anKdaTI27PD90OjWZU/S5jAUUm3b5WQd0HAJBMPAo3LjxRp89V4B0z
hbQ/K7/WocODNTvqXP3+B2hqq+MFsBEnsqgetCMfJ+enLBeleswAuaplS5cEofHP
sTMjqP+0ROPoszwbNNUwlO8Kt9i6hCXlRMg56aPBbhNM+mENSi5rqSXt3rX7jtJg
CQb847EiHsvBXqPVyhgMwC9PpEWTnV2GTumzr8Bf2xGZ/viRsufeQc8hBfIVELQy
WS/7ogl2kJN5uoVz7ohVejeQaC784JHV7E6yfKWrMm4b7K4hbU32u/5ohJdjJKl8
5tXLidd1tVhvVugjN/aGoHu6OXAoU0qCdyf7rxyeMpI+gBi1Xs073kFN9hYIusLS
6cIb8t6NbuQUHblJjiHxaZqZLcXmkY0nOs6S9kTd/V45MTt3qRlU8Qk9unwIFRg5
C4prTqfqUD3YArzems6AmVmAh3+8SEDg7S1lejdSQj0n3tR3h7OAt53u+Qxexs64
F9Nrxt4aVGzmmGTVKqUjWa+h8xrdBSD90RVwALeBuPr3PQPIw47czwllvzU4Latu
hi+zPZelX86zMvx5Z1kJNYToFnXWSuXS8th7MLkNE/+ng0GKxROUqObjX26Fq4cV
RVGnh3k1SheOJnW7KLzW+jo0OgpXu5h345FflT/SpmjbjZOHLDsGGwRyZpjacbUG
Pb96E7jWHASRuCSU8ip5MCmKrtr6X5rgmchwBkG0cpXDlJ06eh47v76s7mqGGk2q
S40efoROr74SqxvRmQT3Mwotj617JCyTM9rhXUxt/f7exyjmVHzUaZq1eX8PjBwC
dK2qUu7+ylKceWCX47/k9P8Z9DFeS6dhqd+6AkPvxDXVoK6bXXZiKAmaOysIAS2L
wEgsFeBnI390w2j9s+lRCvcWWD0Qa4LlW5mZNwLTaueG4+3NuT0n6IL7n+7KFJTO
m6v6FqQvdDbFQpRT1OL5sZLK1CMS1j7JzvydotVqa1Lag5v2dRDxcnEOc2bdVi0+
R64c2f19OBV6nssZnF471EnuwjBZne8rUu1HfNmhVfcBaXv82YtrbMGlRDeQbz/Y
Jl0SuOZHstPPiCTFtMpCq99ueqceAKy3oJUulRp3cjzypyIYcLNvd9EMb26JvgpS
nyKODY/AVW7NaIbSwlkgV5di66A34CzPrUJQcQVgFHEuFI4FmtYMarAGrjfSRrHs
Ms4x5n2iSEghk2imsQE01PBFWcjHMNQeNxzzbGAMy17JSsADruEx3hvYdA9mKuaa
F8qla791/gh75FEc6lPhR3R+XR/KwGNr1Tw49IHfUNRCpE+qO6xf2qAAoKl8ZCiL
MSRMkZMji5ud/EtH0R6qS4YG0KtMuaRv3Yw0/S3luivB/4pUFzrT4VqAlyG+tRen
p2VlwfEFIlKSfBu6XsgRQJFNlhgUZ9CVbC/BXhVnYk6xmowXi0KANyqR1o7RtfX5
z3ClMtcSMA0INdP51WskZUzE2wC/qVvDp/WU0cIbzL/haG4oEPRpTXU3tzfEDsVt
yBvW8DWPoo04uVDISp5anBdSX0DzdI883RHgkc0lSwKfviUfEx9lvgFRW1lx9l8M
/io9u6yB6n+oLds1oJtg5uN/m3C9DjDu9bOQ4cBNpVlaBw268IYKcmdS1OM5KsxS
K2/wtxrUotb5LFzrwSWyLoY1pwTUiQDgV8MqWGsloOlh1vP8kan8jksDxDNrlYVO
r1qxn7n3veu0wjqRAJI81DPZpPXKYVVeQM3Bh5wvUVjC82F7o2Uzqz3wv+CDq9wA
jPk9MVSUQT9/29NavcQNFkeaOfxwPohl7jGEVpRBA7iUsB/DaDuqUh0Jb6bGmguw
JLvLV2SEwOamj6VAaAJCnTF8VQVEu7GrVy+Pduhm+WYyMEdfGXdGX4pKI8ca2lyp
jC9i+4ePOoVn/Naou0l8lG/AAIBnwhohc6wJYqwb18C9I5dzdoH1JTWuODzCs02J
oFQjC0YzfMUQnjz+p1PSNuYKW3xkT+fSMH8+HMl38JpKbvKooR6zQWyTJIjIf22Y
ee+QFZmZbX3lGDWAaGxMSrWUKXHwT+GY5xhUQnEYDTUhMU9yCl+meDQMRjD3jjzO
LqkzxgqFTJLumFTME7MEUchCV1uw/FOgeBGfXILF/iSIxFEZk0o3DWfnOKJWBe5X
YkVyZZ10PHcHqjQZ9ITmrQ==

`pragma protect end_protected

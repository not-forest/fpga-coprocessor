// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
FKXN+B8/BDqyGoa7xK5uZ9brhZT9P5rPcqqbuW5Ri3pmddmGTf/8/qdHeNoG8eUC
+lGtPyqehmgz189dA3ilCwMhIxkq4i/IbWa1T6RXw0VzahnFnjKqLm7CyYxQOkTH
7pTtQ8bJTruHXvPgVRSZdRjUZbifiTT2c2aodSzZrYsB28IL9Yos30FyotYxNKcl
hWhuVlazu6ZPVBIAzpdscowbaVJ1wOx1ZQldzOmg3QoMRQIesHD+hiwtsQN+gt9J
CebORTQVOinBeByQdm8a29TtmZ7NpgfPjQVnp5EyOyd0oa5+nmkhqHJjiv1rTHXz
/AvLn5j3NvN3Hv9TMxb7Dg==
//pragma protect end_key_block
//pragma protect digest_block
2MMfIccNAg84DB730JVa69p4TYQ=
//pragma protect end_digest_block
//pragma protect data_block
2bk/rDjm9U3pYblTdhObLMp9pRtss0ZACDFOWeXfGDURLOqi91wXvp3QYW7Wo/+3
i9+qFYo6YSwWj9qyBQ8BHXH9sSefti0VT9u4LvixYyU8SPsFPUBtTXyHBkiAbuYj
Lr4qISopNXheVnU9cVAjc3kOQ32fQEuCSmiFJXzOGYPi+xkFXU4ux2vU88L/AIma
ctL6bbu9ib6LOjdFBXpU5PvgkPzp1mz8yySZCdr0eiz2++tXyoZThOyVrPFx5mPs
KmYTf37IFvBSStekuMR5KGY4MH5hXwnkosdUVY7m7wnVPurFqRZ5qifWFbyjMbyR
Y0P6Tip6Py5kciWBTRgtvSJFWnTbr0YehPTMiFBYzPN44SCRI/jkG4VXY9BxwVJl
g/2feFupWgDJbAPOFwFcNcYPg4fKPrneka/dRehJe22whZDc4R+LBrCmFdY24BqY
1XSzHxtcDdbbwmcjKN0dyEO3fUuuAguf/rvGrj8ppNubSubarJHgT4/TIulmtg55
D7mMA9zucgdh2FHE9h833BqS1f+NvWeDl/iwMx7ccb4sSbX+qCww5ICpYLw+fHyg
liBnDRi5uWzfEIXcCTfipyuMSWnqIK3kICAAulEls3Zo/ni6wRvAe/5rTCHPawrz
dUfDXEbu1NpRWJQxZDdkKDNAznc97FvHXNCwX+PsPo4U561fBvp1ftuR2ciKbrLj
x0cz/anB5cMNaQKtJhgSZKAtqBxqktsAbE68MvWXx16AnEnZe24zZ4+xpxgcGLNu
FpRxQk2W9q07eOBR1qJXwJToZUjLIM1E2t5unnhNcC1Qi6yNFbKI9+dIo4CAwwHs
y/q1xUEpIHF44ItWvXBROqOz9NZHxZBR+fdaG7ZetYcpxKtfi/QhCHlq+B83BNhc
NAxLlBsHTCbdmeuPI8i7oab3eXmSprKPtQ68xs4TGxHvHc8bTMSJBb0GDTaE+3PJ
zgZlHcQdDPEo8l73T6IjVFm01tvyP3GJfbJJ5QBiaZFfeyR7Q/6Otik7bWYU9zln
6MpPIIDYg6uKKPlmhaMXJg1KXzb6EkC4WEt9CIFyV8x+NcGBxRBWSJy8zONBnRmZ
nq2TqxV0lm91GybOAH2fFwLT8AFKJFdrL8+uAXHBDrvkhSDsxAyJ/HfExl7PH0LN
nNafOzhKl6oMKGCYdQ8a9HDGLbLZ9I0sliKusPpVidtng8iMJt7K0qVFHrsLJXWt
rtPU9d2WAO+jehHqiZOtRpcPiORzA5/kyUqSJbi1P5rRvh7O6fwHX7UMOrMd2mLy
kFShFpLrwTP94Z+c0zPaNOkki9YyMPCwESQeBZjBDdVTCRoz0OxnIa8h5/Cu43nW
5WT+c1ralnnTPC/mF4TtjH3vO/+FXmb/iWWb8s5d2zwFO3PyQZ2votCMSHUN+CAz
XjRQoUPeJlx3mFWw5pKYwljbEZ+/nXvMnId8KppIWz6x5e3fVyOSZhNDh7ILGRZj
YBFGZs7YQdE6TDPrIxEVf5r2UnObn/Wn9buWpq8jRQYP0op2BX1oLQfwmZit6f/f
IQq54HgWAor4DnB/NKGc9hkh5rENfA6VyXC/dIxgGzOWEkIen25ckXnuI5LVMsp2
zdjLumM3f5AG2zRVcuqFvuprP1e5JVpGZi/zewIIynsXxemAYOZM8+/ITO8mOCpX
ehJKodokIuPCoB6SBYDPNRvXZ/gqmsCFbg6c2+MUMG7lNPMyBw0Wz6MyM171fAyi
HvnltUlinBXbKv6UiEDPQk69xkl79Y3k2pZOdRdtOnp6esvj2DWODq7xU0V+ph62
pSOsXpkPX8KYf5G2xRDTSoKrovw6H29dOhGGGNWkfC+zpq7S8u3wMGntCCA5Xjhf
PpwWEQT6SVYB2k16J/tOFo4jnLycvGHag/dwGIzPXE5F52wXCTDtpOrR3/8yvged
dTx6wvZ6g1QCX9k3xsZ75OTlIXglnaT9aUVJjkuaM/uRrNUglEWetn+kWBWO3tbv
TalDBl33OVGndrpDI/J6/zqBFAqo+BBjY66PWEuOtxNfRYBPKhPJ+1V0ytT8y5k0
sZVmaVKjboV1dWSit17b0KLG6p0Vr7NKXhyUF4YFdEuOjE5gCpVXvRrYDnv3FwGf
aQVs/wd8z94wdaRK+tEfIl0X8IEepIST3WWEpQzoHnal5U4BsZZFtFcqpAtD5efm
yEhkjOaW9NB7B8U6SPuG+KU8vUBIjFc1v0oFzdAKA7wAHqR+TjPJP2dSfQd/iAIr
cZpfOfIQhax6Zvbnj8EmK/hO0zJ6fqLsXFNPD4G0J4PPN7nb5jfiYVjuNnn+FTMV
7CvW9/Fm/lcZ5FGxsIIMZNlvqJWd/3MstMo4XW+T3OE9QUnBpttpnEdlmplI48A3
O6RbzFXnqDLYi9fyVfMR2iIdiZM1cqVqmsn6oexO6KUoABS6LmmnkEhGJ/yXjdaD
0SO55NWUaaq/3LtC27Y4Jo0/XM2aU09lDh2+jlgtgl5c3HOkCCflBJt0akFQ4phf
56b6sNoUpWfjuQXfJWkdSMK6yC0gTZfc4+TJ15JIxvwcmiU1MEFR+AZfLHv0GVRN
nOhQIsdfHQbD7TfaT4hRPonpDzIlK89hPFhziejUHo8npYQU3Rwe19YPvRmvT0rH
KaG0SQcUKwwy5+U+7iGafUFu/wS8nnL5X7lS5dZHz21wFOYe7dXtpS7OVib3Td/k
XgjcaSr6GvVoQx+/AwoTel1nNUnA84Y31A0mBbocHAgi5hQHOXSiUpvsHzo4kq1o
bgXZNnlTDpEYabCT2ifofzN2Lz3bfi8m6XAslbJgTR4csN3dxVwaEGY6UNG6+RcA
95q3G7A7GIBER0uyEVBNdARqpvNxLGREBKtwnEbDacTP/ym1N5sEvheIqMjbCWwD
oG7RP7Fe9CkZVIGwd5nbw8C8IUOeHwjJPha7BuKi3kLrd9bPLO5thAq7OvfapQXJ
xoqqS5mVBviXe3NPHW1uA+fMr2+zU7cc19/1QoNCv/CRbUDUMHbPr0ZbekJxfQNm
X2EO62L5cGvslxdzJp/xAArSMj8gaY4A9o/Y5uRH1vuaCdb21aAj4DSh6VeHpG5H
hnz3hJtSF7Cal+1bl19izdg+LpUyo1ny7POHI51qxE0oRUq7u8NgpgG8ja1YPm6i
AIfHuL9GwUn9BsBPQwXeS0zQcojshnt9KXsBM3Tu+I9UwSmgXe5r7IJ4L+aeXmyM
rzfR9nlcUNbvTCVsdoF6FbC6txBW7FED4lS2gbsx41BL8sKaVafdYKhOlthRXp5i
eXQgrToCj81iH3kHgsGm5sYyyHY86GwqzkYuUCDd2oWFCx4t0RzoxGog0c0zG1IU
tx7rJf9fsvEuytqC5x7ZVJ+pjG36lc3Vyf8yvic6BEXv/jzQUd/BeZKuu/XEsdfl
TrEPmxpB9wUUANZpt1wAozGb3K2V/AXZbm72QBBh62RoBRh+yxPEZOM9OsRIFq3c
S3Zzvm6tRt+ARL9M/3Q5l80Fc63XvUO/ypr2sUDsWbRguG33x/jjmbrfNiUiGrlK
WAiGPgiSCtw7Awvq/Giy/0bbnaGZAj8zTtloFkf2BWXE+PYekDHZ0eeyCbGVlgtM
P44W6VBiMeARTqK8ZXd+lLxshHxQ6ORCQQSm5i/x6TnDP23Lh22qrFXKGYT1FZoS
SLz8Jv787oYzhkmeWrQRAFhsH8u2xgmAF4bN4SESKi+hXsAHJN6VGGphU03geASJ
yHvXK+AMB7EzAIOMuPv3t/SBBcqr8nNPdl9zDyjPyS9yY3O1Gw6LE+7zpgd/r8xj
5dSr0CshQRcpZxBZVKBG6+1Ly2stGt0GR00SUlXrbwv5dmEOdIPL3ZENJvtguSN4
3EfYhUu+RLVzAUS4FN6xuu/RsEvgPHeePJwm5PNYwspDoxK+4c+cqB47VxbXPadG
t83UuVvQGBl2SwuLyQ/zZe5b7c5hr+HYk25FY9B80jnMcNYnjyjxH9vw7m55vTaf
MbPTXtcqys6VWc9FEttki1NHA1ZJYkijFa6sDirgErvg1LgNbt5Ctb1VVAEHIbHR
6E1Xs8Ig31/2I8/fInIkP5JTpGaZ4l3jNPbsfeHSgQbiI1MI0rkuTQJBoC2sCDbd
0Kpgf40+YUtYXxw6jA8idKGgxYoM/qQ0wmLYreu+ZGlh814AZL6nKLzeTCVLj9BO
XSiF9fKyxFqMnE3Q8mqilsE+ZcnzgaXuV+1neDOAwC2VsawfgU0saZd/ISuR1uV9
SoHGNi81ll1KtAWbcOlOSyLIfDkxaUrLIWuysiwhs1gk2qX2T/kwQD3movPKRRrl
GvGeiC7/StgCsKgOWJo+mvUE+FwcBzrvNMBz25auHIFKOXToH8+xv1knh4bke77G
1GLLdVuIOzALbnA2fu9FdeIvzS3Ln0wDI5TSXa13m+9gr1YVKhaffBtWt2Wv84gi
P/sj2/YNGcsU8pQCukq1ZWVg1HjSn2iWvul0gt0Z71z0jwx9LrCIiQewHKWXUVol
7cEBlNKKa658YqxPJppbdFDUNlR1P4tHDB22d6aVDnYWnlmrcga+vNvrj/p3TDMA
/e0aHZVoj5NCbfEvn7cRXUI5FY7Fyc7Uc+ebTy3I8kxKPUyd9gMx2w8+p1A2jzTT
ZYyw//sWc9l7A2W5Y7fGrhTHFIXlMkGX5bIgYFrEWf3vx7F8QkNGemFgLhI45lVh
jdkKXj7JZxKP59lk4YOZpzpF0x1BhojCLzJbAS4Tj2LrGQmK4miYNYs3lZeO7wM9
WJb+neBCBJju4INL+xNbKZzwRetHX1A3y3ZtPERUqD185Ew3xwYyPDZ3ELCbkBdR
A07VfKWoXCF0cZLljmBA9PyTp7u/6lcBLBw/j/SsYh8Z1LI87LC83PWWX/cQPXcR
shgb8E+8loj64+o68EJi9vRYC66BQAO0YjE+wHsi7mw01ubczxt3fR+iODrkjjUH
nkwfirUOdxchAHm6VCc5LY1qn/5ulMf1vrO9ozQERpsSuQjAVHWWwunwXQ/eUzyS
C5SnjT1jr5pPrOm/MJOk1+U+HBUCJGhNTnPF86mOoA17i0kCHdzV+xGgqw8l6s+G
lD5uv0W6Q6MGd4jGiJ86q9QgJJhbLN9rlgIZZt2p4YzceL/Mb4iFnzgkS8x6YmMv
lVd+dadIeNxtLTKx6hvyuMxJTya8vXt9l7Ut5gdOTEbWoDpMROLUv9ouTnxA80Kf
11Eyq7AUTZYD+nkDeI71P3Q7YnqckbAMta+98sLnoESOpLDBUllzUdZJPtaMFXOY
nSbYDK9lDMXMWnO3GtP0w38frum2MxUz1k+KVPwvjeWZmOFUa93++MQ3ATGZHg+p
hWMXQaA2XWjBeTXBvQjyjMtaamQM8O0mUh5SCY74jJ7lHd0W0t60ovO+NZQwG0AZ
1rT7zH8F8SIwwyUFICTg4f+YEkUz0z1uawMEII/T+7hQogCFUZXoN700UuiCCjkK
FoWrX8Ofox+rOZ8m2gWOP1O/9tnMJDzP+LGAgODhPn+ekjF9g29cxE/zK4Qf40WD
EVdVjWaugED5cQBfvayTDFKUkJVl4dR5Y6vauaapTWFZpB87ObCR+sbyrAHKVX2l
y/O5vXYTvMxkYp6F7uieHUdNDcuy0Zs9Uj+o7bTp2JSs4ADibqrPCa/xLtlTA652
u5BepWxgtZRkWpRYD7KIA0Vzb9PoLzXdmc9CJSZGuHSf28xTmkYePnuLCFuF+vhe
qq4ZgiAEdE2Xe3zxH1OwAe/2YKqcF8LQpOgHEKA6X61Mf2aChisWST0YikyUB1uV
vdCpYrRsChxf7g+G+YkUBWJ4zJpr9sWaaNfn/6Sk78PlACdhk92XC1uLc7fNfaaf
dCecnsNcXAvlbZOI88eZRagGPBUUlFv3crxFZyaLC/ON6IFeYVnZ+FNmPzbNK2FM
CMQrNRoawK6goa6fygqAlMRTaVE+RPwKuMaeLmZpEyqJanBP6TEj2Hl8GEd3Aslr
qc56fmn/z+Vdr7squi96Qmmap4w2wMqXKmKJ+2o2uztuJ0XKy9rFJO2m/rrkIb6/
dLI+4Gao/auIXDBDz2XMrRvrjZC30msgghBjIuS1vFrgXA7cN/z3UbTKn2sj6M+g
GUsE59ErT5Sn/OTcsvRFsiVSjImB+6NZ3oQfsuHXD2jdGiP2eBjTnhhIV8lU4a9W
KgMIGNZ2G93hV2Y5aZmRucK7WY2vn7BXb1SlBgj1img6TE85L8gMz921QDF8+iFL
T4AUI0q9761GF71ed9vtb91e4Ot/KE5l0SPMSmWjJuNvX1qXtM4fhx//CZQFACo6
Bq+AgQoZVn2zBzUI26L/KJrI2ITW1rr+owMmbnv3lOPaLRQWxhsVfEPzzGiRGei9
IvteGxZvWZvavG0uYh5U8tbsil22/4jaF+Q9qTRTTMmw3ZdpP+Gr37X0yw0OouKi
kyYi8jLBAKf5Enym0d64BjjlPtRoGd7qVkJMQQfW/0u0OK75GMTBv+FBa+ovZUBw
IwcxnEYtZtCCZDH8xvoTlD2UlA+gQny7GC7GCBNtRBA1yU+WW5G5L8FvomkL8p5C
ipb5ke7/cSWClXmqkZCYu2+Gf12pBEH1rSATRWFlBIXeDUzEvI76CIppgHL1aR1m
/OcMeKOQMCXpslyUSRAwSRbAMAZ/uLRoM41tmPUesyXYQZLvEQImePSFtAKwoCZB
xgQfZaABZwWuRQeiN7OJAvl/925d5DhyFuQ7wQCl7D9wIM7+/Hclgyb/c7qenKm8
5TA5y3YLH6GZGPrm/8b9tdjDH0WV6tMSHOzW58FaRNRui9lVmbbsAFteWkzwYV1k
0aQnPjguoaCW/socTJJGgNWXzPzl7oZlxs/RHF6WY092lwaadLISzuYpQcnzGh52
unKTlmuWEbv+6QvoELxXU+2gh0I9FpfH+ymGbuKvN3VkhBBTUy8nDTEOryLEgSIM
kkxncbRdHXO20+aZA+MZKZT5hnTu2l4P75ULQtWGxMo=
//pragma protect end_data_block
//pragma protect digest_block
ofmGaP0hA5S/ch2u28nNJvQGo8g=
//pragma protect end_digest_block
//pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
eQCtXiq6jYaNo+CGggzWNqLyfS117KxQMx8ZgBSw85St2CXP3OdrC+HvA4JbaB5d
BHnjkD5cHNze5HPX6pHM/lV17XLPAgE5K/tYMx2hJbqJF7V8V/ZHV9kkZ9TVdNkb
dmshb/78c8y8qs0pWRlgp/i5sN9M2DoK9NBuzm16i7s=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 7040 )
`pragma protect data_block
mwwHHZLhnYeFjP82AHqP0Lio61e79u8A7D+hfkgPHKwpQg08xr54ItDIMzsB2bDT
Q0sJc4DLz3vYXyOFUePNrUUdv/4V6Mm1YOk4rPs59Nyc+eZ7yXYN6gyCxlqkUmGf
oVpgy/U8E5LrrXZd0wy7sha6lYwVYP/H0dYfr/4Nr8ICVnmVvGsXMR/Fmd+cex4p
1gH2T8FHbYv050JQrrKShG+tA0FihSmR1NET9w3yH1O3/5p7dfHeoF9MUFez/mwA
P5N8GERgb7kjcoQjoFYv0blXo6shSLIKwjkJGg+lFmMFU54Wd66vnSDrY3BtJBw2
BnZCHtkO1nv3Vi9zuf9v5OlcpMMkA+9+TrsD5mk+K5bkFQEE/LD0ngbKARb6zyQT
XjKlhkF8YbllzaPlaBe5AVi9goGaiwPOQhAjqs4jMUL8rPBV/w4zdnqMe1DVfveB
SF9e+x/B/6Gpr/vKvcaudmYYtdhEyrO62Lyo0HRVPQie2Ua5b5pfyE3COd266k9G
SrrU6U8ftS+no7adXtGK5ybGgOmFvM9kFBKOFql3qqJatk82jiiWW31dY83ifCzx
KKoipKZd8KiUKUiCcnIS+1AyPDFyVx8z1fa21JnVlBdK2SVdeQZPZnlD3jU1YN7j
Z2sDkg5Z3EXMBVO+f/nQL+zpiGHjvEa6Sd1mq/h3OwOtCt3eXaOox3M/FkEnV4XY
jb8hqKnYQR8BFamo6FY61aQbJ/Ze8esdE5P0bJAjqwju5xJazBV0O4o/J/83KyLu
9jTDtG0CKZN+04ZqhUU1kAA+vL6Ob3pUK+/z5sHM/YmVBSG8RVwHZ4wIFh2NcQJJ
GroINpF2FCqif4AEk5GrlmulZ+oFI6hFjNpX9JbtS1VqX1LbZqZWB/S2H2WiFuqt
J1g//v8FCkWil3h94cnpvhoCz5VKjROkn6SqMsp4/wstt4PfFTqbjaSfjbd++EsD
OfKjt05EmPFUQKkVlFg3BKEbBNzh/vhkJfWl9ZgThF+WEZZie69sxYyWoPmbM+/M
fjs31Xs3ozqG1NkBtO+G322N+6ou06ArrHPt1jZbf/mZhdAd/52yQRDheeBBJunl
ja6E/jQXp5ek2iCCFix/tJju8Kzn5osSqT1PLqyYE2aPFpjP4BxoD6YbaUlkqW3X
OXtNT+UOvdTfwSWFVYpgRQ8clbfnmIoARyyKWSAxfeNjWJZW59/TbrKTWwVW3xNy
gVOCZKDL8ROFwTZP50pNpqUtPnYK0K2NO/KJ+o95yJhgo3QM6k9FgRvxS1w33bIK
MbgmI9Znfwi1sXmxs3hYQpNe9Kygc+LATMCoUlbybsXgWbxO+sRNAaG9kIgYWltn
IJZHnNr2AaoyoalX2o3E5AgO5QiimDGbVWbX5Jn7iia0gwJ1kFrtMFYftD31fMRf
YLKwAr1INJMzN4QlQm6WV7Z2K1q9BiHQGf7EdxnykwybTPZ4gNH6MBcU+itf5Mxl
I0rIP0yLQ85uLIKgBZpt7RrH8f95Ix9wfqvzci5CMAke5w+RMZkNLHn2nhrIHXNB
VnbaQF2rYfHAPq0cTHZtcMRffS9bmgVpB7mhyMl68ZZXO7w/R7SwRyuQs9S3QGdW
52ru5rtDdtPlD5sLeZP9Qs4lfPye2jSV/qrKg6zFfxAZlppc1UZ4FTmBs/WjNrYh
BrHNv3aj4IGEj+Bvht5ky1NyCC7U+bnaN4qnNj/GMBFyLNplI6kFJuL2SrU/8d/1
B2jtvSp15jMELOhOVQlXlZ76RMLw2MmJj47zT0uZKQCsdtwNA8DOWdOag+ZC/1A5
Tn9oPHgkoZBkhJwZ4wBOO6nxXzhHV2hycmKP1Ks6XUxco4NCCQW3sxAT68aAXfOW
+fuNW0XdIrymfM4NRX/5OYlBbAMueIcdgrtr0SADzYb9nZoL7rMMOrSB+6xKLlOt
9VkJYCKsr79ag9ShWfAnCWRIaeDoY268EpvwJcrAVYX2T7LsATpSWM5PuP/sn4hd
3pG0/Ww/13Z1mq/bFh8glHfJF65BahtEcrOiDt1ivvBVESapAaqDW5i2lUDZN4Kf
LCA5Xwgy3aFKObEzjW6poloOnv7Ul15rdylWm/9q4aFXOAkBEwNUg1SSwYQiHCj/
ouHQ0ibceBS3OR35wX4WGPcpsHuS3KU32BVNA6Yttxw2TwM6WzP3aoXq1w665VJ7
cXBQbvAj4S++vCxJyhC6x7TR6lQ/i0GIYKIjNzKaDHE71B2U5iDI14Z756qm8Jrp
6/U+BMdemr+DEo1l0X7FYsuLdhhjzbsKo1q+M9GjtxvasSYcNL/sxam3Lbkobwj7
AuNXjxDo8UrURSDUeiU0Dbdc8+cN5mzjusE4P8rzj4Pz6dTJJLEJQYGVsZwm8lI2
FyagW0/tqYI/t+fTxejtplBHI0eSSzbMCokhjcuyeH5UaHhMjbBAlcU7JNXG7JfC
aPkJIcBA+3D3sHLQsSdRqyto6fwBWea4tavVNt8dxiFPXRlaLkZ3uZwGxDYqpJk7
bJcRvRD3vB7DkjYwcr61+DvByhHcC5/axfIzS+yhJC0DEmXw6D8qFzwAHAL316Vx
CRlTiL5RFWngMxTo8wlHetzE/v+gnk/eJHsreJDzBODYcaZZF0VVftr5BmX431cY
0wlyTvehh28Ou/EK6miD2Br4O/aAxU0jooDa6Z+WkM6k55Rv9xVT47rUKqqvbw+8
6vSgY1lSdovOy5RIMhbwmZIQwSyL54xXYF+i6LUONLmhVFsD8qgkysxEOclSHsdw
G4zm+M0SX4MdVUxLtslwuMpM/IbOvjubSk+hYYi4jVJdVxN/LqG4in/e0r8ehH7P
67LBekOXsF8r9QaNhPbhKUY96/25Yg6BMsyXIj7Z1Zjvnmqy+ktFZLvNJpspIxMK
MfGsxKFYGGbZQNU6Z8EjhUa+rAw59iJku/Al1q6w8O2avSWxNCORoKyOWzxd2vh9
bTms8oAF9Iy+tfgb/oJ4OBilNZfAzjzm8fqqsQFNTnK2SIVh++HqsgAoqXWNZ+Wn
6QAOJbRnHC1EH0MKYv1z8zhwoZaJC6/d7SCohXQR3k5skt/v3jmPzg1xgRLXY8+F
WR4w/I04j9kzsHZ3tG0QZzRBcphiJ4lIjzXb+yQVt96qhyAlkifIDkQlWkrdiwsU
YNNH0+KU6ueaiXotbURj8WvKCX3aXrkxLoep3LeJJ5/jSs1koGbLBN91gS76Hd/C
gCEAPj+8h2QyaKFeviYTOR9wdDnjo5DM2vV2AP5Gv62AD0DKDjYG+R7FOqKp3gXV
tUVySEWijrGkq7staRppmQxlDGCGmmEuemIVlxr8tQfPYhhLenlpfaPxwBRhpvGy
8yJt8Omn2CPhftGCq3cyF6tY/C5fBTPQmS3OAyT8b0ceie264K8nTn9+Ym4aKpSM
lNHT+y6aRwJvLUp/DzJ5PfCjmpy7FenUnCRZVZMYiBwyGO8E4lb7ss4XbARa18Lc
yZnUq/adqnwcilYhmxiuVx3n80k1pzcWzqbLkWp5nB0UU3E4rNvNXpUTMe4n3mc6
E/EcJKpEraJHxgRLgCLXca/BnmwZfUNFESCj+PQTnFl72R4iub0l5MfoKMknzfqG
4RRsLv9gwtUkOGGUUsrDzEVYGXHBq9fgdjgCbAPs1RoSqUHO6L3nE6LBrv1xdE++
CBbseB22d9rsbyX3isrtUaVmXH3fqNZP/7uwmza8T7eBMM1nfeosS2enK7MogIKe
BqhJVLtJELEFgojZ9qHfNjPMdr3/LsJ2dEFftJ5/j8UlTDXAMdCHRrJD/jZrcBqA
YIrwI/PxQ5ebek9sVdozsa6J9wutzbOzHPz3EGiGI2enLTDhD33UzM8D2AR2/VWE
Cu6LogySPVQKZogKRj1ZcCNQVXS9X5JT0/8j2ne0zBJjRAoSpSbTk0O9RcjandyM
W1IF2n6l6eLRWmK6tGswSE263qIMmdKZELIME/znEq2NQG/SmpwlnKDTfs+hmpin
YI0JK0pp3komdvPUE4Quki/ErKNPykm4OuQp7gtUf5NCAyodYIpjuvPTtRfQFJZM
TDBGA3RQaZudID1IQvhApoFk+5zfUPwLiaDEJpQ3le3zaoTivgAmHh+OdpdW0h/l
mPeny9zF9uAkIVLAJKpjhfojiImUfK8qXA6ow4f14VrFlQKElqzE8arGXOIU4j7z
Dm6vHMti3QtjBQgtTWptAiaTyPFIFW4GtRC63VqU0t1TmILN0jC0gIcGbbl2ph7h
B9n4XFAFP/ctMlFEe67oeBofWaAHYAHonEE9tpZyNe7P2t2zB//lNw2F1z6LQwyP
4tMhLZcaJIFfUIyR99iIgWHWzton97ku+azRwmUUXuPzTS3B4aNGL3CBj/LsqckU
Eyoc6lj6QGA0/h288NTBGdIimT5QXIvwAFU4Dl7pfR1gDFqiStsR8HQE+QHzX3XB
IecW4CjxP8VQZSrUezs+fB6gwUeBaZ1lhd5qzUtMcwFtCbvtWhRyLcuon6d9lhr3
kpyyg+21Aw1fjaqAPpeq2T2SCHMsQxB/9ucYdAPhGubIrLdmDmuuk5TQFLrcWfif
kOwyTeszUT8F1e9w5DPBFiYZ5wZRfx1SdPUukgE+pssctQDlC5ZylMU1PXnhflrh
tHhbkmJnflp+yVNwGueM9HSxq1IPtElnIMNEr31B/5blQDBgru9XCdghE7r6ngI5
6SAYOBiY7sSVHnvER080q9CvJUyRcIi+DG+4aXlhZajYawP39C48IJKjP5jGFrXq
7UW2H0cPAaG5SXg/hByLPnxL3aj+HYUvA/fIJtfqisEl0vjkuNLwIPvCpgLAaK5o
kdpnAFp8yF7yQrfkHwkI84glqZ+1FzF522YkCzmOkVBvjWI5S/u5WkqLk1b5ZqM8
MSlh/WhuSrKfL/tnMnwRbRJJbSDL9e95svRvWD2/uXKiZIaC6DT3871P8qhtkcNI
l8rUwb9fSAon6l/a45cz/g6mREIhcjpKg7Zpe+cvjNuWtx0Zrx8JqX31wK6NNoJT
vDLY2Z7buNQOLOJzRunMxGcmMJ6ECtQljgZ1NETpfPKDpmakxhRFdzPia180xO5+
M+QV0voGYtVyA6KoBnvdKl79yNnIi1wSkVLH5fA1BETupHemjgS1i0BrPRrqNCIx
wJHmYIWYTulH79qowTtJV2mCCFpAdb/aOf9x72z1a45H9XgfjfOc40BaQTe+Qu++
B1bCseyie4K2S1JixTgX+PPCPvb4OAeEYjstxVN/zZCYYHeX91vOn6jeb7BKgr6W
NE3ctcoySO1rgeAzCPYAWmVslhyb0xPA3H7FD4BqfGcBh9l0rGLbGv3tEUtR8gYV
OhZSNFVL5/9jSs4VHRxux+mYWB9tg3zGFhEnVPoGtr5dyakde+yBhFV7mCXibrw0
buajG+ANlRX3laHaWsAnUeyT3XW7BVMKZDKwG3It6Tqx/ugfHyrH7DH+0urcGlhP
xXtQnZ1WQcJ9DecCVIJ0KkWAmz72nE1iuXvbHgGPmzKxqcdMsk3Y6RLspNVDSQ8F
L8ZowWxv6HuPDfH1jKpVx7MZrDI0WIaYChCuVcO3fOgGBLRUeT8IF9UBxPYOarZ1
4kCeA2y1P7PBUYyv/qxR912DSjIl8HszVcP7GrsHUVpcdnW/DwH0JWJ8GwODtv13
+kk2EwLdYr12FDPguRclhRJ3uUemSVuLK0h13NaXZqgZFULrx0V7O/P0Yi3yxWVp
+npLNfg8Rw5GrR+xOzog5OLFK0fEpNs2wXPzZsUdsYxFVurFiRSjNBfoJlFbm1Ny
iZfIS+nMlOhTJxLt27uuJR8zvCoU1spC/j86IN97qd6TXJYF6maWxhHg8M2izEnR
qA1qWwDWq9NvcBPfMrj2+L3YcUvuJBRGoX4GhSaY6vnHAUI7aJaWxXDYGWggI297
xODTk2XntW6IT+N2UtvG4Ma+JKeqBSbwXMqzeHULOPEoW6V7DuDRBg184R3WtTfx
wdR1W7sigAj2j6toK+nd5MUM+xh+T+Yddz1PbKjphR0v7L+evEQe1XKSWMdI78x1
T8dW4oct4oaHdZvD4YTtsLrhekO8qUa1rKo9e6qFLgfYcYcrf8EmVOneeG2KLeAR
LJzAoCliBAoCaeTK8ezZVMgTf4xbC6v3a91S6lyoQEsC5qNNOmw1FyGcEIE6x5Pm
lMXxFhO4v9Nr1M9lWxbsbeaxefVnULExJImhP1CXswNUFvAmrs/LNTHfNt0TL2F3
1dph99DKgtfPLD33aI7XWHR+Fr/i/Q2OBE9S7z0wHQSdmdXpfh4ssM4mJEn3m/36
1++KMvbQsiLLZx1pVsTXS9nF/sz3VJ09Yvz4CmvFgiuQSnPZJrS1aeQJ83KLiYtp
EZYg/HBY8UFAVGldwPXEBhPkbFDqsGh0wQyTYff/iEmF63rgI9g8HaxDC0ZrhS4e
eKYSXy7VlABUjZRGQgTNynP1GfXiOyYiJRYoSDkf/+J/T3O3X2lnpWy4dRveq4M4
UU6LBrY7EDd3vH2PrEtbO9F/FfwGNA1QF+LLhY7A3OE49GOPX2RucVNjA9NeRM+3
GvhJLAkt4SFCG4HVfIthwgRtjVppotJFfLi24eQaaMdvCtVgbYVS8hUm+I40TdcQ
wxbKR4P6U6qSQPMAEgXWEZVMQ1fxTJRJ8mxXO9M13oKdghYY0JVmERVPIsg7iN2C
aPhSDiH9lyN+4jvQWviiBQ82AaQOM3YmbDvqFbdp7KpA59ANaU9HCoR5PK8HfMaS
3NOB2V2lDpAAejeD41xLziDklgU0nQYITmOpr4QaKF74qHYkr6usK0/bacz+yqMO
He6VJPCAA4yWj99cO21YdxMjhMlQtgbBlHiXoubbK1WlfP6h0Ar3IZdfNtEoDCIG
pti5yiyg4GMWSawXJHO8kXjUGbiuY55Z0ScAvnGJ4JI/orqhlRfeCVT88SSRyLJ9
hKAuctTmkw4dGabwWIT+QXcb/q9hy/t6gcUHuHB6278K3+8VklDHBPPDXT2PboAN
QdZJHwJRhV/w3baMIt+/Zrn5NP3oB2Si9y/UKOxqIHOF7ejHBkG3e/qD34sqLfRp
kcllp03MW4v/SOzfl4NfHMNxXGxBC8kjY6bnI9qaLcHt8a/N3sAHQETmCDr0JUgx
i3nlDBYIKI3OQp9fd09QfMAmkFF0qvOBd/zQKVqlLLs0DFsNvM3xflvKC58Ua11q
myJEXgdgliFsffwvsrNAfhoCRNQau6OqIcgFdCm2a/TXCnoJQPXCC1YoKmybRreb
6L+igUZIuY59P1Yv3YO9tSbYlBNDLuFH+mOUmOXvw0fan6A8DxobBe3TbugWyWzO
3mv+kS0NBbLjl4svgWzC397Je/2JtcQCa3Wx2derPvUL26xbDeI4Okb43Cywbqvf
SZsg318rcVgJ70NOdOfJsoTK5V6lGst6D+Rm4lO1AWmMq+yTsozQBQ+bbVdPahTo
CzZmA+/HowdQyycWTk2/z1nEqtNWs3Xg24b1Llz+7yqEk//UVS/ujsseFUV3dFkJ
TvDbArvCetvFNCuyj7fc0nZsqtLpG4qDqn2w+zyodpGtdJalxbN7XppcUes3x/s4
kmN9f8zfiwgyytOQGt7v9BRGdrjaFe4lbWEZuBC6s3eOpcd3cEtHMM3uxX3WJbCB
dMkNQFEtJlouALkQ5Ol8S6TpEO9kmdWSJmmFV1on/SQv9lqZhCRRZeSGbTgyYw9N
GnWwkQ2+lhp9mqKsPzHiNiMq/ABKPqgD548OTGcfgiFS6iJGHDfpiIOYGWBfFr/8
u/Zp9S5FbMFIOsZlOqoj/A6trgRvm9S6DPeL6kmbpm3B8+QLqSpVzLwoaQOeJv9T
PEc7FXT91BDnEHAxLoF/acxvrupP6cr0oUW35I4LxiAkqYN/1IkTg1bRvm7clcLM
RlnpLr3K7g1Jwl4IoxqbfobevPCBUA3YpNtKSm8WdrhrOCEIUvsZTDRfhaHlWdRM
KUEkjDSmX3ajAcAjiiaiV33GAyxqz+3faiBtekBMPQECau4X35Ca8IWovCbyeVgt
1SaEKACINE0L0ibSFZkAv1YsK0ZMpiPyYPjMWW2aAhkJmqSab0h/K8xTtRD4+N+c
L2HefNPi2hHYwk1esHAQr0kO1DLTtj5SkEsE3f/YcqUESnS+Gy7RZAxnRkpW5d05
r7F3iu0kJs46aJYGc4MhBvATCoQUOhjFOcrUcus9B+EDylrfG9tJ7xWcReHbVf4o
Mo0a5S1Pazg5yyVwPXUaWOPp/4bu4NLNWiJhFE8Ls08Hms4/3p2O9B4Q/Dyc6837
dbI8lG2mrNvPe8bX8XncitLenjq2hp/VaPttwwOpu2CNd8wyIQPE9XOj8vYUM/zN
Z6aGwZwRA7ZYkiaPb4n46KlRPZb70UBH9LCSDgy08+VnkUjZ73RcQ726KYYaPoxW
Cinp3THiJyHzirmZy9eBJhKuwscthaa7AkDlBJmeChMpYWnSLZwrSABVV8g8utTh
hDhVOGRRQARH5Zh8xpDG5NamjR/htZYBn+X52Zm76gZ4vt6CfXhzxdS4oTnfzJkR
Dk+Wdxz8AuRkALD/pRJ8SCNfZZoYQIWkr6+rtaqhEcdXbf6NPRrQUsgFWl9K9tpI
e9xywl2qMNGN+7oRNg4X3eWPRbmEz2aoMrnHJl56pM/cyqzSfVK74vkQ1tRY7+R3
xwT9W6xBL5aFCr/5Y2FXzh/ftjuJi+YQKkUFvk6+k5Ys5mEBboQOHIj6/usyEFhq
P5QtTlz620EC75gr2s4XAfd/60D+y4g5itf5IWpOGdGdyqLqM+pikR1BpFJumYek
L4wGUtmtE4x7jDDrF4T1ZwGkixsAURkrcjNS5cQFFYAGAOdLM5o4AsCb4QXZI0iy
rHRsayHbC55VWrj4hNrbDvjptgBbM6cSmAFgZioG9lL1KPKiOwnEnXjNsLmigouu
fk51e+4zReqQZxtuCFywTP0QkpFcIsLFqoAYMV4ds7yjxhRb6iw6WZ5ffx7BsQ7l
jVwCaq6AR/vz8uKX/yookrE2qE/i7D8OSaL23+hqwVmB/+2ZlT1I0ZUC05hahJ96
1izMvvi2/NbDhKFGxZVNyxfn1eT5IQcF/xN3rD3RvfDmDFFU68H9t50NVY2S5khJ
pFwaSDhav0BalaQUlfy1yJb4zY/7ofIYSDoBAXSo8vA/3qJATSZ+d5drLKf9w5Lh
Pa8Lh9kjjqCV+zQcFhYtaRGEclP0Cci2f79XoRe5pMmNcEWL2BqE2Vt9MgXNRu+H
Pp9YGzgoHfjN6ljd3kek5e1WOigQdSCcJfWSoVe655a/ObeBp14XKOuPzT7F+GMc
4/+NS1EREagakg2p6qu02rlcuGffeI0jr7N++w8Zjer0HeoI2RvHHyy223XZYfuc
8EV6+INh5jhWibvgo5aORoMTx54ZBSifSd3Z2knWnWI=

`pragma protect end_protected

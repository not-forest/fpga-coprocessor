// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
odC8GzSKRcwDcw+1myhTG59hE8DOK5JYppS6I4KmybVTb32xFBUDzHLlF0cMksiMX01q8Y9CR4p6
6BZv5pAXm2bl1EsctZ1wxIGvtNyG2ijzz8gROXh7wkYzS5v6NVeeeXuBNb5wKG51UOu0Lrf3ynk4
V8012HgVHD8HIzTWdvwpo+seH5pMxUyKi1ofIoZKVvgKV0zXZeTSP9kV+zATB/iFvpJtg4Pp/YB1
u53lo2YH3jlJcvAMbu4kmCi1kWHiwdX6ZswkqjwamdRbhmknj/pJo4K971YzBNCPh04Xm5g+IsHP
IwISp1/a4eVdXOmATkGvMvTCHyzX1paD0Mrk1g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 22096)
SxsFHxh85EQsVD34RoeX/O2wis+Vpm6i3LS/zAOjs5lAI0/1RYgB7+ic06iRd6laVa+UVlsyJrIn
KyKvb2Z7ollJapkfC2uBR++f4y/rCn3TsjqVkz1vAP783j5yLxPZwNTqsnYFk5Ydr15ANbPQl7fx
XLE1ZFjSxS8r/E3tJztRmk/8rVOxTM0IvxPZNB+hePxp+78Cab9AebuEs/0RFcCSsRdA2c4rXTeo
rhK4Ha7pw4oxZlSSt2hgVgZD2S7ki/b5+Y/zD1XKBmh1vhGbl9+P8m1q8gMAXFA7zU/VjD/uPzV/
RbfrbFl0W2O4oZ45VsqAEUfANt8n5xe7lewR4OxOjIRmQDYVBfQH9RiBzgD+uqF5A48hFkGVyK34
x+ZLRWofFYD5P2Wd5XQQYIUoXKn8tmtjO9FXp6LdIsSSXLdd32fXmn1t8I1SldHlOBD69J1G/huL
jbQmbEJwFZPwSIHh3eDccF89FaYAqrcqPNbmxhtBnK/j+Xl6NX08SxOUwJIbHDcI+QanheKtxEDo
TSUAJyCQaV0VvEVIZbRPpolZ34KtdiuoeHpZ1BNq6SJqMzb1FT4WPPNg9lFRxIevKXpUBsIEndE9
mSBWUdrpm58mkjTX1el68gOacKZK0B5uAc6RGZ6hz1pTO4p02gxRD/AOlN+/2BOwJ5yQlraLYbW8
t4z+I4B+2P3vZtfpH7l+FzIOmMwSH0yy69uRgpDgyGhz082z9Zr7t/LhnNYisi+NZEDOtowtwmoE
YKojiHagljIVoGRzoW06WOc9kKkerQAmZmJq/hgvSM74mZij4cVSV0N28LmmLB1VkzwplXAvPKG7
ySvQSD1Ik160ErCGH5uoWNHOTkOnmBtHZo0EMNpHC1kkaVdWuFCeJFnXnwwI3kPjduZqWpiHFzfz
AlqBbzg/0fJr0njpRb/l51sYCwGOn0Z5hs8jhWnZgLqrTYqrkOg6cKd14aHLHez1w0YDeiFRW1GB
EfQ/wvVPwcOKuflWpZJbv3SHBHO/EKnPkPsSetCOsJfOmxJ6nSH7gV9DToID/6dhv9EGMrmQgh3Y
E6sU+zWGvikt0WGsrdf4ogtr0ZPsGeLBi3/VG1fYXpLdAM+dYTn44//cSQoz9lEazc8eCW21MN20
QUgAL2LENQb5QHeODg3ST9uT5wdyBOiQhh2reOyLMY4d48Jldf0VpaOq6ygTna4xE6lBTBIbOuYo
UeHCkLVdZW3JNqSNjqG/phVmQ+TJnHyqmqVH5qlVwnpTPIGrtSeDX6L55Da+inHA8g7sDfUEa65d
Wyj/riDZLjWhe6kAwi0nFzdlcFb8lJkkXEo7cdyw8YWk18X6tAVsgs1W1LcNF/QtnbafNYTCE/0C
C+GA+FIDHxaYaxxg1NbAkTTlPxn6+BgR8JQshiqLGsgrtnD8YK8BLoQdB/8FuemLYvtXkWkfnY0f
zYYIp3A6p4CrKB7wSqPov/BCQIjS8rEVFLYGslu8eiOiw6C4OnpH3dhtp5/XB2ccXdvYnw0KQ9Fz
I0HPpAcgUN4YfPyy3S97PVkdvut5C+HDxjat/xETAifVvRtDEv7ymSpbllbDp1LW4qSr8GhzNUu6
IC1ikHzkiVBRz2MxYgKspWARCz+jJ6+jfT6Mf6JYASREYNk9GkuDt3L0RUHGvI7rM89H7nNQlYy5
JKTt0pxcdsDkGgqQH/uHi3wYYlWaB76p6wDPmGAjMw2ULyyTLYcfVZCXuz9ZYUsXamqmqVeS5mcF
Fzatw+RP4Z/uiA9SFhOjoGZIfTDXaO2D/vz4ANuQZAPoQjsPl3XklkO4d/7dxqmu/YFII/TB+Xog
/5j7gA7UV61FpLT0yTuRVDPeLUX2bGzFD7dT4HSCu7Wy6LUxl+6ivvdrEdASlm/uCifEW0TcJb60
KAvRwACeJXPOolX8X7K6cH5QOI+zMkUOUT2+g1Uhym6CRiaE9ANb1BPdHPIX+nGqtxdjtQSyFFvL
QT1GqFSORSEP2W9hcXtKSwFMVwUM9ysHIBhbtYqNeW9Ss8rawhzGsQWjz5QJz2z20JMhfYniSCIg
mOD9eSa0mnK8Gf/EYLMS4ILbgYOJ7MPbp9Dvm1qq0dIS3emTs0xW74UfBE+IcFaJkR6i36iqrUTJ
lfrWr27NI8AlknmRZa04vE4gV/6vQ0X8h6kZ+H8HFPaU/usQebawTV9GSp8PoxmxKCw6cFltBo9n
AZ7rKfzd1jp4BM4bIiKprnHDlnp0sZsKkjs/PJKpYUNRW/i0oZ3gXfPqqmwf6LFgjF4H38SHt+yg
FalJU6XN2+mVtiyTQSEf9eINwKBeGqRwZAaNVBPxfUuz050X1vseaEeIDTvZXrd2mxmEtlpaFgPS
aO6gP10bAU8RgIETMkVDnlz99DZDZgf40FGYf/N8zQR4kxVEG7/8YIQ81/RMAx3rmxSWay229Hy+
lBVL66UVIYhhSx97lYDwPPh84QDDGJDSEgm9SWfsmBfj277oyR1qOeRZLPcajwjbaksBNBETWsDQ
2RXhIjyZ/uynWGjtW+XZ0f1U29iCBZjCVqLnlJ40on/aaXReh4Z0RdvlZg9mvCQcV7PVFc6L5hvI
oY7okSK9bX7bDeiVaBgQ8u+xTSeWuI2co0oDXXIwlhXOpMIf2c+IatjL5iJii3OkJvcVldfOj0hM
sSoX2tbBTqP7nlSSTdiY+g682OOrywZG4vpDwJWF0uU8GKb5OiXPK8IwfIA2FyXj8CSqRIvt9b+e
HGGPtWV8Qq4wBi0Ce12Q4ddgSi6rfQfXIN0Pd1ShyakXDDxeZoaGGwPvIa28hJx6l2WKIyidCyUh
v9191Qdji157mfL2CS1XPXO/fq3aLOnZDA2wPLD4Kz/Y9/VqqEV6dAeZz8CSI8gK6fsnjqci7Mvs
YumVdhYIb3bo13UgIsEoN6j6tksJPx/3gJWFlJnGWIW4irAt53pM684as7O/cn//X0JN+B08JMDO
W2jyaOIkaBmsSWsNU9whrbFAWllaAg4i+UYp4nLSwI5AadlnTmuOAshQ88mimKbR2S0JhNu+8RlI
Fxb87Qw/xsqYLfCVVZI/oIYmkIIBkDgfggGe7NuOiskZ//wa9VHsJ9j2DHDbC+scUHrlAQrpIu5H
JF8xWeXn9xvo2YRio19rWwG2UaM9PEWKPkaxwmQ2cYVg8MxO9D4uaGKwAfLSrohggKZ3sQxdVTbK
mR8o60RluCfbph5DeQo80VjsIc64X9xcdEc/NLf5GXnaOIYeEq2MQUvN/oTqQFijgIp2SQsuZLvq
ETDYWOu2aHeHJjQKEPZMisyfMHuKMt7HCub0t7II1bxlp6xQO0k5lSz7F3/o9/MLCZ3LKXi9PwIV
XOk19Z+iY0AK+yoCJp38/T4cQhYU3EbrD1S1rdcswnhtVUHVtWNsDzMQn05e1th2W/RPHTX+e1SJ
19bA9eD508gFNbtZspZIQG/sXANtd9N2bTRvu+QcXtRonqo8nGrX7UhQpUcFpTRds8vv9sbjWiaR
38WqgjMpTXnB9VhnjvQhI8baTHf9uJM/ppIHBKcxUgQ44pZ+KsLuJPBYu7G9hzFUMTIJX3c6ccNH
C2SZ2gyrsZO0LqWuUfybp6yqoFeeylob9QgIQ+AEawJ1p8o5i+J130trrK/kHgFCNGl2ENBLA0M4
bYHawQjTxi3VavsEgk+HKmpPb5WFWiZtRopG1ECON0D9yna4oVVv+gtDlTUAwVvVf51uUkwS3icQ
jGWjgwF7oaqLfHhUBR+RFZbpVVXrR1Eepb9TFP3fcABy9IGScycX7fCSutYbf0UZqBjow8HdVpka
yFHyjickNrbI+fNOLV3jGmT7/DO3sFIqhrL1P2kRbLOeugxvNNqIlgGhhS5qjKHElRBpHR8Vy9pS
R4WeEEMWAFWbm4eBhyw4+wMaB0jzNelVyDAmqpWM+sXycQMTPBGzg7/QRhysx3yU8LOyXJnYVZtF
rPqweIGLHoCBFlXyyNWayaOVBKVSZUSCGgzKex8McyRabque2XlZBlLm7QWr7xBujmN7cSsYNFIh
JIJ4AD+8TEpPeLkWidajNFU6fYjgRlNDZOdXJx7NMKYRWB8vonbV9U5mE072MheXsU7NyfaWOzW9
JT9miRmmANh98nUC7IryrVUVm/ewDMUAyFBdy5d2pkbbojO5OQYNaCE0pUGr9GoKk5OswHlOgs1j
QkCaeNPjxY8jhGoykaZrDzgv/zFRfRQ49IJaZEHAmJb23A8m4AmJXM4LhHPaaLZcJgxvITvVF/a6
mA7gwfMV6nld1eizQs5xZh5Q9tRCyZ9kVr+aRxe4rQk+9QopuwxYvOFyWVOuriwGOvQvXKht1GnS
7NBUYLG8sSkgT0VnD6gaZGg5kCIALHiuoPpEYlnKUmvTf/IwhE9KopIrGY77cIcR+nWot1GC4US0
O64lJZQ53tBQyQWIt1KNpYtom32ul+ix/fjXfY+KeCzyhBS+kr+e/Zadya78smybg67c7R/D7w78
bNx3SZhyWLmnXIxpt33RGKenPmP5ZYWatoZfwc+aeisdE0Vt6bEx2SUJwv+Faa6MqGKNnFlcmqfi
f70SfDJA5rLoz8PF9Rqyy/Gf+CV+DYajlvgyCOwQkegQBtVNOq5U0/pi7K/3d4508Wim7pnioLVc
lWRxGWx4wARP+mHOCR/rVjczf31fLmGxNKNMVmg7Lpgaf9WFHQfclb4cLJaRku+JWB5s+fqe3XFx
H4jTCIm3Dhb+cH0/UboIPTsus/sLXqpJkQLelUln2TEtwsXrb4NkLIHyqCw5WkUdUYUyfiIsa2AV
EZOJYfEpM3z5rUKImaLDFsyM2XL1ObKxpVOLa+Up35j7EZ6HlLL0uLPWzZxid71+re0cavA/6jid
KM95swTC/tMlI+/4ThbUR5mPUFllwqV5tym6C2va9VtBBdH2RX+7cyeOxXLZ2ygof0Zj7tHF3Kyr
UD5L4nRyvXIJ9o1wb3VGz/cMV7DhqID6n6RCn6KsJTeASTZpAKp1oD3DI8TpC8gy7W8Xud5iaGDz
ypx9S6FyD5Fd7Oj4PENr2pIpqyKKOpcuNHaPz2rZJJH1tLzX1QwRg5z511x5liJtrBWTGzVEkVg3
a2HPyNrO7QN63Jx600lITfgZ/xzRgTJ6zaxuW27LdPLZ3dpb8G8d7nU7V5GOxyEHRZ37NdcdNKzR
DGQdmtTZOJcmxT4oXiFwgPCDKtpuBQif6PCetpTYlQgqYYQt2lD4gCRcIPeJaUQB0Wj1XkDJGj3D
bKcsXWoyM3ReiSP9Yzz/6LnXbKPzIP7drq44zfP2Vm1wVJfVb4d9oGibsw3nafyk8fvuH2a98TDH
qXkm5j7r2iUdMy7sgqCDf2YlWowMnpISof2xmpOhpei+IeeDbTYc/gUEo9ARHT481kq1uXgQpcD4
Oaa9101B6ol+YkAdSwhqTn5bNi36QeDCVTlbq5uI62y3MGAc6NKKqf1uTAJcxOPp+sudVM/FlEJB
9r/UDgnsZkz60YoF07wvHWLz8Rs04tMItyEXEatst6MAa03idjsLWHCg08/GTUAd2Z4kH1AWBBoJ
tqaaTI7EZZZdEvGa9TOylVpo+yMW/SZoZgXq6+0mmrXMd+nhtCMhMUVV0yw5taCXsgfpxfOPssa8
NgQYbkJfR0R106wIJhEfsELmQhYzy0iWZ0KVV39KO18z0CuG11ozI0i9qOxfYoc7uz8gYkJ8UTpm
IOQ9r0zjQz21wffTguvhXH70cWqS8qsL09jt3AYG1S4RdxIZf1Yg3LT5ECWVJT+aFKUofbBDCAVQ
hn8DjmL2HOEeo+7BDcgG9tzohqfhFAplqEpZf3UFAJdm/HR/J2dg6j+DePnQk6vbkK+YJCGZzDFL
MJXoXM8ghbSAUUzc21pEkwQmpgvvqhYruy0etikqa6AgbgWsm0Ry9uiAy49tjMhWTlucPbPa34U0
qR/BcAHgD4JhM314I1CV1xWuu8+UhC1PIDrURGUEBLQb2pKWZONgSNGYJtragAMip4qLA0urNR+S
NekM1IT/qiDpzCL8JZXTOjkBr4lNWnDPGfdPEF5t6A+apBTVviZlNSy6rQXM1ePr7iWXv7ja2RO6
uW4fe1tvmMNhZ+0ijhXjvZsHtkiPsfCKflPe5R+t1ZKyvKEQZMzi+ofEw5J4PK0gf3GENy+mXkho
1GkEXLnCb9tLv+o72b96PbC/OUhavMCi3rZKb9B+7vopznZdaY89eVli40g7jtvmFI9qf9TcEfpH
E+vexwjadkbAHzA73F97cNzG026lRRwysaDpRvIDgCO9a2Rbeipiht/zhrUrCDGFaKcsPXoBM0Dk
YidSgXL626rz48fj+RXuqtawjXt2gaayeaa6zcF7COB+bQakKwbI9Wy2F0HbzLz54nJDxImQ9MQc
HemDJCXBCaYQREKYopHzYzYtS9521NsNKvt2VD5EOo+xDZ+tYtEIkiQTwKGd0BbbyzeRt+tR6638
i7QbstSd5YoSNhLLPWmJqls3mB3TLPA6m5dKxexvqyfQg2M7sKsH09hdy7vvtwzPVBMRBN/oB866
l8kQEhsghf8o9ixkMI5MQS/EgWQkGDdU6ucfbtR6/8lUZFEJ6xm66TDA9Rv1lCZsP8RzF2aiFdV3
sJ1GLXwzn1qMXjpKPkqiHRGuLkycC8ifgqTmKZ2v3GB4FsxRmnngrMPUzWnIG+4y2c+uWByUZtgS
gf4RiATPdg7rx2mYOpnshVmN9lbS9PnOPN3eYe02rLWQQbF47xxNpq7B3rhQf2bzDcZV4OOj7RsM
XHk5mdm7o4YNyg3J2YAn6032zNxbmw8u0F9lYW+dbMFKqg6K0plYJ28t4rmvfjgUThzkJqP6EMXu
lRqtg14vAHYA0trXZA4cPzEJ7xXJR+u/qOlRV/67xu6DwTp6QCZVM1X3ccqqK/KBrmd7WAoM17x8
Cmilltw5vRqe/b2inHQx4KP6wDZ45T1pvLUAQZ8/JGMz715t+Imws8LXOhP7xUGTfSjQMGkI74gU
LY0hwcJujeIXUua2cWAHBbKyA+EYS/HOyuKux6vTEbUPPn/SGU80e9w1+VB924kx8sp/7EF+0s0O
fciAnUPxbHy2LqnebwgLeXYA126INu2AoXxPRRGEbkG1OK2z8fehWcyG+n+19QKyErJfjhTbbonm
U8MjQrbuihL0Icmt3WJLC50MpUhyYM3VwGgKTbezuaWdSnkvt1NPw1Qp23IC90ye8BZdCBlnhnwa
bcuRhuz2FjM62KWRQhujDRJGd3Ln4K2niQpY9DqdsK2QBQU4dA2MzoBtgSAxZsOmCBII6hGisX0F
9EdVKIfEMj0wPK6JrdINm7HOGYhuf/3CpI5IlaBws8oKc+ajXKl+F827My9aTgMASAKMAqxlCYCu
Kp2+euiC2j2H5MnlssZvclthjiQceRYAR2cbXkAsI5jHI2lBsfceRQJx4oP0+HdM2tIg1b3/g6nZ
VLftrVsYlSP1pLjPmGkaUZSthvHiPNTgMiJ8RznkNqZ6RBG4iVCHWhFmF2kgp7D1NAX1HAtaReB+
iu13xrR1ZxqPGdLfX3/aPAki03g0vPVhFkYd+LnX3pUQblte6Llbavjwd+KV8HAPvVK6rVrNvm0T
HoW02dcIE+CCV58R9/JEAQ1AbGMFm1hyGb17/dln9rUI+BJwI+5thn7E6yiidPtLw9JwFkBw3Ugq
iwWD3L5Lx2OVBi/yADPgLlJhNNsEGKxNGX7lxcOVjtJQnLW2KvgK9z0B807qBYQG/MPElUh9UdT8
0yh9mJVm56vz2vXOzY7RvEgm7VmbRlN4Z5j4XCIh+JBOM3iMX2x/RuqBk69o4OBIFbHKu10EioZU
5st4jSnYFyLEWGGfwpYbJyc/4FzB1gLOXiArcHakgI8K1iQFmxlYI5UtgbcSz64ZOsYZJ/v4UroJ
lYx24OmD3a9XkKlgsPtdQ8DSLYGDugcnUaeaSSytZPI7xDQgz0zWdd8mHB5ikjaGjUMb90MAUbhz
NtfOSJc3BvzjGYEjO+3lEIwx02UAdSHbUwlIOQeIiLYYyppd28rkKlMCuuRDYRUEGzO5n20WeJMv
vfk9aosv413EXnmrOTaZYDoBwa/B+VTzjRo0xczpabe/nbrpDiZUnPlLAwv57nUaOQKYS/VwZJjN
slDmvMnbTsGrFA1LptlYWK+ZRHraNk1SS95vsCvrB6oKiDUmsRhmiGCLUYFjuAIOO+zsij+z3n9W
ZgrXhkNCuslI/yGRUoGcd4XDRc/0cCVYWn19eRgwhR6q+58UJyzp1M4CMuAu5tuZJ9LfofAk5NNh
2BpQ+HEZlus3SNnBbmxPVKJlv4/gyvNqqkOSf2Z/+m6zNPNMtK92lKNBV7CultH9WvsV5QbRRpmm
9sd05ARszclFkpnrgsQM5QA+mxjw2lS4Hfe8pk+CdOcxBFZb76Azqco/FwlchYwS8r2sHk++JhIv
ElnHC0u4v+D+NINGP0NQUhqgZtGcUeYKhKANFwfGpYzvI7QNMeG8pZvBsiJwFpnsJDpPQDmE6p+h
tFLCrY6CyxA5j9jys8z35ZQRQctBlhzJmF6xON15lojl2bmcndxq6erxnTXbsuJWzlNk6HVnBdH/
EidJKbFosJszO9wD4VYaxBMRiEFPBStjAtk1V8Jq79K8T+e38xH245sGMZ6MBwmyk8SeY+xBGUfI
s32erqdCbLobAMbyMrgg7AqFoTyqBd9hOCzehQ4cYIMmFnCk70ZRdrur3oEa6YaeBaaNXXCEb7u1
EEC0zZyPLBk3Z1+nY87loi0I7i4dWz7PhZMmhzPK6aeV8qflY3vQVkkcxPfI82qHJ4s02ndZuJJ8
hUugaviNYOYDSv8Edn+rOHf4MLS2FF/x0IdO9hFVHh0bsqvM/llXVGgMV6UEXznNxw68wCjNWmI5
i9dJJL4xrR5oNp88irE7aPK2d+AcxCPQwSCGvCZpFNtJxeIQTbhKq4530mkwxjAhBms/kXmgQCp3
xQjAhRnL7ZnsceTitVUqqNX6RBXU7mIYdT5j/RTu8vMaDUDevQ0tKyOVQohfRkjJjy5MtMl+tO5P
eE3wYK5ok+E+cpDdaXvN8B6087FtrE6XucvFtAm/hXBgCl1brhXbEJKoGi2GblrzZRAItvqzjrrV
6TcRnhggxa0uCZyJQ84gEE5WfUrcd+cZ6UDVhY6afhJrm7okPEjaocAzkX5xzTE+1HUYWiiRCfTS
CpfbTYcj6w6OMTOqUhvzYqtkLxOUhyShm0vB0Ma8Oqd5OXtXo6D/LgtpHfhF99IRd3A6FRaVdZzI
X9iVEFQOwGv5NOidCWMHT9l2beG3CMaDkgnK3nY5K3r0hio59/AOpEUqjjq42xgLwJIu3kpnSvoE
QHyR+5cLfYaLDTNP9QsdIAmoMZsXip0COROzhQsmeJyfGigBHImowBEDGlljuwktQZKMGmqcEXS/
8zqB6YRefGmUPGA+6fr8WGZISe0le7wHJTX3PMHssFdSb45b999DWjPzbUW3C8qCce0i843iIzNA
VY/l6/iuxJx48zYsRAEuJrZstU1Z41DWDMQbJX7G30KbEZ72/47WwBBCHvk0u+orUtbWBpDaA952
gASk2wXSxcybWtVPfBtEj4XdExZ9xW1uXqpSnXRFXcj6XOo4LO1bn2+UNRXyks6N/HFrci2sJMhf
ZHFpddyycAE39c48z6gZaJznjXyS3KjI0uz2wUvGpexJqkfb1CTyxE/L40jL9rTJVhaVwBMS/71l
t53Yu3rDhVEq2W1CHovaw7X8m8LYOeERbXUH2u47BKVWjkxLlvJB0aeUPpG/agv8vxRzlxK+ja5v
mWSWfjV3squKV5kqQoG/ytjNJEuvxGFyVrYoAHi4y4yobZo9PCgvktV4Tc1BGh+qOwfHxmla5nji
XZDLzNqU4PY2NVmw3JJ7yy2W5JCfCW4uDft3ghzC5Ij+CiZlaQLGvjtEx2iEdFA3jj4FobXkEepi
DzlJx3yfd3wnXyLM3/AHH9t2ed5YDJGVVrAemW19Nidx9mWTTyXpUGrkTSIMgBx+SkR+VZBXnv8F
xav6UUbir76gPrPHypwFHu4CeQXsyuTbhXwQGpsHgNxI62eMeMJJVtN4K/g8BjhhhtrlATcOwSIM
REiw7knloxaFMGGED5qjqL/GmDS34PWmCb6tv5p648bxIlvvXAsIs5AgBHA70lzRw6SJpOGM7EHV
byK0rRakH+IOKGU6uQ7sZ9Fr1QBSwGVBrcZQVZk4FyIeZFLLEGszE+wMHlGIZQ93OL+ZQLBpd+1+
ZzHQ7OMqbKBNJ2ZxXqr/hjWaIc1o91wylZy5Y/Woo/4cyjq3DOCnEhgdSWVpfDHJ407tei/txS6M
R1zNfxEYiqkntbVf/DZtC1xlP0+03HE1JfRpqH42ECJVNfrjpaKG17Ae9gaTpy0YUMdu4/fH4FQ3
Dju6X/ktmVB2wrpt9sZGFjXeHCn1+UzYuVo3gQurbj7DuZbp+eq9hgyoWb6BX2LveH08HCs21oWk
WQyG666Zc5t+iYzZRinanR2KVgOpy+C+YUMkaOSechai7yxFCQQuw0MHgpEBvEQDALhjZpTiGTPo
xbrybdvJUkpUQWAoDkIVIWUhFHGvu5+qtm4klVas5+DPDsfDkHjbO+SYcPzJbPG8dNzlgEkZ0+uq
/FcphIGwfvgpRMOzZhoZXNGsXE2WeeaEBI+14h+/heFQmuEFlr3BzPbEgC+5fvWhA1fgxNjNVqL9
VkB7eXqdNSvuLqFukh04eb4qTnhZ44t6//ZSMSn/dupiDd2ZzWhQDeQAVj4Wsjr/dXFMrfxUPjEx
/ptqEziyWAyG8w0YB+ZNdBNUCFCmdeEnWg+aevqDDpv2rqDHUqqGDNNCkNIGJUpCDB59wq2OkaN/
1ia1udDjpE+OELsVUHaawI2mAoAN3CBBV6TdFNh9bwZsPWIwglrCuuFQyrWw44jJ4Kei3e3fncxl
11X7Fvx0tYmwdBiqTnwMIY3hnUOc8kurSuA3UfCjgCzLbdFDE1oLStX8K9ciSF5dnw4IzlUTt1Tf
nCyubCG/IO08XzjKlNFQQoEZP0WQUNeCOeR0zkX19JGeyReyJZ2mefEUyxu1xsoX5wNP9F7R1zZ4
Kb2dnDppNSGyKAosD5g/EveCi5cdOF0v5a1T6l7lCdcZzDmSWsQrcV958c+YInN8Prs4PSPovHPy
w/i3KVvtVsU5DWpjquqE6BpvkCuGB1M7zoBhTGsyRC91wo8jOfCdFfO4FMu8YRcNmVXhe5S94YXf
qQNJMefYdKFsO7DlxapJGzLDb7qU/4Wx6a4KzHppD3YrzQ0g9TUJt1bEYyPTXZXZ1C6iv7eXkLUJ
O+vkbDVffEQFyD8/nOrK6UI+AFDPyXiErv+xWYcpks3HJE3syLbdaS39iShLzBB8fEM7QGk5aZNK
mCo5ueZrSLBZbL5JB72wEOMaHb3SbPtwYaPmYLTTJbSkqOl50Jfy7ZqQ9D/GBfuEQ/VPiyOc7m9a
2rWTbNb4hsIaCYaXF30zuRnXDWg+BSqX1wKuYqKUCLhz/A3yKcxg6E0Z64Ua6fL+Bn4f+SZKSI6G
snYjcdlBSmfZlK+yo1dkZhKbDEGpfCCmcylbDPD2wXUUWq7/fPQ7qwS7hs8eysFbagPoChBnXj16
mx7BPOGD9iOhX6XgGgrER8Yp1sDIGgdsK59XwsCsPGRT8zmr5/efGGoATqah7ogvSrdwuvHXOdnT
BCNr1gMvjJzODif2MNTKQiVAKhkwv85r7Y9x/ktfjqFNaCW3oVlfNNDEHD0shkXtUbEn4IAZCupR
rK/Tw1gOokIH7QeoU8crm4ol5ZvjkKqsNrihHOxwv/eTGj0IA4NL35p9oktNo6QWBYfSUmN6SzDp
4krvtZwFATasFIMaVTQ9T3eTMkQ9AUQ9FPdPvFWRfo4lXPcfreho1NUesh0KoklU/cpD43ZwF3Xa
x7PT0jeEw6l7B3Y0RUNw6PnGJfd2JThCYLCSc9h2GH2GVZ4iyhfoem0NUFLm4DvjF5e0CTdhGV5L
L7CWrbLMXEhnDWOBVGSSSnmVXxA23/PNZQXYllofnkD4ti/64q5lV+KQomGR2sbjMtdig4/An9zP
ZIC0MlaZsZJAedBhVgKqRQ1pQuwXHCDiwLhH1DSXbUdde8tjLdk9mAXXOEv5LaXS/NOvGqv8bqPQ
CNSlPgI5iFzK95yzHBrqMxbkfyUEuqJU3o/7T4+mtv3umbUda3OaenrFoibEFaWVtpG/MbJbd5RR
ldkOeFdrzbZubC5K6iRh7go1jhFqsTjgq7M6yeh22YJFyS9Aqx+bBLqYvjqm4QAkVb1CoQHVQbzK
vcPziDGE2gN6E2CkYzr2wrmE02uiPSNjGWgcI9kA915JjucWQpqTU/ppPMg0yCqd1xVi9FcSKByi
MRViLmCqU0Du+LRPPESEWbnKU25f8c36ao7f+kbUUfC+jxI24cY469sVHFs77Jf+Lb0vVqBthEj5
ffoOvf0CE49mPULSY8gMVMjM9lwZUgOSLzK5vcXkmZwTG9XaK2r3ZzJxhbVsRBtissg5KUT+FC1N
dNzPXWOXzT0LBD3BXmgMHKAnrgV3Xp/21t5htCcEXA2dgWQE9/4/+RmwbUYzmrQnv0mflTXDQTw3
1IyG7+c189eVrhoX1Uy6oKOAkUrn3mx18JG5/q5XAyKco0Rtx+rPUl3y11XpsxlTl40R/1YGDPgU
IhAO/DRvytPddWsdyiWRLnQY/G+BdFlWUU7YhmnGIkFwnoIY8E8Q5ReS7W/bQMeQWkwu7OxpVLC0
dFHXHC4F7SDATUh518zFoSm2GbFhOhlBqQKI9LhIFDJDPxUOu+EyIaegyXyt4/O2Aj0LXitqgPMe
4FY9vh4abXQ6hTwOZq/l7tQUb95Y+NZ1/Ess+UaFcB1eDTqCUS2YPxz47J8k7zC3vWHfediHKhlo
D8AQUy+VcUYJCIShtU+Hq7Kdtsmy7mDg/PARR2PfFj3PFiazg/YrOkj8ZWBLkyIYDGPbzIXM4ILl
I0ISC+91YpRpU3ZE2Q+0qewbpYFUn4LOeOjbMvR15dq1m2sH71cDGNBB9GgKuDvSpV4RayQ2Xw40
Pw7lkTYqqejDiAKRCG6rYdojaqN7PP5DpTKt/nCMMG4/klMrXC/2n5U+pjNdT4/6fWO+bF3ayElz
+YBWqYDKcTQxQEOiYtBC9pxRuDLWhFrnTLih5GpOpmoW3z2tpbf2FsvjVlBAoTMFVPTh8m+moW86
RN83o8z3aRnKKAUOf8i6J0sWtizfLrURQPArdSJI5ruu4CZBUHhR+1VcPOz2O376K3gQv544qpID
mR8cFq8go8buOuTVxJSL+fIPFf3pfdic/APYnlbaH87cyIZJY2H7b+F2gKXw587QGJDf4p+GJEW2
cNthTFyc+d1f4859LBhWL34HzSjkQpyohck4ucKpqOjiIYL9ptZHP8KaRK5Jx4pYLFL7Oa4yrQDu
iriBh983Z5742wsoD6PTcC/kmR+/l+PAGYJsEn0YP06gMZzE3HP+waPSl7Hxgsh/2AHA+BUk4hJN
hxBNYl1oDz+SwJxGt5Ux+aTBsPNZkGOgRchc9WyzOoW42aingZjbRHy8kcqVoZy8cxSfRHhJPkku
aOchF7hWgjvLOOAzWXQJahEEBNU2g3kRgBcY6wStHv4hLcQ0ycjfZnfRDwNmO6H3DgvQVXsnFKgj
3A+ghoB/bKcfMBRmwBjcbS373Q5be5eCravSy2D/VAw3JFB1Y7btNbxYuI1ZwIvxf5JoIMRlPZeB
KrhyQDnMxAqrlV0TGKA0f3i2MdY98uSCWaNKI22YuJ0CGOxq9kpN92VRkDZQI6izF79QCXPqjORa
tIBraHCq6KeW8Ie+cUfB13u55g6ZS1+D/3NymxJuMdfkFTpThE6UxzNnqLOBGQmZC5fRtuW9Bx6u
rI4DwOLHZxf66GYReeYYSKznlCFmz+1GXRVGE8d1LMgd240Ki29ZSN1496DOYC6zFdcxxy9G3E+a
uRsWXenUGCYD3EStg2OFQfRm1AL3cPi4OvFKCV7I9t2cO8vOvuXavU4bjXspVmi90K+QNwd+LQH6
5igfTj2vT1wWTc5TSQAICZUVaH+zhoor5KwxPkn771ger/h4CuEQp4pi1g482+vDgQmkuPxzQ2iD
xnsphnRAU9jSdhkIIztci51DlzpVDMCH72Ou+Q3w2qOJzsE3w/05gQN93HUfIJyIPB6u0gS1cHU9
y9NG4+Xp7JKUbNx9t9deCm1kagr4mYc3mSRNL0pG3cSaaMUg0M3ngs45giRxfBrO4k6sAQV7VP2/
UkCijGOwslzcIOrhcmQX0Jyt+AHBHWrcKEn+JCxwOmwLkBsVUp2mFfeZ1eMFrRh07+Y7aV24oQlN
38/LZ0pm+My/QbrCZNb+7t2qaoaIq8lPXWxxksepX2dRqdX36/gn3yzFA5//DYT9w/gg1B+nxerp
fJJlHrYXxCcLrlmZzUhaeY7/2fu9DiSvEGpCGkMBcw5SVTkUw8K7dKAqaAq+ypNU2MA/TmfQG7Pm
EWmH6mF/Y1za2xe94Tou8WKEVqWh9gQXeCVGbzhv1vVF067N/u2X/p6ixqb5obMtnLru5l6D2//2
UEbtkIaPKYDMZsypAWXdO78v0bxCwKlnT6pRhnbnN2/yzPknXkatjuxtD5dJCIHJr55NNMutERvq
7hGDz4gEwpdQCxSYx9eP9KcRNh5SFXx9BXYXe9fwAzgWkon78LRTPbKUu/tkeIQ2hTdDtgG60g+t
OUKM5ao3UHqGo4S934zi9b+40xF0NVXqqEmne7kExDPC6yBn1RqkkjFxyfJvgv4bN6jlH/MwVur7
GC1ULK34UPz71YrD/zoOth9NSp0CgemPUE3WIlElQYfugiRXcglK/IaVf1K6mQQyRaJsRbpMrlSB
CrwhF99sHSOGfmqUcteVYEI3Oze2Zm4b/sfxtU+Ie27nmoLKFwTgLEcY1fqIWA5dM4fQoo07Anoc
VPpBZuihMWWWZbzpmJtTWbRcu/xiy+GaFISy2KVsrAY8Gm10WwOYPunwyXUKnY55qob3nrVuzI+T
J5eT0tMhJnczNL8kqO0ZQVmn72BgHPckV0O1HHTxgsTGcCj14TvK5R1gROUPuU5r3FgqM0wUxu1T
J9bgWQhASKmakhPC3kYaByBOkiEy6g+WOe/yRGNUrWk3YQryucjdPxX1DMlSGwkCWgv74fUDvs8Q
pWzxqU2sOk3kHv1WKYJaODCBB8zFAS+6UM3B8g+rl3dUWLGU3mZmXkjkRmHILF2t4q2ICp2hrOhs
aIcKf6NO5D24Y2RDs4w8rTOg/Am7O4bbX8F/lAYnspyFy+JbeZ/TCaMkMN9870bvSsiil+HsgXNx
JIa5tjCtmeXV2Hq9Eo2K0pA/OgUnPzqyBn02CnLTP4ypPEFDKhFjPQc8Bcj84ntBvRHArh4prGOL
tpeiSTvP5BMbCE5n7A4cXLLf8D7pvkbpH2vFzU7iOrkbUeaIM70NlwrSOj9F1Dmsmke0JS96cH1D
7KBAQWNWlwqyKpwnbpswR9CMr86MViQr/jcdDZeRPgG+9+9Wsxf4c3bwo0nZtaO9cHuBa9BIYT3P
hbPBQbLzge3MX6bqfJopdGcCHfXHD3dWJhzlRoeyf9KsD+PU1ucIc6gl8pOApSzN/NkFfFCxcr9O
KEpnWgy4eBMNqITuUBQuJpvDJB8y1bpOG/GIMXXBaoMoKlE9p760c3kBeTAFiE4tqeLzsbzXCMfb
YKPxwBhFYYIvpKe3FW7xIrJrm+vIDNt4oOLKaldogxr4qgWaEE/b3W+CjeV6FyaXWTBGNl5LRlmV
DL1R0WD5sjSh5lXgp1LuY+Qc/SCGdT/1Zanpa4BrgAISjIp1SlPIBnWOBBB/JCrcIM6hod2EXEXB
MOKz1y2VixX3vK8DPO5g/4N9cqgCNLFIk5tWdhD761mbdMsbmAAoLrAzBO7ow6Nan1veuibmh/6w
3Szs6dRCyw3CX3QZ9pcCs+O6Cl3+gTaGHxRfO8QSOZMIw0bIzceIymXY0lCE7o6vXvJqXkzbK+lN
/evSgEh88Kd6UIdpdM4v1iRRVLES7zceQ+mh6CwdWGJeo0Z/SzNm/B6eupj4ekzEpK702/O2lLI9
u5HNV7Lx9E5PVmJmoA63gHXwNvY7rL9jJrYQbCbVkeCMU023K03C/5TxP9jqMwvPYCiyvjobL32K
7ASZSo6WGrPeCMvckxu7vU7Pw4b1xSnRZ1jzcd7of2cXAWzXWqCIpAkb2zsWCOMATz6ecEspzrLo
0NkxcvTGmvzoHax582HN5DPqbT47VnLg6DtY1QcFclCiMVIaNRYYkzt2e8kZcQeoA2mJfgb3Jb1g
sJd3r2OWERu3PktutgOw+IHeED50Jd71A39zTZIH4+mxZjZcE1mmnKYot9WnKEkS0ES6jp8UGLcU
3NxC44pfuq3vNrEZGnpW6EPBKMP5TN4bF4vbvOCqSjxvYy6SR2+nGwbsW5whQJiQfntyklL+umdi
zyLWjxkfDCdTHQcYTpqYQ/8j6/o8oKAwRep6glTWprkk0a4zvxQ08GBp2muY7qOW9JpQKZLjdgJp
efwrW+ACk/bN+FCUmTWTF+PJ7fyZRHWHOL4O2G7fNoftU/hjIQ0Kwaqj0e2V2W4VHAWvi0uofhmQ
CKd/tFvULXeOW/U0Il/B22MenLE7V8k+eaU+s4GrbNI9LRfK/WzKJjqX1jwiFnGTNIxvl/ekS0jJ
H28e5zy3dn1U7goEEH6ATeIKnTixurcFVz5e4cFL2cOplfdETHnx+jT9hIwi4Hd3T3iKg16V+MOa
i7WMmsZLePGyKn5pStkFAoGbkYESqnCCL5wOPI5G/t57s5mz3r4rL2PSUfU47Zs1Gp3aozoZY6wG
VZIFyNVrzpHxjqyUqy/iS2w7SA7/bTILDbRuHkFgDP5sLSok7ksXEY2ZjMw3WLEiXP6UeH06asJt
EL0KWWSTZKLd0t0jDi8+DxM6/tz5euIp4gDcKKFV/sEDCs+aRfAp95BDDWFpMJ2IjVsJVswUOuUO
OcrpC4fC48bS1PRWI9RFHAjZ5MNS1p8I1wJth9USa7hjfR68Am2M5UfeDaieaVVOnzB3VRKZLdxP
DfZVgVExz5Mv7fJ5yLMQYoMLPPF/GzotrMSeS4XkzExcWZNhDtsRf7RuzrLeHE4s0En4+DQYzu4O
c0LD+bZWojAv4NkZsdfZr1VvvEfBXP4tCcWKZiwvHHgZF/Zc12w6dp+h5ru6bfP89Dkek8mpyCU6
gn6ske35WdSrpSo1b7Bx9Tcn1Dl+baO87b+gTqZiqMwywW+g+ImDj86jmyrLHHZrzObBZ4OTyzOQ
BcGx5Cw6r9cMY5A/pg+RUJMX1xMHNo4rKG3LH93wpQFhl8GI/D7EE9E16ioXS8MucDfsnEgvtWLE
7/SLRsq/bRCLwfJEZkOZUZfvgWXGok1Wx3iB7XTU2dbcbDXrTo+bkKZ79RWy7ooCeiWsXUOnBB/I
n36KS+/xNs5nPpBwhEc8L2AhFZoX7CW1nC9wNmLwRUd5dIqbrNJmNDA2lrpxi8NmpUi8WNcocSvm
BTMeFTBtsiYirTaxYEl0rwXyPfPkNOsXXU19uKnXfojel0pB7LCuUEFWjBao30vp4+uMV8kOGnkk
7Gd69YNbrNpdJsmozLQ9TRJABkv+rkeDylkUSaV+8OZBf2Ymsh6dLe79JkCjjGVW0F8nHvaXanI0
5izmtpZk0sqXf4jBduD528w0STMWinEITo/6EktFxmWwbk6P2XQPEgYJPnWd6kXvoP5sG+MQSvfH
uLNN0S4NVrCzGNf2UoYo/ZVLcFHnRp5SIJa1CRaePZgjyn4Ts0KeNAkiEu+/L10pHoepPicnsjCZ
U4J2gvxsoGdimQ72FBtdhJa98O+NFeey6TQDwkHFNRbG9AFlQ2jLuhAJDVKptgN52t2njSbOWV4j
MyAVNSkkUF2lNvROkDuzy9o2oFNGd6vfisbVUcnbF8/mJfHEhyI7mDRIqyd2vyUm6ZoKwE3LnGhS
gW6D+lyZjnVWeaFnyUqj4Ph1Mw1yI8kkut0a2GpyWN1P1odGJ7iWicwjLPUVm2efbLd07N49Cpn8
G/DhKhgz/eoij4r0xTHXHM0obO5ktgR3Y0bFNnCfwfjN187yBfoTK0ObFdpjgMNiPKkE5ULkNAek
VIZwjz2Z8EOHd5kx+chARjIAu4etCIiiVhiIeqxBy+Du7jpOlAqvy4WfseClwkLry7IoteOu4q54
YyrM1Kzhn31h6QD0YJ1OqxIn0bsjtSdMSFhYU/68/y+1JjfY94SGGdRoe0w1tA8aEgR19XLXS65B
jie/sgfJtKMMb9qTCX1dGoBDlCCFk5Q0BuHE+p9kGo6ciqpZw/j1t4hi7SA8ZC7Hh2CyzaH+1xxd
8kXTPh6my4FeloA4LQjhYp1jnouENmJMZCFtTLI4voS597NJVa0ihs8F3F1XeITyP5dj18qRTlc0
j9T2W3iZec7r5X1Elig/invSwOro4Yz5LoeZIDsMktJSRxQDSJp/sBceiYs6Q/qhESjgyUiOrsVv
B2BV/tpvneqLWcD6GTFyGlzpQcfC7zEu6fWaGLcG6Hy4RIwqiDfe4XuyoTftQLgLWKNbAbo7QoIb
PaD5Ymg13oqWj2/qCP6Ht9QACPeneGY0i1XaqoMSKvSdy/oBqgn8ngSp8oRCO1+8oXFRx42Nk0Oa
ZFjg5QWmCLoDW9R152LAMZXAechr1dVUa08j8SHuzZ0/oCOrlhjPmwzys3hAbpxJU48KiRUufsnr
Vf2UTYNLfqfJ+UEf2zOBwRj0XVO0TxpUOQdbq6gD2hZtNitlLUYZGBZl22cQ45JZd38piWW1DYCN
pGu9vcJ6jh8PJq4VAwS8YTd0CALw8KRI7ndxvyxTeKOErPjMXhEpQ7qB920iwPoSUsD46f4XTO4O
vDzNbiVM7QR11eAouUcFghw0mS2NLiF/PR9HL7jIcTZeezZZcJ+/VT5CwNUJRaZ7RToaL2SA1v4g
oDzeQV0O5izEGvfHr511NNaNGvravUTMj83M5VRmumVdmv0ULVx5kBdD/DknR/dS5PvHP6wB682g
BYmi0kKfLcyNV73u/9Y9nx4a9298IcOb+kvtv8hWEcc6VN1w/Bq9HryHqDDHtZx7nZfMGpem80/3
ndPPBipQdPxKgfVvArn+YO4prHZj+wwQs9a6X9aCaeyHsOG71OK9DVxh+JUDfF936Us7fgCLwxvd
RXDf84muP5RdxjBvmpzgeQz92s9GM3dPeP0a5uCYGqhIuFzXT0LrxKyMP/11ZqdHdrnkW2yUd2dM
M8LZ90HlFCWswF32EuIKrydw8Uq6iKDl4dsIXbINOjGOqQbK7PzIoC7ZJ2sl9ef7V1RvTr2QysXQ
dMi7l4QuqTapyrFrfh+pVak1nd43q3JiwAbZJpAA9qHgin4nShnT2rBPTeTGBH4r3HYfdJUhWkR6
KX7hC4pwOss6t0nWlA4+qIDFno6bb/VqVn+U8Y1NgsHs8/eHDxEdwNflwFHF57GMLhMhBI411+AM
bavbq4Xv088EE4gVThwQ0zJ0YaIUKw9OwTvITXbu2/iJCwzyRH3YVR81z26+ABz/2qG+YOT84EjR
k61bF39q6JaP9O9Q2KKqyUWxXdQFHX2gM3ilELzDYHbCvGgOPp9KTUQfDFoSSFFdeu70oEm2p0xw
vCFpqTi36iKxsFnDhFpShmZPgQSGeKWpJEdQBrVkiyKcTalsSyOWYCfsQw5uq0fq96W99nrRG6TJ
xIMZjxsRFX0FE6IS0dxbK0FLHfS23qfkkXWHdUp2CCJEroM6aMwYXyWZEicsRycQ2xfrQmsxMJZA
cEx/viEcc7FiJttLc2OCe58My2C5UgwjCk2Zu/8L7yY2i7pD1NRpCMMfrx0fuzP67RQgg5Un9FTp
qKmbllt0g0dKlu1Vri22hpSCCtXC/NxrnF/SvASOGupe/pBaVUI+RirTcj4dDsKsU6SmmALBVjSI
hyNSPo/x9tBl4j5R0vjfL5XXJToh876fGptc/kU0H0O6EdrTCar2/HqhBl5ekIddz1i+NN6uq9ZF
gBiSNHZQaifl0/4M1xJ9A5jMUtogiEaFeldbt70GckBuEQc2Ht7ZT0adPbrr+debmsuqMDyOMAWW
bYufJrRqcH1g29nzEKhzQiM+or6fDzw9iMCa479bDlmYR8QNDlOv4cRs1J27YOly3fAbscgqYZL+
7iVH0BpubMduqh2BuZ2hDHN6v26Y3826hYvex8cE1K5Y8U3ovxmKvSOVyFVhGwCbr6Y4Dx9/Sns7
6srBDDVxFb7mzFIiuH8uz3QdO1spmoZBq0KFQ+7q2FonrT4r5MCYylsVFZmF7PDbPJUBpFOJRMxU
dX76oZ+baH2LiOw4153QRHusHv+a6qFdZ9UJne5b4AA8q2PXzKusJ9WePXyIZ6GKIAtUiyGk9zMr
uK7OD01YrytWalGk5c+WRmhHqM67WzNrC26wEyuAIOthcZSDF9PMh7do4swhn4B2fgQAv/BSVlC0
KP+Zwbqzetf8hDswWaPRBGspi/lhw92EFK2CV6QR1Zes8j2VQEt9reKjoeQ551djMlAkwRwoP+vs
YnYjDI/2TVbL8ZZTkfBb8n4LMtDANEEYU4Q54otreh5DRzL1Gw5+qUrqH9nOX6/pZa8wBXdyjCVO
TPU9Im/MxooVBAkirwHKLAFsDhOp+cwq3PC/+pgNRr7HN98Rp9wcXTp8f56l7NeEiMjv/KvMy66E
9EESVXHZm9TZ90taLcgBRXO2Hieyb+ShHLnmSiHpW+U42bKvwlmzWzsbW/uOyVPdFFQn1yygQ8Iu
wLFAcb5rUdEpKeeGSHrkuxjJT4lgf0f+o8sdu+v0gnzcdrmgw3VQKKAiYBzxhGNSZKwiwYcnih74
P/fuOEJxttjOAoo8VkI88O30+Li7Ftz5VkUD22UJqk+yHIBEVXgO+40mp1YJSAoAcCIT1MVzFlW7
bpWvpVgM7IKxp0Ey00TgTI2h0Kf7pm5w875kL3PQSTvvli1FNAD5nJulnl2sCz4O/zuAN2tvSlIg
D6eDvp3ZB9DLd9uRyz6N3P9Upk4UuD1+3rSpX/U9jztld+GpZ7TGb24C6BxDRoMvm/5mKCuR9UXt
Qf1PKPYOTCW8zSM0wmZlbRIhgwhL1A0ewKZN9cmqXZ1U7fHwu8fkHaeeRF6dSELJhXmcjuPHnDQo
RsX3d+FATlGv+QOwW9jOQZ1ogcV4SpBmzI806tncrNq236HhQhF319cXTphunUD7Pg4f9paP80AI
F3GaYZ3Styz3jDaHE5oSBtBRoPD3vbzLJ5L5MItiMxaaspBk/1KUYENgjYj2SCJT8cc3yNQbp1iQ
aKiOvJtxSlUS4SqCFtO/KkvNcRIjLJaPZf2Kt0IkpdbDfKScHh7lY/gVs5B0wuOH1HveWybD4EuF
hkbD2b9d9sogxvqgOPHa8RFApItaYIGd7dvvwmyu2uPo++yeokJKUVhp7YAA6Jw9zPkTUNYs5umE
t/HwsVoD3NWTumr04fVScqlpLA4/6zhZxQO0AncLBWjofgXmdHtjC1sIYj6nBXH/fglMmOiVIAHg
LbMFdcggEca5AM2iWyPCbkp5M51QpwKbvPx90OUkvbh+kF5uig1Is2N7tutMGI+AmTEw4YTPAcX0
y06SMY8ADseJA4KGX/ePfBi7ipJObNEIY24SeRA9IBgcZWDJOO7jXOS4f+jYGFNoU8/NAIQTwy4p
Wh5M7D02fPFFfmBElovOqFDYx8Rm7i6yVCLu7bkQf/iDuSHQAsgx7Ka7p1KXC6lKWS0M2iAa74iQ
Z1FbplOv54Nusq2R98/MfwZAhWjJAXV/LlUdM+hsaR5jZ5KvjJHJfoPRQtY+9Ybvi7FrBcT/VZ88
KryLuZ4ASUHggvgIJV0JIAYZA1Ml/O3MgeGlzk2WNYhyznypCMkvEICm4SpCVK+eTaH/aM34JRLb
Mn/hBp/YedfVS/L+rvHqiIy3a4SVfEza3ZMLDVg7i5LKnAZqQSsS7KIpjSgQ1wBNPa2rGxFnwdkH
6qRVMpPJfowYxWt3Jo9k+9VBw+O0Q89BKaHZvpPK8uiJWVkq8mxrEl/NTUSYBTju4McERP2dpmVH
UrQEBcCHBDkuRWY6ARH8qaw1edH7aISniQXDWYXfH80ltfEY2E1ewNBPTwfOViMtprgIeSKGV4iY
FGTK6p9G6WEHVAyT6EjRp1MZLG5+fE0eBkquakImsmpIbrJcsjKgGDZxYpTYCC5mjBj1F+iElDTZ
5F6z3+U9aq6D5q48k7th+xdTrgLyTboc4z65dn9gAvL/PpnR4KEo2sinB/BhbeMFoKHJfJEEGU8a
BdrrMlKvgXzpuewXUCaVSz68l2wE9iqlwt2o4df/kZMtGtNUX2b0sKpHC4B6BqA5mt6VBnQlQTdn
JUxRUmcw+a1Pwzk0pvFqFV9VWNCJcIWu8yhjoWSfMdyqANW8dUTx9JK2eamrEB7b+UvENlnyF7dI
b6KtnTCt/YT/dPgjISV2B/YyMO01Wth0BVGMpgVRpYK029ftkmENJrrh0mchz9omhznv3ddRNNqG
Rjg+/HzBFfzofn9n72Asdf1zz2MM8xG8PrU6IcnnWTEM3cmkY8nZwHdVBlMd80iyvS3CKT9T7dNA
pPX+jhMDedF19lQy2ymFdi5F3Z9V7kuLL+uAoJmzM1VYQXlYE+0vOqfXCV+fLPM1g708Ea0ZFbrs
c7wUwSoon83gR0oE2+Vs6RCbyqr2xzm0s2h4Id2956E6R7zmQAjUOp3nYz/CZpTMY/tIj3aMQFlc
Y45WeAqfcqYB31ZFQHXWMQxMDgOCg/N5kCytmCKdyzgvRgaVEis0AvofaDGAmh3LMUGn1+szIbo+
rqXD6n6pTYp8uphZF6uZ1gJZr+VO1iQVmUiIyO4C1O11N+KDjDEhUEgaWiYzPbmzdfozR8M4IyyG
xuOGgTX0aoyGiuHeG8er5ucVMKJR1AxL/hUnRnzRKoNjoujW6HPF7yEI93JIWhWJlW9jw1OMeLKR
KCubNb75it0dMEkx2setPSuvoCv8hOtNEE7g1aHkwegtnHaPd5aPmyckVzMpw0NRS7Ey3id4cAe7
Yu4E8ugdHDX+iRS5PNErdyiZ5wdYiIv/BWH8LDeeaDDwYyzuNXcI2XGO/D26DekHUzAaWs0q8mSK
COxTp0sCEVIrQ9OyzKOvAsE86cygWLZrNFr5UPwJRoqDhTWdG0ppHrheITFRD5yhDGIxxnSVy7KP
omyM8HF5xVRurpwJH8COQ+//wyW4kBzk2RftL2nO+weZ7BArsIzDPNOFx6tYkzhKfbf7Mr83sDb8
LibpYO/PCbWwMNvnQnbQh0oiaD2nWCWyBobXbiMEkoteC7fH2Lk5QSxqUeHshlLEoB9A7m5/YLf0
6RAZAF5F7ayrCC808lAjNtNH/q5lO528+t1MpYbYpYYRcHnepQEuTOXcBcoHtEIJ2tgwaSStqUa6
9Xw52g2JlskUDUyngKxC2pnvSKk3NJdT1I0/NaFaenR3bmbRi6SEsSpKQJ3TsUrYc3ViFeXY/kbm
6Ktx15+7CLz8J/3Y1G21HP06XtGvFYU/Sv9RyOp3ZvkPqThJKgV9yR0svHrABR6Z5iqXi+UPhOUj
Y2gJFeBrIp69l96q9oSAY7dyKS0FC3cYr+dCl7fr+s1hDrgCYCV9TFncToMPWvcMBiS3aZaEAfax
8CmuJmc5MpJPbqiuTgYyJkFWfCt+gEF1pTpNXXYbRemmzq/+asmryz2pBq9pOJ9kEWbddnN76zFk
3apqqt6pCZDkvmGCwU0yJz6cN/y83rFbmy9UTJVNeZTrR6kVsGRMypYVzlPvfVJviLUUymi2p7AT
WvpmplP1ta6Y6RZqVusAYJNN+++JWFzMJ2UYcdeVle/xCQk3REqR3l66BXHztVS9cJbIxXmHSjDQ
X/ypXhgdurKNjUExEyM8g5VqCQ+ZIV0GcInMd00FbWduHkBG3rykuEnsyEVDe+5s5DLfkmty7NKZ
ntTdM1HjOE5Qxyl4+CkTPFPcRI0wOXdfZgLLsZCd/hJXKaYFvGaEAyi8/5Re+Zr+OPpNwsQKkdzz
47BTWv+6YsCY4GH7DjTj5yZ0Yw1IHZ2mPHcTSs8Mzo+q5V7TegIjr0cupiTPDxC18Yvek+ZkG4/L
V6ogC+cW2EkfOgvaICR3hF5SNlM9JVX/QIJCVbhb6VwPK7gTFSvLeDEmjwsIv7PIDeVmCz9h+uR2
D3LFSZ/eSM9CJAh0NiWVboVydfpdT2IxOX7x5pNGBKvai3BbLFxzuuSWu6C1JmbCSovePD1s6vhO
N10p8LFhIpLhPmAca8aRf7Ti0BnMG0cqfqHvmYF0c4ETRo/sesQ+pw/BL4t32G+2mmTZJxA1oJg/
TCJkl+0dFVV5GVwdl2Pr9nysvDKaiL+rR6s6aJLhwh4O2XwRznEMtHfrmYRf++3ZZj2MeXl2PpKJ
oaO15+ITbHHECFCBWqVv1wx4GPsCJAxGBzO75Pdt+8aD3rTiNDEYtt2q0nEbu2D7hnmFzHyfPn3E
J5s205gZJfan5ggypq7CWSYuR3N8ajMHqtEHxfkGwDi3eRWww2ZrOQDN4BaQzDoYSFmrLfrXYTvE
dDvgsEl/n0b7V791UEcLRIyU0pyQ0V/b5YblligTf7pf3vT4+FRzI4iXqfxhHimeDtxV5cBNL+JN
qhbqor0+2UjTZVy1a2SQi8YHF+k2I3dR/3Iddw3Tozv8KWeU3PKTllpkoqyvq6wUZj4zIelYkB6o
39J/woIu+y/RSxs0FUWyBUBrS8NTW4olEaEx173Wpu2XAm5B5/Z6SuaSQr3GVuT5r3aQ7t9XpxNS
XMn25kqwrFbnCjnyx7762tmUAIjrPYCo/CT0jayBiOHi2NZ6ndqvZrkaD2cIgRwXidv6usnSsglF
B+M+V+RBkf8V2efvBQhYqrYDwVvAjFH5BCwaFGAr37+pFaMzuD8o7mLCIDOfFeSZMjgG2n6KGGS+
NwiwDr9GP3mvw7Qa8Bas9MwPPrZWVVuSmMzNDEbnGJmOXrto5wAcbwMrxILRM45eTYVTPOG8QxYW
Z4yFobED0zgQbrCI+yi4pvXvjGhE3Pu3pPAqJ8y3Tt0u8kZoloZfIjZ4XSiOLoMTlrELR64UzMzo
/amnT4KUPNSdjyIrsfdg9ZUk5LDlBiZkDYj0+RWECDNGNR92fNlSaZXyD6MBLRrj1H5UMJX6Awnw
65jHubFPHenYcan6I3w2ZItLg9QMXsPK5J+G3UMz4GH5cUWE7N4G3NP9PFpPsx3O3Yw1rp0CJkga
JluxHL+mfJKrH3+qAhw7ziNdzLsEkn9nf1I9rP19JWog7ecpUrJGZj4YIsCudsQyi4mPnbDyPQD9
fF2cY1gzLpbvCfSAbIrluQ4RNgNv+vpHMvrG/vvrihUyXO5NUE6wSmKuX1IV7MNL4QhDFMr+l4Wv
hbdMZtOZubKE+O0yd9um3yQ9c1G6JRnExacIfC4+hh2K5xZmANHGWJtYjkcssV889veiXBrIZV0V
4jOO4f5DsIKjjOTXWxGU3lZ5RKyj3cD04A1a/5/kpq7NpEoC2zoyQ2tL6a02x4xF1U0u1VeEj7R/
mTu855UXic6CAxjJFTh5CA8/Rej0sPKgOCONmSKYzyxcKyZRSLEhboL8wb//u1q3pglesq23bcm2
OxTg7ha7GjbBAxLuH9yKveXauAoCSVFscwizkfHPDvEMFf0gPX5jtscWGg7kadAatzXypUYmglo0
ObZx+DWIdpgJAcUqp0VSYrdt2L2kzhm4ts2obzEfWZ648U5dcgXPyihHmh5MV8p27tSDXy+KLJ2O
nG85CjwQ7ai8scmm2ZX7BTpgO6Krjn7jvhAkaRDg3WrBIV+FxQGhTyeM1LbVRfVYUokFQbpGQP1e
Bd+ucJ990Nqa2TFkwmwn1NFKPz83TGG8tCTRaqa/3IUzeg6UkwYbtwTTHq1TfQMm85eoYtidSRnm
+tI3Rplz5L7DeU4/btHpcmadPZ4ERP2iqCWLuEo4uBrsweZk5GbhdCu8x8Zco7CK+HwKx259q6eA
4+Yg4ld3VcXfAIrj9Qlko+cxzG9YlQGy3csFBO9QNRq+zFz2Fv8ydnbd8oOOXuoV6wuhlZUZdoCl
0dhK84otP5trE23Q2iuvM0VbW8Ssk1jWtHYWb7pb0kPYHJ3YJ3y81ZT6JogxR/1DZ0zzlYAv1kf8
n3EXYfKm2vdidgsxCWvOMO8+7QTd74QwQ2F/eKA6ofoxRnMmblVw0107Q7ZgW1XC5wulRv/JjfUV
MojFA5xD6CPO3dgdxQxZUlEV5ySjgJfN1t25FmERkLMg0PdxrgVqPOnMnhgffgak6UczRy9+GOoF
riQYNcj2xv9480ntamAuv0f/lm9Zh87Hw++aS6YaZS/WXhH5lHMexZ33PRQpkjGm/kJmGh9w5/sy
5m3DrojHNbzfXbuZ0x6/x0FW1+chfA4Ht84rVzFOGTtE9HVocFI17FBcP8N09vTf80G7K1H/zXgo
CZvMo9rWQxPi2Q3x/EdU7Y2xCx+p9d2TFbQdEqw0GvblK7w8PDs/353amsnZC8/nUIeTewe9fsS8
2gyKNXXuFjEV4Lz++YElBzU0uGtDuH2V3RMZJ/8yiCNGzuzQqGfNAoS9vO5STMhyZAuK4WWAM3gh
OL3aTWZJ+HmKBz7ei67Dl+4pwCxmmzh3EB3gpIWZr4XQBp8pHKRVhcpiygVykSy4eOFnZqNKys+Z
ksyx3z6yiGN0+cWP5F4FhUqWmQ9/1hxljNyqUmVUns5h84dgL1zNcDpG6TUBAcVYzgTaDsSMhgk3
yc8mRvRPCCSHUiVBqD9Yd+BtMR7/+8/aW0abOa9yISiwBrvvcA7sPJFo4Z5KEwruzuKE4th53gYj
WFmtBYfP4UTJ2P1iuJpkqhbh1dw/Nn7zOJJIf05FLvllc5rTI1EtghMcCPtIkoDrbYersuNnSqv4
glVlb6SRBm2fx5xSAOLwHsLhuoh6ySj49WdaHigZbQUFREFk9eBk95bT+P1+759JiYIVZ44Kqfaz
qPIPhkf5ZFA1FLrIGkxajt/4enUeancy9RwOs447CBs+7A8wG0WE7VtZKe9klzcFiRSaG3+bgzu9
+aDT3Ls7kngec3w3EYCF7UuSlXkaZJKmET9T5WdGH6hJRwH+6/TyChZpI46xYuw0lIFCw+swZ/Hm
KnockmgNfjcK7mHt+wn90qaP2oXtxfIz1twmIpHLTdfM8Sh5WOMbvwU8zhk2GtIpwkQGBeXjUh0z
gQ3tn1xyGlLP2/rgHTa8k4gHwSjCeEzYlXBGASx4Q6Sc0OnQeOkd4BieqIZ1IQLshdSfT0u+zEWq
9tOgjq/bxIASdMvPAYhhLGn0tNqKpQVHBoJmCDXqf0Gur9RrVDwKqLj7j0Vy3ZK5L7QvcnjC2FWO
2IauZrtz7+zI1C36/MHFCIe6TNiNqIil48Sv5atwJo0bJR91NQymPG0ldMavHSsLebMdNl/Wa9NI
QjHW0WRhgCtUSTJOTwxbYU3Kn2pNv7D6HINlh/tab/unzEGEcmBnPUuAbRdHIOeRXntvEh6xoeoF
HPGa62F/ljj9AcXOIo5Z8MNC4Bqf+FrGxVGwbpAoX88y2Lc5THKmeWC/964JB+VBMSsHaaZ+/vYU
5uQfAcvnqD/EEGTFTPhn/tEHJqy5LjUMIwvly1KCNs6EvF1FsjcZezmPIcn6Z2tQT/VoKls0Zyby
aERTR+jbB8D/FPIHpWpCb3Gc/37Y4NGfbiHUCxw5xp0aHGjVArybe48j1j4/SaWcZ5P70dCeXGlO
3g/V3Lf8LkqQDVN+7wClDlTsYxse+ML4l0xWh3FTuMydcpetRybx9Lz5Sw0u0IrZC96FmzFNIMF8
ZCDmtShR7ah7/Wc/0WvpY82lFWrgl9s5HAMPD8p6ROClLaESFs+Yu5C2yz5iTeQz1UUSDC85MXA4
VwyLpRcTJdakirk5ZUZWdgJ1VXmtZdC42tsX8k3Jjwe+oKwuGmVs9E12hAX8NzImsOKWz5i3M/u0
ZS8X0KKZpA4pXO2rx4KpTMn7bncbjzQTzBjORMNn/3++X9NVNwjq7bcdDDWWmzuHhjdLbRcXNh3Q
ix6IZm6uMUYBavQs989AF50uDSN23Nu1OoHTxkpE2submileZ6mxHTAvcmHTINc0eW2F5hM64G1Q
bS3OdiDn19S5pVBjOvEJNmUVsVpASQxd8kvWsayJOf4roCbJxAj1u95Ynw6awhNVnPo3Wks5cP0x
M7/v/DHvN4G0Pqjc0IxXbuwLOgSKunrG4D3TOMlpoF5qBu+3tudzzR4hnflO9xLyCqGkZI64eITB
fx//gbKYnl32wQPR+orQerI7ZqJfkURUOoOdRua0xOqjLseLCfvmdxo2yLiqz+Oc0et6FikwIhBB
AKdFLJT53GAa9BDksoF7mByxMlLzmivGgr+WET1MfcXOJtyPOrmJGCH+HQyUVacaio6bsWmOJhKa
rRSVdK0BopH5bkB/k1rKu9fnxt3HDj6UIUNcAZl6A02yJMQHV2IUoqNZ1R/jJplTjBA0QyU6FJOK
J9A0ElTUlBdFYLkWxyw9lJl413LcUaW8HMqMpVoE8vNiKyN8WMys5UUVMoKxq9Xl1Y+yzO+i9a9B
mRw9ZeO6zriVhTtwLRNnLhrI9vddsE3rQupmAfd0gVJCqmVrUKm0BBgbZXoLoHpngQEr6tYwSQn6
fSggOl4P9K39w3g3Vk46rF7RlIthABwcTSaKceOYIhwDbckkHDnx3rvtsnx1ukXmpUqndtFOnGWo
7NEoE7y+c+0pXgH8lJGXx7zZuzvf8G8Ejy14005Ow4ncXbrUOEdbn7fMrT0xRPCzMVKoclArF3kB
V+nbK7HW6ZX1I17SHE0KESGYip8eWK2ydXa+T6zRp4IxSwdDhWTJXSRJHxmBvUrFq0WpbzeNSsX5
8igUAcpEFDiDLV/CEmbIyXH28vw2bejJKqT1ZX9Cv4BO0y/S+gI4VsViW0wyk74aXpOqnxkd8SHB
qFrOBBcJMS5MhGI4TjHYH9+UhhuK/uIvM0//hfDG8WiWUcNSJdtash5Wn66Wyu35v+EdHCIS0JNk
8cbzxbqyKmul7FT7IXyZ6vInOXJiu+6uCMeJK8O+vhn652xS3gwJvE+gDQqx/F+F9bmerAlm4jN6
bvzgjM20Ux7NUK87BZUXzwrfcSqiYSg6UvL1FebdmnOjJqkk+pLxfPXjtrr56/Iz+GX0IkfNKCiI
zX6UDXV9mG71jI6wmZZbDKQrfUQM72dacxh8RZNiI8UsbbfrFmjeDrZGxcJ+Hly0CpCRoB2AhQns
wKT0DwUDYOXJ6qoN14ZMWRpIB/I+qmG1BL/qPDG6dg4/N0L+VMWC2sqMugiLsVE4FczJvo9Bxj0x
N3mnbetSSHO81Eg831tWtLkINGAjLiNsDyAj71unNYWa/Iun0A==
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
jh2e92/4dWCFMhweIcarAzbEyi7ZOLq1s1PZmUCHqBMcuD5MHtKWwmuxrhrjCpRP
YCD21+h41FtRH8krqQaZkEa8EoBYU5Q5ceNX7HoZrx6f1bJcb0/HFLnRY5Zp+dk7
SYdPU59gwJ25w7UmH3A9YTGcaTPAYjT6mlHs1ODnAfA=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 63152 )
`pragma protect data_block
qJ/DL+aGBHzJ3XYwu3sRMqJfz631Y8nexRP1J/tuVwUXHI51RlJaAYdRIkVQk5E6
XCBmr/YJRfKBpIoMBSiEeFbHkaWusERu4A+yYKrOeQni0FiL2hEc2FAnh2GSJoE0
sze4ptduIX6dTwsHqU8V7iBnhGt6UcAyotKFaP5g+rkxROr/2LRyFORBoZ04gCdI
PFnFvzniPH7L9sl1p8dnVTJ14PpwAWMv7O4VPkzZdYr0qnB89NE5ZxN9CzV9O3Gr
Ngk7LgXgJZau9vVlD956Bq8T5WsF4P1rfNTbjQrTF4XExmem8cT6AQCP30NgtHJ6
1xTwjItf6Pc1Ied5K2y9zN/zbP9lbPBYaqnzhsRT3ktVfChpLAW0ODBiWlt6gC5h
gUOeuYFjC80k3UexHEy8HoVQ4ZjUejOXNsPFGZHRxRuo74tWtQMIdrTeQ5gzM6Av
NyWvyyEbQKXhCAoY+SNF9fDq3aHkD8FeceRKUgLo2MJX3UF3LX0f8dibuHa22EhI
z1Ll8kgCuw3+OxogcnBz+E45KpIxuhJsjHfhJVSCN6vycu5yKFDUpNYhG/fajAyn
1wRJA/oJHVNGQwIdiPiQaQzuMW4i0SuZjTei3XfTW9skQwvcBSfvVMAfDLjIMmJm
YRhffhD6+44yVb3ByR179JHjG2KiP3WlL9TsTt6NjY/Ti0QiGwWRbquH6d2tDbBv
7DkiLcWwPAp3fW1vljouU+7AIS06YO2qk6iL2AEbHloZWRAXRwG7XicJwnCn4OwY
rHjO9/8+7FZlDN3fG6TYJ/yfLR4L0+Vk3tY+BXJDi87LcNoH6tpC9gLtoJtBT/xk
W5bvOGXWLfCVk/FBn/adGVX3POt4ZZXs3tkZRlU7weZqrhkuwU3wYfOluPZa/YeH
25MS8TVbXAlsYu/9jdcj9ZgHpkriYs0lAj6W80Zu0nnw95nl9p0ZCwv8TyuPAULB
AsD0oGoxOxaGZub35T8ocFZIrbivvgXAKj+Dc1zFukWq7byB4b2iTKJrl+H/mC9i
s1tvdLFHWS+rAnL9vdRfTn9DLZQy0zdURjswcpOmm1MpthsPSCurX6uJV/6Fe8F8
Wfo6VAgWyVe/MyEndN+SPRGqaZUMiMxjv65XIOcNvSXTk84/0KmPZzhZ/dAQm1BT
UK5uAwkHW5AsisPsOhpgdunyhordGXtyqypJYqHfinlPqjq/UVm4WUpQzkfIyooF
/lc95qFjHxlsiJ281t7EvxYqUR9qbsVbA8GrceTPpeGxPP6Cl49TqUo1INJdhINR
JEx4mAtNty0NMb26zL0jDDJboCpew7SuxncVSbIN9mbxbWo9GXNpNknNndKjH6Wv
S+fDslbqID3hGcC4/L+YWVkvym8vNw4i7D4QI1THO23qx5hEySdqVbLBDBlBIu5J
ZBopvlbDk55eTOFDDSyEWHcqMm4aosUZBHoB0MSteVV/MsWXP9KQSTmNRNJc+rAW
AlOexOruh6FdiGUmrlevazC060/vHmcm43C3N1sUlD7wPFai0Ezmv00rRLGhIhXi
QIZaYskd6x2pltmP61QVPGiUIP35GFWo4ylyr0UWUx3NGnFjOKDxaaG/w0gHm3IS
CtnmvUNSZ2PmDBSUAOumpqmcA3LGDdXnDpPo6hOH1wyeIAEsBrj0x5pePlKpFZcO
W4csLck4jUN5NZ3lRp8KFj1FnDIHxp/F50qpkkHkRtUGNOZ1g8PLe36MvZXyf01E
LMXRYak4wAScf+itK2jItfd2rM6S86VpyW3YWrrpxgjI3InKJ9a3W9jk8UsVTD+z
5iSjBWYLonbYeQ5Xz3jzFHPQGWgh1gE52rKZX1ml/v61IZ6rQbOB8pygeSjxqyCH
aRODvGEecoXPDxy8Pe5zyVWZQsA5tOqZrZ/43s130zrUmnSG8y6jtdUWlfaZnTYu
Oo2NADxRE0xv1ULSaACB1YFOP1u36GL2DJCKV6G/+tEZBM7b6L2RiMX9cKqfp54q
z2vPmX6l5/j5fqPtayG2RPxZdCd6riwbQO0j6FmMOgm6lHJelCKSf6mVG+fL1vqx
glhOTPRP1VnbpmMfV5AVavz9Z12yblS+LdzLJfgbgVWHZ3AJdUZt0EWakve5zLfW
DPBP0kwzQpod5pgvJCQivcdvlGoCRE5ZXARYhC2c655J1wm6Ln/1O6yPjJZZkSaM
qKk5Py8L5/0av1rsIcEGEjY3m8XZMJceqtg95pWie+Nhoan3+JEAcbgcYI9TA2Xe
qM9CPnQ8Otmqxlg2CkMyfum+QaIDOw9n4Ud3mWnntrSaoIDS1pHOQ382XXmAEVSd
02i8797amjxXkT4AhF4u19j7EogneknhSFMDRFy6eJOsJarfUChe7q6ScNgwRkGs
cDkDs9iWKImpvti6RInyd/6EPLNapJRQE1pc7mxSSMTfwjCRlb69i9ob9hnnQeMv
ZCiUzQCV56HytLvvYToAVaUXuZXrCCspyyrfhSzb1GMMA9NcKN/SnGUEE5KVqeQp
ePmOkK2EnLCo1TKaMigG9joWavgvxJxTNSyWz9g8S3kDlk0gQRGP9mJ3Cnb7/4Sc
5vxfR3VfN+/leSFzM9k+Rv8X7CVBYfG5ScP8fMRnDL56IrMl8xTv1aC7ltLjgQcj
NVEHbxKfSQydt4T4P5j5ER71tRXhdNv2YM1tNYk1ZE2coWT0zmHbyrPQldKf1Gdc
HKAo2Ok6m6TZldRjHdSpD6xIehaUgiUod53xXMudeGOtBqDMMbPdD+aii2nP39lb
bvQHRFZH92DoiXzZ0h0MRIHHWRku5wpJ788qNJWhaq9GUCLaUE/2qYE67pDtUbuF
wGBR9x3tjrFXg0hv3pJsziWAkVn5vgfzDjlzB1fQ6qPRuxkoA2cL5RYWfeZ13w/t
BcWfByfXQvFftcjxshNmzbjkgvnSnv86ruIg1Pyy3vt5SVCklMGSB0CrgKZYKBHS
XDboQnAN3LCxjK7x/aOi9F3kgT/rUXCPKaUedx0bfD08xWigF9VJOG+swrK7bUpS
ZSjk8N7iPIq4OERKNK4h/sfqruWUcu1tcz8ypxBHe0+Z5I5Ziuk5Mn20MN8MQVIt
bLEq1RBCuS8SLzGt2OBbJQ1OFg5AwBzwx3r5llUUeKxNlMI8FeC8FpU9kyQJfSh0
a2o07OlKZk4iBVg0dAbnXT07xC8WPZS6lhbSWTp1wSMzuqyNPkOxuSDL7CEmO17j
zmMx5sEQzx+MVge/xQq6SGeH5aEg2raaEG+YVRNRSSh72D6Gt8o82nsOAO4bO62m
XHORKWIdYa154AyAVbCocr18aVE5hBb0idkFAdMM5ok0WOmmV6OpsUF0bOBkbKvH
VpyVtHPtBzWI6toZcnpZgMipMyzp43HuTVqYACpMnx4Gl3ZvxGRw4+VgXDIIXLpN
ybC7ZGeeHpuMBPwOh5ylOYdChpSrBaEvT58gHYhmpp8ULAjNDoU4mlHSuCt3gYPA
M0vpS52KkPhEBYVOmCe8VF/hV3+MEvJC5s5s3dFvta9vWmSV2Sh0OksXKUvlcGP0
0V53qFdaAEeO7uzs64UMJSY3Z6CyE28aSLgjJA8yiQdNFKFDk0pbwLs1j/BgsNff
uoJWDKWbEYhbwTLZNhyqEC71voIXMutw9zxj8+ra9DnxWTl7QEsxegv0EfDcO8Sc
egZDbqQyBjGgi3WUyWknkkF9aMj+E6bSkIpFcqDJcfeVhxbkZ2vU3ly7DBS8SM9v
lr4hXF1q3a86fVFe77Ue6z8czKaLvc2vBL+6F4s7biXERgU03NYc23pL+duptaof
kn8HIwZ9SehG5G+waJxwSkVQMGsxMdAjtddZNd4QCEOqrUss5pl3UQTQgcrdKpQy
D8Or/3lrZZ479eY+vB8C55G4nOFk3uJsC4hojvLIyF7pFlaYqiIe5AAYIVSsB+SO
OEYzoMn4RXqLOlIbGh2oGr3jtGPqXVlPSAHayX/ljr6gIk4sbDVq5XN+kdd+IURy
gFSztsvvlB5dbZCfDQdpZBK/PjPWNTXqLHOLcovlG4cIY9PYJAfcGbqa8q98Kv9m
XILVOaavoGYjI4s65lS6bdWhwAs7ytFXszYeOXCpvysuhsVvQklmPNCrgUfKiIdb
+HW8h9AARdXuw9IBzfbJydfxC2iKkrwliXdD5uBiaPBbeIRAk4lQ6x844AAxtt1n
2/TUBlyfcKEv1mAY+CiBdGXcid+UItmQr3ffTcbGFfWLh3i3QDWjPQMR2zohxS5K
5MRya5ocruFQpVMVxthRvhfnABhj3wvSezIi9vZ4OT4vlGKH6cFtWsTqH0h3Kgry
AG++Qt1e5ThNjwKLuFjOhFiTF1wEtmbvFHMj34qAAkB4gswabY/27iRWD6jS/fvn
JhdVdG7KJEb8gMn1FNuJ/c2m1KagYsnC9gcYxmVXNsQnP4qtaA4GIiEU359i178D
RnFk+dEfJmvIKXr61qEfz2ajRLz7BVM+EUl747Arkl9g1I1/DCotTxuk/Y4H1lFM
1QHBfd0CjqdccudpBa7qBwgnD9Tr+NEA3WP5x2MLuCcoCiuTOW5VAUuveotJvlgJ
fJYI+ptFCvTIXz8drudN8GEgyxYAFq4Pa2tZ6e9VyS3WYwCS7f4WjGWv+2E6w+lF
MH7wFALV/5M5yqcHeq2HOVBU/3ihNRq1nZbGrjoj/IDMchRxLwwHWHKrXoVuejs9
rILkfAL0m3kUTRNtSyxohP7XYtdkhqt79MtfuE78k7FPmWeJgRIU7I1z8MCzqtCU
/D6K3IMG8SikvX8zZupkMp7lfTRU8Hh0++jxcXopmCK4UbjhHX0ISAuHz1NoJvR7
CPOgedyfkx74TPQvIaFKvWouU+CUq7qNwwnrZtmwnIO2Luvb5cbNGj3hXtTM4IzA
cp8+6rTYLN/qK3MsN5cMWwDghejK9Lts4SqT3NC4RDQwH092bt+2xSKSYm3fmpvx
ZuCZUcwRSFx/QVlrNhsBeJxQwVhYmHFydOLrrh4CfWqswy3sJvgfULKX5Jqqkkyq
29tZ4Wot6n6eXJ0IsW8RH4bUxMiWwvJz+xPBrkwt8vhudS+krd5i0SGhAq0XNVsc
1wtbCXbCutkefn8VAD84YpuB88fZTZ/NqfmwnA1/cKGmQmDfFTSv2kA6JWg8XKiG
YOC8XAsXNS7cAXWYKwLcy4vU8kM1+T/A/TadT8LUvIQtGmQdX/MB5E0tPmyGJDBB
njGHolE5brHTPKceCLaYI2ZxfuFkXd2WVCeheh3VqoagNAbrhwzlL4p7sAi+n8UR
e4L2OcZ0NY+2gliSMbHN+/exeugjPLSPyCvcnbkjfYsBilDojpsB8gKCUwLnO091
O900RjcJ4qmp/sWtVXQgb7M5tleVdnlzRPpfJy8qgkbWgaxJbgfR4mrKz/m6x6He
F9OhihcPZ2F4aKCxNPIzPzlmalVJUG+JJnZ3cqFS6c6EoG/+uUjXvo8uda7zRPwb
h2xpJR4qdlm71wSbRO07a31f8EGfsgNwqO6kOkDmOC0kHXcr2uqqq1NhEI6HamSi
KM1ZzRO/KHTJLARRmJLK1PEaGIuXv1nYao931UVeYADI7IjgN3aueS6M6VDBvWoP
1Tjn2G2gABXcW1wep7c194RWheg/jiDt/+67FOYElqOGihjGF5CNZkw7PG6oBpnD
i0lJKo6omss+a8SvEoxfN7AYiLaImN/IcxOY9X2QNbLTp5xvIWZ2SaWE4fqLLW2B
l+sZSbE6s+Zlf0ACdg8s25ScdW4nYSj4YCOG4i6DMAGIr18z1oGMbaY3jq1JWV4H
xvx1QKXLPRw6OxkCRM6Cg5Zb2udNjfDDyF3xCnu5yfkHW+zkRIAuvxWe34W9HLyf
r1rNv31+IyxQcBZmHoEWCdgWMx+F2yeqhCyM5DIECGN3LxlSHO561P9KovfxnbYF
86eLGuh/WSduJ8rvvBjg3AqHU0tHJaXCT98JgjeT9Y9Fo8N2r4sJopUy0SrasYDz
1yhoJigEL0M5hMDoQ1eZjaW1QVQHLD5fKo1oud9uUJ2VKI9KbQVt9r6R8NOlkgDW
/5OzVtiBGGJj02sJ/HwFejORwjicLd/raDQEb0H4KLkATl3uGfJIstG57bZRldgE
L/TQ7Fe7Xxzzd3/XFGpJuV5HVDNCZ6jcTx4yV1m4t2xkX4yCNakdlroKtzwQsYLa
QjxJexSRb+h8GSVJzHBD6IJFzrdKgz5Cz0vr9YWCGW/XJTOBt3Swj1HDX+aQ2U+b
H1IEdq1bLLOa3VPNQWGTgl1mvnUtm+bxlpOFwAOU2sW2w+o8oNRvKkVedVOSwr9d
mW8yIQxZFsTftg42qjiOVScGTp2OSlrzqkvGZfXePzwpRVpeS7newRVbo3dcRwFd
W/B/0h6kzxhN/kpGYJEhoO3f2/jrc1AvfkNe5CTpVJBqXxBqCWUR3SQ2hl6MHCmc
JqvIHvra0awWFnoVvQd8pJprIZQNXHZu/tvrxvZLNw0YvgqIUoNSq0t+mQY0coby
k1O50oJ8ncc+wcTWWmY90fNCt9aXyHvMT6HZY5MlPxeVLYlx+FRCluKc8hdkc/nO
lE6L/qfersZRW/taEGMHcJH9DKPS3Jt4iR5bTZ/dInrE2rhKWK6eqnKlOD2Bh5C5
JkZihLiJJOxxVfmgQl3fDEgFFiNNUyg+N9jNnHGWTw1o0NmSiQg3RxT5b79/TH4o
nFbnFrCnBpe1AflI7RGq/I5FvUwnCfgljEp5yyyods0tgqWMLQNt4zYq/syfiyJu
cllAaTZldM6nVxK1B1qjM1RzZ8CJ/xwpaINJYSZOfhMH+Xfc8BePZd29F+9lXIiB
AdeXhUTJL6BaiB/4NAQh6cYFnz2MoOgmaDHjlv00Mq1eUso02Fg6AcvFrJWnY71+
fguFklhAWdMs0ugNkTUvlHZtxNZImpClPogSltUMJaoyfU5GgNUIhL+3i0R1nwTF
1HxiV3q3FS8W9c47sMFUC9Y8XP8Syj8VaFf+iPzhBFYlel1I2aFWgP3+JPpyd2oS
lYq6fgB1KVVzADq6a7kW1RVJ+kWc5NPK3XHsnbEeU4ZNdevVr6XDg43D/hLdd9re
U35Y/O96OHAqUcscfTTGzf4OWSneJNM7EPIqI1CwnUTdkKoAd3xWO6WAdjakmFdP
yPxmqPBcaW3KQIsLhM5sjOBdaTnHXdOPGgLRiTvKxKuDjt9BBbDPv8/unFyB/ADR
4EaihsDc28btuVheLHzxBLQ4QORBdmjaeoL3PF94yc7hcUZSdjX8iMfSdDc+iLWr
rvxtKgegsEb8vI1NmSLbURy+vkqfuPxjz3H5ydw5FrEqfQ+evQmeXtoHbtii2igH
cUtUAHpxy8ZOHzqI8WMCEYjaxZ0mfl2tN4GbCYjdC2JnlaCVlq3bUoE4OyhqvzoI
x+Xqz85p0HtfwNhSADQQksV3C7/uXvkfb8jw4kgKo+Fty3sn+kNoUbL8syWkej5K
i3ZedIVkHMn8jwxE2r7m7u/R42F7pN9VPs9zVXeU/Cl/Oj/+O5IFb8zr0oFXLkrO
I+tttonG/SD98KjICmVRUGx20vz35g1hUhv2YjkNsLEoKeoPRomUFuRePOHjewiC
z8c8SQRCaMJz9gL1P0BHigcyMKhpOtb6gyMU4NfjhMH2lXSQ+JUFJCbk/dVf0UYx
rUi8X8jb+a+48o5O+RK5VY4Xe1gPNLOT6cp4vDRv9HWkNv5mA325A2by35aqJ3wa
XUuv+Ndl6gimdoxyeEyyoL+BZLzTONXA5ACrE5ljjf0d1lg5Ls9K3pBb5DbRZK2V
fuwxWlYGTeKjI7WFe3xiaIkkqPlXS3gSEJR411VjOEquOBDdkk4AiAYB0fpQnn4/
ihokDExACohSMRjhDeHmhN8+5vNBPrtzM4NpM4Otfc8iAOmHJb8JrGmvZA5RHZSY
DvGin90ZZqmC4K20B6Z0W2Bkvs1XvG+3ZAkoOdoHzEomoJ2rPXdfH7ff3JPmf8zz
lHNVOm/URbtX9xQEYHrvhvjc/qqbwZ9aUxJ5VHZQEgZe4ZKYRDXx1R1RGi0x81E5
/5ebA5yzJHXr7Qf6kQL++Y3NAlC3a/k7yQfynMe03odTbNV7eChfouCs5apXAWf2
eTsy0OT/Vk+/TKDn7/KXo/ZGv1dkOmC7zwMH9X3OSofQMdnRwAWP2Ba5d7/xa0TE
2l8xdYLpRgBS1brXU10G7ew+0rqCY1tVu27rVDb8h2y3R0vb28cAAsvs6wNBG9O+
Op236QqGb0y/TY6EOI4RV1Z/7tazEzJmjI0VrZAcFm8KBecEoMCvoFma4lwnQrN7
KXEVUKrFgaS40HlUgm3CV7YJuhuRaU9VVwwaijCqrKSGhVqv+z/cMs0BkK0m4fES
fcCcABmtWxi/ERTJDsdZrPEDYHAwkCAEVxJRy0dQXn7/jhgedUvQb8uigFjQ122c
8VdiJnRUhxaeE5eM9zNIVeiVMPPX8LbkWCS//0yTnT1dfcz1cYiMyEQVv0JS8ZDf
fTpOBMYNGHJVYKqe1qkUbEY9S1OsPMbGYDlA8FZXfxUD7GnhV48jKfjpBdOPZ6Fm
mKEqeFTEJjvOvpXa1w3a8Xc1V5jUxPCWoz+i8RpS4TwVLXJPDMkfTMekXg4lsC68
daK2o7Ts/qUpOdWMK9TZeu9h2kADDHUcVYzOvGAqawBmreCrxcU6/FyphUmBDhf0
qOt9OAVeUHYqbK0ge65gypC3kbJ+UBk+JNPTmTHjZwssVGuVuJRgziz2avqLiAqj
gt1DzIl8q+Te/JHn6hHmxetvn6mbeAni4eFzYTkUl+FLrhF/eP6TtY8WlFPt11Y+
VRidAGQzB45NdJF4Y+5C/tj6n0+bWXFTeTCYtYr9PxC3Fy/CkWeaXKMASuGOq8W/
6ita1PkGGXBtRFL1ktO58Ixt7Igeso46b2+x7T1DtJZbbtQdW0JPr8Xni0dysOjv
cDWpfo70fv+Q9EVDrmnKU1yP35gSEsRw0SawOn9mriOT+v+4EtQndXD0PeVTq1ru
ZBg7rbSIb+2T3bO7xcbIjVHO1TwxkVaZ/U+r2raYwAmW2La2gqbZpzm0O9SgRzSG
ZgCKVPKcToQE0w1eAYJqTKVlgMfRS77F5takDeHjDkZ5EOvUya8opyfLxAs6Hb2E
MBdWg47aUqkSMn50HraD9ptlWIwl6C8GzL4JWFfn326YGwrVzUpmf1BcPi03iI7D
aCSMS2JJkU6jwMxq22qMBQm7rA8XoiA79o7gtcjBnZhvfqJai56sFaDfGyRCQy8a
dpOiTNy70YeUFubvyH9TETxqrwgtV6pQPvJkYdF7fUCSkTfo07JE8uj75UYKgiSI
APWzMHxl4qMS4RwdP0UgA/bhriOW3vwlOVMdviYcSNyeZ3VMRDn8MnFdhp/WiUJR
Z6SoqM6KEzTxrH9FmSlYiLqR8Flpt5E06mxFMMgjHSEEdumTRn2l6iZaKuRP/nGM
00YcuU7xZggH2gr/3pIUdGcBdQ67mljJVvyxUuvwuYjjhUiFQYFlWZWEIcORezK1
ixvgVDZ0vPii/IpFXSbFCeh/VzWNIVjE78SGDt/Yw+QGqvoqXHd6pM0okSVUUd7+
QPq1vs+63jRJlOawr9eVDYU6CyxeGJbWI5XQ2onY9xk/PuiLml8d/CftFl2oWAqG
/Fqjww2DqW3euxVia5PvT2X8aa8WuBIygmmUBwyH7fob/ACzGLMrItnMVwSDa0AM
sGbI2EnwfhlJ29l3ZvGdRCKay9FMWQIO+leQ3ZIsSV9nOwnlX93X1jCUgNIt1/eR
Od6ULsP07b4QGaCDFigA/xIkgHE75Zsmm7T6e2nb1b0o3zpe+0phcq0OK2iktCN3
ZQSzGsZ7d/9mnRuLtrHk37XwUmpQbRtqnRxgDtKLpsBHB8sWMZ3adXMcMKhCSW0G
oYBjIl86khvx2jT9uGcroCPD4x8g2ax04VMnstHSwMM8g7fxGh8ZfGm9+KgXphVD
Lt45RqDBLVN7dXlOn6BuiGtpk2AOyo8PE+kZAr5awZJ5whXz8+yGztYwC63qXjCo
89HNQc3Flr3A/cbHUEb+XtEoK/JxLPJB9LlMXJAJGA5fLYJ2kT2y5HjibfXOqR+x
5ABQsqKr06gyRKE2BNqZtNL/JNK5dz6wSoOugFwTVG4/SHDezLBYHxofnn3qe92Q
LWP0IA9PWN6XbxKdRSuJj0BkPbjDPdbx67L6767lxhONL2WtDVU6p/TeDNfZ0HkA
jgNUrbXX8FVaRMunqgS5hWyU956ZUfiVZPGMDLbSPY/T00JdRODpTCJf4X+Xk8ha
wEMGkceZ8bnPF96JO5ipQfurvtf29lzDew4BqDWWHD1ICv4sZ/ldZRKVEqRGrACh
RwnPQ3aSnsU11ZyA6fnWdtri9yjUZhv9FbQKj9MbZWduOc2sRo40fyUxBy1ArOE9
lxJ5h9CHPyH2ecSuCfl1Re02v72QYZLHTHZCg05OTmTdBxZtKeinncLs5KWHsSP6
BydrF9EaN59QctWLCxl2ZGUNVZ/bNI12po5evh6GCDqZBhQuEIi9VQeSjXrB9cAi
S4LnPnIWdpp1/IEpE2Wfa5EjFUlCviyF9y1C1+XudkYqhdtKAVoGRsiBiM0aVaQZ
7RLB2z3b9ke7AHm7rfUpJC8su2kAXFiqctywFavKruvj+0gpAYefxWfifOMZ59bt
1QOj9JfCIOTmvfDLIO2PZBF/0DwGOyqdCmkVT+h2AQ8LZP9AbkI6wFRN4SKPW8PW
yW7aDf3uBJi0Lcxi7OvNs44NXk3KjlV6eOpwwMRuz74qo6vwo6VOSXS7bfwkP/o0
5g9hQmTZKne4qnYcYmeHzTuOb96AQC9pKTyrDgUH0xxeCiD2zue/ReQK5PPa8iUv
vNTqzmw7OeAWTuPdVj9PymIcgqMzBMfzrMa42jQjfyCJ1EHu8p69BvnE0o1gnoBU
86xF/qU23fLAWNd7oXGkHDSAWvPLBsJtRYzV9FreWhHMjYS5T6t1gVh4e+W76TYk
cNnNG8Wlwsfyku6uMl/mAU7PURqAU0bu0+K9UzXTfA1JVv8sr4D0uv9l91M18HXZ
F6C8Fo8FV8TX9//yRKAoHnaT8RpgpkUpQXB0k1BNQUTIalxxJec+CztmEz3AEkMI
Oo93cnYQmr9mdZ0iM1fHafwDdxXVvcwxyIHCuqFCX9r5sy604JRaD0W1YGm0tMh9
mgAo85+Ito9KPAZjEzTtXWEcL0rpKopAnaZ4cl8qMZjbGV9JMeJ1d7jgISoOGYdS
7zeo1wO5FgB63AEnpRhm6dnIY5PLlGRPsKfQsBocKdOP3n8n+7CEhw56XPltvvA3
HhlH/AyVIPELmuTtRZmAjpWUqa5ItR6c+Alxm2rPwfiKMD1Vdz0gclQYSvSECoyo
frhNGoRlUhaSN3DGcbb9LvJgnKp+lkMU4MXKbkVmbrag/HlO9A4NRaFNLfc4PKsd
SAc+SudNONGD5jrVFToQ0S5wQEQBzMgr23iRebSDwOOPhweWesJSqMJxu0oqiz7J
TpiyQiqjtV20cCUd+mKwQaVCcUTWmoBWbW6jKuhRZ4vcMpnlCULib9ZHQz9YNsIY
kQC+fxNTHLRgwVx67oRP75ouoR0Giig0yXwRmHofnls2AKoTyJLd4lJPLnzSEr4Y
FCu0xZiSIRrcZ3Ir8BDJG7vWO4x+QrvITifphbL8botOydh2S7sJ8/GFo0kazwt9
qBP6CYzDcIm0HlUbIiNlh5DlQfTlWt5MNrzFSRy+X5ygwhoY37Qg4DYqJlVcBQQd
4EUEOg5frvGXsZJl/lF9uec8+9xZ/dJS07z50lAJLLSoaf6QoNZ9C9mZ03mVB3Pc
t4e3SW04Gh3nsSzjwc9lx9wqGbBrqmK3qNd2mg5GePDJNGPTEJuyLg2GOWv5v7TV
y6Zvf2jIECBAlA6wJMKqFr4llyy5pm+plBnKcATlLLwqi0PPlN6eP1xfWvW/CxeD
zYvRXdbwT0G1Adpf4zKkIwihy1gOGfueflVc0ItPNGlVRcJTVoH7GsTCIbpsAvcR
PhTjRS1lcuPiAcyV5/jBdFS64ut/BVV0gPc792PE+w4GP4DfhlRsluOIZV7vgE7a
Ex87/2k7REz+hAAQp0j/HmUd81bxIEPKQAPp0HiWfrly+BuaREXoXm5wJuEiDw+h
Am9IiKTOmxKmwHDO0DQzfPH/gbo/TBk+5isHOGu0XU2a0vWAriD2XhBWGSOVIqXC
FKkgVriZcg/47uvNBw+gd8kv2CcXCmIMPpXlnf1d1yEpD5ySRHhcp9mgX1O0z+mp
5p7NrH00HJIBpYmXeYtk6sLkp0lE4//13W+s3T2nm6j9N/kI0xJznvY3DFudFtTT
tydMERS4K/Sx/zoQYtthzs0faBotAb8KdiyY1g1hDenNQ1OGFIhoSr3gpidHtDMi
3KyrHWUKTwfEOH3zUwD0qlSWFPXP5kw45+F87PFFG0WSs2NzAfJOQkcpaBwX04kI
4iHVrIZXcZYOBJ0ukWxDgS2fYscFoSUPUNM6/ktn0iGU+EgfGiED34wfEXxC6pbR
lRi9VkKgE6NepsmQWsyqN+tcUpD8usz5iyPC3hsoeIm+YTySxFLmZCTLYpPpTCe0
kOialGjZWKWeuUt2Qn0ekpBZLT/kdXhfJAUR5FYpqAnmAGAZG7bvBC+205Sg+Y1S
1QrBMVhSq864+1Yvwzrxo6553ondCraJRkaWjDOdHFkakRvbHyJldspgzUJ+eekJ
H9NUluZMbO8f3GuqFj5RRDeeITcIlcXa74cKXvRlV4iu/2/wFQHVO85DhE8G3kWI
VMv+vrhCUECuTe7+Pq/bQIhP+D+CBGThMyx3DeXGgJ+Ptx2j0vJt+GCsYwM72qLQ
MdLUdePKs1pGfI40r/FpAIY48wEFEXLLua0CCxac+GY9ZH4AXu8LzDH2xSYa3mNB
hBa8T0OIzKs+Z0tG6ehRFsT4KVsl8C7HinQr8jMu1sXIvaH1loJBGb4BxffWcY2A
dDoHMls2K25P8dOdVUqCgXMDk6+ZNAJDLNombBBEN4x/sQDKZyhIN8zSeZ5Z/l3V
cOPh1Dw3pYDD5BCZUofYPyG2sfy7EaIHWsU0+MKWhBl68JXBLVUyOk4BsaIQoRHV
/yOGzZ38fwFWWOmSwnwEDL58ZAragmlupRZgbalsp4kTvYqLHzO2O8hiMRMV4km0
Wl5/nbxZSRHL3U9esv51Ma6S3VsEdISFPt5jZRAGh/jRJ/c+tmB3q1D9cz2NxRGG
r5jJ+gOYS17lhZEdxpY5XfksFp7nVMSFbHyNVpVvk9///HZFgADuKow/w3WD/4xM
qQIkw2N41MXYkhh2XmvJ6cCubsUlFcRdl4ZG3aNA/k5hUS5J2LD/jWoVDznJ5sJM
qtgQf97nUV4J+tqN5mzSM8A1LEg8L8FlOlTZQMzOovVfhmMdedoPxMgOjqbPH3VU
t/uCbWa+J0wkFYqWbLZjcNPkbSKISoJPr14p7mNLuBKHgN5sY7K/nAb19pWEd+EW
EZUMu2YR/JByquqxGIMOKaL7CM2UDeeNL3K4JpsTgILasz+Tt/wOE2kGXXSRjg5u
xSQaU3WmuAXWRR9hRyIh6xV9dfvNhX1PMGL/nTJFpg1eu4hPxm/0DPINK2YoDlLx
8paVIhELBuimRb0mVSmSphPQw2WctLZJVPJN84Tjy5U4A1z6zGFpyoIBYB+LLhrr
WtwETNCdd4+MkP0l0HQp+jhZ+qjlXee5eXrXnRmdXrr9jaxaLlIYbQjthx2VQooO
vahZ5d1Ct+rdGO3zt58Dfo9+RjqWrt6+SWKzEqB0bnfHJEBC/eAm+k93+Ftp9Ee6
wLrwnbEs3aFMHPomRZvFCwIBCnqrCnqHQeKE4TqwhjyYkpKGiljZCvKRG9uqXvNK
a5PsyIyhiUtBNWPR2FpgWASaEGac0mSabMhG58iB9+jiPRY/wxHSpI8Nd5mzO1ul
Iqa9aTcm4cs/CFGc9r6VT1US5s2e99wttAnTwri0LNGQo/YRUdR4na+JUQdZifi+
hVmTxoAnFZFbFFgpyEjcabCa8HM1CrYQI1ZZE1J34f00SLo5cnEye8WvSg5iRc0l
rRM7XnAoQ8572/LBPxOUAQOCgS1J9uBukvWYPDyIAd+TWgAh5H2G2V3kIg73QHgd
HPe3ikRLnHJAPf1Pj3pKzPNCBhZecUS98hxwrZ/UI0+TbHnQm61r/1mUIvE6iFLa
2HuPSD7U7E0k8PEtVuAGj1zRZR5402qEvyQ87O+hcoeXFdkiXvLh0WKxcJM+Mj2I
S3lhIr+5J6k+twFcIATG62fGOx81jN6diDfeNFtNZMBuhaFyugiBvLdADt2yF4fW
XOYQkGIc1cOOl3LFJcccq9zBsfXqtI96hlSCed3ZHd/2XfN7Fi+mtsmhJFfqCM3x
GqgI0lVNXkKSv8a4L/uEihbdsYBR9MRkVgb145WjnEWmFJV35XW4l3ghBn77HfQf
nqcqkqeUDxzFJ6IxlnO2MR1M0BXbWypGwbgNdL1vXcutKD1b2ZbEfh2yWYg6XcCt
Ae0yymwk4Roj77SGqxqGD/vlAsC6Fy8xeEprUAW8DgMPWx1QmyJOrBAeIZfV0y0d
pi7/nHzR1VXRYgP3aDx4sZfTSp3DBfxxei6NJOfa6uBarejIW5+kJXb8A4rPaGJx
/xzM3f88+EiQGUs1PhzsQBQTEEins4znSokTwhPU2o9MciaDcJeuuwR/TGIIDfvD
DsBCshh6FFR/EmeDHX8LEWqwpuab8mHGZCH7ijkssibgUSzISOMVLOzHuAJMxk2U
xfYAbCRPb6JSFlae5X3HGg/U9IfVyfhOuv3THfPNDkZN6J/w362EaQ2zfJi6s0Aa
OreMC1EzkhI54LwfBCfLbBjdHVr7Xkr84XtBvfzVrl0YKasvXOJ6kwoWyydnhEbz
IcIpQbXX2tWIe5yigpvA1JuL8/Vr1GxXpDJ4+0AsZwhTc8eVmIs97NiW5+mb6x9k
KfrCiDQ7CAmJh5eDM5AUgjLEqVg51avkPUAMXXkf/jmJ34Y8mY1RC7XOWLTsPgh0
r2LjEjDJ01XkwHZvA5+cwTdrAf63BQoqufXlz3qERkFmkN5/l8P2Uu1Kp8S0iWkW
xoGKt73PxK1f6v4OyIeIaegfzOamcFR8ZQgMVQcegzyXPGw5i5wZzGYVFJZHwRQj
VG0FtU6dFWuruG0sLyx5XCluCFBDeb4tau448uaTbp7N1Q4Wzj/QE3gXEnlFL/g6
oiSHSjI/rYAIR1DYN549n32rati4mUwd2FV7sLQQakdB5taPmdYWjyOathEuK7ke
WryHVHXVET2Ok7JL/y+ozE/hNLcEA5xDYBf93AtiUH8TDXZxlfIulEaeQ8bX8VTL
uJEun+ichTZyzr7Dwb3aifmv5ElC798ru2AlLqrFjvIeKp5eVflSKMt9m+syVgee
aQVvKnBf7ISD30sca+6TU9IzyNhS1n/9zlTLJdkpfRWgiWB1/XYdaUwvkyD8pA+q
dg7jH4ErDtOgkLUvMdselO2QJjPeNkcNtiSeNwPNi5Iactplj1HyRYsTVnDyycWS
dsORCL3IDIM9W5xnTieggHKN0eZrDY4eAS51k/2VfXXwSv+H5ajb44W3T9N46eao
MuBILYGMjis9WRTY0lXIX1XZ+HFi2KVrzLvM/8NzCqjQ5v6Z17dQCB5ZX8lP591V
Mu4X4rrzdZCSUYJlGstKrJXOcCem1u5Jg7fQE1mnLQ7JiOTvMfLKeBHKD1lB3cKR
i9fOqxQPp/7khcxvDlDv7KHORte5UBoVk8g9+yAyrlL2APx6DQLpVoIe+QZJ6f3o
vYQNW022aFp3P0QOYFQ/I0S27ycf0b3jD6HnwemA97U9nDvVW3MZmar0sQLFszG3
xn7/6ilkPATYwfMopnBfm3vqWZhB+dgN9W5NKW9w3/5o25D3fQIT25lcYpUdZfbo
Vq+JrIsW/EQn39TkRvasbAcwd9KlptvNUlV9TgaP5Q/gFJTvP/Nyzq9zidq7sXeC
1NR+c04Ckcz9iI7lpRtMmH0XEohm8ysEBRbhv8Yz7jHXuZdQbgW/5EGG8xPxLzUs
nQi3QCvAUoJnDlFLn7o3cLaejZsPfIQIbi9KcfRgHWpw/JwG6JvNmUIUjbZ2nGYO
/f9YAZzBJowlBP5v+FEtiT3DukVI0ZKYFpHwPS7Tq7FdLKiQC/rjgdwbebM05qeA
TZ0cuP1dJtXoTmFzlo/x29VSB/ePfyCeEyRDtKms8vhii1rm4lYztMmBD90cBXZk
HzXbWTzRvThwsoEZPT/4oV+Ds/QuYdiOkXhtWgFY9E3hA+j9Ef5WFIet3P+SaUIg
PkoCgvbYWupvUZzgTw+yzPYYy/X+ntXzV5rPpwK0TUvZ/IGID4GokOlHWfviZOX6
ECy3E/D45f93q0yFKVDuhJNU+4GS661P2VRl4lj/zbgUVsBZyy4EYvcA0csBY6fM
4SbX99MOnPcMsnU7pdDNWAT2sy61G6W0JG7pV7lmbKibx5nWrROrRBPEt+TkijVl
HTRjrGwuatQ1J8t1710nS5gVniPGpViBjs/jgWt+cF1WLgcZT+R9EUw6sXDUipKI
XeEQOljBaeEwy9Vi9nuF6ec3CZhmVIPJPfqfsCANYxkkA+2U7iNPfMbnwHCjhwKE
oci4aGNCaAsO3xUI0Gpx/VB3muh4hyXDJU9s7fTV9KNeyj1Va2Ai9K6bPPO9BVPr
K1YiMIwhI5dMH6Qta5KIYsrR13BpBxP5HKUG0o8RjAqp3sl0ZrkjeuH4ixHQaVMn
zEtOVTLq3kQqvFtf5OjO7jIHU/a55w3e3LHHlDE5BAJBrFcltvJxbwc7cNwnf1E5
qYBQRM9K/gvmYOKxNNpXsXc+uB7QOxK2kNxBSmkOSf521iOBqhZLgzBIgiVuEyxE
FDt1TKmsSYPeXuv7qqY0hsF2VuI8RuNKs9pfaesSN01+2kEPwC4jflNDBIJf0uKh
o7XEVr8LrPVfuWzrL4gAcEwIH5Vf8Lh/44+jYD3wDNVE9eoyBZYclD44HOEfehuE
W53XXX6GGkCJOM39G2JKs0COt+eI+1lXORNdI9FU0+GxnsjIzJSySHk+TZcInsrQ
rySx6+PxIOTYHwgR03kjqjLDfjj4wrmyb0QeJO07sYxs0sh5ArWLbO6UXvIyQpEh
iKSH+FbVZQycIHE0cYLxJ6YXbhoPPxDVQUbEuHPKEeZv+WjW7UPl17hSWCJ97J4m
tThn2QGdi5RkRoSgcwxKDJgXSalT8OqFvja3E9QrbfkV8SCFYxn9yN+2Vw8skSBT
wAzPGv2qMOXcPyXc8ptu0JPFxDGtKrYLQz0ejtCWnHc2MW6CG9GMVXGoZfo+UVGW
lMIfEx0ElXquqi+l+SJP+BBejwsqKkTEe3cZJGhIZhG4rCT5lWhzgDzpupV30mmh
8W9aJV13sfPX/DzhxdrTkFQixpoV7z4Kr5QkulWI82NhGLOWXKUqWkzs1scBr7xA
opN8wkEsote8DzsVs5CKeVxn5vL4f0dgvcQ9t2fxZc0Ue5Cv9tgNtq+bM1XWbpaA
EOMipPD6/1b0Xs+umMUaR8ED/Y0llzSWWZveO7XX62bs1t7JAmWEPhuXXR2FRoe0
oei3kEq746L7gjVmsJ7Q0ekzqT+sNLA+CzJSIgR/FtLeozm4K6F7ULV5QL/PgeVI
PDrmWIR2Q669HuWCiyRl59zFKqDKpvyaif9F/siC7/MVvRJTzpcgywK2Z9bxQbet
5xwVNblkR9nYhahb4RJh0S/wxq2OIUdQiD3i8o5ASlu7+xoYyjLlv/CnWeMcoXbG
kMlZMK/FadXNxbaYPa5y13lkLPAJMEMzQMKjIXF3E516MJscS08SR6NXKhBffpAO
AjtTjb0W1s477EU846d3gbxyk8YENBf8veo6OB0meak4R4N0KdIRCteov5twz0Fs
gCGJ3nqGXyJ6TS17DgyRuu577lncn7QgQ2v0bzo/LKzx8+2v6V+emwkVftf05NWy
ePZ7JkwjzJdc2ayIXq3ijQZNF8CzDpiTDhgn6P/8GLM2FjAabCwF0LQLLG5zQ+qd
CdJzS2bfdGRskkEkzXvwe+PXiYmECoIwBogIkc61nQML8roOi8n9HESyrTkQf9Xu
v+a/gwAX5TNPVzMSiKc+8Rk7NahmOQItItukIy+mPFZvIKPUE8lpv0My8T6ReXt1
V10ThmeK/xj7piUrqKaTkSI8rhV11yzq6M+yOOFz9yfc2sJMpsluY1Bbq1t9EY+A
K8BU+fGWh7jn064w0T8N1EWCbAAkvDFmorrzU0LTmxdeNZtOJfzzw/FWHjIpRKEU
sSgoua+FjDMGN42y2W7dC3dS0enFSJG9VDm4rnOwqtZMMb5O6DYhbGd4q6YUL8ST
QtVVYHHUdR90mktdRxYXEX8Rg4admSmxQSO0omDne5frVxmwHGUT/OWsS1q0znEH
kwG/5q2vN5g59IrzQ5YPyKuUjx0sOA2yJbCPgoP8wYaw4u9YMPvrkQQe8I3LJGbv
nHwj5c0UzP5BdVErORnAa7S7VrUOEZntr4XB7Rsy0FTWNsJO0q7H4St5s6oc90gS
YDjsz+scTXsDUuFBuIEywieL6GL3lszv5rZRh9KgQS0JSGzYj3sh3BMaOgtelP0U
nAdhfRo8PE9Ti8TTD4FiPJAeQkQzgI83BVbH2LgChCBx/v/vCKbln6v+YQ1HV3jk
eqzK0782/jZoyd8O09a0onB7jQH0IJKrgEpaOy1z82AF/lD1agov3Id3LUMUDvNR
2iPtWV9DSBx6FE0kzpDMAhl8JfcKeTCVlgUJrh24/+GWhEX0Dkco3Q+IBmuJnuVW
KYhvlQ41eU6dFAxuKZigrzsPo52JNcnMFTcDyrV581rQ24e4X+yPR94yFMoAL0gg
vXSNfbJXHOtJ+vwB0/09u1aYF+VuNXkYYih6UvhCGsedzxVzxwe6hzQ5MASwEFIB
vrMVhxrpxepN6S6gx9Q/WXK05I+q8BJi8x3Wkc1Uo9l4zhLPdD5+fAzwP9xTSbWA
rIwzAZ056/v0t/DVatHj7KqltNGgQIOL7oU6tYzwVOviu2jZrKCWAH6O74+bYrvW
r7tQWT3b4iWktTeGqRUbS8EshRFcsgzhrW8GyoVzgg/wZCFKGf6BX0JgIgD8rEF6
dw81kVc7ASNhJebjy9TH/cKnRqRB6uM9aCgxP5HgeQtXmvvEWK5TL7OhxnlBrCbk
+3uXVuzS05/Ib+AoQ9rwtLbkh9ysN7NHDkALBXKUJX7PkRIcEP7vrXBXoR+Iw2S1
rfEOFDJjzuoDsB3xJ/MBH/TdLVVnCGeJHWmgNpcFmFixQK+2jpmzUd4IwKE6OYtf
KGKXb7Y6oCVEiFoQp4Piw5brTgrXSBaSYlaNWg/ylef/LTgvBt/2K2O9opmngkVb
N5REA6roe6uUtbY+HaNdF727rUPu5/4OZpTZ3ZEbD0xVSzvxXbeB9wMYrmSiyxxz
9h/ahOdw5t+94+H99NOoCpI7JklpSlP1TdLsxmxV3vE1e/7uU0+Ziusf5NyPunD3
y6ryqj0W0do1TaxOoNCJHhzpUTZ3BTqNwJxFd2qKvVNymXEamANrKa6s8j02pzZB
/qfcUNX54AlMWJ9sp+02HYBStUuFdDZ8pgTcrxOO82khHoqNatPFAzTRNobBAVvo
oH8yZTtmWHpTv3If1qJ19WWfca8/KgPHCy7RiPsxSivRCnWCtEAxg/SCKxRvojfQ
7L9ocPfpRBT+a5fWI6dq8HgWLthYF/k4cA9bEui3DifSfoVhpDOtAPqf5BuhsfvJ
XgTOF7Sw08CmXcCH2ExNJ6CqZp+p/SeQHghq7fWs8U64OEaoSXbPMlhNyPoazBpC
KTRu53btyMn6D2R37JH3xDrmSinaWlBBENC3le77qPmNDTwCQvNdTY2q952jq3Za
WLH90XhpEhJ+Un+Lt55LthDcRHH8i3eX2UI7hBGP62M6YY1W/eUMK3owD3FrrbpL
W9LIXPEjzmwvhnxgRpoc1YEeyAqOKth0sATqPF19J+kdopGWmmXvZfa4zZ7KKYag
NhuuZ4JaBW8Ru/KS58+sdCerXGIcCoT+aWFAmMeQV8K1e5k7QBYA+A9yrJo2DyAF
vaBj8s+yiqwMOb8g9IEmrG4GUd6Z9SHbfgGdRybVj98NmuWNHRBkTkz0AA3zft0O
36yjcvvzLWdYf3nA2ROmzmNN4YtZDzaibNdbIvhP18X2owIldxhqjWa2uiupJVdQ
QmxHA+VVh7AfZLYkE8zjdnqsabFPf2YcQZqBUM0fBIkY48IRV3wKbYpxKi0Ah4L+
Hqwh9wqR28Xnl+FMNwMCrZLLVW/DaJ+LSJgJjhsqFCwd2bymCPqM32zlkDAS8ftL
V7+pYHCd1xtQ63z2FlJOYK5xxIMTF6sxHioO6e9AnAzpBxpTxa1Z/xm307SD8xHh
CoJCeoJ5bgmMd6P5hPC+EBsxG5zns+Ng+5Yj9yfKaPloxDVaet7BOnZZy1Ido8gD
RobONPscQE3IwNBjysReDHMEUmtHgd2j6hJveEDX56C48ftqb0FHDwMoDvecupQh
NF60+6XUZRB4/ZqBOiyMdCJrl2z+nQCuIfE+xbDHZSfpg8H6BiInrQJU2LG3PW4m
0JuGSsGT7r2ZjgOyTNR7WtuQ50qyBeYrNpuIhe4KzrE3tTtnBtzkF5ePriSLTSEC
N7RyWQ/hUclBVEX/JaN/Nm1TrD8yD61pC72c8A1GhSiaC9E+0bTF0sxuVKeomPmx
Zvasx29vr6nfk5F3X63JMaEw32+B0npnVz2atms5T5XVm+3RcBCnD+lmP6vj4k2+
P+z4pDAjb5VKP4XYT2FvGDNgMYkHa3RaFFssQNJZUECa8Q8g83pQnohy+XY1GTjR
sBMkVjo9NclxpTEtIJcsjJaqhPzWwfUOwLnpAp/eNDzqkvZX1xdzXnuhc3az74QM
WjpKakChzR2v7PSnwKNxEGVhq1a2sPe9x3uwQnxEMnpPzFv8SO0Yy77NWWgKtwrV
p0vOP06l18CHnuY7ok7V5c6MwP2zNan5q2bUMEXw/8EbNlnItUXRDLu6hGNgthoF
htGRSLtZV2oVPgi3XshNPGBxdVRkjD/Fwrmn+IgSvT3BmQM7oXTJbc6RIIBO96Bi
8JnOCQihKL3XYmIN1hK2uiYZNJGKdDdNYufCbGYV/tXC3RnLgG9oPcGicGBfuu6E
pKY8/eNIzkuLBdTMyalIF3KM+98juqtvAxRv2olTQGo08q2WRuhPXdrJvl+5Zoig
Yvh4CfMzcCDYlvDHRYr0l3XSe59sFY+k+iLHaED1gCRyS8yseUa6pXDwoD6VT28z
trs8wmFYhU9QDEt3manqE6Dbpz7WTBwRAxMwyiwikmiiouJbTHkAtPWijHQr9laZ
59CPkXbw0RKJoOpzUI1tS7vyTdRkMOsOfGYgtE5XqJM5pDFiaoPT0h9sE2hMRtYJ
OqsuxbhA55Nv4KwZCxsudIklb1oaKESwhP+IJZ8Ujc68KPLvTAl1K8lUSWvmBCrH
XYRlomoMZ2PCGMluYJ296kh9K4F1O+3o5W1XcZwL48Si9W0xHSLVpyGdC1ZWCoDc
WhoupHp4Wl5HUemXT5gqH46OcRi1rZB79uRZYIz5ed2ZhHJWPE1mOS0ZAsUC0p5J
3QuMbhn3CxDpdyk14ipQaikQ+Nzv5eRi0f9mbomCosYCClouIRp299q2QCXpoZao
+xk/WWCjfAerUIxr5FyTbpQfOj/TOqSgDk3Y7P+Ec09mnYPvSQeJTbYLfV6ihtHH
yZ3M/0dglXP6TRdZjNgjB9UF6yWce3NBY5vmYIv7OdExhcGqk2rno38xSaE1x69j
Ac8aqK27XjScIy+3wmeX0wQjIdsR8AYjnsNQb9GokpTioR2Pe1ityfM+wR9MISC3
C/PgmHfMggYHxfA6TL1lLMQ7Tzv7hQCdxA3n7utOz4FBFhFENyDdPDc1NopLx4Dr
NKw2uZJzTWsHPbLo3ta6/izNppt2vKZWX7vKFzqxxrsBCJvbfuAFFDzWTxnpLLrW
C/UvdCRyx6SNSrBIt81EpR69T/2q1w9F6tYJsZJ3Bs+jtheBgwTk3OlpupMoqRgh
osIbI5a7udPdvEwEfuDc24dM2dSMBaSSZVE0avr5JoI9kP16/7YRiyLDqxzMENAg
eYi4ugIuD8qHzxd52d63EkvJVOqeahfTJiHmreJ1tlRiyVLi23E1mPT7HbZbeDka
ZysA68+cSfRwD3Bxyd0xq6qS7D3NM/UnJ5cAcwugdCq8Ks+LcxX2PgR5wf5zJwJN
ZLUAOCZ2mOiGOtyTt5/+cxYEwhipMWnUYz8TqIkWPr26pTS1d06ztKG70R+OO7Ch
aCtHH0dqyNh7K6or+A2hDtC6jOyjpIU2Eb2io3jHZDqrlv+7fYdjBVEjnMR3YQk3
2yrtaYFwv0Prz4ZA+WNphsl/mBtnwzSAs/+8uZoyRsZwDstJ7Fnw2O+saPy5fBIg
lvozb6Q7skUTKIn4QB/jP5KSvs3hoOXCOJFP1EgO25OMY994oBTqDehrTpeFVVd3
VJGuwCFxxBk04RHIlCM0/veRbB08d8mfjmd4RHBOytJ4T46Wo4qUCTqQpbjNCyZa
zng+4cPoA2foe43X+FrODizI9UUufO56emMhY0OlrLrTQi/nmybxgQTlwh0JFUdu
gH1uMoXLrz4HZ6T8viaZD0IhdV31UtjSZdLmlDB+y6SlpK9mZ0U6mxI2LdvfDZXR
4A8PMfGitIU2540QN9B3C0cX5oeMWgU9XESviwH69I6XUGZEq14YaOC0pEyoBGES
AY36WG9sRfJLRy5T9LOZ/aODRw4k+Xmx65Q5g9IeNn9WB9LU+PoaYDupHvSmCgGd
7dgQzTi0F03PUHmD96LCCCGqUhQ06f4UPkv4QQdK59MpMk3OIKgJDAjZIcZ+tTqO
L3DwsxpyLf5VYvOANwYqAq7U0KdNNJCfD1HYkt9SVuP9YM2xjoSp6zAVzFfQCk0o
B5r7WIot5SmCgwGLEkBScET3e3NuECwKXjHJb2AfJUiwYHsW8lZLF/V1NVHZJIRh
PqVwBz/Hv2e0PZU/6qJjBkum3yBQQdN/xuHvERtZwq+/SDtGxWAE0A684MBY0r71
T+uoRorMxWCzFECU1Dn5UukJva5MGv79VbwRZrDeWk4tF8ZKHgS+kQ9DfhyR/+oD
o4v4xwrcLRPBcT4s78VhGXO3bqPZo3AfTXqCWOHJhwAmhyW9sPQNdyzAXqIlKu01
0wWqrOu0uAlbfFiVZqYQ5hFoYHRyFkHAzwXsbEd0GVFGRYzRPVr951klQmpUutB7
vWldZF/ki97LY3wzjT49EolVs/gilWeMeHLn1Zaw8XWTkMiT0BCtoBfbpGJMuKCS
C9dgemqbizTHFYmxo/YwETV0RalvES1WRjFShQFxsv/NaxzZh2WEg6XBASL2FVEl
ed5VVwYRDc2nLOMRVp22FF1lB33GGlhRCaXhVBdQXSWvgFUpTXD6dHbHL1VcDh1d
UVI2Ag5g/dbvSZho/TtjaA9LGZbjhtKhzkUrZyQq5svsv31L5A8mtGp9uShGoScj
btCBvGOil4iGt42spHDEcU+tyn1zk6cx3oeZqSZVzNLIpnmBPVkD3IVDkTSOoElO
FNMelsoIcAWokIcI85Qlo5xqINfj4+ryVlWGNNsWUSZsRyO3Q+D4V8x3pKOCoy3U
vu+jrBJQkP942VGOywqo/CmL88YqZpew+3T565cHJSQ6u7TfTqjSwnkAjAdG7y/k
+TklZfnJQ7pN1dO7Wa5Nc6EYGQt3jzjIJjugGgh1trGj/xRTJt4zXuBY8cClmOG+
fSeMynzWFt5Zr+rIOvJpZZ7Y3pJ6nHiWFyVq3EbbhICKL5Bx+Rldl4p1QzqphOmC
FuYhG4s+DLTmKZXA4Ef88Ho0B+nIFXtOvNPurCOTXju1hUYeoe4McoDs4KsQ/d5k
OEfrYGdtpX1rO4uLgA2k2MOv8s40gF10pvYdAOMV7J+bOHYtqBefSdSMA+EIHnk2
s28amWkSZ7aywCsvvkVz1q+JcuAOj3d/MXgbJrzYalk5GzHjUySz1GSjHWsZMMH9
Ik4ysUiIhcGdAcPMIiPmjvnvoqq6YGfVRAwYxNQBHXEfLEzy9HycPcK8iyMP+6yu
Y0XrpdQXN5VPSNtHyjL3ixDBAvTBgjHpvbRuxGT8dEa/glRytsPMAv4M0CvhP0CD
43Cy3O7sO5bQwgOda5B9t5Yk4JIOJTxzmNZB72IeNdHYLyn0h2AtElwGx9ZZBRHI
iwCIo0Xa0bDJpGMaUZ3cDssDUrAD1EwNkYophrjd8RNN60WvsDRIJ+5BPVZejHHX
wl3/3Wm8jF+huYpSUQH+aROAE1E4IokOm45vGRTIYe50Mot+CArViijseBSqY/tP
7I46aHmgcdaS9OXQV+/Mvcklye7KmZWShN86CcoxoICIX3SHnNA4cgLcID8DkTUJ
SCI6JaE93uR/Zby+xjoYgz8iyVDfi1+SHt5KBQ7gOaw2wc37jPG+uCbqSPGjj9ib
flS18lABFNq+XqDWuQPIA9rowFRJ15PJKz71hfslk2HuJ0v/EyJAcAHxRonDb8fB
VdFX7HlLijpaRikn6KepGhafgndPt+NzwGC+kSmZ7hjKJ/goXWJ1Gv1o0xDKjpyR
aFAQfSML6YWQLkaQ54owmHiWuhusZ3ZtPRpTtICIgmALHaPmWdtGO2P25avy3eP+
uVkAW/9wAMz7gbKk72ZdKOMffD9DSYA64NGUG1nUKThoY/JrRyOw4+4Qoc8WvyzG
an82QpJvJWNn7SMex32ab1cNQ9fD/VAiZnmXAUPxeSVX6p3Xa1xZWOIQW8NyAHcn
o5vw1a8516mrPfcKbhYDBpBWgEF2FcqNF89QmZ6HOz5ueTgiDj1z0Vyl7TeVG/rK
eAA+0Xy11lmVf8+mH3zGlWY2J6jUJ34IYYqOwpicg9nD1zAWPToWjoH+itR2YB8l
E6FRaHYyt4a+R6IrZt1sMrahQJSqAQs9fO3z46HEByI9mT4aZe+8oraJ7s5DECIO
r1hAX/tNDAfPW0DQOzjtGbr4UyCYrop7FwOjx+JZEIS2wyFb0NP3YnXLLxhSQX+b
PgPrLxRRzPEP3zBn7c2/yRPMeDT1FjkJb324OrvAaM/elwjXArsOX31fqj8TW59C
YZMujbmBQEyTFIVNy1XGuWBpaTreQwbE9103kzKqT+M42wYiYAz88L/s79epek9u
V5KxE2SgaK6Nobkv/Qs7ss7i9IWFaUjvUhjphaXUAzDzCO3UK2svfw9Wg7mAOvnH
+PNElQQZ8V5ODQiL6wVtiNvtEHNH2P+nqTm8mfDx3YndJT9RQf2gQAyf52jGdXfQ
AGKzlmlxwxk5WpcY0K6HrlvaBdE+2XhDbe8YcT1H9aE6+NblVWkMyykPjpdFmt0f
eIU2YxZw+KyB3KITIoE8N7oqwoSyIfL0vfzUVNs3oMQN/77VWljFvVwJMC/YlCjF
xxdUW1kK2Y+wuvONPYdXNsv4irnVDOlXYOQQ5XmQ+wxvHbgbNjx96I0i3Y0JieNq
35U2PjCMId9LYOzgSGKz8JYAu4ljDhfwqdZBrM69DGquYAaS+/ypuML7uiiTXolo
eDTys9my98Y3D/KHw9hp8npjCZMeMTic6mN5TpZkEtWnHR0EMCU3+bBeLM3CpEIJ
qj97by7PHobK5chAtEqR1zjrYX5mmMsQPcgBIe+48Smg/NqMVZATO+ExSBWdpGmK
lgB10YdNWXF9V0iJbRwf9pmL+NSfvoAhfG/l/FOavGkjQKeozA9yiNZhU7YZrL4X
iqQDzEqJsNNsOGHsAXVTmYpqnbLpMucp1VsQu5qzAG6IcfKjcmPCGgNh7RUFXGRs
BAAOMC9QSxSl/JH/eC8n7oKc2oD6KOw4g2iATdMWCq/h4qpIh0K5Bx3dYmOT33lA
KPblMOKVWcAj3cB7B6YdIWvBrAwiFG67/kKsH0jK9kYBGq7u2CPGMg4XHM0ETTxW
xaeRI24ZL+RbjLC+ar9WZKYZL8ZLvDY8ZbeRB6swxyRes+b3lc4VkY+jHv8PVeN1
LrmLmXu42dGTiZkCBA4ilTz/3C0wg/73kLDvGfiLG4uUfkc2o7Mi5d2C8KophMmK
obo63XWSiqQbB9L8A+5XI9DHYouHMN94Ex452E6gQeDQjvoPVNoutWojKP0P+JYg
NPMkmF9sxfx/etU9JltY4FiKfOeSdJaQc/+ODBA6l4IwbpQQzt7nUoNBjUo5rLAn
zxuhFLTdzY258SumyZSzLBvsL1i8PfplIjzKHiiNmdmvS3bG2KOQHkmJRwan5sWZ
raQpF1onbEMtAtxaZpUjgBTzGQdBI2I8CWZ2BbVr6HLVjuP67dJLlN2mni3Ms+MV
Icpa1Sd4kQVohrQVc0YrbTtpRv+VKWtDwfQpHWcbfJfsZc7oa8mZlp6JdLiU1xo6
0Avhmdq8H6Ya0KYnjf/6BznkXVuvr8TmiEo78N1jX40hQiHD/OzBNRlD9d1oHah2
oF9FRsufS1jcpO1GhvamHIfdM70URW87HNUgRuiEvO96CHbMr2Zm6Tyss40ET+oe
HuZ7Qc48DXCTTC9ACoC9OtA5GIntXLbowPfCLGzvqu0lj0uZgttMa+n3+mgVk3/y
DM8hzfp/E11cZJqVOT0ZohOD+uwkbV5jXQgwMNp3PqYmJEzk/nI+5XduKqwqN/EA
Xua7YsjrPDMkGhPeYuK+xooCOXxnxQFd2aYTHR1ZA/a61YVLKl8N0Q4+xL0eYroo
eW/XHHGOox0zyrEt4S+gF7dIeWmlaQg+bwv2S9JkaMbLQbo8NlkpEcNXoaU6RotC
ymTSRKrvkv9H5yoHneF89st89t2c1giTtRI/8YZTukxFpWkccqvIfCQfosgE0RoM
oM8d787q1YnwWPGqSHQVgRIX6LGxSg5ZZMmSNCfZzwTq4TovC39Zk9Mv6VSJ/KdT
9KJGJrVnzZS2mzO74rukVhtz8Wz2k/ln3/q8OtPfHpt5Kh4lxzhfEUbEFA8rU8FS
7TvdGgFXHI/OULjzVR1D2xZO6dvNydh1l2nKj+GGvMmu/fteHdQQx02hD01YgEfG
EeFSOeKRwOwQM+5xGtIfSRkXs1/DsrekHhssjT+Apmn/jIR+I8HsnV8VjJtYuQX3
CHaJKk1DWIcDeiFlH92WdnbFW4HETxNanbACgCOGDRfrIxc3uc6mM+y0Hm+WXpqq
V+/q/q4vzaV/+akLc9h4xlrS3dTL1iJkCKTAKQc25MHoScrLpzKz4n2M46Pemb3+
qhK3znQJnq8E34i4QVthiPtxp3GgcJH3YMHojYL06s0ELmCbTFSiQmJ49hfBe1Y9
ayax8TzAA/rovk2ebZPwqFSNKLbDHPaIlWY2QtJfoYlvv53AO3P8jWZeaal3RTFt
7M54OStyohSZYpTEfw/+5dVB4y0SCgVgyRR/Nx0c+0rDH4CwBZqVsEMaZxPozo9Q
hS7RCkR77ZLuXuctDwn9RmK7h7FZ5p13ang4eLtf2njAuvVHJI5EUodxFnkh/rby
yxVzy5w4uBK1t0LlrJncL1hb6L9WcRPniRLxPIPukUIxk1EmD1isb5pQeFB0j+50
v7ETX+vpOKMKg1nns2PyuRa1W/X9cBjpb+Q+Ek73hIewfWIWRXCvmVYNZFHnlbvx
NIxkUKE4TwoBEZ8cUvuM5a1pl9b+zi8HCnn9Yl7ynUNivKA84bDKx9CbYkgWEH9J
eqi7UZ59YNn/b7or4N9S6u6oe169ypiOVB+ZaWuu3GjUEC02309jxoxHGD21O+v7
lNU3ZP5QGd6eJt8WyuuWPwQO4s8XpigvxjB7oeCVEBuGshlyq1tUJ84USFaV3wz8
TI4Fw4cav2lcxJkF5DPFphV1wMsBsYxxLoL31HgIbzXSCl0mdeMg8vA0u2tHEjXS
wlZa0mp7OaXoXpNOYsUhtXISD6YZfY4p0QJQEjkRvDPmKP52fqVxWZqNRUAIBBrv
H8iwRY5YXW4WE7o6pn5+UevNlk2575jHERjyg67sMGN3E2ymv2JLsqEHapqH21k5
hJQ3wSNbUmJjOSWDMX0uovOBmUbaIZyVTMkyPtqPxJRw3hcHHMete2RgBgsGT0Z6
wHZqedaUty6eUHGWwpOmZxRIAjwgWtYERiOce28mL7k0dXU1Di4w0mSeuL9mJA1S
E4byJoszdh6/bSskaGf0UWetpINW6jlLVUTseRRjwogrm32lQfmYqZRk10iF79/+
r/KVxrJUi1NYrnzgm+VwtD/h8XuFe+99cgovGFb8GIgDQFMaFaf3GzoZ059aWcC5
ZwDKRtfZmbDSDRQEHr4QF0OFvk9fYokPfbXKxeQgwTnv4ZgD2w3kNEunVfni+Vdj
sf4sb2WhmXhZt6Hn0XLRFMhs8++sbYngQZYW6g41CaFTdYV1JEg9OKwH3BPTWLT7
wIVifkagvUzMN6fbOK6AuVT5zl850DGwFofGLQgKOepUiRRk6SBR11bpDBf/ALFF
W2iUSrLcmJFudMccJc39Tsnyg7YbnQHMjafXZ1I9Nz8tPiUWDCJ30x4y6r9jk3Yi
0gXxCly7h5txC3/ORDvzYOQPK5EftrXjmz2FLBOEKvIOP0rGwbo9E38CsqWzztpH
Sf2SBJuHgcXkXKT3w6j6UPhpHl/ISUbpmSIKYiCGEUsrrfXntJ2u3lxlDzWhxVmY
WQS+sS8ZrshSLiaZfR4rW0DrNI/Uj40SebLWai0OfXQOrvderwfVVY6bv8ZeDD1D
KKHyib1/BjccAbes9yPr6vj5bXB5zVFgJhhcnBv5w+2PxQG3mUdCrgxdllo1qnak
Tzoczs6/YZfFawRKNqIVvXCNztEETyrBR6NASGu6qw5KZM+OmIBJLO2acG7VX35F
F4W7O+rObrg54KQu50qpmwUNJBmKOXIz5sRM1b1S0d/mhv+G0Lpnh46g0UP4ttSj
ZEIgt79Mc+I92QqgYjtZFsr5RdTUfhneoQecvTF13yyiOSUQea+kHRNxavquXKAC
uW8XM7uM/10uVOI7SD9CAfDqGB4SChJaiGpDpi9zFfnM9aMugZbclp1f2afNS/Hg
JbwwgQVknImdgXkh3dqGjU6SQOBYbcUrPJXSVjhxWNsffezfjJM/gZtfHeKU++lP
6r410PA/vJsoVFvbmwMwj95lcHA5adv3SejNBuflHh3WWiwZBc0xB8Bo+hQnIZM8
UDOFBr4vmP/SWkhJKniHOwErqnN0eCGWOW5WxvgS6EVjBLgagsyGfX1r19g+8Ath
V4V7pPgRub4QoqR5AeSZpohMKeUjpTxOCBviGclBxh9ow9yrAbY9c9b2oZkEzIuM
scYrA1lxzWl96+qIXePkdxdETI8410FcHqP0B8wZyF/VRX/vM6izcH56c4NnJkck
zOOteVHuonf9KcNs5jMptssCmF4g3KMMDYTPRZ1lZJtu6VEswyuIbxXVSwbreYxW
HpoZYi6Xsvr5CWvrHYvZ+d3tKZeph4ZhmjkntIAWb2cjlserqDVQLtsAmyRSQ2Kx
mi+c2thoiyfK1iaM6dWxbVlfXDYo1j+13whPqT9Hogq8JhDLGnSeYl7Mn5CYZdgb
jlJHndyUjDK/66hGz5PeL2ObW4v6+KxmAP386DvAloTE5ct1ZQ6qFMfqoL2zfy1G
+8muhU15Egr6gvq8LqFaojJ9bmqUooMUeWKG/AGn2NUGjF2zrg23ou3SFnzI1/4G
p9/ljJFg6JDj5HYordHPQSEOW19ubmF7/d7hUj9kAAvo/4k1zph7ivmz+K8QwZ1k
sR2nmmhYT9dEj302RzvdHiZo3N7VdwgWDXTQqvMCyX22yqLX87izqklXneSj+jr3
HPKNPWssFi2eiJgtb4xjGPiYfWDvOMm4gGknmKiVcwAoLQzk98kHpZCOjAO5lzZD
UfejW6Kl2SpzzSyTO6dPy1Cnq8EXGWI3c2TzMM8jJg7rhgVl/LfBqZnGLq8eYc03
F5w80MQlBmn+TZW5d0glkF5MNrfMjx7nfUefXkdGs6C5FbKpaQYv7XG118WbXoLo
+PbgSWMQbR3MHnzHCrYPfwjOV3I3iyLqpHTLcuKH17wym5oFDKZOAGRKhOPY2N82
w07I+szrzAGiGVq+LMXnWesO8sfvHlMqtKsOQlhN/vXB8KO3268YpKUhJQDRHA1e
euRW73aMKnTRYAuj9O4+tYiORzkd+V9nLrfoRt0qeiPbqinEdZjikusxmgEOCMUY
I3OAECTbkgCiKwtYwxC7Cg0z9Vg9MvQocAMahM5ndYJykMjzYqiKWGnmlzB6MB6N
JnqM168lTST8wZ8UYTfKruPZZaSsO6TVvzPYEq4jkQiuibUSUqY77zGu2BLNDgb8
aeF6S0kSsGcmQDWTsXE5L80n4Oyg4IY+8jY0gcPLvx5prxUOiOtpNKqN6sMogfB5
aatpQkFYB+EgRpHUktDjIAgStpLpRQa04rwW8twAKIVjAjbwJi6SiLk7KcCr4tw/
oeXBirp6vr0pwYk8VYbj/U5Rl54yuxw8T5oH5KK2eU+Nra6MNjD+lEVHauqcrVRl
1mAKHI+lrBsiabk9h/AwCX89g2vSgaYL61r3poFRAg16okbaJQTiDWr80iwD+099
QgbqE3GDeVP0LWCBRxyqQm+bJFIWRkK7y8QesWNu614dDqGOu+t+BYHnpEyNk8Bk
wDZh5tqgD/5x8FmW1JB9x8R0KUZBJ+ss+L+i9Cyrv8r02r2HVjeQYCwU1HN10AGo
ha47csyCItAty84PEJdRFIAPvXhTpm41bIIBCtqjznhPz+NisNG9TCYo35/8T1vA
qZq0G8St53b66u6gKeXyjBPGQ5l9GdWpz2baOA0ebk1p96B4ng+i2pGqHJxVYW2g
4JvbJlTUogdyrZuzFVcuh3S7lpSbDh/pmmjjdmkQC72e9/FOPuG2QxFs5LmEKwhq
Izwc1I4fzilFFrhK7zK2buriWwkrejA7eTBySp8iyL8At2/exmvP6s3wx9DEmEg4
vB3+UQ1YZnFfdnDp9NQQJe7M4WrzUdT/sAVoFwyiPwrXGJb9NJB2AkMgrqnVoj2A
18/00oI3z2qdLY+SE7Ie/ql6p6XTlsf2NgwPsXSbVb5H4G9So7ZXoAY2YRNjNB4q
EoVJQ2Uck+7aXIhj6gxb87vClgAv2iG2LMWg8QYz9Gb58WsDEcsGD8zR7qn8Mkkv
6Qxth15/D8fG9f1MODZwNvZToGLw4DhtfXpaH3K73NrINJfPRFn7P3PoC3HZehsh
XHxNIUlW2jW7ccwdD7py/lQDFgB3Tn9QW1aQE3MALhlyZzbP1HOuweoKrJm1StWg
3+9jfDO256WG7rbYmXrprj6oki6cb1G+HaHTTbr+CxQ9136ugfIHKYdX70cCa5lI
7/jBsCN3MA0Jg06Or6fhgsdgMdrPxW3zguKSwZfHrli26w2xJipWLFL7B7+V2zzD
ZpGQwCS6xWBywPzELEMRCyRN2XuvpH4gkVBeLZF3UQEAPIe50eUZr/4MBW9SR2dR
Supg4/1vJQj75VRSCFqT7nQ6uuG1Ad886EsRAyb7hWr36/CJUcB41Akt9j9sQiv4
vsvSDBIm4G5CSQnS+y7SFz0vCizFcFbXeYB70bbBtsUgWzX9tTT6vqfjRngZja0z
YY/ktIXeulBV0cODKOA8rVziyb4aPoeIF+t9fn8/il6bE5CbVDBZUYPU/+3HKNiV
AmvCyMLUEuzsM0UF/iGCfZxVdvPWq62X5cJdFvlot+FIF4UWRxIDdDxxp2XBnA0t
3EoZoqGLr1i9tFddhzqVLZbDwoPnY/ieh9f3K9In5Edq22G1GtfGWEKjrVkiELD8
kkBYrJqHS8CovjSNeEFsyNRhE9+bBLHTDd/Iy3ICOgEkktRlaS5KgEvZEOpB+I4Y
4JCjBY3dWDZZQ8tEatrXmdS82cOphGH4dZ8MaWld8srIZbg5OGtrDW2vhPc0qarY
ah7fZ6eBa4f8+JYXQHKhnnMENHp7UAhn6FQE/k7sstY5wDFR5YBlafGGcF+n8UKq
1JSny+IEJg1n28ndP8bXRXNhRRDm4Eu9VAiJekCJ4PZlwgGDl+GjyVvh6IERcLjU
V58gYqdsBRXK1JZ+5is2I2Jp4xfavAEA5Lo/6T9ID3BOBcmVmbKIrZyPbHBS/KPo
zqqHBbke/K1Ujwdyakem7xIEWGrr1DYM4unrx/ZwvmuXtIrKPZ2es4h7ax/q2KHa
MOUYpxLgBQGKtSCrk6SPsnO0MyYu3swr7jVFe9ZQZDEJ9p19qUVhLpuQVXmOUws9
VhQEl8VAvnII/kU/8s/qvT5yQvCBZTK5PTSYyIKq/Jdlu5lSooI0VR69lF1Lfh+8
F19TO6QVKrt95/I7+6EwrIw7dbsoFyWBVwYjAiOcebRm+BMEY4E4NJK7zzDC8IHL
EyPLn29yWP+ErH1fSPfRJO5Sl2hQo7aB/rYwC6h7Ab/xzpNe4cu1is9WFNsEfhjQ
FbmYVmoIKAz7zwZIClMcQ3oS7h0le4+wKpgRupBshh/qzv8hLQt1nuJpYpB7rkSZ
0huaQxnrx7wwjZeeWHyycdSDVLzeek2eaS0rUz6WlEpQTz1drCPZ+slIjro/PqP2
zyHxJOmd6n000OQf97tXOc9cBeAGyD0DMT6h4Kz13PfU8yHm1qT2dJbtOx/v9zzY
+iTzJRSFlri9qkIO4AaQs2ni92fsIvAn11hpWb8K26Z2eevJXSbL0VKsHJUuskdG
pnyW4gMbwNOdo7mNgNm7VSnNlBr2YZN1DYO0/B3bFBS2hHz84FZQ+vOPQ09nViw4
CVZuo/MpUyZlHFjP8k6HZUelcrYXkPo5/WWUudp4ot5/SDNiDUa96rYTe8yF12n2
hCFzHKLQ2dWX19kw09QnxQdyVNjk/cotcZmDVcHiaSCDgqfA+RzdmUTHO8q1Fdbk
1qODPiupBg91Vda6eRofQxtp2z/57FbDiyMhKCJx1qSTzIbi8Odv7mdqmzsjd1gQ
QhHV8o+3xLd52HvBCBrD/qDdqqv7HUouPVs4wecAl+cZVha/S6k0LAGtv9kHkiSc
hWxvZCrZIhRuqoKBEO7/s3YT3VHXtFS2FhRY+7mx5KmSLRsX+1aZAI2p2YhLaY+O
tGqvzmktnVRF6kb2unfuSjb3K8uR9aX0J8nzg7MLKf86jVYopUy2rAEO3XVtw4za
tBAZA9Rxckl+qxs4bCnnQuZK7/TW5GegkOx2qP2YEoCzQfJB8ZWPBwVnyKFr5/rO
R84g2Wtd+7Ok3yGTUx/6B+5u5K0d4keQsr68JIHYxCR2uVdmWiGhR3Vf9DKb+BCv
C1jhJuJzbn7MfghuMVQWvDcipwiNuLuOCMQ9sEhXOHjS0Qsf0XER+4GYpQvNPsCj
tTyLo9mKdKSL/Yo0hbIPy6UBCRYcN91tijYQiqE3bDWLvLF7k22ObjuiqoPROIsR
0SYCH7GBnBXCUpt8jp4VhYXnYOedLoasPv5qYSHepb3N5PQpPjcDmvXqM6zhx3jL
Ja9yF66pDtU2pORnTZHtPEGQKiaAZ8HG/w8YjUcn35BUCVg97ZzbwNygLGpapZVG
uAnyJSPJfw2N2i5v+CCO6euvM1oj+IGbZgBNqkBa98gLJRs3f4jvNHkKX4QVZrqX
4mHZFYSixBHEZmRvDROoB+CnhVxnntjxudENreb/IvkUJ57b6uC4StgybZCrmRnc
DfmEaLNVjGamiRLIgDCpL5cz3riq/NunUQmOsbr1fHwUTjl0KkPootE/NXFfQx4K
uy/EsMIYC+x39Rub7hpKnyMRUn8yULjK1Dzquh7hO3ZXkhHlTDWuUEe/lmCR+Gzi
AdP37B9deL2iHk4vI1vmkGBQctZ9Ae/G+Nj6BPVJE+Vdkg2hHlDg8xXRMhVr+5fC
YbMrbAJlj5GxsuiFxLWAqPSUd+JbxnxH7+GEU13d+DvzIUSFm3iiKj04OCjYaR27
GSX6lL0NhJU3JKhl+5ZVQ+DWZbXcQQZ4jwmtE9XnGARJPoL3rJKsgEoXOSfe/AtN
cBYMmDkiqsXZTLDUTcjE3ODl4eK8DOR9A17J3D8QLap/85ZDnJuf7aGjS+bZYeA4
kRJAyYAq34TydQVr/4HAVpXCSY7AArMvKldNZ11rZRUx+TVRgV4tE/xBTT/gyTcL
L83A77rrE4KSUhtEoZnyxgD+8SjqziPZkF5LdKq+A43oWKpF24+pBilNHB4gk95B
OTR2S64hPChIMWVHrArlQAcX/uzaVy9qc0E2Y2/zinZL3NFs6YcJb/j3PyGIujNw
Bqd31KLWqN9l7ZGw04+34BXtzRgdFXPBLc1SSz2m95UiJp4ooPOZfm2dqGsOmHSH
Lig6DDZNwe6uQ4H27St9Un2NNIMLi5JCtXf0mzi+N/2AJmA9nXKT5zqZEWc6xPZO
o1T5xG8/wTMIQFjmvCMa6tmokZs2gJdTPo3LZjiS+nspluHeNLwz61IXuBZLDsGq
ofBNT74JQHtbZsvj+xoUBC7qw6TA7f3pAAwW5nHjMxhUhWyhRiIVYOqbIoraAN+h
jRLtYfn9hFy3BZR0+/XYVZNimBZ6Yu28prtNTdAr9m9bcRzIzhI+TOI3G97eiQKv
nPGIOqKyDlYienlP7zMfny3iIBBegEfsEjRudcHsiFezKoqAKkNJjCZ/Riq8+fGN
wCWH4E5ojvQSYWd8E4lrZpRkOsReotUz708gE2lWK6XBcmIIXqez75FXI2l7vXOC
oRiUEiOzjAJkQfUUI+fu7dQRSLZ9ImYWu6arQ8I2Hj5YL6JHopqbwJDylfmFsRyo
ESJxyXcXCPmjpUqjeu77XGxx3Y8JyP7jBAcwqWK3T2CIwjHogLEbjRySDSzYUhOV
w7FhdiAac60UkZctPC9oJEnkYIPsMyMM/JCXPO1UwrrP7lYOCZoiFCBz6eXRFCvH
spqpKBrQpxSk1Qh4lrbvEcVuCs60VUkYgqSjh1m3hL8y8iDYlX0YUF0MnXNWpQub
lH3RUKHBHQHDbOHmdIOhMFtNxRHh/PLNWyplLFQa19TH9iSBlmME4FgQ7EjzrkRn
T6Q3M8NpCI0kOTVe5HBy1j4J4rIm8pg46ryCwWH97FErpii2gQ/6SOb2nt4REaij
/fEUaWKswxgbuZES6YfW5eS84EJg5sz47trABfsercIQzJhU5G+nxVwMXoQSLt8J
QEcG9M2GNvrXohjCyVuWYloq3ookNTyghTAxJXPhAb04kY9vPJ5RSH5QcOIS1jBP
qKHRnANX5bqlwnkW/AzGMHQyhc99dq08E+H9ImTqrgLiYOHeslF0jh86taxNkjnw
SQupW2VgwiLdd+CM16/OtfJAMmISH3kklRf6qC6nMSx8J8spfE3BLZZPe5FgBbP3
aOomZKrSR/+Y+21Qnuo/YHesBTa4ACG+BSDGJdkpKmF73O2Tn6TPIXWZ+zi+UosL
Y9vzheO7rtwx47bpfHP/61BvUpE6uxez9NF+OkOpOOxG91yHd2BtFjiWw2BLcLzw
dNrH6GdDuYspBBlFOQvutwwb7gM/13UNxpHT4D9krXo3AVccSVau7jUh9fwVKLwW
MQVumRFRwWpE8Y5XXztKufPim3HfsizuhWoBzIXHbVsM7ZJEHYDqQKIyuJ9MwJAe
OP3VSDBBQ5/JTaM+DujAOdX7JF82AxnhUJVYG1ZkKUhwCitvaz83NXK9BIbaxOcx
UiS5v1kMz5eJIbY+bpvlf0qHOZwTMsFTiecZ7Prip+I5TK+KVY9UEWMcpv6uSClR
wIf0RUL51d3ZjSE8JfTv794IGZ5TZHaqLmllXb1kqMZ5f3EttLVjGrrwV+48PZdu
m7K3O93N3XCGG5iA13dWpHkFFWcqx8wR6zm53LGrsv2vsmURuKl9t+P1LwD9iQHv
yeihpeO+lp5Jtir41S4nvd/uMC+8Ic0c5FNRGsuib108q0PlPnSuSNxgnww1rliO
29fliBIvvUxxG8q1fV1DITpmjJEzgxN6TrWr1u6/4eHLpwqy47V9ZhUktPqr1qcF
gknDrXeR3VgxytnyH8pCQvKIuO1fnGbfswiNJgzt27uWG8rlrWSgKazVA59d1I+l
E9EWYYpSFe6HWqnt4unspdvhEFxuoexA2JxuuYlwDc9YaddMEiYJMi1/konJtOQJ
3y1oyFjANRPIgj0L2JbWatVLDCk5s9UKW4FERoL13H0a15OZ+eHvoCvD+B9GcKlM
4Nc4UzUzbAP5cJdIkg3meGlNyfmoULiRMxL1pkegadvDrPb5BeGbbBex26z662Vt
pH6dFVGEO+Nj/imT8cV/emD9+OuqqKbu9/6Dh75zunDvOvfXnn5Zb2/AfLC9t67p
ewMWO+tVsShH6gXrtP8WsJgWi4TyUE4onD2KJ/XeKlAJvbMUVnFsg2PUdwgMlCDm
0cEhiRoUkjvMC9GTcnehrrpjBr8FynUiFn2Oz/hfNIY7Ho8fMr5wbm7REEx+MPKj
AI9JjX5UpLRREW0gxvyS+A4RghFgQztsRcnTr1WKSEsR0rz8zD5NBYtpWP+a2r/m
84KeGgqv5vMyHYs2AAIaQlMAMgHU+U2pBAswFOcto2fwUAPdU+0OWN8bDFA03/8o
4MLw+2qoM6OjNSVNOQx8WzGaNUO07jPR4zF3V+Y/ZaLNvK1tn+oQmmiISd25g7fS
MTVXlcpvhwXG7agYlusQoFDGKU1G0CIE6EHAvq7olYv3kiap9qcKAk+x8AHk29lO
HndIDqTtF/m0PqkkeTCqYip8yUvHz/MUrRoJqhK1jFv+rE8fZBgQB+sSMVLstOue
IRQqZWsONhxLkQr8gHA+L0sltv6o3UITi8y91dtxj6GOVgtHGN/4Cm1Av1En7BV9
PfeaPq26Biicbm2Iq3pJLrqxOV2UqCbiUpRa9VYw5ZzAbHbowUzQMYxnICUOsxDk
DIQTAuGySslqFzOddcGe91JPOG50SMsajm2Vnin2Vkf0OJZ0Fxv9HxzdLusFX9mp
k50C04zgm8kuSZx+1YGiPR3uOiN7a70VENllXEsG0JMmVa75e514OXK8tQfrkYmO
OIGYxwnpxSQG7/p1msfLfjjDXScS75tGaVIALxQqXDZ5PnuGqlQcGoyFzSraOEyd
Or1YGrbP8Rcz3qxJerPepBd9rl59q9415CAQjYxq1HQHennKF8NieQf5LCEQhlAD
aE8FNtB1Cr/KkW8T116nt6kYNV8S6W8S1F+uxo6KrImeltAIGj8yjzriGYF9OGHb
P9YlKnvpj71Qc9eEmmYQPo4hMAkBrD4t/Z+T9opy00uBRWLJ7j35v/gdTJl/2v8B
SzuWeZqNTO2KGfZhxITkAbh8EHP+jYKqqJaTfPvO6I5CDV2CN0rOPz9RKGCPalXZ
s9pYeUyRhKkTYS9tJIG71JsRrE14pTYZf44raZOc+opb4u18xoumF97B6+ll3Nvv
jofxvWsp1wZjmf4MzRggPHAyRQpAZhD3rL3SGSx18HXtFKLEEhre+deObXSyQBHs
UOayrpVPhR9q+n7QPyG3lkNLZXsjejrePpBt8Ux9xouZ4xfiui5+DVcnB+6s0CVe
u6k3zAWvSULerncVDJKM6NfxjOXtRkyu/kFx74/Sd9ZCqONE53IJKpqmy3FUbPx2
StES9i0lQjQ5DixSsdZQJcFzzTQRuy66C3RPqeQa+mWKDmguH7s1Untr2V99CyTj
sIH+VtfS/WmKnLIXFlLlMMSp4/CC87MyVGy0v6gTDQI3SdMtzU0Y6wjjYSTK69Lj
8Nf1AuF7xIGKDhB0aSnRyjTtk/JktjGbRngWN2Xlb54oG8QedNQb5VG/0vEmBeuY
8Z9eCbq0EhRP1bIJ54fSRuv25/PiFGOHyX58kLpqFuzSWE/zHTc69fegCis8gMI1
ZW2yQdT8gopcHNaQ9Yo8+Pp5eSmmVGp1TMknXMseGIP1jA+5m+iMs5KR8GLLrAYc
ZWgupOK+OTVL3E0eeYjW6DrurjQGhFM8Xu5VitzqZPv1jNyLg1E/P2tWbcGz317x
l0ykDckt0ehR85fsS+f24ON4ggnC0H52YBYSB+/ULU/Xmtk7asAvuShY/TSXBlmF
P9fftck1QPjul+UONyQWwlgkpZ5rv8wTL/ExEwSb4d8qVljpYk/rkD+qR1jWppqn
e/Za341VrFjLRmT7S26VE820Idk0MD+VT0T8ge2kers/oje4R6PBr2PJqCqUTDho
DlbgD8MtL3mRjUtYrHPHU+b6nWH98KrycLuOmjU8ctsq4R4GDxddY4bTSnVbgq9I
dB5QZew1yhJu0qbyKiU0NtwqxGSfeyOLqRSFgDOqKp2DR5gC9CADYo6ax9w1thvL
7xihQ5XbRb+BiPabYia7Skmkg6sDiDTZplihD/89U3/JDu1hOvh/tQ8bbIzEKZup
ZadFMuL6T0YGcJRzE832wnpt4BxwApsyRGEwhQ+iVYS6Hks/uhZWgl7Wn+UxXRQ4
sYXYa4KVXVbI2Ldl85hwDpsieSB59F7IpxAgFZDitKsEQkDa2gOBLMCUMmCTIwHQ
1qGnEuV7oipOIBTFUJlUdTzWx8Hym2Ub1/XHVjhjpX89K+aB60zEKYPZjBgG3zMy
fjE6fXYIeZfsUZS52AxvG/zWYAftouD7h/LLscPy07KUf4XvzouGB+ZEyKoBAwGJ
+1CI75r1N10GIzkpaTazCOGL6f6/YIbViDTNedza2WEIzAa9smu+1RehaA/KtmvQ
3Vdfze/KfV3l2qI/VJyTrnyuyfHWYspzfdvGUjR05v4tydze1BXF7xXXMbniNzFY
sHc/3ZlKtJjsVVxO2ATMvs9t1RAVw36HzEDHO6VwX9BCSECX1XHvtEhDXP5ARyBN
ASLsjSVdpWzzwdqVObQYyspcB0m3avz4ZbXKnCgIT67WjxMueEoUTJ9qqCI8Gja1
ga19DjeqVU+YE1V1xKh+Xxb7+I+oKF3K3xU9+0LSFEAPhGw/kjpq4Jr1dFdd+Ft3
C9uxdCJOAj0FkFS2j0gZ2erLyz9rIM36GvYA6kjSU1DX3SyQwSTMXF2NWeh3TdiT
YGn33X199mMCIpbCVyPLzan0AvI3KUVHFFgF9BpBE03DIaSJDlDYcrNnZhe9iSl/
KYaOo7H0FBbeReGW0+g/kJ/c79y0KFL0BVSU/X83U6VNcrkbweCtdDzxia1TDuE9
9ne4tHNEfC9cwUbXl835zxMEKu4tvPO8pN7blnfSkvj3zgurgjymZ04eglNi5Kyn
ecU4CMYlD7t+Sx1g+IfbO2N/wN5lwuJZDIQ85gNKy2nFasMdjIzou0E8Spk6etaH
FIPzLz79KnXr2jQ6WjkYV2M2q1mtZaK33pHzPVkSOwk9PxpkaGnrbX0KwOOMyygI
8CEjMOGMbNxCMFt8TOT5JoLPLMw1L8u/IKb2vLjXsjKGxBklEpKo3qTIioqZx+lK
UqZ8FnDIN1XsaRkCSul1UxQt75EVq0B2i7X5+T7/uSJ0KIZWjt77ST2unGTUmoSO
Voqz+6JDYprKOhpbP+izfsNmf4fr9eQp50CCvI//pVtgsLD2DJRPGvS87A3wougZ
b2QaSSHf5awxIDJ8zrSAA9Rvq5vIYzam4ChltT60b5ygkMrJRMn7u3VAFbymJtif
1P0yVcNFlSCdgbHZDTTjo8a7EHx6/sOZCb4s/EdQ34Q7qDmV+M1ONnNzUgvGLKEx
q7Mn6PJlEQHJkgUbbiLMGac3v9TleE5PFR6MQyB9qAACGuHFORyqNXK9ewoLMjwY
69tA6E/ftYr8dDFYLj2RmfFger6GsI7Id9OQIT/LX7D62IEp6acjG/0IrUqU9/WY
DAY2/9sjBNl5XDeCkr5MXrNnR9y/NwawG0WkEUU2O/lpd/1JOKC2f2GDO855m3Er
Hq+Yeac/A8ZLXdJImkXNH/KdXgdKjIJBaXp1ZdkBfCcuhN57ivC3a1DA8jGIN29u
IqKqgiVLkvggPLbof6i9JbXrTCEl0nfEekeozUniDegiblgKqz5pymXezK6QeXVt
dPeKQp8xH5MCXnKxO3hbUReig6Q3iGqxUTpPw7lEKwaR4HY2ksbfkMyYncxejLVk
7LPpIAZV9lue99MRVXcwLRMJjyfkmyaNHMVEXSUjqb5fpcmMeop5O8lywpXhJamW
MXxoxo9p7hF3j7mniluNbewENazMjJRDQtZJ8GR/HauczlxhoYoqpljWtaSHQZI/
EyuEwR8vNqvZLLzIsPYx6bEctXDpYK12z1VJEsXdBmYh1r1EUjJDflil9Gid+dAa
VBPhLgJppPMcHdM1TdTSBFN8sif9J6rZc+iablsUq/nrUM0YJXGD+x2C8FtbSfV6
s9RGjv7STHbw3ZE3Jr73VcsjkvTz42YELQ/ffI0e7vyy5ZWg1wyzvKM6X9k/FiKP
AiO9r/D8yEldV0CKE7gJlHSHZgGQ8x4CUqVMjIhvPQMMEkWJv3mgApIUcqn9KkhA
PV3v7S/9H5imIUDTh8lYswW3hYQ4VozH3HpIFBqhXDeBP7JyiBBzkeloSElfQgaO
VigI1BzSIx77QvY27G38fKDbGfzw2aoTLXUFv6iV+9J6MYzfjV1/38ugEuhT2SV3
fASoIhShEpZzka05XKm2Pz1AXJP6f/7IAIxrzR8AoyF3LRIOqHkiL6DhpbZsC5+J
eUYUZZ+cuE0kutAqOCpLAuNjl6mHF1Aa8CCMc2u3e+dks+nhYyOe7idGGWE2+osm
JFNCbsf+pBCwVgSBKQrkcrZEeePr8i27AqL4hhU9L944D8k9qoy9X81IvvPist9F
ZgWc50eaovpNIrtOMMMz43QtuclqVQSj0EwpLdodcCAzov/djN40qDJ6ilWtR0cP
IOGfkxpbOfUP5zdbC3uc0eOHQ2faQEDmgRlqgGWpxssn5BpiKj1DS2/Q8WqEucl8
tNHhWCYysSfkOQmB+kOCyJ4RVAejRjsMhIt80LVXr3A0bXcxBFv79EcObjt9sO7Y
gI4KWWT3S5fBlBAlRsAtBN5C0SlibEsm5Y9rcMAn2gEoi1sRMWOrz3C78YXvyk0S
rvA/1uzAeNTfU/Jlz0y7Ippkqe1x3An8tNqnU0XTa8w0LLbVvpbEDDQQDRQ+0oY8
VWDYr8f3eP3C8ylFSOP7nntghaL1s+lCmSNRAGW60jews2HDohH6Iq8Uo6Ix8yIz
R9/LrOTcUsvmSVC2/T6mnujoURbenOYYNHBKpLRa9je+JUH6TnELJk/2GWOKnd+e
NVpOLhZeBJCY/kaZQBS257B0RskTXdPRgaQWxwd/KsdRoXdVgtV4BkZ05gPppN+Y
b2565XHqh9wLQypf/Q+jV31YQzwAF2NYPyE/J+vkaEH3Ch9hbLDvSfgIiMMKIAv6
fvBoPmSzxW2KEeui6kP+rV+qUCWpM+Fbg9LK2hhBUPlP6QcZiPgSm/DTRcYhXZsP
pmtB1GYtdvGi4dJE4djOazER6o1a17a+wTAB+4tgefdTb0OOrNHoyfFBLxFdW1we
c3vvQSS2Sf06r8jPQ10gHFhDMrXQHIEgCz3VY1bY78otPAL36Drlm2/0khtYrxuG
emv/sLMHR1jSwRkwmUAmQGsl1T9xZ52QQ8DQWvqTkZtTeoGVmrnlFpOX7LZdbvl5
72mZCdKSZ2Sc/ZQRKvf5yg//9WV2nZAfI5ax+t60q5G7LqqcmC3EBbZYSHK2GycY
rKmKIgEmNUt6HTbAo6oCmGpX8rJCo5Otl5AHD6OZS4pnrgjpGYgqez+VypvAYspj
5dh+eKw2bTnAFc90XiVephcKqvbbxWClnSfmvZPrxIiUZgxc1ChqnA2hQtJpoh7D
p6lBo1+hB3Ze8fWf11cskbP/V4YuFf0sWEDBEVMqKTf0b6nlE3CFd2Vli6GydRSD
LiaCPn9f3QjrL7uLT/OqILOYUrMxS2A7svKEVVjnKnofWPluYkSVsL2ue297up9G
DefjwTCfrmOTchLYl6xSHlPxPbcWLwXGMfxZESAgjRnNOxeiSQsLBw1SYuXOpyli
BD4kthKjz33cRG9BrXGs4rhP/JZC2hc2eXuGAVwvp0bQaIC3dU3snla9x6z2E8Ku
So4rrkwf65hX5Yujb6lNg6SXonIVWzB8WgJvJieRzoFaVbjNlwezRjCjOsbfs5P4
TtiFM75m2u8/cIJeOxKVFcxLegMATKpzN233wKa9YoMCRA6lrrZAGv6nxDhPC4YZ
Wb6MDbc6sxuyzEP+XlvQQzkn0N1EWTNu7twmJBLxOJeyCCuY2vJ2UdxcU40KGCy/
DX0F51/r1Ucdh0n1+t2Dd7KVUK17We3p0rNYTXnEVCAf08itu7K8oVPNsmk2HUCL
GY1th4kT85RC+ZrtefTTjjQHKmA39U1L6Au6FUl+//HcQl2gA/ygCsLYI8tc+D6y
HqLEdCpEVnh6AlMUVESIs3BtcCn0I9bBvuFxSKrn5x9AZiqbXInlYF/fp8dqPdGJ
dEa0+ziY3KkuEWAvUl68TL4qQQLQ7P878Hgja+q6hZHrVzDnyQpTe087quWoxzRr
PCZnpcbyMT4awFIuRAM12H1quRBnuCNot7P/yMK706+iTOBrUcz/k0zinLM1eqrr
mquvYo6/jWLe7te5ywxILFujEzK0t9zALRU3fgD/YQM1EBjokTIv2yg8N81/p/B0
GvCDNqoxzw7xVzwSA6st4rGthx+HwKN9tCUB6ZuiMfGkv1vDxhHC2j16Bx7EpUAV
bdxUpcakeTwm5lcc1wfjJUkhdyFttZ9hK+OIlb4sShmhefTiIr9V7GoYn3++cspT
e0S3eUQcw3wdr+C9MYNvYl9LIDcE1ThB0Dk10HgyfrY7Qo6EQ8VN1hpfibnYQWQb
Ftkq33UIKET3YNjsv7y9VW58ykXjr24YtO8BuTFjaa7yXjk7rgQOhCuoAdn0qiXT
reeB0bR3D7RMOCCJpH2EVF9sTFsUuwiMwo3UO1b4hM81qp9p7nSHLAyLf3XMKDps
7rJppRXeinJYnOIYzKSz5iv7lLmUHe/q5qirfgE6774qFXfm76z0pG6Ef9wXvBWQ
Dx9PoivY6njJ4OELgjxBj61F5HjqSyP2oAsZYhu/XHVGMx2NzlDuSsjneQq9bomB
2TgEF3JZ3rqmOi3hm04+7XXtQ27NvM+rjoUGMYxO7Za83ae+oHOjC5nDeoQTL/wh
hcMj3mRrWDiEoZwvczKVgM5NX43HvXTt8ahyuX/rBWFfH5BZZ0BZH975nkrUxw82
gURP7Mo/Aj+yayZO5vLFknA249O6QR1fJI6qXeafUzYzJ1YhrtyvkPz9Hs2O38ec
t28/AnVHQeS75Nca+Zd/jwLLt+rrFGIkcy9WnVX/rKigQMvjN4LQ/fB5SCIIx74K
ElFPsqA5yTa6EA0SeHjnLhPvV72YyHgKmMBIP0YMlDqfKiPRl7NacpjUJ3sCYkKU
5cUH2NscvyHLZnVDVRif9G6DuoNRBG5v1StyGgG6lgZ19a/5aBydop8xV6bsTkvS
0wAPcbHAfLSKgwIQUfm8Zrs6ZIM+CAQZNb3SLao450wwa5QrWvAT6FApomP25+3B
5fPH3Z8i6Zdv8vlLD1OaY8MMn87LXNQgNeFdKrEBHHJL8o7d6/j3ztZzCBle/gDV
l9CsOQlxYfu1vpGOFHE/0fdbmdLd2O60p1lVFUq1DXVxLR2rvP2niWJqYug4x16h
qjh08Pgka+YiyWyKNfw3jbx05tEK1K9aVgh8iCYzhvTfjUFr50+RhOQ62UXKwGSj
y47JdnW7au3nzN2MNxDTr6TpUVGfBBEY8yBZT0/sJ7zBqadhJcTihc372W6zFX0M
8E7DGUMR2NPU+mF5l93Y63wfqDjn5HYUD7ghUfnHM71qWt3UYDhFPnsydFTIuc/U
zjsGAuZt4nm2vVn8+B2LIcOzwlSqq5Gg75GNah5tcjCSvhgb9yluSanhdMC16TLd
hwxmdIvUzdN8f7tEccAVi9ZL99JxMTlK08V9t48hlatOUoPas+42YyDmDSa9QtLx
XOCRSnbQQhZvote602WDafpoX+is4alXnYfCtIncX6u+6gcGJ/2EmO/XG4Dn/sva
PLUX29+XRx5ja6FxE6Au3h9YajkmdEx4enmrsS8bVrFS/aGKV5Y+nwVTTEWP4EF5
I25FwqodmDKBBUNuhG/UPpxgUPZUQydjbqjGNGF9M0wi7RnFPx013fljFbjOPAKm
Awp2DQIDsLkBNpb9D4koQh7GpsW1+gdS7tQjdIIhe9LawxSE/ali2vNzyY60LDAd
OYhDrybIdO5VMQHTRaZxYYAOq7NfmnXCdQJ7qlgb5r1AExtZbGzyE7kqXUF5qrpB
bfcPjmznM2s22f+FBUirhBxgw2GYS3FuxCN4k+6J1UOorw8BHEJqymaGt1jj1GY1
w7nRtjyEi2tCky8IaIOjDrh21iZ/ce/LqaCIE31bLR7e66XIk0Y9eUhn20kKcBq8
MPlYHrknp0sGyo+tbcRqqJGGi51a6LAr6RcrrTm/m0S7sKdmd/bNukcuaTGChHzk
ENmXloTVBc7ZcPPUHE1s77Vwhpz9zQGDEQ1JkmAiRrkWwQ2VQZEjdL1lclnEe+5q
ssOD8I7BjWWosAudqts5ikwZ+jnoMltaF7VoxGl2aQAuhBTYaIcb8veFXvSCfER8
9paJ8zod/nXmk3qqYZOYLI8aAioD/GVbqAsffhG9bQeMbVFtPMd8xjRSyOWPlc/h
lfsO2afdgcdhcEeShinkjmAb3gd/g1n+e7194X/oBJYpNqj8WqcIYfWSQZVakDtU
fo/R+sO5Hz+nIcNWf1mLmkPi7uUVsUnx+Hl75Tjs8i8caw4C0Om2TWUZtcV+gWGd
XF/MHg9Xplm2QHSv/IkNpuAkY9IkXi44dFvmJALhK7mRkMvi/+pwROU9J5oLc3in
cZa+hMAfWwXy4H5Wqwy3Oj9jgcNEMlomwrENtqM3yiop0/1/mIW/BkvhttMrJpx8
PYcyOn7xXtjwkFLNmaAGkQFSgKEQOPKadNTmQp1unxqHK1htBBJh5SAgU3e0n8nf
lyZnfIQ4X9rK5k/EAKN0uS2SKB0hMEAZCg+hU0Klwmz6d/MAn5TZpPiaTiLehuPb
0d1JcyYiowu+ip40ktEZzWWQE2648s6jSlZuH/yTOHkvK6l9Ljfc6Tn4iMSJPs9d
zPB6qubzC2SJ4r+IRCY6kf7jnV7u7foaIhfdbFIOfo87weE5Hy0q4Omq35Fesmok
L5ILa9/uPOYLcpJT05a5XMYc590yiIMDRhzrFylG0iSYDTO//+afA9SkUmCZ1+Yr
0yJqrHWWZndUGGdr+b2HZjGj0VrFob/rzufqxadzLsqI7RsnWwakvk9pzt3rqEVG
58GE1nLfXl3ORK79u6iJMd9+skQDb8UTO1xNYeskeDoZwMZqoIGytQsjpcMobryE
9u/JIINNriYCf79nTvNmDZtBwfO3tB2sR0STUv9SbqQiR7DPjnYGVx7RmYDAelNR
wIs7cPPdnKgyF81yHsbQhAGiP6tee//ejqE5XHYUZM700NsuC8m9CDkBJ/y4cM2I
jqF4e4IcCcH1Sypy116h2DGCbMPO7JbX0EeFNFG2TsXY5P5SgKSOIQTNHAi6aoxL
doe6pwLJnGGYuLFxFUuWP7nRrNa527CMcalZc4Vdk7tCmkPzpxPTtN1JomNogFPs
xmHUulMKpQSQRfw6+nQKT91zHoK4fGsIEjnuqPJm2oVM3TDv87777+SAUcuiI6jc
nIrm16bC7nHuTH6JJACPyR63gCdj9td9tmm5oiqimVMMl+0OWln80TERPZUnbe9C
9TYENggYoBo81zbC9d3aCMyBEOHgrE9o4Tingvr1DmFUSgubxsa6kORod61NogPa
Aju/7RAw2okjKgrpkkfP8IfNbeG1gkixsesQY+GCWBvX2xk1R7NVFRs5gfZDkEs4
xwOKyORWAczzXIfifc7NB6CX2zM5j2r2mSQoky17co0MR7u3SClKWJybxB2y3RtQ
gzssHd+zuwr1zLTFbDVOYQD65uMfcAJXACqXtOwks14IZayGkGEck01xHR9Zex6G
ZvpGcZ/M/uv100LPxiMLdICNM601Qy4XKLlwXjGg09SZ2EvMuJH0boV8mRND7Bet
qb4sDkOxyloeX2HdcUwkjUHcdvCldNn28lV6/QutJ2fYeMrGgoxehbVqCxfZFHw3
9mZPLCVyt6HFsGZqZuJxkGOi9U/kfcvO+P7iYxNiXMOdVla3sSeME4jVFHEfpCS8
WGqb4mDZvDzFIHwRAc8XJJTZRxZfXrsHoYQ3ZHmk9CO8MWFzj22z9YhXIW3jK8Fg
yEgyZzEOmvxDUTEIAsz2FdeUPzMgkLOkLS/8LYEKgUlQQsm22Hy6MLC2hslPwnn+
e+LC/I2gdsMZUgnEG9Qal10CzZsznQ5+UzdKgyrYRLrCZM1dpjeNdUGHc4qoUS1l
EsEdshFAyLHzG06TNtsdZVCFvgtu+0gOPG1nsEEQDD4KNjAK/02quRR80bfibIqw
F1Qfoq6wnH/yU/4cKicC9cWNIPCM1PWAmM0WzwcA9GjYUr8mQkWUYQmve5SdNftF
Alvuopoj6znZ/UkY6bx9fTyWAmwKWuCBEDrYlmCovcjVK6YwjqaFi8FUvZfztqYv
s0hzHBqH+GXmzuD5wIIIyMacwPkNsqdF8Ven6pw32zJEPVYG4c743byaZL5x+Xtw
IQIhv845nn+XJ/VuQ376HVcavAKwhqFRoeafB9Ck1ZwcRbiIP5VegKRM7sa1oY00
IMZWNqcgphOTH327b16JExqScReaOaiyU9u+EcbWwc+Ci05ZoDXlhBPAuYSnlnNP
baniOk8ZEV3jsyaUv+MSc/sQ3LzX24+hiWvY+SvQFBA19jrV+FcoyzKqKhJaRtbf
a8SxEtCKDuuYSahtrF8MytndtwUc7xKYNUdRnPvYzgW11drVg3X6Sl2lLiZMmrlG
bSVqvCtcIrDW4n4m6mUALcNcODTGaqKtllPG4Jy3BlaT83bkea4eB0P0ZKAVwx//
CNrjlBIWD3JWIrvmTq/1zrukRoiLdHWBeuqsUmdrykTOiEDYzZ7qwxhtmDyjfYS9
NwIvwihUxHPAPqwfQHOlcweb2oxOKk2LE8F64k8U8ocGyaL1fX/V9aTS2TV4tcWT
NSof1i6UG6igYvrzDfvm5WAXJ6oATs2e883i7FVTdVDBvmGmezc13fDdyVJOOwZf
7aeVwB757I+Kl3JRjXydIi4RXZP2Mlorsx8NapvHpmmNx4wFSIi12YpCLubsSlNN
UznhAV5lZm2+sBnndO6wLLyW387Jvm5zQGoygwEKuJ6vKNxqZyb3WZZzEE8aSvwV
eKPRtZojBPD05WkIfkDpeHq0/A81tdxXi59WErw492pzYHv3c6XAbPhOqa9jcEW6
c9P4iXM1J5ShiFaYPQBuBwUbjLxV+zVMKtoSF0pkT/gKBl4MmH/WF20vmNelGkxr
dkYdrdIhArAkqLGn8XRPtUT5Eh+WNCrZ2+9YrVXYv+SRKrdEOZxzFyblSBk1Rh+g
IVZTX3TnuQ9bnRKg6K9jM6WwKzTCliPRRclv0dTKjcDPcJfo9BBWLTU/9Apvlaot
E8U6A0y7oHspMM17hyjq/VEjTFH3UVy2//W4lnggHNOQtKv9lGTf4D1WjxzQ9lOo
B+W35O0PlFukDnvpA4aDn+BWpyIaO68FwGMy40P+sW0Rt8fNdJNyPRzuAIszwak7
Sha+loilXzQTsznG7Z6vd/41xYV/Zr/5eBy781zH9Kfhls7GmA+oi0Pf5fH45g7b
hYhac0qqbUPYklM7n1qwazXPISuMSR0j3rIqncmeycpflaUEeH51RZb9Xnxt+HBS
D4XZ/PBAqe2ap0F5UGv5ypfEt3XhiEf22SWHhveeYBkW8bn/b22TdaMbFEjn4fpu
BO8pIUNB8qZasc1a/96wTlLGQF8EFb4iXz2RC0Cg//r4MJIJJaMiodwQFYSZYpFv
k2LnmyGd/WZALqccLjV+tVFeIwvqK21HvQfzFWYfjcGfQo3nc2qwCFP4QB+5tcuv
KiLKV1XITL/K7MllYsnproF6l+dPR0yp1v/Bj+5gRuv7q27JT9RWcYIHabBPtjY8
t/ZbSvEMmkPX8EHd5DqQDTTwESSMPC1mEdRbL60oKgkK33vGx7eLy4fczMFpa4Mv
IUXB48GUxXkV213pNqGBZAk5y2ju+i3yDq98VSa0ayyeCQljNsNKxWuZlwd/GgfT
LKSBPXDBScEY0iRcO9Qr3TAWg3UNB60bLfnn9JUBNvchY32zevphPbiCPkAgQeGu
PZW7ZZTfFvDvUEGbVzT7AOjlFBwInC6NODFXKHqlP9MRGfGBXGSoIY49nWt2oTaZ
bD02DFdBbUQjQmw78jDTuR2CsegFEfgDUrXM5KgUPaZAS91aB3LJd6pXhGfrFy1X
uvtiICM+LqBMMYqe/gHTLPrGWnje8IYGcGZS6PF0zU6Zd7E3DUE60vra7pI0P2I6
Jv25cb5AR4Mjn1tmnWon3yiaslIKQXgd7vD8RZWtxUxecP7ZFs1jE21v30VcSnGN
C39swICbAERaX9QpqDNfrEaJ5Fnc7xY9Tq+tlQwXPXsw8/2KpHWDeKaob/garIYI
yOd844ZCTbcqgJM5GftA8TCUSvn4ev5bmneZlczF4jhVtjQiG0OoeJ2l0oCGpM/u
XxL/PGJAT0XySWWR2u2d2P/ElVjuTvACNzzpRfMfOj2DNzwKfKtvyZOMapZwhM4u
PSK3IjkctwWUwosAnbidPGloSYeVmfE/IkxLHEhGjuI+JSCcwo9IbDgO2g5KIX3n
NwbF+qRwSZUb5ZSgQtjbewA8Pyfgc96l5W73BTGco7J2IRToA/iVtCjZjdpkHGcY
/PsQ18CPYPB+Q2KObngzdPv6aKG0UM+I9O13Sci0kJBtsEKV9Da5WNaWD7qZbeSp
XK0MW5NWUtVk7AMEAKCTq6FMolCcNKGMwh9y8ZrUaL/lBuOGN6mOYYIqH0CxtA6i
KcdBwUJHoKTqsehRljO72L3wI0ud1oigDP2UfB1i9PHgXz3OtvazKKBRK02e18B/
6Msfa5gmU8c5fRW60wHT9VS/edo5WZLYN7QrxXT5WcIZUZrXxcT4IuLGe52adsGV
GTdyFoTC0qJpSBognXAsxBbhWp1RUT4Z+ui3fTt8zq4nUNN1LPRrR3EgQ4PBJ7Rb
z1Y/KGskClAlJvFggqHEu60wGd/+GGNgsgvxhU/6z50NPJW/mxvi+Yp2S+y2r7sz
HzLhH24IfLKXuT65PJh9Ccw/Ou9Vo1Anwq2gOmJ3DumTJ5O53wPSxZhQ9hHt3LQS
C2qIIFAgyR72nh1G0f8H9VcvGJRejbsRSa9CQ8MyS7DWwa0qY/BAaV6/kqPSTG0v
auIVzullBRj8EDByjf30jh/SlT7SJOoo2NrmLmSUHyY99e4cM/PEJFeDmjil7Pha
svFkgEQpA/IqfVglVvzbNey4OPrgK/xcyEhdKMgi/ErTdZUqAHC5BSUxPbllh50v
ob3u2/CfUsPXy4qgPK/TEp4qhxvESI/T8jZx61umAXpAgE9CS0mzT4swXfvbAr1T
x5528pb3o0OPhHlE7nqWMHjQKgLu5hWE2FL/s9tlw8SSOT41Pc8qqeosOt4NV2yt
YYe/ZcKadw0DQI4rWKPkLWJhMVRZM5fXL+Q5LKY1QJIZpC0KTjka3WAjPvfssYJk
iWxpuAo7LdLuc8kcWRHSLp82qjpG1Kd5vytrN5X3iVpWaZ0vlmQUN6k0QX2C8equ
vJKftPmcphkGPv7Go/Wr3sLNyBGjwwzzBl5zf4/Wqlgy0ihXAulYCLL7+K08xE2y
00yj7q3OJXHTaFxsqwyaNzSE+hog4n9OEr+b7aVkEQGWMk6hG5y1f2X5bYdnnUxr
dmM49IbjoF946kuZ6Zk7LoYfZfaHtMVpi4ipZabJsIn9A+vMyE+wMcMAFKMa4JeL
EVR1TesIDZ0C+1RUUodXLM3nP6YrgdtPm3ptblrNWKrjudkTjUtlL64jKwe2cD8o
VzsRQESpoGWqHYuQdJdbVDwd4HnmyN167YBZtIsG/hUC5hMsZqwdfXCES4VDYRiv
9kiOV4Wz6hGjcVV0RzLVIc29T6ykF1tWBTKY6MrNCtn3+361iD5KTvFGybabzqE6
Fs/s2AEq6yx94SwwXsAG6OOZ5j6xTks0Z3VOzeF/b6wZ0ooipaZLG4MCCF9DIqT8
Rqd4YN0ci61iqhyqSv8PBnYC1azW4nogmtshOU8TG4GGuwt+PfEKhQIUpWFp79bH
Ry6GSL8T4VxsPDdKZyVmPEEckXSa16pY0GjHUV6+ZOBsN2fyMjzXTZahYEYiuxb6
w1zUPc6DZZX+HqHChSv1RepzfGvumzfsVOeUmnzJCglgwxiPVLySgRihG5O8+xUU
zrzXP4bnKoPF+W/cqR3cn8zz7xg9v1EH/+S/JWw2+ABIRt/UYu8o1CwDlgtV9lco
6lf9e12rJARsExxT4BXv+5jkU+KSKiT0pkWKuTCPsd0ratbhuFpIqtYMcw413SXY
B8xlwingeHAFNs/VJLuLZ2JjZdtqpYQmb5NMGaZfGqSkqXMtbjyLQvI2gfONu4Ar
XEIvqnB6u5E9atqSgJGfWOQm9LiGZgw6hpbr+Gxo9TSVK4NDM0yWWz3MxZKP7BC0
fJzkmH3fa+4f1fm/obzVkr6VcY5+Bg/ppkkBfGHwaJps024YknUj4OSfNiZB9r1u
p7fcSLZ3TE1/VsDO9zjqZNXSqGF1JUEhHfVYKzCDDsuKN60Il9TwaeEELwkot1uu
EuFJfgfHrEoqEx4GvV/VldIjB2erKANRzqlf/pRzTOXRCbD3T8UbXdyB/zGP3ZKr
Gnt17CIYVoxhIzMB5BCwrQN5KcpbCIRHP5hmuHQ6TiBqQu2UbCKBTiQgq5CrN5bU
4sxMI10wx7dVqSx+yoOVP4jTFDi9aMF5ZUApU1DoJYdnhohFXW65NdQ1Gqy5q1AA
YQPlgMbkpVN/TFCZFa6U8kBCEwrCBcLZe6lRjlgAc7XSvR/n5oP2uluS0VZx/Dg8
SjIeheVF1JqdGXBOxoUX60wsWty/zVa7JoUP9mgmPRMU1UENLUiaERefeHaPmcAd
HQWHSsXtuDILWWuiQJQ85Doh3WDiG5CKinpLQfqN6Vnrm7YZkb416txtas8g1ZSQ
hr8LeagX3NKdN68nkRwbhflbEuUU5rKILaBXxgtH/6OW51Q62zZickvrkdI7Is+P
plLN5NPaKQQLkf9Uhj4Rp4UvMRSKwbI4H/hlN1grioKj3bPZRoLl3ioMsowqZx/S
S5XN4kIlLhtADQzg7rX6um+LZO4avcv9kL7GZbMDTniaeOVYzEK0ypbNibXo40CU
0bgh9yN7o4Ys+8Fs9eECOkD2tdZ+1dG/TLeRXykJLSXYpEXE1m9s4jp96xoQnjco
/1ENTVJenEaPHOQ19lGTjCt5XPjJxFM1xQ1HdqKGK1nkFCZAssZ4cHsD/lShXQow
fhZCXsxj/XkK4sD88XnoEs8Nm2zK4uX/+CWdXMfF++ou+RDGKirv0hXSmEW46lzM
SXec8EDtSrnqXZKtjlgvH3UqWVi9p+l9Gy6ukkTgq29nAAOJ79PO/Sj5c4D3k8vC
C9MkB91JESfa7KIzrwGKohR+gMSkyDW2z8Epl2pq++y7T+Y1mW9khX3nUKpOcZ/G
YSt6pR8rWQjXjSJ6WZnFfem6YKdBgeFjdnqwaEgo38xlmHgxIRqW+D29IsPy1H1a
Eg5hL4P0xAprp7Wc2MHWZ6ZcWCV7VZU/JSlfWS8fx4Yo6f1FnEKb3+Q8nRMR3q9w
sycHEZ4E2PjjHdBCPaJ6TZcKZ0WNAONngia2rYiBlqWcnIYPjx7I0Udxe5oUAPDR
vOuEor6jT5W6w5vT0tsvXGLKdoCFsRGNrO6vGyT3HBtg7QO/XpKJWQPFTlXxrbB/
i3VMKrrVDLjFgQNiBGJOzNhEd8PpIIl/C+Zwk1cw/Cy0axJ6+L1Eyi5JBk66EteN
aKz8rqs0vmvugqSXdMsUI9QuBSCMSO5CXwrBTand+eTYSoPsuILrUq6KDUMmDtEN
WyihwPAZ24HdHObD/TMiHGQItryIaw6AmUjXPwnOrIutipBJh4EgO/r5hO3/99de
dBABJjVUEIMNL+vJkqdoGHvqRsV/6RkP7vYq/s5x1T2jI54qZb7ecDXNLcjgezCd
xmNfNOQ/PXMHZ2aSubOTOpmJhdCidYgTry4v7a9JWHIIq3m8Q3oO9E0I5wwNVA5G
dtqXz3daOXMrosMFWk2fzq4RcOA89zby06aS6wd3K/ekI7b5cMGBzPjiZ7h4gr8L
CyaL/kbhN9/e3GLUo0Q3HgtxVCvPTWIaYuZ3hxWy3zM/nhjMAf2xM7rUzuBlCo9s
lCcPayb80O6ntamm9zuSJSjaAbD9hQ+Y6DCnglfDTxu2/N5TfiNfKBkLYFUqEqFQ
ywK8YfQGVGHCNnV137KkD/dFios4l3aZgPRTBuOxRx8td5RKd6hus698R0Pz+TEY
azWh/HoVYiYxWV2ZotOGNw1s73wiAiXaug+V0x4prA0kmVGi+G6i2oQYkkKM9cBm
9rHzxNL4gBIksFniOdOPfLTBc0ZUY5NMqsTJ6yyC8czdGwFhk6Ezm6074cTSa9fF
k3lEo+G+gcMTpMEMBDwJTeUAvjc9CUaZ2c1FuqxZG8EyjMEBWi+IW9VgSLiCPBkp
/sdeEpeHOrCdddiUT667O7fbb2qPDQOrtL1EO7nPtXuPY3pLHc7jjIOetVikeRM0
Va9Wcu+JHWmyBoocPjQ4ui1c09Iovbyw0/7DLjqkkPDAOZnaHTRb52wOuZUG69da
gI1NxNK3yYBUkQosz2B5Ud0WDQd8huB4pwEjUDfdHgLyqZLonWvA5fqC7+la1nQQ
PyAMOjOhhfCCb2yEsolSQIiS1h72PjgG2c1kvW9MvvcHHh2oKDNE1Rbu8+GK2xa1
6M3ifV2CvOTcNfEz4cj+WgmCRPhVC6JkOTuVCTi1/MKAhQYB9K2CAUSppgptaifH
2nnMUYCYgr1pVvaWspsPPt3Hzal0QsY7fDIKnRGA2r5Kmka5cCfwi2q+X/KChFqo
Mtztakc7QY/dkIq80Oc/LsTcQFg5aCgpQEM0z5tglDIZvG0/Zb5giiknFd7X3Xxz
5hKZ3VijQLbzN63QzuDvv7/9/qYUbVSNXpN2LKTT4r2OvWtVBtg4nYy7bxEtnbCT
neaMyB3xqvuC+l9QjzK1SsqtPHg+dnnrsNMYVNsriB6EfVfL/rJD9w/NO++bhuXI
JA5cfU4pKGbKHR5+aH4+pLUDk8yRSpm4IdBuXO5ryJbi2bTfqgO7Koi1nR6/fv/U
32yHhfjF1VoWzve4piGSNZmj4akwKkY8dVyz0axj0rdN1KwaNMu4Q+p8GZ3EBeuu
IBWYilGXOMCV0G9+yTps6Vuv5i2fcpXw9gg/70N4ZnRGxxlu0qWZSKPvP34JZU94
z/CSyUIJBgaRrC3egnlf7NHcXkoGfasUDXCFzp8Xssqk/r1x1FqzVrCiJn1dfVIR
zugT7/s0Np80q2LNC3if6RtMTdkvRHRKUkA+RVCoCZ0cw4t/GK+vLMQ735UEXhGV
ijSZcnEHF3XpgxVc0vHqEMJHOiNadLrM8iwHF4SdGikzWeC3jmlJyqnjaMWosKmv
6qIzoZlMFt3oZea+hFqo/Cp4WBrpJoFr1jwYaDeOCYOwR1MZZQtR4Y8lMlzTxYr9
84iQckm4kSsaZXLPWyLK/WQk7qS9eFm23J3n8qMCyiaWp09Bv0+8pPC2upGXQqrU
Gk/GS/71mKKUZoKEcw2+t0Mjb9wNp57jsKW2oxEL4RofdGGUm1vdTY8KFhUDu/r4
LHYja+xzomlUig//WrswI6/wyjnvBqoyvnAwYkCr9zaaICqJg1KPxysH5dmdX5Vp
oQq4Jtq49dffL8ka4bf0RRgWwcBUU6gPjKnZL3jFU0369fxQpufmuCVnuPvExCpe
Dq5T2WJ4AH4q3431/oAIq7cICLKcm3JQe6zIDtcaFgfUGcV2Yua7q/lvFr1FxcDo
IYzRaE+iDNbypiH3ZPm6YwsXgYcgy5moF1UQt7NKl4s6rxxX6M0it2PzZkyM/hD3
2UBMeL4FiNm2y9R1rO1qgIZfrvRWvbOMnY1T4bJzLhv0nBwxaFtNQQZrPcofoSDb
lhi8HgjvqrrvvSiHu0sVR5lVpXE5ogjz+4yQD0pXBlaWPwW7jo25r+MNBeY7kxvH
I2vspmck4rpnkRQ/xd2eMj62TLjf7kE0boRqbaE2loflWmP1tPp3IZePH9mG04Wb
y+5zXHiYAQDJKOnpC0r2654rV2cjVLhHXAytJ9CK71nYaD6NAvO9G8T5UWhMlvBj
sCgmA2mXPg9v3+Ffe7g0J5EfXiPSrl4ZED6QLgza3ZQB1mUHNc2wC4iQ6LQmRBEO
SStK0o4eW9+JEwb+iupMVA3wyFjJdAbNZLE0gYdO3iYY3QacF45z0tmyO751aZfQ
516nFksPYtsK1g0zOXgvF5NdXaVNnNzggemKWIQtrH570lmiOHxIY6y/7tR7GKZl
rPQesZe6m14ARTkUiH3gYBi95gEibhIFalUc2uf7vbeyS7zewfa3AB/muo0FCErY
3xWmayHYDoMS5bKP9A7T1qW+0uINj7+lpwJ/7TtHGKwRODf9MYOS3fyDqCQAXJZH
0TrsGOw+BDvevtPDOjhqKU/2+cQvFm8IdjNwVPvKkuKrNkI8Ug4OknDXJrYBMJGo
85oeXtwTzmq/WTY24g8KCiMd1yvSYn1J5VN7BR0Kr6QD4DsG9quFZNTEyqP3k2+Q
4tVDCkibGT1rH41JCuaUL/RxfCEZn8WK0WiboQFubuPN6F91nLZxclR5Kkw/ROIZ
U/Wynr5FQfD52d5K2f2U5FxiYerEO7MPXCYvNk2CdHupJrt7WBE1+sQeNuwAkeWO
xGVqtZaDCWbfIzPJIOS/uriUGrGJo5pxBzMCxESsUyitt2o6ZgWvf02zYpaG8Ziq
5dnPkr35ZZN3wpqdD3KSmW0eNjTM0KuVXPDPllfOhGv3gzjSs07NTAgU/er/cIlK
owEDacghgcLVjVu0NvQqWusfjl9CqtyUAaTXgiz6JqPe6y+wMFmqssDcHJYpOn3W
sOEoDGf1Gx8ZRX2n2A9Ib6sBmRPNRrwmIeNNm2aPEsbZ8ro81OoLz4GpDcxV+y1w
jG5zeBrpbMJuF/gI8LiHhWIewqJ4sEtIP1Aml+bQ8jQKUKIy8Ulon1NesHY9+Yjn
J2pLllo/j8dlu9+cgKrq9nCTmJuyee2BswDhsv1cVcPl5VLYObqwGh6JlAsrj/vw
pgo52RNtoi/pCRXFPT1tXCQa9fY6BtZ3qFJkoK2CNQVvlpbd4IbjfEnFtsSvTCZg
nZovwe5i/jat/ro2xtvhhr9cKJOShNjchSOQwF5KWda9YdKFmd3vCFWf/o6GTUm0
DaNwTP/xzWzqHHjE5Wl9/0/DlWxpiRaWKWn3PBQ4n2SnHK/7zympAudWCXfqpsyX
SDnbHeyRa5CZL+9eZGTBSMXgm4Efc9JvVcBvmwqOqaVpvdbeEQzLB6FQwq8i/8Zi
iQTnt2BLcxwBnJIf41s4LBiioTla+cftT9v7PLpEqdOCEyU0gtybY3HRDOaJKMCi
UOvDJhlxkb/nFFv6B9oYuEYJfMhJOlynuTGj5YmfcCfTQIt39SQHb+b0SJvWCHKn
9b6dryrxZzUh9EKJgqQQIVp0x8gdXJG+Ga7lH/wkbBZmNtya0uWRUWDzx9fPV3TN
NSRD/z+Q9uZhpL4KnpM2QJ4cAbLl41Png0suIjPQJdw1972zzYP/duetZ68zhp4y
Gs++Fjlsj1Kl3NBpGF+8h+tKDZR/A6BF+oaYL7LoNFJCJBRZBsQbjr+U2mq2xiEw
Plysw0H6DZtvjqv2PHkJkdk9ff5f60JQ6CoCJDSU1B0mMzG49YCOhYzTuMPfnjM1
IMDAtXkGfjTx30p3NCx+60d7OYnlHbJK1+RCDr/gCAFiN6THLQRPdinkITc6tTAc
hnoX7fW0ZN0IIe3Oq2FWSv4OZvf6REvq37GByCC/zsNNlEaAcjUlXCSixcSOn6yM
Wnk0KvzjNY3PDKqO2RZSE57EWMCsyxDiquqXgp1mShLYa880jogCYO4BEkeTpcwQ
9PhYCO2SERAtTAR9NomSILSrFGgv8jIL1jCC0rC8IwMZOQcIVLQT4xfs/QaFFc77
zl2rSnJNm7t8/bMCDc+8cqy0vDbN81X2adXM63Kn9DpaQXTr1tZoQBR5Sx2uMbYx
EmueOZcDN3iK01VBMe6zPh8ycog8W80AO7KMi8vhl2Ot/W4ooJ7atUeaH1yAT1NB
itV3t+VwnxuBFt1Fbe2CHWBYTuTBFM8qmTaA9nTikhumEjKINRMTw3xithQrOs74
ZhbEVro3q/NnPCXKEtumdqxx6NUskL/+dRN4IQF6dn9ouepuvNpK3EaCsroMljbv
/ybuaQkqNgQhucslPXYfv4oj5vnNUx0g2GDv65RkG7Vr/fi/mE8MDsXti0NgWtqn
q/AefAT1ByQs9Rs/iwEzuVmA+eQiSLeaTEskCjSfz5+T7tvLszvtHqv9gaPvq8qq
tzNzq6oARLFPq4VdcUxaMH+CtbiqdKvCHqObCMl0Hy6znKiYg+GXJum2zVaj+hI4
LL6zE4rlM86/UOxPPhmydJe6WgOAyQ6Kv377vzmaOcLL1RQ9vwz8vjWJiL1bSJNI
5ZwzReNEgqRnc8frG7mfl4Q50EmibDLDKNDq1iek19c8uFhlXgYtTqYIU84aFt9U
sVyAo1F0VfgvvuzzelFUd0GvsZYbgOHBAgRhCxTczk7RlcLiYqjVPSS5ZGiRNIHD
2/aoBVTsm6OS3hI8KE38jaTNOybuDC74u4dRrWjUL4HQX+NJe9NqIImrE5++Q97A
VjAud1wIqARJTw87ntddg2JtOsVFBV3RhX+YCVlQM1vOJtoLvCmaWUg8WFHaB39J
x9lR6hIojzbgWMyDcZlv2lxbI9l4NAs9MZv1edLAQdK/S1cFxkB7v+k4B9hfEkP+
FgurePzPCp3qOvceARQ9LKZQIokADJ/GiXukH0wSXgCeLK2jeH/Ydz/unWZVPU3C
JyfW1rjezjWuIByxWt293370JmacRAg5ottEZ8Pq0tRB05PZ0zdhGDBR2Pp/qh2T
fzCYER97Dru+KTFhrXSwOQYn91yMk4iktYu76GhyRCUvKTDlOpYOmhBii3BihXE0
64W31i++e4X6LXx3WEeTwT94lDzYEZa3imuhpyw8kyt6bbcfY7r6qPVTnD/w/nxJ
9jf4XBGKAVts1i45lrzE3isjgBezxFXJZfAMLhJgio0xmPyIHcCKpFGO0QiSbyWF
sG2HxeO6t/DG0t4vXdGyM8eAPjuqAlds+E9nNV+eRNxqvG6+h330ZJ6wBLhTMry7
iHsm7ZPKs/qxbuf/WQQhKnaeEEUdrn6y7a00EcJnHUNjufGg6HMmYs9TFVXbt/9T
42zEqQuTL9LWStheHHO14qcsyYQSKRepdhzQt0nCK51+b+Lns0DvtdqL/nmpfDed
SB3HLiAYeXKbeu8DSv+6Y2/6cXSdNC9rL/24GUOraHFQW3OggYxmiaoyxmrPTKiB
nIZ0BaTvVyXV/O7iS0HSiWGOB5zTuo0bJpv7I3wJIn2utaCd+2+8sirv46nGJU5c
DdgxtfNAhNQtu6qAVdZCVlfQoF5GabA+m93iJGZw2f/UFEIlRB1MunS1AKgY821/
ES4TOmYlg+Xuwh18ZdlAy0aG3TpUdyvLZQ64l+C5+lkjKa2cvnI8CIs+jFWN2sv2
Sp58LqBEv0Hb6fIlNdMwz+6kHi1YbETm6gpaxZcC9HnfFGIheg4MG3sOGN5fxj2c
LnvCC7syoaHLgvld5slmhqodY+nY9fCSCJRN6dQ8ubJf+cFT3jjJyg2dICJ9iXqq
xkmvwvhWL/LW9BLhBXSMnvMZqc85tYgEEOaiNnQcZx4TdQDng7S5US/OPGWXj5Rw
JNQdFWaRO9yIZNl6sTBB5jIIZO60jbUapE9DGTWAqozgs9XF5Vi+hZ1/dyYCxUs5
tqwLt+aucEER9mVhkCyeLyVYjbXuXuFr9wdHZtr+bNYa+YxYY/pyzAf4n/2+2Vrr
ShFHrPmdG4nIukoyyyqFyLtfmhFtm3bsPB84QKnbkedV3gtHDi8nqO2cDJJ2FKyO
UGr1vQOSu0OKZp8TLIvtU+23EUXAjXxPGFAado7x56VBrz6MkszB6GQa/qQrmzQP
3Oofa1WU2aERDIIYs09FQR0Bm5n7xNMd8K17BLNn75iQMFPsw/8I7hNOzhTrF8vl
HYgOiOjLuT4mMt6twGfRwNpxzmPa1rAq4v403Zy7XgXkxiXhLREtWpZlh50YI8Tj
Sd3CQ7leRV1pkL/GprxHoSJb2H1TrK6BB8Tp/lXESmTP9nTvdw2T5CxAJfi0BcH3
jF4UqtgUvduSKrcgrFNLDfhQli8QXy8CrSx+L51UFWAFANiHoyIcACgU3lh/fl9S
ilReJ1FGWhxzmdQ97EL78JDhUJgkaph3sNbDBYqoTOkEYzhEsGGK4pW9asi17hgl
qj2cbBVHU/lOmIyEI3BdapLk79tvfA13MstqYTLIO4MWbq5Wb+U+WHMTeDkVh5It
zYhyVI5i/EPDVB/Dwi32d7kL9wx1HUmmSN61Z8TvbIF/BQG04mKQ4e/YGOK5MjZi
Iw0mH6aA0lEniXQz5f4yCOq8I1wVJYYx4WWFz8lrfGVvXWq9jYUkGKu6LTGopHs9
3kve1/tcnAIpa+8DEcCh6KbXBtzJpgiCUqAOTMB7R/w5ZCo70BOGGjubwh8Jbty8
R2C8Y/OGHGhyxpMkBgAgTQGfOqXg8J3JZjXd6MIt8gJtLHWCIm1TmBJvApBLWJ0k
C5CkzL/puDoJt2lz0Fb/WK16sTfUf8lHk21VeeWKhkBVfNpgt2GChiiZKu6coMpV
zbxy2YPzpqBaUqOCo8+SyYzvpSzy0YsHxBHtrFTmoMSl/b0UWTs+7KdJTamTughV
V2XRsqiwtFBMIj5h9XoWy4qRlvdy1LD6LRKo7QHBpAjAJaBMeNmZTrc4TjdSzrL6
ZILRMzbyfiBzftF/4u/+pW9jx9RVp0F/GNeydYIr8FWzwn7NbV2BBV7pqvXAnnuv
5gRqODDelwD7GcQpcUMTyEoGLUwqKaWDPCWfVoZ1qiJg+JK2tX5zesdPiT0HNzq7
VdLFT4umL1AEHxRTuo0gsJuid/4AFsnuVlbM1H6PKgDMW40pDwwbaCQCaVj5qLWv
RsWqHik1ybute54XM1290NEON62kSvZy3yaPuOFzaIuRnOchJi8saaZaXsEmSRsj
UgRskbxgrVif29Oz6vL/1SzTpdRn/o2kbqaiDhX/FA4fkCimOZ0z1ZZjC0qhKVJX
4Eq6LH37S+59S4gkegKl0p7Xdctui1uxlEdKjsFUizpdOqcldx45A0mrCcni8ImI
/mfmK0WBiL14pMD+WHXseXFbPoEP2oKtZLDAc0B+57PofKe3g0XQRNxUv0xQKcTH
G8pUOcfKZycIZvFXowrRTkxvP2RaR+QEYH0hh8+DRCrkY1Cdd5/3YTv6qF6M8ufa
Z6mO+zE8He/NPJ0GpZW05hkoaPKrJa7Cq7bZiST/+vwYTOEbq3GnedXVH2/VM93g
06+SGBzUgOL60pSG2qWSmBdCicIqKCjXk5XuBNcm8zAzYWAcy3a0igYrpSlQVWlM
HoIAl7ygpefMZdMkaOkb9pdV+zX9n1B9d2gef6OHc5BkJNPi3hy0kGfu9V0S+He5
38PpXxtKYWWIT1hKo9s2yIorRf20H3EB2BDbDuYrw7PQJApGxGxmLBBO8eKUx8fH
9Z4tEsBy2dABclmCy4y6FdKxgEuHn0HdbXLTyLTt3geA5pwQCLSaIC8CCmdpn2Wr
MDaLMp5ziqD/NPciGLdl250uOuDY7E0EUWy6YpV7Hm4G1g60uJ7A7O5sPsN48lee
t5/EJZQCSLmIayhcH64m3ZSUngBqruY/cxnktLYTzQ4J9YUgtHENbNrH9v9ljsPz
j9swMipfjTUE2W9n6eqnqNZn2pdYw5R19MvaKTJbdesXP6eJvENEqB9wWkDCZzWn
EOFdSoI2NPqfRlShRsQuL7iwQ4lG+Wzi544oL3BfRCdtVx+PJgeNhnBz2rsv1s+p
pDQ7aqjrGepMoB0rJo+fgxWioBT8kt7VRVsdr2Ticv+rX91bgutaoOCEWL+dMFH9
3G6d27klRMfMkhLn1p0L2XwbfB26o9TvLj6lwZS+plbOkuj0kta9YqRTVmxDRscO
bw9Y7s7k/FdRKdHEARg/XSPHI6WLOrcdS8nqsOQf3tIwD5xNyf6tWpVlp9H2TcRD
Dgk19uE37YSzsi3rQOiAmJST1A23CIGEwNZuOh2svQ+95hgncmsTWGy/TZpRzhs6
HnK2jvytb3IXrFE0lsX2U0kCCbznxF2ydD+SbhSG3QL0KcXzjt+mE5isBx9CcK+b
ZD7LKFv2VcFGfCoE0WZmbLDECoyPpQYCey28bK1f1S4Ng7Rrt0F9axaCq/KNUX9M
Pp2LLukxgNXFQxf2okaDNdusnL1vortKqLztxltBf3U0MJ/Vl4Ee2M16RGRlpseb
VnHP6ewSPFR6SZvzjzpqjsKUtg/tiTi8CXMm+aPpAGRBR4TdNIQ7pwUmI+2PTzbs
zdDXCr/KHd96aMnQnhQZ8CTZtyZrgWhty34Sd5M/EHcMCXeiZE7bLrzkMQSBYdwQ
I6pxinVmGWf3Q2Nllk4lLfBpfS+3b23QYl6aQhdTuBKV+XQ3oyCPyyYj7XkFKjHm
i1YlUQvBD/mw2C+aOSFQWprg3Q1dHYsVYPPa294mQp+MzW0xeqd+ly43An31jqjY
ZIpakhlrtsTfORE9L2JyjPsllGXZhcz/QiAUTTs1U5fizs57Wrj1jb1UsU/LHTP3
ZvjE1svCB7ElB/s+vvzY36EmMA8wlDGCQdnaM8zfxeiRzK+LBfLe1qqaXO0UfSRy
qr63X+R9EAqU4cLGjK1UYLhwwJjywiB0iFujCaQjy2XB++MXzKY0h5Zi9kPYHCkN
K+V3xL3mZN4j6vgYjLXuWnheMK2Im+Fpk+5prsqtpuNvY+SQveXh7IV1v70G5j32
pyrW+T+E5Vj5GaR8DLA4P0nO7Myhjl6vRa5yakbqI/G9RAu6Kxc0SdgozuvQBDkF
3hegyqxejQZgS+rkqDeZZjjLx44sbPfSKHXiMHwOUSsralCIVTwGIONNk2pofJOk
MOvmfo84wSH2APA1r2Oy8VBCxLY+PIdCJcPM8MwVaInHUHYENFr+9J7YCp+XQ7gF
ocNHiduL8xpOVsg/X14DfuycbeMDNYOPDT1zd0TdDgE0KsNnLkGCR/YUq/UXiwjv
7bL3+ixFbG6MSaV2Yg2uhQu3nY+FsaKGJHPcb9J9Bmw3oCkZq+YwUYvflUmj7uz9
yR+VpnmIct9N2xHj54k5vV7U+Sc8JJLUtt01TMVBr0HfQwvG+Wr1zsDcaOEYDoND
xdrnyHdyiaZiY5e+q0RH5XHN2qJMjcQkD6toh6xGNY9L4bJvhNPGnKaeme6ltArC
xrKDk6J+9TSiIX/L2CDMbruJhh9jp0IUem/dqymdP9oeYeEx4m077cqoHQCP7SbS
OAudDNZMepQmbQ0gzyLHquQk3D8Kugu625LFukCae6+CKmqF1TvVTXJz4SKGfGXA
R6JZ7FzlPUkOkeTBA4Wme2Op1Bcb0EZY8htJ0s5tIoYKYV6e8Ku+2Lnkp8EhCd5a
pvlei3FG+aEVCWbX6ZVKLdqUO8QWR1KZEMEvNg3G96P+0dMbNfXeW5tpd/T/mQaE
EpCjfRwT5fgG2jn7zBVpHuEe0sIldqMQssdH0Ftzjj3yCT87V9XpyuIyakLEFk76
92NhD45sA6ReO9agrr4bd8yamTqQdEXzYnPI6T7DiK5GdC4gxnw8tAqBfcvKjtK1
4NFZOafPpHCxmhG+o4qhy4SGZKbGL5spXTjhbwjbW6UYtyzC9v8yNkf5brkWoBge
VRl2J5GMorMSAnbLmStj8J7Wfys5oKDzie0X6ESpkjl+FzTFttxox8Gwg7e8bm0x
nN7TgO41WLusC4XHw59Eq51N3tiOiX5JZXLy9PdVYgd6JaMMNFDIW83zg/wVIoOE
NsLBLNrq7MwLEFhMlSwPSwi+iU30xXO5cY79kNb1Zq+kgKTlngYJIq3c1a/8ITql
EYiUsOy+lnKSZGcfElBKn4JXdyGURu/Nn9GgRim0b4VZKL9ZK3R9HjADUQcwmal9
bkKJRHN/UD70RR6BeM50UK4G3kzGWdUK16URvTkuqs1t4KpFEVPJSQZFrpjHkYfl
0hr8bUDK5oLmtuUMoAVdSTYbt6aydJe79A2TytgIVVzyhMTxOpXArifZseRxVDgB
qkDEp1pEfIrdpdI83Bzy88C1v4od/hva+nMm0L/eEobd3ERWf2m5aPDCryy12fMO
6yiQ9EctR4C2Z2J1VPVTVIifQpCNOW+46gDDDkbePEAI7trTVQjdfICltGVRD02A
Ca5cpZoi2BRO3wk0fE/ttxWQ/IYLwGXserVvmaOjMTu5gAHzhO0kFEjYvp9WhByY
jjMf1vGsnZ25ZeGrxjVtpM12nwHk48o0Vq42vnv3z6fjdeT2Vr/dt+E86aAfiKS0
lH5PL0dWe4XsIpoBUDDnoJzljrKKoK5rjJB2PAE9Kvj54/VMH9QkvNrvf7a0vEpL
GrtudQ0IzR7l+Wy4mu9bUZLt4DWVAvM1JwbUS0I2LZU71wWUy6x26ANpG2NUlBlX
04aJuANzH2h3PCntb2KIynWqmmKBWVraDTTyuME4uNKW3wcJuV168EeNgE/S21w1
MJOdlyb27P4TfRnNnZ0Ud1azQ5hLJEOkhm0mtbJr0L0A7alS0oFNXfvhHskmXF70
yt0OTz+hVt4FKk3pRz9/pyJPZzM9VizJaqcoPwQSS2GZOvYS2M9oErxYA9AE4RR+
lpPNN57LhMJt8cfYImjNFvpaKPEShwq2cAXP8vrFIvAxH5F+pAZchgXonlkJDwGU
ufhZmzVhEPT+Q0V2h+PQWGEArYK670UFLjX2TIi7pPMoiGq9LtP2ZmoFolBr/pJ9
uS5n/E+Id5P+puK4YU+RUNUlXvbCmg/L32Ol9Xm7lXhgsiUDB/UxBlviyf5iDF3f
R4J6SNXDv1K187KxIoKIkfJYhJB+h/C0bGTvZALIfOSXuY/rPizPfSre3MrSOisN
WYf0EEBRZwxYNwcBssbDDt34oYI4HN2No8oYGu0Z5+8has90fpqCHysx0Y7F8bfB
ztGzFidtFWqoewXa+Vrl8cm8W8bVxUFnFtyhDbel0gkNLvJoGFaomhrqzVInL0Qk
xsYfSUSxjdnzKWlh6WFDtNfRc/LUnDl5JlIp4QszFly6Zz3A0l9omDfyElklOIRa
XZuqUobarG3L2vaM1piSaNmvErvBZyprAnQNtvYERxma/MInBJoK6b9Xrbbs+/Kj
A1ChhPLibVT+WftHFEF5VzNftlzqvnP1dD2tMZy2ymxNnsc/UfwTDKMgoTeBAyaw
1iaHfsZTfPe30O1hEyT9MT6IM0gg3xfLnKyQw9997wvGM9sWMPaMwg2s/eWa4SeN
kGFQInWWRrfx+bdy1cU3qrVdqGVwvCFYJ34aO3Wwua5JMmuzWSEHZqRyuivJS5+X
4Ikro8YGnvWfOVcz8XVTnD9XmfnXRa50VhBoJ2z7k3BAhixwstbZjwENvaIx7Oa1
qCw3oUC6ipEAngvwNXskmO0ykozDsFpW5J+UmJC+RLKc8oHUCLlGx5olV5AHyqJl
8M5GuLyi2Ii5roxBdkHWt9zYdH+yqtZMuNIiRflnMQGAk33lHAbaBSfc/0CdRzb9
SbkflGSCmMmxtsm36VgryVlTFQUH+g/vrnqIiM5cOdZPbAUjwe92AC5/dHCazzEo
759RLPuDi4jAIg6n2eCS//KfyPfNrywtrvHCeflP+A5mLAAb/Md82hxLSSsHQISN
/ghyHhdz1cpDtSL3A1kIzjHAb4A15bB+e8LaUAdW/P15yj4CJS8/lN2koqlV8X9Y
dv6ZFFjCcjaNDZiDhuFM/eHUsiezkJuS6PS3a1VLcc4w7ba3def3yBThc1SuQ855
ynwkNGMPIkao0niwjOxQsNISTV3b0TfqnJzCDA1AjW3wqCcYv2jWoJ7q8VukFJi+
bQubrJXE7g58nVQz7ZX0/hFS3fG925K/rm+7+4CA6mLV47hj8my20hLmnD27yDSV
oLT7nUBJB7kr8aHHvx+VeKZCqwdv5MaXhzv30a666/JV9sEo27q6GGPWy95QZVqK
pKbBEvtw5E7cMRUPsOlqwyJcmmw469DWnCagpwO8vkZROTjMOVsS03Tnty/xO0zM
Uvac/1ODNhsV4VEglFI2vEVdnrdlGNMB75MD9lcE7kvoTWa9A6dS3Q6Qy8ujzof+
2dKpSOCtpCm7i1I/YECA+n6ZUlBHpbFSz2HbQ8tqsONit+Fivqu8wXsdZRV7+PVR
9K0j+o313ZX6WXbcenC8pzKeLlEL+B68yDiab0TE4lfKr5J4iupZgfQbtZNgB1eP
bH6JuyjVFSEmaLN3ETMker8VBzlN8hD4nfol0h1rrQkIbT+KnQRVrw5+VkDGb5SG
MvefaTeqtxVsSuC1xRrey6KgJwUUnRuA4W2ewtPHfH8uDG1gABThrBzKguly/8dg
7AB/KchBJiLWfq5U9OlsOsgYSMhqPKxSfMpQSfZoI/1U4ZTWrwioqmu++hGMC+DL
59r9PvrA74lV/ZTJEemz62T7P83rdcI8A62K3ev6q6rxrwlg2DRiGMDCOle4L/pm
7I0hqOryDAyQ98+7WcvmLYq1IJQsLUzKKBG6tPidd09AebDDshsreQfH2yjVt/GY
zLDOb3m2efE24ecS5TB+Np+gbfwcc1drnPqKxDkRJnoJbwnnLIR8EOD34EoiaffK
GyMuFDW2iXkNsL3i+ihCkyZA+DixSfF3Gq6O9jD6i3a0xZ9B0M3j3fCeBBkqAt85
gDaDENAZDykwiis2YgAaD10qnNy+zyJzN1QP1w7xAHflBgB/lYmvyp/pl0iyRj9G
MZ8hnxtW9/NzlytekAbRN8PV+Z2I35ccyuBDI+PtQazpHFHxKy2+hZqyZ87Nvzwk
y3qc9c7IBjAcChTiajs8GiDq7sBOEERsxUIKn0t8GcgI5+gpEzcOrrn6dmiVzQAD
8+YuvRCNz82Fbj4OgQcQVlQbn5ZsQK0cRdOPk66R6EdYqtyLg1bja1nsu5C7SAtc
Bqp5XPOPsEMBOEOvGGh4D6npCaZSg+cElHBRO5p25nt7lsVzVoDX+WZqEeVXTyRZ
niIlMxR2YhPbbPwkSZJvLT5daS7Uqg8cG3L8+o8y1Yevn8L0qdDv6cXNAycc6I4U
QNtS8xUxmLMKk67V0bupkLqa4hWsVPJEWEUNYVOEf8/xQ2vkEq82e8Rc2/Tq5Kr7
kf6tR3cD16uLkFVVXFTfa4eS6a4JhZuKOBuXfO2DFovBPFWMpUvx3qlwnh1DWVJM
MpwSAJMBljxhbZd0bQq2WKe5i56UonLfiTUw97kVDEMS8hbLzwMQbH8/LeS7PXF6
8PRK6+4/qfbinKDtdg7W6QSJzsFCuNiTQjYQNr4cQ7y8mBjIU1zZP7IIUbGKkcLq
Mo8925XUOIZNSnFZbHUb1+MZVIvhOtGGFuer3VRUv3hGeHPnMfx5536sbQ+8NCUq
WQ1z/YywGI3B527nkg8IGcOG5T95m8Go/8I41tzn8DzRwjxooxCUpVAyjlWX+sO1
xJgPyK1qSd5sRZfQQxBdJ/U5Ab0aA0x/HiD2VAgpU45p3BIKaEQicMTlOwFVAqy9
VgCjOt0YoKgKJ9AqP+fHg8vTh3iMfHCBLVsOBPAxAXj89MOEJotgFWUUHQ3BFyZb
XAco9FHFFJf++01oDf/jD8ZRh/S+WgHESdWt6XyQBt4X1X+PTnTT9qyE9Oi2412j
d7PlMTQWs7W6TTGNwzuxEshik4r66rY/IOB7PfkG8O+B4FqbECTE9tMMuS3K1ysI
RrHxzc/4PHvJB+KKt6KyFgADvlmOYmDz0GVz6LqWrxc9czkvcW0dhwfcX0s8Ha1t
813UgE4E9h78+WxB6FQ7gG0qO/VIeu8MpuWKkYrhNf8lY5gPHx7n0sHJPvZLLE3W
hicQV8pMm7hXPP1ZCsKgAJHv+UhD2gn1SsqzFvyIjc20zfg4zSsR8E3mswLAjjTA
DmFpCXzifwAZtVjh4kWQffCM7MZAY3ZdwbE8md/WzatNEkQ4q3pj83nzQTHqDSTv
qWOowhm4oIyIJc5E+8M+VEq1dpU0H4s1bHLSMGzNsNE5cZyB1XiYv7YN0saBK6zF
E4CChT2HCCRQy+7IG6ils4OsrybBhssmwbOHJgpx71Y6dj3yEYa6IkidhcYfagMR
qkQzv1UihhMrZbi/fCGrm9c9ieonZI0fWL7cfMRLzu1Dl+zd1ab7WOY7x8PHJmDI
BTEs73ww4O0jujqBT4VjmL8PyKlZTX6PWhHg3KNM7NV9yY+p7WUK5BqOSCvvKb7N
fwbILndOZwTx6+5IXUU7o8Foqz/SxJCCwU1xJefIkls2unALhrDFNn9W81KdH/RR
QNu/cQ2hJ08tTYaUkTbOsjadeoJ75HQOArt9dhGzNFITgCimI0+vHTyCRnZEkPsi
a/4CLARb4oseos3BVairTO1FNfE7Snido7aQsTnX5FaZZV4uPCAT9PUiNbratXcZ
WcSHerI1ceNtmtHAbRSmfXBq9nDuTH7qGey7vALzA2JPK7xusv6KTLFE5db04kUy
PxStOepxCLmrmO164l8jhj5kvHEuzXqaWaZETVMagc7S7fiko/3e7x8MuTUxXs9s
QDOBvcz16u6z14RZfqk5fD0fDrmhuSsY1rqkGW/avxlSDcOggMjvVE8ekS8tNznL
bBFJWcAB2FUR689gqbYn3Pc7V/9BZP6aPxfi5Qom1BaQfrRsWOhRygV+rMSTlhip
5h6YxJKmudCj4Q0l5Cb5wr2/HvKeCAsv2z1ssZFS1vwOoEY61ErZOsDBnfx99jTw
/vE0zmPJ+5ja+8a9vLhlbuBNzO9G5L7t3gM2Gqm9Mx1V2ezWCyo5A9FdNipcVtQt
8aoCsFa2VGeFG6oevVQ9fqbNabGuGnIv0EU0/V3t023QYMYjgogpbxCUyT8XRkq4
zCmZRMK1krLtcIZMkFVAw12cJie7+M1jQhSxgFflz6bWftiJbcb4Q/MQ564ft0CM
Rk8AuRsuFCL9n8dPVz3XMbPpC+kD32zm2x7gdoKOB1LWYl+/MFm35xEIEdgSZL2h
wWzlW0vU/6podSJaOn95oQKioxM5RoMk/y4WAKHRdrwowg29Pk6dcXJnawsXGdJG
oOM6658cKh1Y4zv7nKOOWAG4LfoMr4xiZ7f/ac5EdL8lFBev+sZ/k7RgIBQBN/Qd
NDdp+9giheLXv4mpuIlTp4Evb1978KygJkUAPxhJqG0bF/cWvlqPd9/TNb/YT/oS
8jvQURu7dx9sziMytn7Yb92VDW9FJNv+u+ATMN+61fmNXaJAqVaMngRyWBhQuEsK
sm2DgQPbpWUvmuE9IXKTuIZ3INAK16AjNmh8YftWWanJvs00Lx2PopnReHGf/4QJ
jZjd9YMwkwYirzta2gLtcISQD8Zae0vUUFJcov5hma3qYxjtW98n7ZKwCYVNJNlQ
RzHi18WiTMJIwfrWJXOwYxvyoc/ROHrRt635ooLfzhbKU4k0OEDzX8CHXEE6PCAP
B7R8w229DuIlZt5WlEyVcR1633N3iobEQPE6IMbbjV1nZtneaOEpi6byr+lT5KzH
58FHADlip7tPGPVpt1bYhN/Y2pDNWRjRYj+GJ4YkSnspLzxrC8DsAsWcIkvcukXi
mPufxAhH9ppiGr6IigsNZKf+NiAiMro3Na0BGCDuE1I4Vq8gxvqF31r6Dx0X3y/9
mOVmtgli+ugwa8uy3IbQzdBv+rdYA6e1fT87uQA7kkqT1DTXUHtV9EwR/C98GMTh
0j8rLT2z2Mg/dVTLBphZ9wxRIqcW0pJRtgC2vkup4+v/LdAfe807VNfgua5f6hCy
qCH+Z3Ttevs0D/FMkHaVXMD5+SC597ppnYJwKmQjB21q349tdvWtWgTGfQEGdVkM
VNZbb0HpkryScqADehoLQosV7L4gi87FGy4/fTZTbrWIrIWEuv+gybN9QwAdkhMJ
ewHGxnBea2RrzxJvyRhM2xRXvhRd7+OJC9dIZSQ58yJfrd/sLzrM03Cml+JGmzId
a4paiaSG++NS6Jia1YcZB3oD8YYTSUhSAy5fMg2rG0GXmRoLcYDtwpEHy0VNKger
PyDPL3rigX+KBVBZV6CtCVeh4gclPz0G3AQfrL8yai7KJuAOC754AG+yAu0fTVOD
ZouEbuKFx1oL48bbipjqoS5YPQbfXuscWuZQy0duymviG32xDHN2bcx4An7m6GBk
CMN+cr0rPIV41Vrv2wOhQsPO8VYsfbVGq7U9/vKTTLym1Xy0iCP4dY+NrPYTlxeG
LPF+wWBRk2kb4BPUQdCy1zNN7ge4xG/5/rtNLd+Oe9tc3uCjAp4a5ovaFVeFkUCH
uyxR679PAouGGRbAGbflZtiftTnFe07IwI29siSL9Xl9xfkrAP1D0GzjdasnAHyq
vbMw5y2wUWc/6wuOEpZaQv1EK/eB4bmMn5Edab4gj66D5FPgAargq0nBOx7XHVgl
KFzTArLB4IdPHAOu1QlNPgTL7Cqp6uc0QEqw2jH8KFrLzWGW2KVirkQkipN8tPd4
Plg49l0l7O8MeHForKFirjHpX8s+k+Hbd57cafg3xUh2VpP/8HtIFoHvBiS99239
MXaXnsmNdVyi7AL97QSSz3o2H1nu1x6hAJR19r6WFGP9JzWIHA+tmajDJ+BABacE
JOKBnLFySyNJjI281rpvcRlA6fHx2tiR7Wzvi92MmcvaSOWJNjtDMTuxklOwHlHO
1quIRPA/sAOWyAg5e4gUoFAfv8w01sLQKre62kZhjIJ8gS2GzW6FwC3WbWKCGgC9
7lOlI2tFeaGilQSd65xLr7lQkQGYVrLzyiOKxRQJE+WKAMICMhxwAZOCAN6xjWC1
XTtZUnGGPmSrdUoIsPlWjz47nWeZ94+fvsykhJzTHw2UKMLklnKnz+1a7wLS4Xoa
7bsRXis8VfAW7abiphDGDeO2b5BJrGknOhMDxWyj/y5iq3c+TOTeO+jtQ2kuIXEC
6P8V+Rq60AGSqjzdXxvqIBDElC1tF4MGGHa8iTrygju2+0Uvg3d0FJ2yLPa5TENe
VEC3wQJmYNgsTEHmDmNUSwbG2N/ZHK7x91jgDcAtep1+qhYPYikK9nfzDywwETzT
yuT2JRk993WFDDIiUMil359NOJKDtKnkjSyaGB+kzp4CzoIAjjsBvokVPk1MK72T
uT+1Yg6EOIrW29rAUpoj7bt/WOi2+Ymb86LFfxnWE8QID5YjkDutl1VuAqyUheJB
H090zrlih6paE3GfI6jMOagWbHZDP0xn10KPW5gHR1DhGZnrfrEEspEnAzApptbA
dZuhL3C84YAYr8WtCCyt1YePQieampVAnuWZWqdWJECaXELN2rD14AIr0WreGL+0
UzSth+VWD6xK6+ZqOB5kvwZFANWj9GFUWAJuQjKknDaz6xvqsISb+OlAC+eC7lJy
Jc5+tRD4eMj/u/ZtTq814TlI6/mw+99irL6jJ6qXgeFXsQNp88jzqvkGrZatUTiV
S7JqcxNuIopSdh/M3Oo6AXYiTY8oyC2vXsMlcQPTTxJtDn+Ie88ooXdxW5rjC2FI
cp2vKsyxTaUVuDClDlUbTkwHrmkWbo8SuTDKraRC1D5aLhfrmHHPTTueEiGrV2/0
AN82ZNYJGN3Rca09aMUHXk2Q21IE7fO+fmJ5Ks0MWA8MBUDDHCjIeMJdQDDeET0q
68DAu8353jiB4/KUjo9mku1OHbDBX2Exk+25DMmtR/7wsmy0iCIbk0kinMkXYjzo
EZpkhGZU0UZRAFtQ2Dm3c0v+PZq84qFeeYWPeEg/FdBwLJDs7rfvFtUU4rc985FB
IUFIlHCQABwFP8j1KLuk6AjLCLyCWPtLaMleQtZcDm7rdv0HqWJUveAytSjL4iDb
Xvgvh+nRS7+Ht4qtJ6yVS545diRsfNR5P/aqwyRZpb5fK3vaNa67b3bJwe6exLyL
WFQFAyNivQOy9YpTBbZoW+PpRnlGGSYmRxvS6zvZOJb8vv8T8W2utjCwBRLNnD86
YoZenSsK2/w2k41bXLEt9Dmc6q1yoBkV+EFxTH7UpttbnGnnj+2c+Nz+z02ggXUX
Gqp+P3BjkBV2sntFBCTHuzFNO1Mm1tA2EVFXm3FA+n0NO1d5P/xgCL5YKSULrZZh
NfT2dp+TdNHjtIp/KeLUq+3nIgTDNmL1tN5UPKtFcpipSJ5GUo06hSlRhggoSpjJ
nJLl1045rCV8n4hCtbkjfFSt59o9QSPgUFNHWJQjKcFJg/DA3cj4+m24J1STEucG
y3f+6otBlJdz2qi5E1CH13jV997ML1POOBAI2XJnAPjYIHn20BRUokxaVmxZvkx6
WtD8SA8UX/MK3I/ilkaCDGIdwHXHqin3XkhlGzPpjRrHRsfb9GxyAn+y6kMSSAFd
g0TdI6aOa7362iocCHGNe1THGBzqXjdx2ydUIVENmQkxJtQblCix6joQ/hA+jGaz
dhf4CykzRsWmYGH0uEVCcHXlexbHrE1NE/hww0qao0VpAGeEwm7ifQuna4heUAsN
LEbHvWx5Ux0KxINJRBRJlSfMdc1tjQFVjSOR37060LoPsON8Ic4px2KirBQ9VNBq
UgQy9G4x/qvEjU3aVRjDFy2qAya+EtjQGUvIjH+eNZm1ObLJwKmn5yz0NohDGWZD
BawwNDSmgMya2ie3S1qGbJ8R+4UICC8+6dADhcX1T9/URtOai2fVDD4DP1f1v5cK
uF8kfKZqr8nLzHbuuWODRjRCnRI0oNlkBRqEIl9X7b093SW0OBJ/OerpWWteKv6W
Zb8MbWNrpz4aYXUn2y1cVAyIZ8cylYRAuUVNK3fahXF/FTwXUkZQA1gi4ifoh1P+
/WvDu70lrggA5vSAfpOlsizvphy7/44D/xxGNfnpyhJno1e7WidBfSf8ZmnZF21R
a9eskq7edyDCia50SoCSAzFyadxAzp2OdkQMaxW/HNEOd2kDQbveh/Yw1rrgrjFK
7TtenmdnQaVbTGpx7aKcOV4gJWzBpU0EpMkkl/pUeslHyFT5wy+GqThUzrxGybku
yJGzByzUvQbAjH7qFfivguweLbndwJYn0Kaw+LIaw7fLRiGBTnozVa3Xu3/SHq3j
QRQsTpN4YI0RSbYjFvGl9xrW61HMfE0gxGfOQcZBEispDGMpy/IZJBoHw5qjQZit
cfIoW1Sgp312GQmz1a89nPbzc7ZswX0HwptCSYnIPZhKEKCPLTJmVl+MJY8xo97v
R0gAkU5pGFbM9eLKuoubnALtLYeEonTx/Ivu9FBoSz60UwXSr/vN3aCW1Sq1y93+
phZjeTdDUUszZi6bcM4hKKBApGGT9yQWBdFHm/ynn7k9p8r3S7NWyKdlzhHL6uDh
JFk24u6TJ/rybzJfksnLGdWnLEKpH6dUz75IqSnEGqKuub2fcv3wvwQsWfwSXtya
YIUS2TfNHAut0pqKJ9ShGpowgl7akeX9j8j6yuS743jS9p8IV4+ZikPMlu7HIvWI
CuPe+XpL4k2zBBxdgXY8GFOPbbWJI2NhmmPHsTn02zvtBlZfwkfRHYPV19C/wHjj
GJCkk7MEVh73ukOZWle1ctzo/JtLR8h2/gVcVJx2djS3VgyCL5mb+HrD8Gw0Jfht
KVKAUn7H4791WfE1QNBwBIeNj9KYsTI8ea5K8NhMDFIE9Ldts+Vstx8ZJLWeWTlu
zvVx0Cn1McEMUqTUaidaiiXDwECtYC8GworsvcnTWjuCD7vm36Ar7Ey1/jDQpc2u
K4RacHxceBieRBGdmOBy9uuYOfJU39tHKYpGG3MwZvGEIcuI16o0LAeoadf4dUvZ
YYZrFWBBaCZyuXBxrTaMu6eoNgqVSMiJBmsvA0oA0rh/w3eOPv6M6zQ+QWEKKOct
dSzUujys20Yu05z8w1uhI4Lh0AyYbf+NZ3Qc3rUZlxk3eT1mvT0CR/hueO2c8tGl
KuwMXS4stR0P4GljTjJJmLbz0mz6YZeN+kYgvcypYDIzlL2RsapWY/jHhgAsQqdD
yyVl+DvPSeWIA8ib/4dW/agDyQtTRL4u5VST/Yzo/wR5GQTDHtAS+YrZPlz2WuJC
/exOJhMfsPkujfQ8E6XTXTeAELw6AQ45kvUAj4hiaT5dFX1evSI4uSXbSL7bECd+
zVJUa+f0pvs0b6j1n2i+x9f/RK+p7ymOxd+jzElyIgK+qrgBTu8IVLLyqXAHzCQS
YdLx54lx8JctduNwbDl5iQFe8tOK/D61NbdhTsTrlbYb2tsxSoTYaTTP9HmpC1PU
9k02XF0YNBM4kovhMZKJddebgXs8qLs4WwJ77xpLSUnzTDAWpbt3WB5d2LB5j4Kx
tqIEnMNiG/Yz7E9hcEyW262IS8U99q6HU5kx+1s3KeiZRjEkzAH3XHwr+5VfIPC6
FlDC2VnzjiH0EHjAuZ2lUNcEJd52CcSVelUOy/GXksw0dctGln4tHQ+3trQ/YFhb
XQVb9lmHPYsKBTKGx52EWf1pKWzN1pMKGFNAxnNWtGGwIiWUlJ9sor2iSTgHb6+5
4EerEIrXSdwjmw/7tm0ceGh+w0Oqp+XXOz/l9fzJ3grtibtXqWkSCloEueEzJ1C1
iJGhncawcnp5T1ALFrbuE0NDuYbHRIArX2QQYf1eZ0R6feXWJCuHRPLrp4+rdH5b
AaggwA9fFRY/hdvnNcTc8/cGHPKWbYSVFbVc/HmOVZE70Pp3cv2azTzHUeVLQABD
411JPagUnTDFJxdwerya4lKKR+Y0H9g5WgLINgHksL25EXl6F7Kbkh0OWeq5iKpV
Wj9PiOX8Nsp35z3GD4A/UA8j1nda2wMC7ivEemuzwQim8AuXAD+3PM4cSDkwoUoc
4+CuSY/v97x7zCZt09pCWH4aj+xGIOLSkuh+cdRPIIpBq0gnJ7DzLAAwv0e+QTWB
Is8UGDXq6ok/R8UBdUw+RgQ2PtEMIigMbJlN01oKPB8j5g5DcI1ClAVtWOaFieUj
oOrgoAeElmzIZFdr0hiMf87fR+Z1+XCmXHyOoOH5qS9VOcX/YP2v8jqBSG3eakKr
kqwtap/IEkESuUA/Yls8+/bI76R698cCesJ8Wo/mToV0hpEDkRXORWnZ2QKu9xGC
//HYSW1pbyI+PBv5gCWTiDPLiRKdAfD3Sy0rqkxHxf1SfoH07DlmVO1kSOIequ+T
SBoolxSgP1M0z6KZWiYmDg1XtJ+E31sAyLwLBd3myZ9hUYLqw5uBpwAuqJAnXpQO
/7wP3xQoQDHHUt1LLFejPHNDFbIBp8gM5+pGWjDUTrwjrY017pQUpH+XEXzzUGvA
ZLxbo1Nl8DcDc0+BuV6Qxq3wHE+XeZe2qFJ6AA5gVHIh2/8DyfE7avpkrijM3ZNA
ZwTQ3bOvi5DBsM6Xrk+mG8yjwxbQG8Hn/uNB6nLBTxtFgp1s+Nloz4QVpdETXzi9
VUP046IMCFCJx29yvPcGIy0WilNlad7SylnOVf2xJ12r/8ib68Rrqsarc6PyFZZt
ZViO9XxsN6pfIm6UsRyBGU6ub6iud4YIv+gIz5UP3EIJ0FaehV/AZvi1BHRvnKxE
Jhafo2iPgr9do9KSSrmvfBoDlw5XRmKiRSWJKuxZq2Viw/RLbmkpJEpxCFqSKjRj
WQi2OhFo+IpbvzFk+E2PdyH6gRgkDpKHmD58fDM3XtBsoTrJ/MuxDiV52M6Ccnvi
kS49m+1nrgqmRncaUqls/bKGwfMV/msGlSQIivWyOJ3qSGDHLC/lXqiE+ZrBDWJf
3wgRoM2DxqH5Q+4pr7BvShUaEgQFaElz+ba++Rut10/rXWNxZJ9pxKrS5JBpjr62
UBtjcgS3K+4Kr91nUKphhNzCrvrVfBoiGZpII2105dQiCPlg1WEKqpCmSAs0eB+P
1+5l2zumjkENRK2Xu9af1q29q+QBHAZ3+OweSppTrPeCfIe0uVd0CqG+naUtLO4L
ftiE/1VonuLafr0NsdNj3wxuZy8eLrGKDyjZj0Dy6lNZ6uCUIseeTRJagdjdpRcD
0y4KMqZVYgdnPXVrJpiekqKqiW1bG5f9lyAjGSKDoF8NknBlBl/myKLBJXBkHj4K
CZ9VA29X/7xJRyiD2Fuvb7DYNRM7MVTpfIJ+JMi7rHW/IvjaxvNBL3rzLsPTaoV1
fcjnqG7Kdir4dV4sf23qcF3WyZ+RpYgG18UXnHKeHioubNutMTJ5u7zyxVfPC91x
z6VY6IafJNuDYTVm22Hzt9UBT0sKSyX1Il7K4emJ7Kw3F3V/XHjj94xoJDfk79+c
8GP24FbgVal5dIZVenIPxGYXAuceMcJmGgYBvwxm1ljk40YLCCaCiuQ4RMqNyi6c
ONjefZQNlIXM4IHW0cT0oz/YgwUoBxWx0p5C9z9/v/CtN+nChXQcspl0t5iXog/P
TifOUq+umAehumsJeoTK4Ahig0le5cZ8SVLYgAaofT2UDjPs3G1/lgFv2KsDzkjZ
yX//bID1pBAi2cQnUPXHBHNfokYHyWc8HD/5MN58YEJKPhMAg/BkRsDPUo3Ojblc
OwRmb6DgvPAJKOAzDusAzqZ7CTlGZP1YxkRXdjOeYzUJ1kzWZMVkiD7QTfzPCYn8
pN5u2nUvcPCjjgtcSgv5TMnXAnHIaWKGbqZ63R46UZ6n9ZelFf7Fs9/PuglSVbMy
5knHMguAUG15T7CMwBgsFTdZPBn9HdJZFSTC3iEaio1IfZUeB92fVnSkb4RCXjxX
yBQ43dIr/69Oge4oqgu6dbGigQjfyswJ/kCPbckrK43zM3Pkp+YFwJevEv7x0MfX
1NF+OnD1wg12Nf3jzU7T++HQymG1tIooOVUsNIAoGle6WuCZZ5E0LHFVB0hxvx8h
yHL8Tbln61dXQWTu0MVxkfNIAE3ABjvQPKqrhQ9n+KWVj1WqQ6y+V0jH8+oLf048
lekuojFPTs9SRmOSMUjqiAtPIrO1iW7HGCLJuzhbq+tfsWd/iUzkTQpzehcUMm0J
m4AodkLSp3BL8a8FBxLpHsoSAZNP69bSHeyC4J0xvnsDR0mATvAqW/D1aIVNh5N1
pr5c1Hms5PH9RUMBSLJfX3iJo/Grq+fCClwYF08r5dAVGO/lWT4K7BnHafqqcPE0
/SpvHwUUwjmBCuPqTroeJkWML9nnZKFdu/4DhnHeAbgFCfwgoOGOavUFnKJUs9rA
r/RRJF1WOv5N2LMTXP97m3zP4HSQvxxPBJib6bqGccICb6YC1Sbr9IU9SY+we4jO
/jUBsLI2dsZBNOq4EeRfnEXMcZrGtWVfxLgEyCD3+/5fO/VKXoTFsmzsPee/fP9u
DbssaumrogVqv0jdDImeJzuSdZZhcudPkeJrdko2SXkbc7mEa8B1mN7FbF5oYe5f
M8cLVK7KKLN5v1mmIRuAAJHGHMVLTc2JQ91DYBGQZmtOeW8vvUCD9rzwOG0+a8t2
qAKGkHKApBynG9gZoaqdMkSoExa2RpxgTbR9ZLQraWIgNn/Gbkwksqk3Ab/vmyEi
VqPVJFL5z06fTzRVdwfqueG/YIuWKcPUf72ajnYVSnn8VhOMaK75vr+GkRv2czwA
KL2DIMxzGNBUeHzG/tquOubtFFXXP4Om73CZfnhyEFZw4zggX9JScIbal1kGuHnX
d9bilb9JnbEQE09QJoOcstXTEF/kERrtKUltcfeaVf7rTCTCdB48mO2l64QFiRm+
ASLv5BV3cW1l0nAWKq0Z9XAr7usTbpTXZbQ30TLVo5m+SLOnsW8op5LlYWwkIdNC
UicBfT94oXlGKOhrPNI3b9Qe+lPhA/R3Jl/9TZrcKNWX2C0qPKruZVgaKqPyw1h6
zIHSMLQP5Pem+CFLZRO1u1an3GlV1mST179l3a0ZjeoXplI7sszAp1UzcrIcfP2S
bvw+8vWcFf4DozbKiVubQT9DggjLB1ickVd38whSsCnF9KzlC6oB57maUK4oC2x5
KVPwqvwc09aRxKJsNjzg40JgMZd0hgnIhsRLvLn9sHSM0oHQk0p/vxRzm66CUR0y
BBNZAi3YTHlXI9vVSCsg/LVguc6pqO/CeFENHnPvyOvP4D9WiRJ/CA/aFOVH3r6U
OHgiDWmtfISYOheRfDWONNEuCbQiU+RjSblgAaLU+N8z+Y37bnDYZvi5kUEQY4RA
ZVBzy99LXuvGNixysiXX5h0mh1YhkNtQE2XwmGwDKAgpt1ZFPQ0J73Mr8cLJm49X
KWcHGuyu+4WwA6drco87gknOkTQr0ey1jzSJ0+Dck1rz5H9BU8WTmhWur328Qa41
aaAY5GKeu/HYxTePW2GzzS1I2qRhXEVEVBTvLT6stbmLenqojvitVF52JwrGf+Z/
1smTsH4phF40hcbcQOb/qQ5HzLL614Qka1M//rcECHk7EX9tQmcBYOeJIt4FYeFY
kQbZIHa/IgRZPi26U6QWq7GntSE2tG9ua13wF3HL24Fw0zBHs1agrDNoLlpOf/Wa
jI/vccY6ZliMcP6uKUvrGUJnlSthLGFMZUGoCfFlzLSbFz3lovRYTL9svcQphJ49
NWRhBkjq3FiJjFFGa+Pz4JJ3IN/vIBVnZdSHc42sxuLD/0Ljzfd29uION6x1+xv8
aAOLO/wvY6oWhr5+KVdUUo7ZvbJV+XiLRnxRp3aE8hFHYtpG81hfjn3oijFS6b6w
50Dt2odYFrpIw4tiaJfYLLiyrMc4wQxOV2C6BViGFhopq0+t/+jyBxNtD8ICsj/M
+bLHLJKVAxuNp/4GUDJ6MQTlAAJ2+GxhCAle2V3ixiv5MwrG676cAiRrDmMEPbxa
hs+CcTKRJEckgnWGOlRQm5diiqBSAmuA4s5K9Ilqx05/cErNk96i/jkSccCSLCAG
0+7uDTdwQ/IwYrEFdIf0KaCOyWK6oqdcqxNdlEwuEbWIdY8psUNTdvq/KABEDeWv
Z64MeaksG0HBi5xlrd1eTXbREcbNwbJCvJFdQi+aAlQ1TP9KqPabIidzRCsbVFC+
wI2ultq/Mpzf7cFW/EFaX55BGW7ukBAqliL5G6oO4BSOlcL5ID43E1c52nySNrrP
ir7t0Q+v4AkIb+a/r0MnEq0/q8PrpvbsCqpma0ZcrODx7gdwC/MIHklClvng5rrT
LuAA5nMpUCxwe4qdptBTdXdpCfBIEjYdSzFNLvjLaub+UbAgfwjS4G9xBa/bnG9K
BdDg3ilhO5+zFo7MYNVI7gPb2lVNS/BsugjTamETbsfJoI0hlofzXLELQ86YyvAA
LUXkS2g7tfRSmNQu+mr4Jn4tQRBHDYAN1+J2KcKuJ+YaqFRn+2dNh5ONnFpjiGAg
yhlhddAFfUJtiiDFyX9pBNAywbJVLla8HxtNVXSFgGOZ7waxpdLEfuNzy4vU0MX+
mlnQF/pR7DAv9tiM8vPNEOKtinQDXTXPqRGPsKussKnaMuojxAiJJ2t8xCUqpIw/
MKTM8PjiOlz4zFvkzwhzgBMd3EUt6gnQHs6m7XuHxJODHLT5ksCsDxXoSNCT8tN9
1K4VZv0mYs5fjvOY7Dv8TO6mzsRhdXkGBj/X+lraNQUN3AsHuyd3o5xzkX4AMdLT
3Gnc7fTYPSaoGM5aNvmz9NBqiBwXGYuztVFl+cx8p0H9m2NYs/CLN3pH4+n8DETz
Ncy3T3g3scAW7G2v4VbyWASYUXGkF5hPOy5sN8EugqDbaQxz9LjkdU719rzyxpbx
9T/0nKeIO1rJca0DB6qyspHd1GvjbkSfPCllZISt242MVva2uNqqxyWrlFxJwJI0
ljc5WxPxFgMZe5FrEHQn4DdtQFZJg0SJxG/UpD316qxmVYYKQWxc8wru9ejWjC2+
VVU/OJg8KxExhp0QekQ8m8aA6QPuJc3Yla8/SpjndvVMHfpck9SDHoufGwH56VWq
U+1qip/dDVwktGAFhXuIjltkmAi+tGOp/X5et5j9iZoGHA9upWamKW8IX3mnFAbW
SdALjsReQms3RkaWt9JQlRcQrdjsEOZb7VW90eJtWLmzIaaq7z3v1EcmCiWk9MM0
0hhg4yD2JrrTZ0AeEHKXJNcP8eO8rm1UK3r0IvoPHDb3g2fiGE+L0NIQNnRDIPQc
SfeQusbao2xR7ttPW24hQRAGMN8MTOYWy9qaRH+Uabu5Bqh4wag8CDQcffQGsXW8
ioGwx0wrtxDzWKIvXQQ5Z+o2w4KSJTmfrDpQnDCNQBAOmFpEOq53Pc/0LDUBYsGd
CI50gdc8cuaXAH3dg5+OMvo8mjCpSwJYPALuoo8lR8l49hihtPqnvkNbRBGZrAAu
axpcw7flzMSQ0Xc6NYVuUHfUerPpYhD5Huhr5cFG0Tn0K4UdvQACM6bFNTgALo5U
HKOlH3+TW5Bb81xzvNgOhAk7AaRe0lrOW0GJrrfDF6aPZR8V/2znxtTv9l1WfOR+
5JOvvU29+hPRpUVxeTF/AKRzTNvOk58IrG9g8DxMyjQsAciJKNcq8MVN8Siuwfpy
/h7DMQE1PuiYtmEy/7NiSZHPid72WBFxsOI6kpdS2pHsBCxsySg8ivyGTxMogtpJ
8RV56H4Rgz8TfexPdxxvg7gINui8pGtg/1nCCR6MO9grOG9ZsaUqrv8jrtqRqqRD
kyYbqqOSS0dWp+NmiN2q+40WYeIuHb0fOS85a6OeRk63efACSkO0hfbJ5MmMdgK4
P744XpF79LR6DzBcTp19cMPbZq64sZhZLgIlXmzysQzIv6DLARltW+gyBSuw4nc7
Q5NpxLi+ASTEc8oYZJs2w/QpdGR+u84JvvPTRolgv4xd2//eUOO92fxvoJrf3iIl
7wTRmFBgpBBXPE3FlrFFh9U5uYiuL21EvlSSlub5ie9F3irnuXpcJ7coPNVReiIq
2yc4huHK6bt8f2oajfdom2c3NNe7CrSSIFUFsziOkPvB9bAOPq29pPUnGjHecnl0
i0DlldfdiArQs33Y9sBeH2sP2/V7UfLxIiogZjgfCLa7iYU/If5MnUlAhcvymhw/
SRTkHTMyLRwNQvioe9zg7mV7aEJN9MPKQFhpXE6fph3+W0Jec0utujd7vDi0q2iR
J32eawTtJZ6DLZ18wpqmgM3vl1su8AGDBYp5sRYmk+L4xpgw0BTfWD7F9fdRg9W5
gQbcM1JfKbjxzwyCbvpDU5yXm2jJaAVG9qfSJjvu+T6jihpFUvUtzELyVgxlKkpt
MmI5NXhIEtNEgs4ReSC9NEBYD8Cw4UzSwD2Fh0cB0HZzES2405Ydwf2BKbya3Yvr
wX2B6s0E8SYeJE1gB9PogFzWgNaUxp8UQqwyt+Gfuu7mqp7xPdk18vGbGZKegCg7
FuzcVSypp0ORsikNmeEBjbvZh9tWgR2r83rdu/5dkAmdyYEfxqHsbFW/I1BrYJ/A
Emwp9OWfkmEKWYcnajtytRzLCv2wI5oy+6HAGcolUV6/wXV8OWDtGb4Xyz176Icz
AJnofAK8aj0bn0q4A9Hvr6UfbVaCA9MFtYuLvUVy0jMpYLIZ5Jw3jrTqwFbkUfCI
LccghhqIy/UK6zAOrCSLXsHNxrFFCb1INF10z8D2o3oIlk1mOWMRBbu3jgCjcnLw
gSaHqAe7oX++fTsGkSBw6CkMutAqImlPdm/7rMjPDa8L67VzfX5agdmEYLEJGsIc
en4dp13m/BaKtI/u2h9DcBC0ezoYCR3wNXTPlY9aPI0N+5n/gzWEFioBaFCmIm1W
N0vIMWqsup/myreQa17Kz18+gA31eXSQIsB6Vwy7V6XfH9vEhYXFpJskvllkG/6U
0LVRT3XLhJ4wieBHs+VV80nO8wv7OgsCE5lyH1VnKRs3jQLzd5nliBqtwOylNEiE
hhsW1//Zd8pv7dhSQIxvb23Ad2uxLQui5Du1DKNO2276YmU417ojZfGbls0nj3Di
9FNQ9zeft2cXH02TBw7BdXyBAARj0Vk7EUPZ9dw/8Hratgyp4Hkn/DzGTkoBn1Nm
cWBzRbpuYzOacAvTSKTu2dglE08dTjlYZ3Pg5sAlz0W1wmUdq1lw1c7Rc1foUsWH
c3fTb7kg9rjKIIBXuHOjbmm69nQ+RQ+8x1NFiAQTceWY3nD4NMsRx6YyYjA442Tz
M+8fBCQZJ8taEML+Y3pdZyHki1GSz1rgu0y5iaD3zAVX9K/Q7nVubHI3xm70ZRF0
VxlkdEgN2l5eJKXfis3hFo9Zviejpb8oHZG6t+oPHnT24QZ31K60HJwWHfK0eSdo
PxjXq59pZQD4Ip3cvXPk1L1lkFkNUhZcLssE2ckdv8+OrYdHBUIEc/ZTGHiVoRvC
VJtPC5TPijF9t4AHZwRLTzpbbzKFK74SDXUy1OC2kGgfYNyoVQfNChLPnA0s1keA
y5yFQdbHWDuJp7JA13Tc18Qk6RM/V6V/WZediU6I8CtBqMAO42aa4GRZ9+LMzUD8
sH21yJ8sPV4Fksacm+RtLo3i47T7wxqk+SRuT1oDZNJJKZ/2QC8qjziBTfi6ITLC
5wqxEkLw8kwvNf+MkzFiwne9XOq+sdjfYpKixL60AaxHlMdVoax7beDEWK506Jva
Zg6Oz3gNI7RTO44+wqIB1qAkooItPgPjxe9B2PFg7QGMavEgVV6Dhh8yef0f7JNo
heQ7+DObLQqTs2r3hgo1lRPj41i2ATcYh2rv9XTaZaAisFch6Dw8SXNk3ZIK3+M9
jJz7PDIC9810zgi9j5dnxluZTjQWB0erSWWKdKTvZniPrvs4a5t0y0zzvBivfIAT
/gz/s/cD4vVgs9osreoOeqKQOSt9qI2tDbZC3yH618bk6i+4O/Gg1bNC6V1olnQ8
cS78EM8OSaM0iix1Ph99VUWIcr5O/2U97+k5KWHvivFBAp8G9PLnDpEjQGl7NhrV
F+8+9rf/6yYyMvTIAxDpVRZhO1pjft9ViONnG6/9vHX6SR96GDkBsXXTPXnPc4zP
v7MdU1mc3+QsNc1TMlrHMqhX2FoKYjudG0tZg7zQqj23nxWeWkEuOQUm989ci/pg
C7xKwR/dpnJTg4xK0j2n93QAVQG/U1vcqTmcx7wZ6Ex4tzVm3fz2Yd3t/1nXzNBz
IUZfRLs1hkx+FeYbroxkWmbzWiBQJfOKK7+CjZNAZg/b1aw+psyMQLMpDGtwYxNe
REROQlUj0/uwzQv4e8H9M0xObVMLAf04aR7K96IuzToOxXYiE9MtzO0EEX7tZ7hk
a4eCWKapyjXLqEnWEYjwXCSJPGQX1Xk6i5bXgu/BJJYQnkWG/gnkXnZEwGTwrGTr
DIw3P2Wg2CwnbwrAD47J/h320xYSqkrZ9MvylV3mIksZdSDOS7MRCFY40GmH5asC
l9IwWrla39c+CnsoRhSFQ9qzudMH6Itho6nDwnW0y67VV0g1+0wIQ2rC5IS4XeQw
RnmVkui3m7lnfN+jmloxkysdXklwxYvsHvf9QK4KTkFcc1r8P6IFGco5ueE7Nw+4
54OBMqqwv8m99zxtfZ1j+nyrMGAAaV4MkLVsJwgtCiUY9NXxkwcaBn2RxHEFHwXm
iO/AzoPr53n95CDuQHoNaf/sVHjSXo5+JHhYakLJxUZHnGke53W5oewUJNUcnKNK
4NIj5Dp6Ijtpxl+GCrdqrmlRqmSEgDWf5Y+kTTeR6UQ7u/DXesG9nHTZvCbgPq5S
b03gr0kNa0mjf56HqWFNmh/YecUZVfW+MxUhMuvrwl6jwlBtO1n1zg9Xpu4u8ATW
zfZls2Un+SxD4IssUQVNUH72zASGeIiQ+BahQo1sjTSOD6UAwXnBLkJlY7tzLvaS
DlRRFtJc7nnA1WlAYvR6TUc2WlH3QI2EgDKWcWRiVHygadHDWlCdOvf2OpjF8xm2
n5rjsmkajFsgF5VOLzNWuqFDWJj1GbwvlClbvv/oDU039AKPPNidSkshUcaD7b2V
cMgiKg9XXnwFJq7fPwjgRRNt6UDNvL/Q9FGdAWqB657wVolV9/IMNgB3GuDFqjXK
81xqnDUM4Lt7154aUL7iHg5xgKVXjeLdhNO2nbgkzH1u7tDLJE1FLKhSMps2GSE/
vpz91PL6KRLYgVoypdLjLjJ5DU9Qa+0cTSFSV4GwaMGYXFbrgVVJZ4hoJlSHAXtC
tTthWLpDlEIj863HDnzkX41CKS6DpsLEBKe2b5f7BMEXe2Ivmay5lC9hPdxE7osG
318AVKEETuNkI4STSsyFCC24Pa0O36WRtOFS/cjc5d/WMPOls4/SFGZgBmuEpxDs
IcVewAYZEWvH22Z9Kg81GmQyNBHnzlETsvjCya0K7FBxeOYHEOf92Aaaln+ByF5/
laWfcRUb/Y8Fuzj+uDFuCFlb3/X8Dj0CoyPMIU8gohbwvpbW3RyCyQtlUNho/xCq
w5bsNuoGu7oEM8s8MVEVATAsKAD5WZ8g78z9wDjK/MYY/PKyCuYbFfxPh09pjS66
2puWTCNDElGWKSHNMpxxY5/yCudN1/VOEoQJ/N07Gs3qLh46F4dRS4aonXuNa4Zp
q+Onn9hwWZnanR5S2hcZ8FwMi3kTm9ANZ0dQNDxLj7zxGGjJiuTlhM1DqOG2wa0k
rMgo0PlHKZLmysWhhPRiE87WXVXLNmOyAJ9nAtV3ajtPq+E6nZ0hMbODLVru4iYn
/aJy9q3Tqs7RWBv6TApwdw6q4YVSQjpDvl99MDyBcel7q9wu2iDf6y/WrXmQMDyq
M91fX8xyutP9oBbVabTS+YTSpgodtvGeO14aw6jkpOC/S/cBT2G9GUi8wgi473En
uBd7VvI+geb6R7mElm1vAMo2ouvaXM8BcG1CPWg38hFtOI2zo4OpOHTNGUwa1w+M
hVi0w8Egod2V2Bm3TKn2UL4usNfjrAQLNZtTxizX7+Grvhgpsx1UQXti3h2L2ITC
itFM6kNj8X2JtWZKYocH8tgU9RxMcdpbmroSesjUH48YTx/+f87EdJPMJNIfdoSq
fn0vmprB7YL/Vc0IXbDTwwD65DaXzjuJDcly988auS7c2XAd1Rd0efHbrN5KsjPP
oe+e+Hh59gzwLIyg7SzH8ZHVvO9w1dx7sjYbM3V0MI9g+LVRoLbUTTN4PF+XDcu5
APLQtA6qvCfMlQXmn//cDxNi7ihhslKN2+KX7mHX0M4wFhsopXBHKFhzdUkt/bdQ
qovSSYRXp6HVz25Yaw/GR52fsxbs1ScVtuDdf4CjxbparH/7zzesXq4dcBvaDwlQ
Js7QI5W0hQ4qq1lXb+ZMYy8qoBpoN67z2xljufNCVrM7bWBH+c2buvGNEDAq/JDu
pSgglSWBMzyMVUybJmx4QxXEBS+PPxK8nCV53If4PhVdgkcz+4YjKTGnSKbobxBw
vS5RiJ6LsaeokKg5/5mu/w/rjfyReE/L2ExV2w2VU88OKted2wWjLeVv/ekdN97V
wSPhgcXKmQGbIvKd3AgG63rtRirkN41xQP8uLSJQhfyceo11NIhvyjjEyOuvyCju
SekXl2YETDpGKIPuww68fu016BFaLtMChzTUWGoO0WNTavoab9Yrbc7/hoiDceob
rBVydfiqO5yacUT/Ng33xyzv83VqcMbRsphO5uxtRVFOZg/egKkjpDHtb2elBVK+
S1ohn8vLz2CPtT8LJtlcBEiHjigUh8i36RCa6uJqLF+jIDt160+0CxbmMoMlLvbF
gBN82OjXxX6ij9OhYtdhFQeeUAaA9s/68MToWc7nceAW1ar9yuQvrtc1rV2XN86x
ygdZkGJuHJJR3jyYky/pH6ciHbeIxGcZmomngL6fRdxHgiPiZ1A4LpsPFOXle8/o
us8aZ8lx47QGD33ujDjKwielKcK3SNchx+rEjo1MKzua0aWJslD8O7f3k8VsFacd
RuU8/fb8jHxbXOvXdLROJaCMPhJF3aFDhmawNMRzklW2F65g9qpoQhN+UIrkw9un
yijyhZD8rP91o1yiB/XgA6KCGs5j58c2hPLWaJDd00wlGNcUVYbVf8A4Rl6ZHewf
q5QXUjPVvqDs6P48coMzGrfY6iIiuDDk2sPv87sLUfIHO7WbMH0Hn8ZyaH09QEEr
ekhmy5ZNQ9ITHZo3pYr5H0xK/tRJj+5sGV3x5T2P8DyTzlUzD1UusB8yWK2kdVVt
CFZNHBNixKjHwqFEH4N9uUmK4btl3j2LeH+TXSdqlUpTGbbNXplr8uzDRYhCDUy1
lwDUroWCXWvFO+cttAvlkv7Ux1mzZ8xAY9TYCtAa03A=

`pragma protect end_protected

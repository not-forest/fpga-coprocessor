// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
F/X4O4ihUdPqpfRfHzTJkfs2QxzT27LkP/q4DFrSlfiboKHbwQpc9NeU1sEYVKfCIUfnmoNHUnKi
FakZa+I7JImSG43IwmtXXUB7aTfZXuxMDuIhj3pWLEmrynto7X7OesByCuxztL9PYVyqTwZClLSD
3KhuH499DOxR8riSQQ55Wz3zZRL9m3AYnaTYfWrNq5wBe62bTllIINYe/dfYc+3ogjz0be169GrJ
/lGxXSIbU8KhPyStQc4A1uAFFS7kQ/Yd8T/tXb3xhwWLKGm1cc0FC71lXnQM3xiXV2yQ9FLfEox9
IaqDAIZJRLx7iH+RcO+6D3WRV/0d/Ntog4/S6A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 6128)
vENBdWvqQ+FIjgis1StpzgEW8qXbiw1OCNggJB5tAKDp3B29f7j8/+IHST0afeOkutMIgBSCZysU
KePQE6US/FQjleJzvdfe1evBvv6qLjJBo5XB8f7khCAkqEcciHyiDHkx33a181cYuinSnK2+NzlE
kvNY1LgJfFT0RY1XJpNE2bfQ2bOmv7A80QDkAwiWbG0lKsW2EEnPvv3+fANarHuVZGsbJnCg+PRF
Pe8N5hUWIRjJz1JXJ01uhUaXTKUJnhXB3nPACi4KQ7ViQ+CYtIjGh8FHjBjPCnnfGNoJmGhQzF52
fuAAFOVnEFZu5eQym6FmZMA98mL4Bwl8BViVKGuwwvKjlmCgjPhQ2hHx3GSK/BsPy2iu9ScUop2Z
wo75dUUlObaoyR5MbL3WjYAqIOvt2nwI4gjeil7Q6Y+VA6H/8riKkTH8ePZtWFURI+TC7Hdz1fDl
OZ9N7R2hJVcPMw3Ur8wrGrsdpGvJtm2OiQ5zMJtnlxs+xLgwryph1n0j6txjsHL7jGeG3eX1IkJd
Xb09FLHnVGoxe2eazXecLKh41VZwpEdSZQnrZnsFtA4dKerPM7bLcWYulLhLo9szgnyt76iepDkB
uZZOA2aweGl2tuybCl20AmqkuGXlJyYayR890siZRePkm1y9S71902M3PBPdljtAloGoz9295GHf
Md5OYFgg5ndOfuP7CkrDIqbzaY3P4yM3UK+lGlt0C0mOLmTHCHaYB2PQIGc/2dG2C4NwoO6HlFiv
AVlQ7sn5hinO6vGYZpc3Q4EshmgTk9HZ6WsCkckdkQvj0bpsN7n2HDEvU2jcyJ4440Du445pTeJO
8wEj0s5UvFgLWWWzPACG34YfGz3bYUgsF7oIU4K08TguYa4XPJ7kiwd/ajJGWW1sXE/Qs9AwT1Ad
qsg+wP1ILDDW+XQ8BeogixNSNrkMLBXyIoUdii5yS5ALOAj2pRZjgnzXlhyAcNRQA6rxOf//0uh5
O7MTJQN4wd3YGTJ64ub9r25aN5OLJkpNG8SoVGGODo7XFQYLQMwDVmDh0yj+jt0oFfjF4EeAmCLq
y/FUuXaH+AZKQeztw6kTTmPjHsbpJOwOE8opLkRTfcey+GHOJaeIuFFpTwjSmsAZ7DCXOsNkJOh4
HG0e1faai/UMVJObsoEQDgtRRlPNsbe6/zICqwYsWwFuH9RDqSVNcbTi4XlrcwAkW9cZeNSU021H
dFCBkbDGznolHub+O+XSUjGAIEw7gbe5BZk4QarhpBtF0XI+o9Nh6haa+VulD8mpdr9UMmxlkf2N
h2W/KI9Q3EehxHHStq3j95YR9hD2RPtCru3cjZg7kM8ioV7omOuNiYiM/ZlcFV+exCnXY2LrDjMu
HRsoU5UgkeEWPy1PXeOWhl5BM/fdVPB2epUD5fqepjqg7eIaqEbNNt/Dwgk4mo6sNRxOSzva1Jsn
Z+g68sQ7aBVHKfKkTLf0aoxykc7nEK+qyDMhgJ9v4fZPtStNCA5tfYosW/SM80XktXNPDabVCsw1
7HYCODxjpzUOF9oU3Y31I2LyeMSi4F2KBqBQMVn//NJqav8rQJZ44sHTMWQtlNSqcLLII5fbAjXt
MnhpREukq2amBsOu1P3pL44VsfDlplLNanbtkq2LA6OL4j4UuxXY0QA3WVa5Nl/IwXJATSQ+tSuI
QDT22SyBJP06h07VpGMUgie0EGrJPF6QbNCBnInQj0zqlV6SWqyXqr7uTVWIaKdv1ogtAtAsrJ29
Opmrn5H59gMqPxCwW395liwPc1qDF2qpwXLQ8FZqLnanqOHoxMCKfsedbDM7TQGqNLkVRMWmDb6p
VQz1+W0Mi4MQIp3GrJalRE3xh4wdhFS/EYVK82WxLXS/2vYZIXR/3HbzLjHCrQBPlBfuMIl+cI8A
kp8jRXVz6NxW6wLs+APxe1jBTWdMRC+NTHSuLx60mk+zbmv3zlGkP3dwyhmuSHH09UCOlSbW1r3S
Pwuy6zZktD04eW/QbciHrEoRMqx1XnbvExXtukvsqqtKwYAh4VqCi1wrqhofhL4ES9IHLjLpRsBa
qUou0A8FmWdZuIoH4gIYpttgx3+3SpZ3muOcOWaihm3wtaIPYUetIVMuwq9YjnzFORFNsE/AEq6E
8LCKnVK5xWT0NanSzsi49nFBeORxsfy4qoXCpC5QWgBliXna0AmpU0VHsKkxx9AoaV7kuCubKnGu
LtrK6Jal1fzrlUxo30kHASz+6Gb2agGstd9YsE0kMcFn02DT/7gKKvOCyNjkxig9kSmfJvyP90ut
gIsG1LYDo52+SakNgvsQpa5heBnAIsAuXdAtwoPiQaVtHs5bCJ3p4NPnsCJZ1+sRzX8K7+dyhEV5
kcSv2YyY3/lDspn7Gr4nDm5/JvmGi7P74YVYgXXc9hAKCuj3pxH9YnSTSbHf/suRQIGAdOMnDF/x
T4y5iAXcf8tPKLa5wsndazFVDd5T7Sk25EWaDqsBNA7+8s/uPXKvTOnTPYH2go8QL7VaLTWAtGtp
fFV0S5Z7zgdvQojJIPJDSzWd9Jvcy4dYemXFSzfR1N/uw7rl7rCuzrYoCx/ssS2STT0aBLIZUv1G
G3b40c8pzXum5AUPDIZehYfajRkE1ZbHPfrIJjf0P2mT1N+5egPtim/ywWEPo+ypocS2Ss59BMX7
c1RBJW5gDdpM6RqsZkeBPrpCpVopyA5Tl/ucMuGtJEgG3LRH66+/HWphsQDimcVC4X8R2zxmPjE7
XIb2aLeJ8P7apAoc/LR6stg3gYTZOQrZD3zH782joXVX38FsweIBKFhhYZTtLeLlo5CHymadcT1y
YkOmwRpvjND//Bt4aqob1tEwDXcZO6vfJjeA1HlsjN9zr8+o8ZnurWomTUY6jVNCwJ0Hg2PbeVFM
VnphRy9qjRZcM4RZLGlPbtb7x3xGWHntOW25zvI5Zjw5oCHXX9Hii8gxE3cuZKHZNwC2le7jcAac
yfb8WOq4BZPQ+jphzZWNXJqsvoqFnEhLatXVurQlppTa1g2x51qfsp3/12gNjyBwtS9eXXdBLmu4
Zem/osYbVJlOyst80btUDSn/OJsU3QwbteARAsjsZHypMrGzD+JXgC3m3nxAUrFowhRZvdQ+od/z
QR5AP2qIxn1OH2iPNHJGeZ3RNcgpsKcb1GxPFOc5+dJusCw6Or0iRqc81rRKkONC96PbQKlBX9Q4
MFUt/bd3+IR5K5i1jpAmb0fTc1jW0EhSvwGjChwNsv5SE32JJqSW4lEzGxQ50OiN7ZKkiVvQU/mg
hxXoU8tqi+CMWc0FWY+8seZMEGeoUs8WW/O8Y21HIqIiQCR5/5vU/SUPvhtIdo1trhKFSrfavVBf
feMmquj5RbMt6LaXB2R0cvD87FHGC3GCFOz7xQX8wqJN+Pg0KMH+GxeWQ320cu99jIto1TUQ0eGG
K4ww/abMwOA1OiLBTSqJNNhvVz+oKMQVkp40CLJo223fAz7fU83CTCJFEMCU/f9Y8C4JS6L7XdsA
dG12k60//htxs614s1GYtFnIYpBpPSY6Zl46H6ELJ6hLZcX9U90YTgMJnPgORFOcULNuyzn9KQwb
Q47eEbH0G+9wK9XyVFiyZZ3IpwBL9NwlIiXZAI7JzVMnhUXYUDbnJeZMRw8GLmMLYRxGRZXL30rg
gVdZsDpqTokc14cd0qJ9A+jSbIaUPkoEOaZ7057mORV1kVBM+37B/RSuJ6drrjj52+767GZ3nXg7
9HpfI+gftMlb7GYJJQFB6bL6W4fmZKVZd6eRByb5EfvQc3SKNToMxuxhOWVOQ1ZcL3N3gDBI9UAk
bpvnEQfOWELKai3TU5ZsuIj/Tf6/7UTZ+6/R+F2V3yx8QLgMJk6izqaMllUhnc2CitfnhsKMD41r
Jh8SWAX8WCq2S0LDY2XvQUuTXAr2z1qIq5cQ0eRVWf3MFzKETxvep5APmRb49alvfEvTsheqfQDY
C95k6hvcTd+mg6i3nfroaDibZSjqQJjBTITaADRnuTHhdvC3zEqxSwGP92h3Cxs3KjDwqD6sck9k
4+iogb8OB68e5OlRtcARaVOdybin2PEYbn1zwtbGAkhHYOUxJ+rehM5H5rOrv6ihCEJCjMMqZ7bh
42eGUx+DAlxjOjxLHBvdam+GncgORipypfAdQVSBJVvYUKe04a1Ib+EP+4UbiFps+BW3Sb+/3q9g
0/M/06sF/Z39zNacffFF7E8OrpOgv40sTaXoJH0Rpmmh2O/5vQ+Sqzkr8lVq4lYri1niUPm87A/i
3noMrLoTUd4aLTF0kBscSXmhWFEAS4WByZmZuYZiDomWl7655eV+ix4uqhXTHya76r0HORbheSW4
2/Id6kS/2spqXS4IBDWIYQuBy7jK1qvw4mot5CZfoeRLueJasZDd7JwYxNnk2Ks80pu0Q0Vls9Rt
HwsgfwI00bJ6q3wR6Q5XY7hlvgIwxxHcjxYQxKY8huNhzOP8BBG7h3hl39G9ETQA8R57ChBPG7en
aZyE5a7QYwb+yAtICVfEqx07PLjLGE+BpXxGZp3Rg9GypTCJoRmlNIPY5SGFnCoBEs68iENB2j6v
H254WAgNQ0OPzpR2T2B9oFPPGCNs/nUYA9hG6sJcUTuZkAO8bbeIqkCocgnfuh1huhbffFmqaBze
slyq2F5z4ASkG2OBBPqvt5cBw85jd3QWkIsfShc/Vwg6MchZa+nrfGDXHkNUc+5gyq6DCOIJX76j
8IlklJ1td0b9mceqKv/PqI5026mj6b04lFME3zas/aWyjf6Jtl4QB2jG/8FB0CPRLQ3jf+Jtk9re
jtxNnKC6d/UXTrWL5i1oLAHj7LaGhMy68zE/uiWIqMhmog/g1/1RjOjB4A/65781uRuozrrn9Dbl
IfjPcNnSVT2UAbPw41EXMTBuKnDlhBg9PTAh8ph0ty9gJ6FGznBrcyQGcNoVMZzd6pGiHjMHPHZd
RNrPFbjSS1P7L39pSc0fwxdyFRkE9+3rBgrZWW3ByU72eT8xxkr65gm5jeZov7/cnYRoT82JufTc
a52s2Xu4sLDWMbnIZCiEDlLlMI+gV0R1Kfku8vIPCCbALqaDiHD+y30ycgfOPPa6u3SVec6p/zWE
P3L7NnxZdl64BNFVILrmj3Lc2oqjJ/CjHHWpYh23fYbLshC/2wipLNNeRKYHPQMUkx0CTQj2krM4
VKcj104D5J7JnMYTk46XDX14oY8MtXoWCUMxnuxNBE4bK6rISxkft2ISdaKF0kWqlscW3HqyYUIS
Xh5eoseMcaiUUPBc2Q7MhdFOgdkmdyRzDV6b54Oik7RZFwWITYBuH399cYOnjhzQeNtmiI3bK6no
2Tq3Xy7c9cPMlX4hSUSkChbRRT7mW4E2Mpy+6+Bwx2dngIRXkWQQM3qaTRY0ZqFOKRC9qFzpuuO+
7rlrR6c04/AFHHhkeZqIWUAYOZTjP6anHm8XMt9MWSt3EXtL7CgPi0klJQPskDwjs7rWtf+RaURr
2BVwvKWy0vp+m9LweHyELXos8dxEx3iVgTzZIPo+JjlARnH83zDncxh549/qYqxTEzJlDfzKBXBZ
K5pp6wUoFIwPRN6GpToiD67El+y6ONlxmZ4lYsNtyiUxFNemAuwLeN+WYwmyl9wBc5FzHme3yiIB
r1mbqJHSsUIJEoV2tx1/3BFOTKf9G0RQ6j5W59Y7L59kgJGMYJF0ZumQpb1bRub9Ro1+d+Ox2aQK
rw0odyK7L8hjSUlcA2xHJxJsn887UkkdZojuCeAnpkls+39wppEEHLQG0ShwPT1KO/BaTdMGac33
JT3LgKbvs+8tawcVckdyrqvY4EfhcN7xeQ3SiqZoIx3+HNM6azXzN5R2p6OEE3FxsYXooB/ciiqc
4gaIH+1BQZpsCe+RE4LFq0asyyRfOXge2pYw/tK5Uyx9LFz/Yrc9T70exZXEtEsGZshlaJXtI1Ma
h3NzueyxSa24iFNyHXWPH14DxxlorGiclv4k30K4UsMIBSsMlxho+0SGd6ehtgAaMsJpQF5R6/HS
4+H4G5IryG9ggNw1vVkYL5rNPp3TMif09Qp4ojkTUgdX+HuJRMDztpIcpFmeJcW4OsSZ4Iuknw7w
01IL1fpRC79rnuOwdjdgVcCbT/6qSVmglhpfuZ83xeCcO1f6S0Tz8iPAqp0SwXW2MOVfIrEIS4s7
jG59je3NMqIQbpRu2KrgiGmgG4QjEYuoz94SNA/FOUdZ0ChiDlhEge06jw/miyfmSX86Ih1bMtvf
gFdzJQNWPF1i/B7Vfc4r6PnxjHfMge6Sye15i9O5WvlmzNBqiwFIHhm+5X5zGfgzhxVcpKYMtq9c
mmGkxfT3s1oLv/B+NuXkynZsuX6HTn7DbZqBxWyY/arNBBjCHpcP5JHBLGXoEfGSIFrfNg0HjpgC
h7sUCvcYTYMsvJv4Vl0amyrDV4rfU2kbMQQP2Esvpyt4EWwBzHIfxOUDuBSF+BL20P5wmQYPBnsL
fHWDNmfFpar9z8s2aKl7I1zpj5lUErFyRM03jwP+4EwT0HCMaPRtOMJqi+uZ/0KEnGsE6yEg+KfU
FWWQ+uRbYYoMobXMi8rDsRHBcmcOoKkv/Z8qcycVCgOkZXyQkmXTS91jtg31vI2eTvI9mtXmLPjK
s3vjSVYqSZu3bKcgR2HY4znF4s//KuMPSrj/gBDt9W7V8JeI/al1j/WT9q03D5e/bcbKnMbdeQLc
STWl+wzMbMmnuEuhs7nLIuLriK7epQBAqqcexIk6EkqUUeviNar9Op9/2z3nuNovhrHENe160WIi
1xE5aZVOzaLf06ixaMoqkkenuU8K86ODINfRwEIRTY6EEmsjeqcwW8QJNgVGZoZwrwyNiNskMqTb
mTXjv6QqHgeA3QNNJAZ8orQeEKZRtPgIi9TS2Uh15eO6bIXsxVPusEcUr/bPaY7T27fSGFchFXvA
ORqiRJq8w7hOmU2Y8v9oiLXlB4WVPWy9rGPZDvaPZsADwL3tdvdc/I4AdLJTpb8r8N1Osw1578yo
G+YK8LuzC0fdFOUsck2dOhXdsJmyPoUspy5S1L6+1dsX9RP6HBp+8YcstpJqRVvnpHATOfJlKCT1
rMTVlTr9UP0+UgzK2+QWcVp1KoFpr/dPgr3AQMWTUcu+tGgZTpPluYfi3uBHWukFnFyWZ5IHHLk9
TF4Xqgy/D8wcqWCF79mhWcIjee5a56zLp4zMwlHDiNs1tNC2tdllIl+YcIoOGfOg+7SwwOQ8p3Vi
55o4/qAZCBXebMG+LTKbAciNSvvv/qftd//lvOIRpg/sgSP1YONTUrFM4McgJJ2coQfB8Diu1WvT
YoH2YnsuQZr3VUXMtxaPUeAdO/2ijx/6bpDe8jr4gcCFnMkoQlfTGsUsZ8nwSr1xqVzBhwsvzMfh
H2mAz4H0ykqQDApcyDeVrlq456R8rOXuyWRYQFKJrqJEMUqozKQpKnD1vQhUUVY1jOkd+qFAFP8G
n5JLxC70uVb1FTnycF86nPrWjWNVz0372rmtbUDtshajwgkrTUz45B+2lyPtYdDs9b3pCjT+19cP
gZFPEqDcS6/q9lWUVkkrCYh3JM78maltK0YdhIt5TeF01stvJR7DDOIf8eCyHybp6NUrttmjBa+a
zAFijkB2v6n4KYnfmwHRD/6q1UgEJlZ6RDH9wrCE92dTVwGMLIIkP7ywsrXuhNRghSspEbevFQ8G
wpioQO8Oqpl7XvSh/9KfiyzXZigTM2jWmwzq/cV9CXH3UCH77ltLQUnqdbF6N0mh+ahXyJ0j5HpK
KU/AqzM5G9sivxv1HTgcdmnjswok+V1VyFsUMKYrbiUJr9w84ZtA6tdMVnrixAYWG1ht0TJQem/6
ovlutexXIAE/AYrgrPzk2DOaBp22fAhlKKKXCyf3+UnDyQjS7UoL+sC6Cc1NsiQ8HiQ4kn+IX28V
XgHu4z0u7ZdhHyrqyhNP9YMHBrKXPtEimlqCWrG8RZfoi0vPd1QYWIBZ7k78FvRKEPcDdocThN5P
AGKrDYkzbs3P/GnAZIqLY0a6Yr2tiK45qSFzwdHfI42k3M3WEuM7vWdFN/v2q/eujk6p2NC89C7+
kIdQRyyyeEcrs4YWlZykUFs6ECys52vVkDoJwWF/Y8N0uLc3kJct75xdUezi2gqZ6E1I2zVKhYiE
Dxgdp3nrW6uiSWgufQSIFFQs5jBOKQ/ISKL8q3M=
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
BeMmAgFnW+7/D9c2QGeRwALCjxAok4rYiOzLCGd5rAi+j+J+BlmTKgLW93EycDD0
8wpcIP7CErrDol8y3zs1yHJ/DfwJ4kSWTR//ShsrslDdvr3DGG7zzOpbYu8DC8mx
H7Vn1F38To+STvsjKZXcOH/vU0cP+QhWlVVGb5Kj6FnGpdbV5kckGTTXBGiNUUiX
1oVLa9cpDyzB41965w0C1RZH2yGbmyBS//D0LF94SBLWuolNTZ5PTrOm9YQkWFUV
R5fJJxkrKNdkwBKaCoAbMZdj2XpTv1P+TuWCGcMVdV6jA/KREE3UuDlZIXyPa4Z4
YTF1dvnTIWEcUKhrZ3BhMg==
//pragma protect end_key_block
//pragma protect digest_block
XZEWsHk0BIL5eXjVSQyuUQa14rM=
//pragma protect end_digest_block
//pragma protect data_block
0iBO0HQjRfvfm3FSWzGqSYdUbtP+dr+SWEyccef8yFH7JMKsPcMhd6LIfdA8o4B4
3Fe17fPOVR10aARnIAGsqQADFRax0HQ6kFTl2ikEs30pMKYy+JG+gcwE/HYwQGHH
ZQtd8L/vZoE0w7nUPR/3mm6rRghIdkqRdDDXRE86utQz3zqMyQgB9QBL03ikNpiY
T3RBIsUpkDyKipkiHfnvKmh154OvrVyLobdWPe2WULYp3nn+1x7I7TG0Pt4t3iyq
X/QAhJ0OpT5X0yFD9v6XOpSihI2O/YAfGtTOD9fOttBtchUGbDoR1ptiBWVvb/Xj
m3EUIrPtFxkAv97kGTVc+jpAh3AKfsDLJQGU4qVMjBNjU8zoigzjE/w0iuIsYdFV
KNp3NRHhhUwnojaQTQxCfjLi4qcHsaJj2ND2dXUCNu6MZwc4VgcNCFXpBSx6WXNS
wZBHaRfWxUBXkZMz5sLINUKLcIC881KuOWIaPsFircOKbL04AblpABrX5UwUj534
yZT5SMGgA29hLST/ZADoo2ZrHkNSCmj9t/A7/vuSb3Yc/T4i5PV2EXjwKWo4As42
j4fLPs8mUp+Ayk4fjXJ5dob/AZzxT6x1QF9RWWilNrcexMEkLZMDlRjNJJHGBVXq
dbsYo8ovMsfNJvji0tFEnbALkYWotE6+tBHpv/SfOtjbHbwg0geRSJnII7xnCzYd
hfPPu2HOCBGwyUSDedBMsrV7L/STd56E6YA+xuHJh6EpCFkRb+IGH6qvBOnDZrgo
1h5b1Kq9lNqL+T3hH921TuI7E2dGvT3BEkzZQ+SOEwHOeFTLZUSU0JPtgHHKnG65
wB/UTsP5WSHCXQcfNP1J6Gv/LciAYXdvzmOEWgiAirPAmKcuSBMS5KdgL6GsVgKi
UcjktiWel1lBgqKKZQlkZxeIdIM0xkOd9addaUPD/Ruw9gioDfg9Gk0NFm2ArmK1
165JfFEr8P+4GaUF9LBCBQLa1mLsqh3XKLJwjRvD9DtvaegyNUSkU0iLNDqk6lwz
bM1/Wm2yb5x4buSdNvFsLkvFR7PpwToOeA/L4PaRl/E7b0+rZEdz9Kd9KlHSODjv
3ZgEyxZpmBElO0rrRoATL2Zc7rgg2PUhrCJzrbNTjRi+F1GG0HIXcBfaSu2GoTxm
wUcPbIaqYICFZiSiztFho0aSNjWc8HvoeIBrwjZ2uKrKowb67n/1z3MiWRleZY7V
7X9usj1fVGHGCBE++lrT584e/hXUWmPDJ+Nb6B1GDRI6PQHRLus4mKTNv9T03qhT
pSHJvSjydnK5VWEdKWwIMvj5JjkPs3iYSGXtw5GxkIDT9wkdI3KvE5fmLk0tXWqy
buD+HEdHJctM/miOIMaj/BVtROojMTvtlGnVX8hDWL4DKLnHYGyKY8Kufq33UcHn
rWca1I+jaNg4X6MiPFcyJF7ewnsrxY8UqH7SP3EHlFdLJLTEfYsOsOZZgU5BklPj
774C883naE+NoOgWSwEpkLXPFnH3NOiNIpB53pCvG9mWXmYYxlZqUborpdJvDGB6
IDzoEvYCtdLo/dKYmRua5AHOK+kLRlJSTCFd3UaqUXWzW2PTasBU1GvXfgATiAXz
ITAbQiva+F02QmRUe7UKuiiA9KVpE5ipSIYoL/hTevE57iUo5IpTX3n0kaASv7F+
dktGqcn2dZak6dRwpozQUyYL4ef3a8EOZYmMnKubcn9OEYlwS4ZBsrd6SUfktAbL
kk0QIvAPcjjd9lcAmKrG0SVtGIH+VQbdwupxYncxUMFHzHAUtlMmH6Q2wTIQcSZY
SymqHFmBCoNisXbM1gIcDOxg8YKoY92kkJt6noDXPZPNObcZYqqsAQCfo0pFdj3t
jNGZQ0zC2VhofJM5gLyYCbQue9lN7ZBX4NyfELzfoxh6qjpEaTVZdL3PvG6qzcqh
KUjOhClyU/Vg5CnadOLF0KgrPBOHKE53n7wiidScawXnUSMbyEAVV4uLtKR4oR06
VkA4Epjqyq/j7F5u7IOy0jFdobF2MuPgINaafOa2xHJiiOudT9knNjq2xFikjdpA
JZooedYiwq4CmRWFFJBVgCuFCIhElGKpDFq4vpk7zelQ1N+3GLo96RWyR+za1FgT
Ei1ZAFQ51DoR/KTrrCF0xCq6iwNsdWayqenK+mHFQCxZuwfB9Kg6DykS/rVlwYry
ii18nnjGCdjYjuQtc+DG7pFBtBun8cj+4Z83nxtGq4KPcNX1lhbOBs/viDqfw+ik
N55dWf9qe5FmeKEfzk5GVOFVQk7ur+uZ9l2UnBCmAZtfIopizPZ8uzj/vmpJnIPH
OTUsWiqu2Q7kKyKQ7162UYGxYftrPFcgdCEm27XCkD/z7EBzTGkBB3zHG5zmCcm+
WOV9ZTtuY/5OEGD/Nj5quX/0833MNRHXXC7FGfFws2TolC1HS5zQBO/pFdzqrZeN
FKJY2/gjBfiCrJJti9h1dZaTYkZqqOq/jdt6nIl4yOn2eJLPq+H9dv7vBi22KcU4
0tRQpX3ZHY7G3lCyVsnnKmwrRnoXhQCvn0SL+6XmuJXjwuBTC4wqZQiB/5lH/MFr
xAT3HaBWvvtboZtpuELgR6du09C0LbDto12ZoDThJKNGaUJonriPe2nA6VxN7g9+
qowER+7OdIqBFllxY+mKk+XSBYDSdDerTEgcu65/eCAHB1vp3sl2jvlS4ROXSuHI
upRxFp/MTpb1vv3j8h+OExq65Fhlm0rAgKQfmiAqflQuwMdpcggq2/KC+r+eZO2f
PG2dczQo6elxKRuW/hPnXqGy/E/xhr6S19DTNbKXxNALkeT+tATfXjoYA3zVEttS
n3biydQt9GqpSJZ4zgA/sq/MppBlNbP9oKUQyWjZW04pu7NIF4GUgRv6Kma6FpAk
y6Fbg3dMpwWK3RkDVxs5RM+mzShjQ2yA6XJstksuOcU01E1Nnsku5ugp3ovHBg/o
RE8HdKBrOJnQNuFr3hvidnCcEBORkTXSmfvnm2ydfaX2DsZ3/l50WjuiJAO8+Lfj
d7EzQ0hMa3PHw4dyqHYUzDnHImn725sZ5rWZGWCtHWem8q/ftje/kW/V8OjN1dS8
ZPa1PgXYksQSB3HN3ijxdjQqUIJ+vEbXWvJhwwSlmJONXMXcQglo3JqZIBGizvBH
1H7wQeaRtoWUR52YFyWF2tEk6hEKrAPLNriGUIvfCxcr4wKoXiLN8MqbWCydU3KT
haQ0xFz/IrY7zqIPuLhymfjGtfOosdULmfs/ddJLquB2VPhyUSQZkhnpKVoOh90V
YoGSjRB2ibBNuppm26f4zIaxqE3ynRvKoCcIBwOcTjz2z72wDv+aZKUwbwRs9vnk
050ynxpYrDItrjpxpF+T6DjnhyAQbIpx6vs5d3rCcSfRJAeOZa0fF9sHIjouwbQW
1dxoXiLdYT+COvmqS5tczdwHSytRaUJDa2Ondzl86yHBAZCaDvwr2BA2JqYEnjp4
SOwW6EnUjx4ic0zNKaCUqv7Se1M7OcwFfCbM8CQED7pEyumGjcBIbouEtMlL5wCK
3dx35TYnbyfFNE9QPcMY9uSIsNVN6TwmJobQjWuyYeWzrO0ine8SMZ5SjBH0dATm
eMVVgckNrgIo5/b3QpSnCFspBvfuZ9+m/GPAf9JAZlWg/n4utyNQGLSJIBWSwmnf
XnUiNV0XFMnlBs8cvtiNH6/qBvWKDj3N550PhGBkbSin3n48/VxIe3AKN//l9WO5
rDojYMMtFjw/DgAV3CYUdM3CwGvMOfU78lRlCxG0TLvtNpJmh7UHEIlInx6qE7ip
wQVAe6UvtBqB0Bew0dHlGx6qiUqq9K2Nc70WHqIUM7SkwLoprcjBBNn7pX3nZq7x
SWSqoqUKfI3vdghmHT8XH/37b2pLvtlwcRUirARxOsFU+Kce2YMCmpT1n6Scvsv5
Qqv2tPCLKiyc9pZczqjq3KnJ8257ywRP7zESb5Dp9w0DPSr0T9oZrc2uTmz38NZN
6WkS6TRDdRCiY27u2sMqNoI1BLbSsxDy+j8NpHN0NoiTqgU0lH2oQ+oTZS6YdlZw
5oYqQQ+q56MRFp+e00tYVcOLobpxKjO8bK/yarvwcTSAn00YW2ZjQlskW3+5ZfqD
aYhmnn4TKc1ceBSm9rLSw+u6Hf2TujwWFuCVABygwRS0ZY0hdPVBAHCiJSQxlbkT
mW/U6KjAdiyQRPxgkiY1kHPWS8q5w8GvKufFzXacFB6Rch6iD1TKjFK7eRTsWtxH
wglz+qzsHHu30/0EQBzJMK4DCoEiAsGD8Y9/onmwSnULvKbB/5O3dJ1fbF8Ypsb8
Ns4KFsX3Whi2PFac4WNRIMUZmT9UwOpeLazxYBfonB+p37O/MrarQLDpHuGVeVRM
nB+RD59U6UHg1yKmdmz4lM670DuRHTp7WAitVy3bQ5GodsgRqOC6owWBh0WbS07l
UZXginux1JiqNyDGVVtSg/SDBwhI0jr6qq9wfggkIeSE+Hm0nHEkINZwobeCXcMO
BLtPJIRVikbECGFaAC/w57EjgdzW80CxSkX/pm3SQDFrYqggul+XuGf1EdFlEcUv
lJgvKvfX09vftTHDyOiYAm0d4KWcsADCcVBjP67FpuYi/hUlF59exEALj4SsiPvP
Jvow7U1tWArxKFHn9biBkj84a9yxp5jfEGrO5HAiD1QAYzBjD7ftqW/F/8IL1FvT
c3EYeJvnkTMUnXMFMq6MEO24rF+BEbS2Og4sbAyeUS+nBNKUB/8dY4FuN34fMfj0
zzz6M/RtZG1XhE4hucQyiH31GbEvL28w6FXBDQBZ789qurdlL+9MXWMMT8mrbE0D
iYrj+24RAGj0mCrlvuopCDc1m2wAQKckbfk/3x378Tj6hPk1IItV/pFqai98q0zb
xid7Mq6DCAHLwNH4agZARqQVj7wB+cyrCeG+025aItHWHV9Ifa3XXskDsqF/Y7q+
+2MEJOAf6h53qCzzVzb3rA79KPYSAO/2QyaYQhTjZp9dTC6OYlkBEdzxR+gYP0y4
mfJxQEEvGz9yGbHoG399FkXG71BA5f83qMZUTZB1Nq88xB7Jjmc0zT8DEjWOJvop
fZnnBlJzA3YTyQk9LnTDGF81sEHPLzI1E5stnOG+wwd7FSpU8gdDHfYufdim8+g6
MUPSua3rD4RYaUS0mLt+226/qK6IrRCVd8fAKLM1BxOu/wkYoSQf47IQCLUG5MQs
duP66m+/GMrz2XaCkWyTHGjldH7AWtuDJbggSNwxzxsZGaCNx5tz8uU4YuWjejGl
329WOeUAbqGHCMB88Rj7dGJBSMtZP0Jsqfo3yY1jLVu+MgHzR8fyJWYSQ1ODqSWf
AJDosTKqNCD4hKiFjl6pVerZCKt+x9+LSudBMQJ7rB0xItkLKPv8EXqMKtRpOIvl
iZXry8/CkYUziv4BDes8Sqc42TBeU4+qHql/X9nzK5n6L/rDxahlPEtHCwH4kpcY
A05HyGBMKyMOdy/SJ2xgneg+tVVBy9rcDQr41hYrkaW5YVMvtoWHoru2yRs7EANZ
JN6D+itjprc1HPtj6lpvBaKkqKl9ppNywq8CiDb38NqQWVK6XFxAmoxgxLCVYdRO
o5Fv6nKzqXhjXyWqodunmt4hZOZUsmppE5L6rhnTydBIjwkqpVr9OyR/DG2E12qN
D/mloF2Er+pWxMm2THiwVEhrzgwbH/5uMMcqSwWGBxvamqQC0u1VwR2ibStn1+ei
O0XqSufNZc+eauD+Jf77/frGH6M9e8DeLpDD5TbKDA9ftX2nfwqeykS1AnwGHx4U
hdfhUr7DNnq6Bqq8Zmx+5p0Uxtk5rvXlLC5lks/zFWpm+NEBZUP16YX9my6xZWEQ
le6ticB3ikS57kxGadpvlRNUdhtO0Cc1Hyb3lKthF+8IbtSVsg5hW9rbBs+jmWSw
l2rv0iz8xJvcVLfXohKWvDKMffFVdQxXH8nPCPA/+e6yH8uqIFtA4gssBdfPzlPC
lXsSq1pPHk6BUcB9XXQGpVLWx4h7CQyy6cdS2OuC93ZiO1mK/pHU/bJwu6swVhsd
AlIw1OmfhCRiZAeu6fwsF4f3KZS7IiF86x7lGKoU/IaDJV1X+7ljkAgthUMlx9cT
r3USVOgwZ/mO4CczeHAv6ryCNs/ER8XYD2HXIPUnRgxawKIzwpIaqygl2yFh10f7
/Wm1oEVIH5POlnQefUfE/LoJTgez6mQNr6AKxD9ZA0E89qTf0KP8oPIaoIEVBZKq
38bvmA0bFLJCAzBGwOGSonBx9M7KoN9788ZZ+6sD2wDPA7WydkTmWhYkJAZKyxOv
UlbU+5jDQN5bEeqYENAs4RAW4h0jc/ba/lRXmbnE8S68POXD6DPm2+bFn78cgYOG
opuxZHqVvCxV1sftckrl4hrZidbjHHX8kxPdbSOz46OaltIn6SkNzNYTgU6QzYvb
Igcohl1i0aenSX9KkRcUSKrAHSEpyzQgSks6obkG1UkTXB77R+Ad4QSOHDqxZkps
jEXtPVBe9yvgIFwj6+uqgDd+sMHej1B6iW2SJ4HC26gJ+Yrl6rBQvHDJJY7DOJ6Z
8SZIE9/HSCNRDwc1kVcsWDtCS/CNTbhs+hJVNlRPKWYCQWNCdr5ktn8OQAfIDQvX
nnou2BQLQCqgoPzrs5c55jMIP39SVOWPGEDXN4f0eODw+OqXkb76raVFDQRcjoH7
dOslC9HeKn+k52d7ADqxf7lhsMtSS5GWc4C64Dob06nVU5rx2J5VMBJGLsxCjwmr
m1nkiIaiT7JP2wRaHQoqlwlKsdTp/q8ylOLhPjxLhN1OOEedDlvpgPXTX1Gbi3fF
hFtUHOFTxozfUq28qk7dnEOqHXMTfUO5viR9KBJ3wy+fc89CJieLHjdAZmiT9pVH
6pZKSNZmGiGUvNfOS+hWQ890lCl31MPR/tLKED/jMceP72ITjx2pQsnEjQmmc3sH
GLm2fip3qEW3PHOw1WLAdD3aAXQQ1S4WemTsc4sP6oH3P7hrUQzFZeXrjYeb00rT
99SwIE76+9wTQUx58JPFcpA84O41/k0inLNbqQ7twmYWnS0Ju9VN2x/73/8AZ09w
PltlqQChk+9W8ilxmMb7HsX1NhuGIEXt9CztPY27VWpKo2N3Vz8NLVOm1L0VpiMs
mb4d6c3PJ+A1MyzSrTihtU4bhgrRWVyhPlXH16Xu+wC77IH2Q7QUoBfMkgNwx2VA
WwCjGZfMjYa0yeyRvZWOyfQ7m9dUjSNCmjwMdPT98lHqBROqhnN9fcQkGBG+nAgW
lJPO++GDkBRQz6k4aA6gddRbuDMsHSwqG3mtT+iLrgQztBICcuuVntKNvKyTeUUG
ZtJhI1LcnMTIf67GtmtAlOTIDFUVtpjGANYBmE6O5VpU3q64++yNCLH1hPm3bPJw
ZH0LBVhDpw3He6BPu0VgrP6bdozME2RIi4KPi4lNepVygQJkIRyGWXtuGszKbUV5
iaBmf7aWFpc2VScqos61Y/EieZg2Q+3ozbrVWHnSCiSLCq+e30ARXgiQ3ENKtOdi
2w9usTrGbJOZqPcCSKjuzPExTtKGPccnk3zLxrnrrHN7d1yctoq/CBS3Blyz7GeS
Ueg1Fq4sKxVgq8qFx0tW5cpYNDBtV/i/t1spdoLGAcJCrKBQtzennwHh7gd2A3uW
J9jjkux6pRm1+ymEqIEHzqOOmvySeheEops0JpNdKetaYTkidNt6gRwLL836zDhQ
91AOPAbKC2btQ2EGNkx7bWKTIZO5guG9PVZUcZ55vZb4b+Y52giqOGqEe1z6KKCl
dZuwdKQ7hmzzT+H+OlbIQ7uc4HsBPbbBicYYS92ZHpkDzo7ls6niFSJwAKm3+hqI
gx281Me6nUJKFUAvEdP5qB+qO16Pzop7Cl41oHDg/Jew+ZKxJLVtpU08ZBCIG+SP
/U0aeoZK+mWV6r/EW0BQne2j8OKhxVzyEXyPtWEv0IReTA1El2BhRheuqCWY+uJL
tipVrE3Cbkb0jebfy0XbWAAFfgKGfKdBwKDEmqudbpIjHXDRpBqUQRJ7UZKgYtvB
sKsWBw7h2PV8MlBAUy7YNKbchWwcMiS01z1YpH5k1cIaAUT5ea8h8j/m3NVGZbCC
kWkT/ZQhtzPDzjYTKSn9roeXl9GGzjOnNd1+N47sq7kC86Z5GDJ9gYT+Ont1xn7S
md5ayc2fkbwuHovNrQx+2senNsjIvvUQo0T8nmDP/taXRUFBcYRoXShL9+5SuEO+
DrWeLLUK4LY/pOSpTGVLnPK2+FMV+tEXrF/PU0/PS7aSJc1pYChpIgzyhR8iKrMQ
xvlj8KKlr4sgSDOzjIVNGbdgPbPOwBuq5BqgJefo6Wsln7aYJf9FDg0XcYeo4+57
1nNuSsrwxiv26VaGpwOE0mjRjEUzL8JrQ+/8MH3dmxZ1qW232dvCs6gAzdwAYQlZ
bU7vdHpsXGt+64m5Sg5j+YmLlLn9EPt7rd+U/9/hBH1M3OWk9Bkny7xMHNDO574a
9iigbM7xvRTI8Y807/kIHRs+fqcEeDpG3HmER3uI2OfmFmCUr5EwU2OlcQIRl6dF
G/Ys8OzNgs7AeXPAOBVObUbfGKGNTM21GG07nV3bfREiWhYLFkg2QiNsLY8p823d
THLVNquhwvBm+j+WPK1cJQ4aO9V625IjTz1Zbm3dkelMbSEI7AunuQJgs/6t3xfR
dNqEg/JOZkv/xQ3RagNuH2qwss3Af1CQ57dgc8QA5CF7616hZBgXRctqZ2C4ZAiE
SdP5g4JIpP1YMYG25CYy/0cdkwsMAQt+6e7geS/0gdE3Drhas+kxybCAqknMTgrc
Lqfz5dDPzmD64ox/+nQx4ZmbWcM2MkTitMAg9c622m+CNzepPdRrksOnmdFunGTb
9RBNfjqgkHCLwR2eVIz44d/haO3FW7wTjbx8A60f8Vm5P5yhdTq2vrK4X829PqvE
J+KVXqP/WnHEORaPsb0flaqqpmu9hyfp2xa5vo6W6Z7KJY+hileuGHT7xgidxMaN
JDC3zr6VDsIj9EgMHxI5zQ00yWYMpJ5MeeFV7eAIbufbt7fojkgsuy/efRnS2xoP
XFKXwKjK4O72arjZGrED5CSt/pMUCQcJD91oR5ah/v34pGxRbHRriQXH+veXWjZ7
3Sg2ZJijw2vSrw4WsZzjyZmk0KSt2YqOtRKIUswhI3WvcV0ZK9vt4f7dXmk5Sdgn
CDN9TVMGIXAsilYS/VnBzPdFJS1ftL9rtwiYldr9pJ2M7XUHCcPw/v+9W1Z0QTZp
04lqNDvV9mJpGoFmj8EQbQIwTj/yl1rk7MyRfSe2Vcq/Cczlg/9fh2bF5Xm+XuZr
vEMdgMVif134SJ3ttby1hJVHlEH47dHjj+sqxicoDVfyDfj9EX4YprRsBQ8Wa6pk
8xsTHbXrCL17FsDmaviQjKbdLljZO3wIpsMi7zS2PPD1vhHchfojFdyOaJGre/Wa
yUSIXSQXC9ZdDDeNk1f4/vI5mNPA4TWlQYoZadu/9N1xRgWEg8AxSqb4TymctWNC
To60f8Anvs9IELng2FwEpamDvqQxpXpDRIrELUFqigwRJ4bb+NG8sGzEk3PBBnOd
DHmrY5nfTtemhiWkPCb6+KqTKsRSaorqbZzysjVGYARvrTzEttDLET+Bk/jrEAr3
4UmnTyU2EUVcsjUyl56fuY2z2qykXxV1k53Q30KOjcNNx/4KGDwiwg3AlEqbYkbc
e/wa8rMvxsO+mLd+U+X/QD+DVJ7Wfo9yt/wECzLytrmKsNbGDJLiUUZ5Tj8t3sEp
2gN0CJsezT2WAwZOu+QGETYvbvDGGdKT5t/dJAc+drxKA+tVezGz/Sh7mfFTaNEn
+XCRN5BzUSCXk2gNvgxmB8ouW1id2XOKa3BynDQC0oAdmDjpwS+hY9a2/sDwJCv4
GQvK3toVxJOELs6GgQbNUHtgi1thtdKvKifntRujHZSFEncfgB+smvzLm9fIC2Yc
ZnQrwORh0EbEpyAnXIL27TJAxskNUyZZvW01Nro1oo7OC6TYHasoaUldqTtaeyVe
if1oCGRA4kQlO73MzrlPnVf+aJB6oUvuahXaDhLhJm9qq9IKASL69k6G1B1WV3PL
k3j9CRZRv1U8WecPMqQJM4XDpae59+9KTwb6L+rjUTFqpKBE4hhFk7LcYAG9X75t
ts9JbXaw4tc+nAsDn7hNTMQDE57poXE/koOI5iQXyZXA62Elvuq0qXukXYBg6qWU
2eeGxdRRcXTJ5atmNBy3Zq5WBWxWD46BChtuBv/Wioa3FpfYjtln7fYF7FpwXEbp
IkB8eF5CxK42yNcT83Ltn5mjSy1N1CuLQt7bbbbyGekdvZPJezKXdBilE8IrkHfV
FVl3LM8i5SAaLUP3GRDgymqR23gMYcwlB0DzpAtcpHTY5rnsXRkTFJIFcoJ0mPZn
A19AlZNAUYh83HrNqwWuvlwuWMa2Qle0A3u61DZRr0J3FMoloCmpTnnpn82S4xyf
2I1bNE+xStzSsSZn1gcOI1eKgW0Pq75CG6bwdhMttwh+vcMFNcn6s3SRou6DlRAk
24skNehVQMufQqj3w6aWox4MvEEb+lR6EQ1MixZNGbQx5HMGHFEexS95w8m2YLCS
ijxm6Pri4/IgGMvJC2QGK3KfWPQ7SI0NwOAO/Yg91iLRrfyfMg3nGnVjtRnGu8VA
N4d6vLHvXjiec3bAbWmMrEnG+uVqqrBWeVF1hC2LzSnpJNTrOntk6/dOqybTVOvu
9cavdEoHkRtFB+XrTyw2iN/sd1m2WwJQf4r3I2G8frtva2ENhMYgopjoFzIaFfCO
mw3ynyQ2jOsbydgVpnMuCTIydYS1oy0t/W+o28ADg0qM9nWC5nxUbd4/1mX9PPPq
GO4rr8tYgEZDENCh/5cZIJsk/mObBB2BzSK4V2beCOpqzU9GRn599NxaVByhSalM
YLDI+6/HllmvweuAsZyx8+eQpsgbTNMahPRhgFbNgatygAyYd1ej+PY8/WRY0cn0
QvzM5S3T8qtcaXDUEyqRQRJgYcK+8sLl5JIpyDF8WUOgXJmYRatNfagjwWaScMOQ
sOmBblD/ZaLhtnwYNNs9PIJdlDa4F0/mq0iyiWluoXZF0pnNMN5tTdlW9TTOFaJS
hdkqYGmK9aBMqG7mTHkurVZcaOWMQuhuYj93FvUNyjGdcahRkqmZwOZ76XhjrSbu
0KuQsNgOEgzkYqHYpEmmZucDuXP/xGdlbO2i+pzYXZM4OuSnXUl9ohdW2bL2L93C
4YluUIeC4myrWJFKov75jociGdC+35YjRtTuv4GRemrXUFtddddzCYItEKdXNF8u
So2Huq/r7gn0eZr5otJjUfwXEFGx3LiPNbDexNyS9M6cwflWsH6YDnpHHwVAeFns
nvdgYtUCIJaO2YbfpsLBz7gkOR/OzaBbtEqaO1F9h53jkfD4v/4LM3cZqG6y3G1B
HbukEOiMhpyZEnttEiFhmW6ws+eA/LQKwj7RAHj7Mxprnajhv1pEtwZEcwldP2QI
l4m6D9SbPKIeeNqNdKsbYvkHP0LgtpqnCFzMZOnKCQu07ThXNHjzQYkQ1aupMOsk
W9IdeVTu22Q+T/I4pWAIwxZk5Ykl9Hyw6/gU0j5sbeqSnrku71WDbECtj3kOu1kH
MQbvN+oPQ55zRUmHLdDMaK3P1X3ANIIavVF1pxu/pANTnzbcRkccwayvkz0uKwqI
gxLXPVf3XmV/mlncONCu75OPtoEp+NHnipMPa9WdsqmX1P4y3d8I/vyo7y4L7U3P
+92hZAYcyT776W9czP3foy72RO9Ls6duqQVRcfGkRzU=
//pragma protect end_data_block
//pragma protect digest_block
3redTrmtxUonpib+MpR0zpeHVEk=
//pragma protect end_digest_block
//pragma protect end_protected

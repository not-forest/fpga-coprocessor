// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
pXEXvYVarblK8p3TolL2rBmFFGGrW/WRMr2M327c+hydJQtIk0N/wSBfx5iEGtHPIioklyGwm+3D
dWorm1UAwbqzcNh4L0ZpXD/ZilVXiOxUMThHzjuk0o8GQOILB8K6mtqu6GxwH/08dZqOaUG9TpMP
jZwhEoDWQOKNDmnIn1F4bmvI1Xkr7HuNfu8mnZ2pFU+oVCdWZ4hqCWAGyfhV407vp5DvP+cC6/rX
YOceLRpxUmEHafWVCOp4ol56Tght8/tapYEvLFnvBflOr1gZiZpKqBhd+E2gfw6tQ/RuKfOGz9iT
VH+4XDVPvA+0m2gCrQoif8Tvo3J+SYp15wI/IA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 7040)
FFB+9nCEvtpPEnDXgZ2PbkK8NE7zTbkaSV3/Bi/7YGi8agEY09stlYvTJgIqT2j5AZ4QWwTPU7Rt
j4sRtVgqxl3qusMYL1rV4LkMBuLANavRkDIhaeoHsxhf9B/97gl4rp/5fnbG4lby5SZ6g+F6udgR
wdZRPiUoTr8Aj/576wluknJhPs1Cs3HhPTKhD8cj9EjSuA2f3L08No7H6cy/zTwDtENOFf9XWq0X
Z2KZrB4cvU9BAGEMazDogcKBrQZmK1XolTcFMbZO8W7LIxdsndzXoPZsj4W4WUPQiHO7QWq9so9T
6rujZs3NGYy7PoZ7QwLikLO6fkRQLN2wCLxJ192Zt2QAr2wry0RKI/iHeBChfHyYrXqo9Xj1o0OV
S7WhMAHmOpmL+Zl5v2Bc3gsNPbB2FzBNUJAVkTBPlznrAAp1h1BfvUf15k7GC2H5pOXNaSdr2Zi6
lWcosv5n91JkszQBsoam81pL6OHC1ytbv02VNJpAxhy3CgXN89w0FeKG6ZD67OfUmSzg0zb4lpqR
DcmnlIhAduwV8b3dtHKOrV/ZYq3At1bLH04pkXxlFh3SjCro/dVeqWZrg2gfItf5jRTkaA4DxE9l
nG/tam7TXj3AbnPJV27MPGYIGmQyLtKoyRtmHlenMCsOB//PiSrTimxyppqjhf9pG403xBbWlkGT
ZhJJ/VoubyAVBYTrblu8N1Hm6ZqFm4Psy32rxnyVsjEhoGactXh0ME2drT9FQo6r+bVcxJ6uSYOd
7xQT6azgvtOILP45dvT+YQG5Y9MTJCiwsIuem5yPletTM0BEjOIqTkINKRFUOKbD5rZ/Af0K8RqC
w2rEVNZM/Yb2DVHRv3KOR0YLZPK65X7MgOAGWqXoZW6A1/jS10/IIZ0ID+HWIVvMlcMBwBPs0qy4
5aCyjp1FRE96Fxh2zLgc7Nt3B1eIlEssj+ev8KMR/Z086VsBNkJc6gPsrsSXTSoyn2s69emj0Y9t
f7AQ2ukRonm23Upbo94pR8y/4ApISrh9nD2yWFpOILpXxYLhaSjcYdiit/BeUgRUrVOQqefZ7EA9
5vOOpa+GkiE8q3bqwyvs4IShzQjq2upmbb3Bw2iXnjyyvVKuJiPKDB2zydzwFHguJkBe+3vFPuyq
ddBkOtNecaYzh15F5qc9MH355+VghyaYiDjQUXY2OMfoHSPjoU+1fgBDq3506Y7iOSxi4UJAjA+g
qPyjsmDRPIibrFK/h2EiRP0qycg4NY2OmSGVkU5fKvyUhq6nMaL2SCirmv2lj1fQaxp4lpnQXMm1
Fr4bE4DXpVzwi2Qcc8tvGIZd6kfYWio0fuCRN49GGz3Ezo/sGhRPLMMw0HW8+/kRxIe/vFTk4Rqc
myTNpqidG4Z5uLHIKyIUUqENwSUlDXat1A6yzDUpyrHLvFGB+gHuhN4rwaiRr5u6GODHEery9Dyh
carfqeSoVAXHwi7ApPfWhjLXeJBqQp8byYG9wDmUWJT9jpCNo60uMvOYkZhexzoN6g1OSfAbXtUV
XXDFA2bytPA8szNAoucwU7vMXxmrYI3IxMqnA26ywMh+B8aQ0ovrJRir19w2Uo6TOpBWEqjT+6vF
hg2hLjiDudk3pnMGPTMEUPKiBpYa7XFxUdYd8l89SiZ4HNa4Cm8+dtY+9FyEIgQnsCs7nrDOW33l
rrjLNYHtDLPuf9+IzwRk0Enp2RVpIBdi6hGUh+j/FZVRY5GG7mL4slxtHKUXugvHNUITt52EJGv9
dt8j3mvqMWJrxa4YnUBZPT+SQ3NGulmdX+AYgqGH/05wlQRo+JzCYDMjK8iAwXZGhUmrOykdpEb5
ZKE9Vttw2DMbbzBrHm4d8f6++jBH3RYpIb/8Na+ru1C1bji8MeRtJSqj1tTTzDYPYKS0YIYnmz6y
4Moh0t1reZi+1j6jLL7gT0i9cup66F5MrogoECeU8JHC/QnIL+xMlrxv5a0gfaS1gIGZCL56ctqb
jPwQBcu8ooWPWG5LkBrOsI2buGyfHpFZ29bPrWyLh2Sogs+h9vNw9z8nWFhN5sKGDZ7m23t2X8YT
ct4h2M6fmR888tu2oVspaJxQAIx6RU19r4DQRfsVxQaqhzEyYKEh7TAdCgrsRZbgpuljnyL3AoPz
Lz2M6gba0SDH+YOQ/0Bx3FFNyjpucpwTshkGsv4/JI8hYf9re6FdEZ6oHhMGZh9EHmxS+nQW+UET
+O9mrG8kW2gB6VFJSjUt5eZTb2PGubNOBgrchVubZn/AHkkpVgn5nTkr9BdhCPzpSTR7Tk+qjsX0
bTJNHOzFCd3ow/Co2skNuIhdT2puuuHQqR56bN+zMakBhIn+wVdZSmIuVLJbzYgp8VFgzI6fGisb
ulkNUvj/6fiYinRqmq3/2nUkCBEjYtY6+n9Ek61+L1zeyquI3+35HrqaX/Ugs2fSkGCdlBCEYLC1
rHcbyVJcjZ9v9Up0IYBYuX71Hs5qIpxMLbD13dCKHUflp9NMl8XuEhEBmiRc27kcb1ocHTiaZWen
oXD9JqlzgM4/KQLQ+Rigj8SWIcVcwG3QQ3IRf51zbzutIYKQVb6z/g1QDfn0jCewY5XRksH1zCoF
XZMWMe1JAmjf4DDcyEPkELAYGvAnuF1o01Pu4qlmu93ax5r1dI5QXCi+QK6sr2nEXU0x5g8Uk9Xr
mpC9NqeCDmBO11GSY/pTYJsjP9LlbT76cWGAdGZe0b335cMgdRma0XzWaU1ijAmnAMVSJ3AN1gwk
gZ34QiQqsjq2dHWPi3NFb/Y3VozSAkIeK45sLnfl6aUx64Vlesn6n9jE06C/N7e31YCRjNgITfyM
1it6ZzcIP/952eDoMDtIXeJFAzSHhbQ+fT5lXWsBmNvb+BTnVyPXxR5SGnrKuHRQcUB0WeqQ7IVf
gQ7KVLZdEocAd6eW4Zpp6p5vhPSsbqPKG9QKRVxge9b8gmJ9Ka/BsAF5JVT9zH/fmNV7mNecnUpm
e5IY2kJFOnShV6CCULhJzPjq/O4tPX+sA08FRm1u8PzgGEEdZXBYHY3sxg1pAOX5eRCDbsfSYqyE
WCOh1EfumxkwmCR0MEcWbF6RAIe9O4iw/0bddIV3FiCuMOwp9FWOBx2DUBwQo/2MdpIcSxrS3TIU
9Wp9G3UsLARQIbCbzKibgRT0UMa9VaLp/0XTfwHRq7dc79QPP0uv31mgw+AGGTrWemHSG2cZ12hG
2xEfOsNX0uosuSWGmN4D0CZRN8cZ5khd7/X+Tzp4o1pPfip0Fwb0zQKd1wq08vCZiNI4WSzNOjbu
uqgX4cW84gUbDLlJDsQWqu2Sg4Wh+G0d0ZYDn9zcFR1FvCz0KrOYP15ZUCszL6Mr4gD2fpYglthL
ZhVMEa6EmtVQS3CtR4n0BrarW13dDsdMTXjkjlbkVb0IGZFaxU7FaKNwLLyCFXtT3lp3m8glbBHR
Vy1wnoTOFXiyeUa1hpZU0YpmhS5Fjs+4l9VNQ/qnPA3/WaEqMd6g7MWjdVbPEa8c5zaKNsJa6z9v
PnoA4UK2v57lUT/3TRCtj/f5IwZwB0gRGK6B8S+syAqiT4rghu4bIlIzJagsANgvIugH5TkX/Dvk
mFSRZRsqej+G3/2OqsCPFxxUKtE7R0URkCbEmD+keAVa9M6fTlYx/fVkPNheXnao+31KrLS4vfo8
wTKh8Ey4JVWBwYLKA60R8qWMtEt6lm8lWE6PFuxlO/8Rmp/dcCm7BMUd+jNXMZy/zaazmI+ioAHi
ycAZVx5X8vmzyIfeCkLbLghHaWDRykrDUiESljIESoKcIWcnBnQbi/QxnnNWUKV7l7t+mI2ZkEwQ
9uVchyasWMM5bTM96ui1jdFmK2dx+THuakaG8seEz5m4NicHZFSPi68BOKjhk9f+7eBuJ7AOyPCz
wSPsnbGTnxUyoWkBs/sSd3rHhTZOB3RSAwR8Ar3PsrtCwKfFKAhR2PkFILKk+ZbQO0IMzn8YCSYh
UujMu5hD842o3oR27VkY4+6IQ+eqiryrFDLl5stymfqN+EWIOPc2AeVszYyqH6HhoXFymu+jYc7v
pyXgPG1/rVq2DAX+nDlrOACEtSE8Mtteca7Ui1w/LWoDXXBrF7M/QpuJzZAT1YAAqzPCX4K5UlwB
eHI84QPxOGHT25g5Ep8Jh/oe9YL+Q/4z9M+LbC/G18tVML8XvIMf9cnVWMo/S3wGu3F0LcXMaW5i
8OZwBhrORw2Uf3g5/cf0HOyyxS90kC2+UzcIQsxJtAbTSTJ/sruUEaoWjGiVSqTR61PSlhoeA7iv
gB2wyr0Pv+9xTqwYbfXeQnBXwQcjU/+wuPUqr4u3miW00pbSZtozWKEK+Xwzqsch+EO4Uy4K1xAR
S26qzE9+3ArGlSMBTQmoInYLn0FmBJEExWqztXcvvJ8NWlXFxKzlkHrB2LHSPeAoI7DhCYm8n9wB
xG1rSq6id9hOgRWb25nAr6sjDF6LpaJwcPVF39qfzAVC+4KAXDZwqB/aUdftdZORJjC+XgtPCU9S
iUJFMAA4gQadjXx0qpYOKatyAigf2gaLCM0fFwmfgv8hwnZ8iM2SjZ3m1SMlNZI/FwCvDDVPH4DR
sU8cELDANArp4KhxaYCWRg3t2zdxpbSxr9qX6etwb/uDKwLzxL22V9Pgcb0vx6DNKYLWoRaYgFiH
GVcCgIvobhJXTobZW+4e5gULmMOsIjpoqAClNcbHQr2FnhB+/a+0A8fdllfBTFd+phu997raMC6W
unc8SMfOZdkYd3owycVDPGQZ/e0iKAD3sYjszkVp9P/VbDJmDITJw/Qtu+h+06zZCUlTXnPGI2Gu
VXerjmG+hpGL5Z+w/DLiNkWB4B7jpRajZr5MMHk+vj5buZJUtJ3Gbn9g5ezLtYN+y1EorGp383Uz
EjVpKJMo5obx+mm5tr7gSyVeSO4efLkeAJ0+uvJJO0xWHpX93TkMFR8P0LSvqymLbnZjRueJMXs3
KREI8pF80AH2i7ym1y6LkmKiJOjrLLWqUIAP8IeSeaUgMpOb9BKaB8CdUJTpVcgZr9Cn+mZNJyc/
s0tBImmqKAFtM0Y/YlxIPbrn/rubKtA2GMZByGgdqrQikUtMvDtIuCz1LNZDP8OVVW3OEn9I3cah
mnIGlLhvBCSBCScAhTAtbDIEVtu08ckoKeCbG4jTn+C2v/72ET4GC1MaHCHOyLK/FpiwSo3TO9QE
GXE6VyOhVec6XH3Zn0p3VuGSJGyw9nVjb17tPc7Hy77NM7uC42oPjKgpFHzHWaw6copHseZV9nrb
OaafZ9/n6P2l9FAOqACkt+Y8LCausKWePxnADyQF5SlonhMZ4QBRIcNA2rYu0g+zAcp8L/dl+nIa
frwPjqgjRz9fBsrOFqrqmIksrSxhkl9W9xIj7mVzftrLpOaDvvE/4/HoBxq8pHReU/37akWGWx3R
FHD/Wnj29Q0JjF7ewerLWH+2ZaqaWnkK7pP1X3bSOOrVv4GGT8mrP4bsoBrW7jHyjxsb+NWSuqUs
26WZqosoJ0pQ/IpOZLhTRORgq+w4g7N3+k583/fuAm+IgN87ZT12s8W2F7AU/zPOU8g394+F0zVX
HoYctHUCCBz8zLL3h+2mdp6YqKbJO+e+zxZxkQKufom7Yl2lfKDadPaA5Tuwo6H9vyMahT4AjwTN
axuOxbhWkMaI56Ba56+lpDYUCgl3WQSfgB+hU2YiThqSEb22yh+5+HWo700CzFCAhSbo0Uyn7zV4
KIZySvmm0TmflHRYQZ/VnkkRXevZb1i2JT7NwxahgjuGJTLtmAVz02o6RUucEUsdbRgWMySsqnAE
X4zk8/tjmB+DnFRu7iKpLA5yshyE8/wu+3byWSG/BuxbD8ttao/dHF/UHlUAG/ayQiQ7J7XeIXK8
/BheZWmjq+KdX/dWcBLUL9BgRgCn0QaTTi9VenpHbmqJRtrUqr1mz2+8asTDtYO5NC/njGee5UvB
LSR3zOLktv3cPcr1OVQMZPHQr2bhghPWrS7qpep9VKmSPfvgTK2T4mH3qh8i1PzNiprjIxpqwTS9
CY+H2T689vAaz856KeEatQhEIiO6XJAs95DGoRKhayZtnajqMNd2zgEz2rEI5UyubbppYlj9oAhs
TsblJVNNlk1jGG47f9Di1GLyDc8KngxSJEYBRxOZrQsjz7VwRYa+KU0qskuDwVq3WB5Xbi9CxEfY
SjT9026BRhRQRYT6B8ba4vn2t2MIfJmcPrsuDhmziiIgmU1YNISZ8eQIuzEyWXUS1sgGT4zOdwhC
p2CELUNUQdhOFgamQ7hSEzPNy9o7DfecZf/3L9l4mh05C7OjNzNSrjB8R6hbj7IFS7kXYyvl7Aec
pBweBuehK2gKi4H4gJGt5Bdg8Ty+OkZWL3Kta9CjddtV5K6/Wyeod0AfQM8FdyDFjQdfuhxwMoHo
MAPt/TYvqqGe7ejsC5PfbpfhoZ/7XWW6D6AOk1HdWPHkjolWdP70niTG+OWln7N0meR1B8tPI7j8
Lus+MiWfuS3HB/cwb/aXxPkCzaAXpxBLYa92+Epy++pdL8zRAgHqKVSCPuj9hNEfvozEKDNjZr6C
OtaMq5fnjnL1GfAl8aPyN9J1UTbi5KZZpygI/lZIqz0Agip42lZzT7Z8uHF9GNN6UxA4BH81Hd0D
4UH092rvwGOfx19z1Py7P1aeWV7q/X8GsLz9x8Yjm5Ae7zTtIiexMIEZn2Yr07zoMI48KwZsp5FV
aiwnOY58hXTeO2jZrxQo9PTx1x27rDLcVhhccWDIVS1TiTtmvFXUYrZjLvV+FmGoVJr8Rwo3Qb5M
VVFSerc5LN0yY8uP5lvrO2WyKsPVD7FdYV/xztoEdma1C1MXEA98J5fm9nVPtVoox/L7HAC1i/Jz
8ZKq0q/XYOlA83hpCQHPTUre+CdAyiLNlKoF6lvZVh21ITto20Uzv8z7aZzg+ECW2xmG2ZcYFkfu
HHhhd7j6iaGP22nckzlL6N4F3l228w6k8klkE1MoqFIg65Vc6v3Em/4LXyce2lS7k+sH3qrRGs6G
fU5WrUAIaYvCMlWfyDutDJkuNLzsk5b9lRzu7cpFWarBeXmBNhMpMEYajqrYlojRRpfuhiM4LVbM
XzXpEtG4APSIjG3t864a0cfrbNPWm+jMjrMxFNiYJ6iuKjmUpEE91j/IOxzEhUu4G/QLH8rYYbLU
+jtOc//6FQC7oOJN7/dI0m2yKMjcyK2tKOOt8/JksnA9UxP7mELY093yBGrXr90ic+By0rDuyPlY
xM8K/9WZvDqPRKRQMTwUNoGGZG/sPoS4iwHn52k4X7nSDPA4CDznuk0sAyPBVIBN6LQyB9rZbrcu
amTeP6ofA6kVBIldWjK17rlGEQaX+JoQL/HmT1wXIfHZKrrkwPWd3/s8G9Hyfl62OHeTI1C10P3c
5XacUkAzxCp7E0KeBLaypn6C6o1N77euJwbMK7+fyh2iJvGp+obdRu3a81g3yen2kt9xyaB9HOGG
IQoRd8ILerUFEC6+bVqW6Bf3+nm/WjIISi6dRlEZ6AgbGF0fJNmsWe53KXSnpmOlztt6rsKCJ+Fe
UxbVbgeS+yeqKtNkGsxFETEYkXG0y6njxDuIoRT+3xBxvMEaYq+NyyZwTU6bjUgFgAk1nBGm1eOc
gg7HJYyix0h0hAGt8hARWGm1CgHRdUIdGhFa+mYslaMCMjFL52WSGz7qGwU5xLMyn/U+TO2sV0Iu
DPeeGNg2Z6JdQsULcOsIuQu9MVsCgrzmaryQHEeD1GTVv7Fv8Mz71I0TXShSEAxkwTNO3YNI7mUR
xFywHTCr9hRaVdWNW8DQyhbh/vJ3n1fTBb+mPQ2KkLWRrOqvDeABT+Lu+ws3F+cg3Dh00B7YN7nr
DzFltQqClWajnO9wIiXVe5jetvkyIFwIRTrhOwH7apO3V1NQi0ZopSO8TOacVb73jc0y7xJ8k1GU
Qfm/JUSdDRNr0GeO8M5KNQi3vVnAvbc2beHckCFIZ1vN7tdw1vmXmiHwsj2jro3VD/V8sxkTyF3s
Tbv4cv9amNfKB5M0n6PF6gUMsCKPmCxlq01wmaGOdllHoYrkgmBZEdfBMFuY1ha0O9/i78biwRBT
vgPOv/botMeTe/72rnm6fRXckOls929EeGl+YfQvGXpMjctBgH4lECTlo1sgy7FeASfJG9zG47a/
oZttLYf81Wr3wV1sfFXNEvGgMJ7hDbUX587WIGWFg6n73rwJmAX7iImZJQQndoSjgSHonAlV5hO8
9BDv6yDVl0O99x6PNMVsgSiokSKoeSNlJ7IYBsFFGwkIRQkAf/EYsmwt1Uzi1tinLt98lbjLbekb
3c+hA9gaxWIJ9CEcHcjT6T5RIXbXXD0GAeqjc9nUy3G0KiJyVbQyAcanTQmVkGV+GPViGTYdlxNy
IkZZjLuf5pcwQs6t+9WCNdCI4rkE6iCpDfM7/cTrMEDx6DieHN92qQDXEdjVVMoiEwGfnoWBSgQ4
QZeCS51JICHNfx2Aw6vs1OGNqkvin+nLF9nOfBcWRlGnltPvFlPG6w8x5PpCnL7iKC5ZO4r3iCUQ
OjarAwrEK7vyZWfYF6fCiyoNx0qG/GerqWg1X6iIxq9frU5LItt1yTM3lTG6h5scgSMenIyCY+ng
s+vltVawI5WU9ckAdJOVk/9etPs44Ic06StNjTRlpsq/XwdcMJ9BgskXpE224tI77695mSyJ4+kg
uLqp8c7TVcFzB9gL7Qqp5/8oBYp1qlYyvvTWuT7/IhGfC4SJPg+p8xpKxkdUd1a96BXuZxXVd8X+
hV2mcOxiZ63NdK8UJNuh9zYCdXtAAfbJAB2Mx4U5ykHHWhsuW3i7tR/RAwvDvoTUDsWAAFNuZSHI
xCJ5Z/feWD9RI5iXDJBb9ADxZJ42qBUDd5F6olLWtJpncHFyWqi3bEGXzBIwTdkMdIgd5TmWvv/B
vUeQftjKIhmLh2ZGfwNqaDt9qQY1Dow4u/U8pj9F7n+fuuDYlM4920x6lpsZ7FwVKcLJbfNbMRU0
0PI7Qd4WXtZGA/FLot7o7zeNt4rHPK6uMxbg2kWZWc3U07Q5WrmEk1ocAnC8trAnYov4SMUa6CSM
qZYzHnQZRVu5/WC4NeiwCAPQnRwYJxc9OW9Z8CxA+r40aVhrfTytkQT3bsizq4QlbQBbBoAWKvTF
gfzpdFyIyBu196Bzt78h17vv3FqDazvsdHjzXoqDoqA7SNVyUOEaEuPnjXiQr3d1dR0y9KPgWjqJ
mAIJJyE9hhSqap2/GWLyCY8uZVrGsBUvkfwf82R7+AijX+VxaGFIDy61kezJnfPwWVtK1OYoMoHG
wTYkQn5h9JTTNYvgKQx5SPaz139ZL8Yc+2kPGIgSLT7F0Jdf1xaAyHGCjO1alwVf1Sp/kw7An5QL
1CNQQKwnjTLiz1L3P+qrFlmFaRKUG9XE9wPjpK4=
`pragma protect end_protected

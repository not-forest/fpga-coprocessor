// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
B4bLAgvotonVAPpcraivh2hQMNoV/0/Agxqvbx1CXIKEIGPxYUZUybsbgUMYh+Sq
eUp1mwaU5Ztoruix1zlMyFK6IOQRkLPAxpDxsbmsFH6vPA6PKkzzGFXOJow89kYk
py1RIwivzfmCe3aRumvz+inIJdjRTMhXE+oZBbvpOE8hgQ75Il5z05UCqEDGvePN
fxNh9/1yTC1zmqoJ3/j+DwA8dd9gFXqhmnwgltmuf3Osa34kPeeBOXZ0aj+gbMSV
/ZsLQhCT+0Jl1hsBFkyTft45EbhZO/YVESSyYOS6Ce+oLSiw++ZCu7CZfDO65thM
2J8vCkpAopl324TgoM1w8w==
//pragma protect end_key_block
//pragma protect digest_block
lXrPhwYjyfgghhUQMX59Cv1k77c=
//pragma protect end_digest_block
//pragma protect data_block
Y9LQxYvUscuMMYJsTeEJOdzO8OiIqEygELj8Ks9AWoSRGelKU0NDHLQpEO2BHqi+
K8vPegGLmAMxr+wmo+AhkIZzuOHIQeNcpi8YMJDRNPfrBOK7/FidT1cNNTJ7+Qnp
/oqe6mVo0+Wa+YVlwY4l+5AHp6zW73t+ikiq09kNGa3F/ZG9p544zeLG0WnNYsMK
YD933L1uc2uyrNxyIRMILtRCD1UvjzdPKPs+Ad/0O4BI4ge3R7asvbyu4L8DNOPh
5cXvNTg/R7JKR7Dg52K4QmdOYmBPf4ihs/To5oYoP0izZMBYnl5y1+XXLJqkAZuz
IOgi+QnVclAe6BxKj/4HQf+gT2V1VEx8eMr3YPEfDv3B1Rzl9RixdlZ2DCJ4KqVL
lkWCVqur8A1hdZnn1mfHfNU2oguKuCD8eu53QHIdiyPiDDs1gZcdWPqayGmdZGWL
oRYOuMZXyEEtnFGIHanQx9YytxYXuFNJ7JfQ3+K1iO9eDPdz4XY3ykQgnI7CLvkc
PZpZb6cd1IfdsTl5/cH1+YK0GPXTnsp/d8s0GDhIBJ4aw1Ksq5Td9vGHdqWrmIbu
1DeumEPFC3FINhZ4WnJoviVBikDmzF3D7lcjud0zQaSm30eaGqIuFhLj0ZNiBz2j
7grlazIoCt1m7CNwzq1U9CxHi13Lr5hPKt3AYYDZrS1X3BGeNN/vDPtHaBRt+hzk
Cd9d5K36JblBb/ELzcwDTiH0prZvIaKXC0CJky9ozvgeiIqVNaMzhXNjPgGMDlvD
GsJn4XpCoUjyemFbf0EwqEYGi6j+Jl4m+B17cChy8lUkgchC4aF/Xi5SolatzCFE
OB1jOETEbKvVTW7hBVn/fqcIgPehDLCryqPzztG14PfKeEvsRBhALQBEsXAE1myQ
IrqJJp+tpWt5Yw5Sm4xaYCx2JG2MKWHoknkFc+K9AReRBAKFcS8U0yl5sOKzlzxy
zHhNIFupG06gWJCtzsCLml24IY69JbgED29AyQcorhEQqsI5s3uln4a0KZUEkHrt
EcLptMecpQ+gnyiYRNzT+jDymRQuG3kwjlurqMo3Dta5f0aiXTdOxtcH7cABX+fz
SRtg4oKcTeBytTEIN0krl3k5w1uDZZonr3Xwqsuqj+VAWXdYoKYbG4dHy9kosoLj
evpe4JoGADunxa5nirEM+e2AzW04NU+Oyfc0Fa92DTnMzidEJDBVxKreUmJAMVim
YbXWz8BWcJvSsvLG34m7tyMkkdcVwiV6nAZ/ju0dp01NhOwKjmv630ZnhLnRpnQ2
o4lePzVNTr6rLYVe6A9R/5ERyPvjIdQoLYyMjnvXY5kFDFKa6HDgLaBDmST2dMag
AKH37oNjZg1BdN90dWj53cY3cOmsQ3NCo8F/y1RNDBCJwG6o3I3k90ZDc3KyRT37
SqJp8m7qdGI+3XpBx0B1bFsseYTlvLF0dCER5tbjSaWZul4K2AZj5dlLtrA6Ma10
j/NuVL2dakM7/66+/FQA3p5h9AmwTfeu1cykAvarqIWGoKmKTSqUPBZYcNkg/gZP
iFND6jrKSyQpw5Ge235NOBIo3b1uyfV+OfJlZfA9s5fK6YT5Ger3YLCWjxDdBZgx
dsTmu2wIiwQaADCh1lxgrJn/6XhOnRncRCFzq+0bG4MEOEqSSyiUP6/S2+kOaQW8
ieXr9Fwv2ojYlzk8TLbIfk32ML2rb7dcM7K/011a07h2jpshTZKtrVyTBKwg7U+j
/bv7iJdeNMtfv76RRk+dA+ufLmL9qx5yRZNbdKV5RJBl2+saG85ybfSF46pqBQGr
BksjVfkdHGc8vu1xMiK0eiFuhRL6thsuV7GssNaeGF//hUma492zdHkjft9d1+vK
QZmZtKkINkswPlDdhIN1ifdNgOUXQsLliJB7+us73Ts010HfQ4saD4bLPWRF2dGH
F9EDP1jUUNJxcNioZzlWFIi8LzxIoAWcofoq67Y8fRHlskfuMcWXc8VkOTVdFS+6
yu97Pn7PvssDN3Pj1i5mq/C8/n2eaLJwRxmUZZDmjXHxME/BJWhLHGW47HP7Qqpp
k2dC8+lCMxQSbiTMnl5hjc4LoOoodQtv1VgPS0x6vgjtdDx/6kUqqO1Oe9rmTV+1
7E38R9DrGSli/lfc9KBy/SGHXltGI7XcXGY5lDoPX7lySLB+L+YbPkk6MWVtTKiu
sDLy4/cVy1Q8WZFTnhuu8tUSBcHXFyNbcoDOrMsc8VhN2Q1p47luoWfSa8Ky677l
QmtQvLwUGfKcu8KPUNE+1aOwCPkDycGTzkzt8ck6AgDvotXIs7cNdYDwT6AgqS6r
43xgvGL+8bHfwOnWk+9KlzduGV/1BcmlCNIglFZHNL/uqL4LP3g6GV2k8KCXluv/
Hb/kz9iarLm7vABiTXvo+MYDiriV2GfQD1XfL92iXggyCPjylHQLuZwijxCn6fao
M650B/vtQ8EAdwxdk8puU/732nT8MpoEbzWgoVaghkeM0rnBJSZkbp3jF0Zw9TCY
FSPKW4jndcsJA7tKU8YxmwIdNHfufXcTEXueChluzW5y9dQ8BJWieKFc5O5EskZb
sKZAqM8XqJwBiHHnGptWRIVqrL4m0iI8pzZ2U93pFHzUT0I8SynDCFKsg0Jvjh48
9jnJay1TrLOnF4VXu0PPRtJ8iKdqacdHntfM44FnTPGaCCY+9F15//+xc1aWvyk8
/OM36faLLCSW8ovfSlBvTchKJU98tYILAelyHD+UkNINudlBbpspaL7QFuwUsqzC
U08tNTyURpsR3ylRgB9N4jDFQ8xdaNiOvEaT+LXQqHGPIC/cl+9Sci4/vhD8/QkJ
CgEkuF3/UxLerdvZ3IvPeRQXoXdUp+9mFIlz6N113OCu8TbvGcuL96pjQsw1+33e
vcjhrvgxc9R/z7+scZFUvN2QqqE7z7O2F1khwrnT/0w9YO/JIOM1Dyxrvn92IeT9
McpJ7eAz6waZFp7QfVgk5clEYnZhBbc+oylOWxJDTChsnWYOddiu8KdypOpsT4NO
+t1Y5y7qZ7Lm1NVdClsNSFQKFHduMcMObkLe8Ha5wdHKJCWSAMnRukge+dDDfTTM
A1G8yEprU9ecZRgFXhfyNSzZBmbWdEMpaApuTTddKJJU5ZqV1F4m6ocOE1AtfStY
pbcKN0nE0BSdWRw1X13K4mz3kb7XZbA9dtvBjUT+bX62ha5jsw5T9Eezh9sKFJB6
hMWCUpaPgOspTvF/pwgIJK/zvQ50O+1Aar74Idh+Fo+aviBetRDQXbZC/mZMm0oa
NfwV63M683iOee6yQwY/7sDEYVYkUzT1dobe4eISIxh7QN3CzjpkqtwysOcdxRcs
psoOTRZFpFDuAgjCyXzlgAZqSW0SNfniqeLGugm5OIf1sxCzcX4TUSVz9vUW9aXq
E6qsquBUyXy+1eZ90znLHRC2kGZQbbl3V0ZzILlZT9Bhh8H0L9EQ0vAa6kUZ3cC2
hM874AFK9GjTLMgWWZ56E5Rk46lAvOtEDKYVrl/+O3co8g+WSlZ1oU91rT8iuWE+
JJpD1Shh447DK9kYOXaOKtLVGVniW8v2SD1e5G2SKrnSKOjLfFi20TfZ35f23Jkd
SjYNbSZdMqT+GGiYy4xSdxP4vRslKmmFO6uBw9hhlkqUsBXhFVSM52cwajUsQmy4
Xet6tuw3X8NaqizDK4MIARuAqV2lFOR9S1cfmajrp6atl5boULoi7beT3LWFHptC
5gBVI0NFrGSI7iYI9N4r2A2AD3nFsnwq5A3LkJ6YE+0N/PQr/9h8g30GYEOI+Ipn
QROd4XlwKcTFsJmsWuWCfZUQOqlI0OEgpiJKrNYqX27Wj28fkFqQdmKYs7dKpS0H
nSzOppbXqZ2iC0Q/l2jdMniSVnw8BXU1DuDjDR3bboeKKPnfgg5UoqqbIeLMxcMx
Xfebq34xtWQFEVOSsSJlfTvRfolKFQI+UTjJgtrYe4cm7lrhki1NbHydidkcj9H7
a5edr2RXqpWJYhXfF0xPog2dkhEDiOXavKKX65JhoCzovr3U5akmUjpckrU4GV9q
sEboIGCo/Lji9cmHs5Pr3ferLg64dkiVjkWciYx87gGyEOcx7JwwjBPEa5fZCMJa
ynXd2BF2yQ09AcfJ5ggB8IRDTLSsKl/YGuP6mwh+HSvlaCjCWB6PkvDJhuLE+GCv
0lwIx6BtaxVcBvuQiIbYQQ5KJDfO4esVbsMdpqe/K4qyvtGuRRC0r8CWpvfA1u/I
2gl93pUR1mFqQLpEG4u4eCt6Zuz8ol3sWGL3Zmw7cK2o0sHdin/8gyKJbGcxqheV
WaD0snpqFbsipFp5HBp6kyjsUmtnqaWxJ+HzCOVzpkhftWxHwSHqzL7NsyQEEhVq
xikJQcH/G4TKCehDWYfrYTkdbUiYQDPRla3tCyWxFiPBuq7FNbNOk7Vk/JOzqN4o
4ZDRIjRCsPUW+zk2MAAzdr+m+LC97KwQxtw0VZAexGmfcBK6uki0DWx5k0U7zzxn
uDJJ7ZZCshwFpAtknavY8JtD89J017FGltrofHCaYcTund2Ya/uVQs/K4mHi7m5u
el1IIq0C+qK3KzeeQaMY+5lFpKBm9vajfxDY8+Ab1C2JtpqOAV9EoZtLpCKt9eTC
SYdeWFEdl2fELXRzfqWhsrSE//qmcGCDURFORYR2QLhL+qNpwwlUywdiy6e6lCsj
/9duLGm5XROKj3d10rdHFMUpvjzLDYYtTC4fjLzHmFqgZ2qx8F8jaVKZKRGFDoFA
qUAJOd1mf28r5GEgW10nSZ6TrqbJrwG5RSyZlvaSshoBVzK2LJsyxrQMWy0ZtGVu
UGl56Mom9luJqEYlSQoWKNwYU9f3WPCcw+BVz1NdES3egvi5mtVBYWRFG2635Nzz
3b8h8caOR06Nv8afBWXJgxbzGNIO/6yh8tLYagwsSu6qTia2kB6drzl0ARS8hURb
bN6Q+gFNYRAOk545oHx0G9zAzngYpULgxCjesrlbIC1h2JmSDc5r3fF/TLU3SuxC
gRsRZWpWeAe1BV6huOp8EuBpQuWFv50WAM6v9eRc7AkosDKZcV7Pa/XBzCGCF9zk
COIBc4oqKPLuUCsnV225Qpzxm99PcKH/RwwC/7j8oITVTfS/xYH8diu6Ma0w3ZNR
hDWpwPJP8TMcwQ9TjHofxfM1uJDbHlDht8osLhfUEtELFnl1Bso664sXN82R2zzp
vzMav9+CpQ/t52VL7weMW88dCB92/+czh+JgygTT6fh/jmdeEcQ/9V9YIpQasxg3
FCOsTuIwQ+M7sXq9wLnX7/r2jIbTKFwKCXkxyhah4rWnQNCn5og1GDW4WtHS6tA5
LevicJD346o4xLHejGiNdGNX6WN4cXiQpuDMxR3xvm/tGiWWVCBUXCDgw7usu3vm
41qyZ6/Gyh4Tbj3LX2mctAKDed4LGidDR7ufg6ANV6XDNyYhL+iQ11EuCNNsEi0X
6/WUtaJVVGf8AuIDz4Dzxu7S+daf5HggRU/BVSN3+Bm5XASaQjzhtNj2MgHMW6Sj
8I6hAleOTyc+ElS8da0x3Crg6QLTg0R//x+aoP9NO8h9xBBftqgz4FnxjBeDYpb2
wLmfl1WvJJ+LCbZs4W8ZYO9FC+MAT9Qo3dAUm2UqEKCBQjrgtCYGqdjP/YWDgGf+
dHeR6UlwLURYqlsdQRzcbkD7Rt+Iq/zUxotnj6xpida2pe5Hu7DmO3YlLscUkFYp
UzTs0AmQ3i10GZ7C5BfX09ojkaX07jhrfpPc+drB+8th7kvDeHKFKFKUu6Pc1yY8
DPgmk42KE4nVhchMWcEL/RzvsRIhDDaUUmjpIdMWEca177NKXLXyJBxXzz8gkWEn
HIzDnRAIAWsaNkV1RtLWzUTvbSS+l58CN6+Wo59JC5tbWXNhZOxI+5M5jAj9z5S/
zEB5pjzg6+45ezCsczHqGbFINE197UJTxudPr3TWxC+4+X0qQccCJbQQv0/CN/nr
eV8oM48LWDpyUeYzguvTI6GmghIpru2KuzN+aPuZr4PVjYripHyMopiiyq1p3Otq
tQAM06FhJR2Vv5/t49ZU0v1X4PF1rTyw/Z39jwvhN2vO811rt3WBJpMd6UscPkcp
vEceV/nrmbdKIzL0f2YpUC+X38D/Kvd7PqSuzisqIwA6b9iZixM1hTmjMnMIt3/Q
2xN416Vslmfa2IX2BnpDK1wwuGa8C/vt6ecMHRiIRt5UDYA9a7h7a30MugFVPuw0
Hgqv/E8u9si/AFu2CtkMDtho5QNItTguGxwVW/jj23C7ZgK1LXjPxRzoLJXxdoiP
vROl09CCCtcNbsIX3Y1ZDWD7U0glsURu+ekIH4XbP/emsXgYCMIPl+F6KjD6avpc
AhQsqkWi/D1ZEIqf/F1hlLOFs2hpesBnoen/zejohIUH3RK/CzNQZGNSX3teJgkN
ax6YNgfMOSPK5o4erFr4E8i+d4fbfk1S3uiU7hhG8FeT8Y13XsR1w8w54ug6bU6q
tEthmFfhH6xbffmoHVrhWK5Vtm1Zn7f/+3jZfZRHtj/2RDuZi8eq5WkrD+1d+Oe7
1R3GSz+C6iam9SnX0WF2PbSJhN0t3bCYbba90dss2Dk4CjM0s1wlumcqreJ8zd/u
Cprq6QpIVAtplXlobEBXBgt8UrZ9f9I1t/dtTt+y5uFlJ+gECO/bfJ9C0SOdQiN8
F66UQ8yEMgijT6ff1rjuSlBh8LP+rSQzH3AnaVGzeJ8w1bsim+5FwRiuB4tpWAMt
a+wMf4djftx0Y/mKivapUDV88NhlgrtLNrNt2ubJ91CXUZaFObVpOChXRXArZuRE
sohuPbscBNz/L9OA2DB5oNhso7l43D1L8LluZlXsZgdRSfqO71/MMhXerlymsmnJ
YaJ504RCfIU0AuJo/y57F7bzxUdPQGN9PNods8hSiDpwmF3codfqphAKzTqcP62o
GmaAeWjkPZzi/VcfyxUUuF5jP8zNkTZpjipeJX09AeZ/mxrp6lk1HE3bOwRiNJcM
UDCpEUp95gVc1/BOfWwa6lUhDR4KI7IW6jfXoXpNcJ91IkvJoq0wpSO91VwwOU2g
O41+UOgVlvoj+CHFqA7o7DmhPOdb7bQYEpCe1ZufR16pV9kKpks+xd4B2/kbtUDL
rU9ISoKuZl1qqIUq/YrbcbIJA60M7q85nq+6Q94PhDj1Gf27+aoSyIwpmyN9CF/z
6NFaxpz+QuLcSYNzdugBQJmcwnpa/ouCLgOn+mD5/ScvGYjeK0Gq42BD0ryX0OLN
r/boUwinDpKgWmczp4KG3CBAwoeCivac00sAc9JXnZ0bem4vvODMDalyqPwPBxkh
JQyXrchcx/rpL3dK4MARskko9KuPGr5+msr8rWQRhko8J2d3pgEMzRmWHpiKEv+9
J10OsGDsHx5Uhg+qbXaGSG9iUM+cutofbNiC3AASREGusIXTiowdd/wmti2PY3Bf
4Y+Iz1feqCLQIADx8jI2iCMUq084AqIXcCD3Dee1BQEVu4wQ7j7q2xSNCErvMKDw
bPyXwlIYEbpusbYt1ER3psm3iIJCkWIio9f9FnbM/EP42Qv6gvGX5l8LKTXMfKiB
0I5/eZ5NRvno1JnXQq0EBOz17E4aR0VxssKE6qWMn55e1L6sD0nRkR35AQImuqzj
Jxsy5U16meJcozazXSy/K5cgy1bU76ZvRgov8eo7b5TFHLEuaONc4KppqzBURMCK
j27tlCt4FO+Mqzwk7OP/UVI67nkoc06eJSFDSuexsZLsg3eaQZ665RErgX+Ncjrq
PTXVJIDE9KdAQ2areQ6NdDGmPADSRh36X+yah3jTFWwKhrSfHWveUdT3Nnd70txR
R8MK3JzEJxIFTvw0PVuXWXgwiNiMZ0UKDhvm7qS+jL5nr4XayZxnRoJ0G/HYYhlp
Dc/ymA2C2uhTqLjkRj0QG0W4lInt+wvUgZ+MsMAcjxdgZzmAOPrrnc+nMHZAr7JR
71mLth94RBjLuJtXQ5tisxHrVo7PQu92TsgzqMKaaRNnGwLB+1Qh+7NOwkNOHi2A
noqFlU8h+B7lz6jzXPqQ94vhDypm0J8/CEsaWMroQaHV2rLSsROrdyH4cGpyqurb
eF7U8BzWKRgOa7ScOaPcfn4YR+x/qqAV1OKSjX/EDWFDw6Ih32+2CymNrOIeqb5R
Lz2aMx3ORsHZtm66qblV5QYwHnRkfyZ6aHrQQImTTZk50o9YdyMdmHAo8D1bfEFC
bWfVZetAsZ1ALLgQJ/uj5de97Ib3Gl/8EwnauWGVtzzZCNKZD9ecHr0xuZr1PIlz
uzYF6Dz+HvV4a01V3xyDAtlHgFfc0nvo9jt+DEPXrChXGDswm6TnGucesH0YRDhw
/3qF32Wv/daNx4o6oaRLBBjPbylMG2FS6VdjE0O9+ukQ1r0Zo8+uE9h17Dk8d5TN
8COlt4sTBkHN6X9cpe1RVB1ycVEieOiDpfmUC4FC4myKcYvMRcpvjf2tJ+dDJ0q3
KZ7FRQwBe+TavubNWmuRnXdkV8YAfh18SoTWMSTObGLmCANvVlpxh6JFR8950RLX
bv5uxIETfo1KuMaYZnh0clAMFw2qv9/wXMZNZwImtC5oPD08XaDFTb83zkwmQh9Q
j+8Wkbg9EPRFyaOFoVKoV30qxy3Q/XU0Q/wvRxtMHXlriDpKVw4MUze2RCwjfk3c
v79r9h4HnPNEc4AIRqUoLoFrsYqJSaQ0VR/kPsk0BfLo/3BlsQRPq4PlaMiWkbxj
PZd3nzaGC/IE1Ksaonm9Mhw1WCUhypttpr2LpsXq3daA/ojEmu3QXwLax6n5tq8g
sIKYbw/5DXFghtuOZXb+u/77vYMHV+GJ9Oq9lX8s3RTNBPTNPdKGY5k3qLdbeyy8
0vME+alVuWNBrPFJwzKKhMXue29Ekb7qqo0iZEZLI2tWyJNf0/8Qq/VmyLyq5tWL
t+rrDP5LEifMbGNWTkiQfihTnfv4nHtJlmvo2/mA6vQqU8DIDxHaEm5i1C/d4rtK
QD1I/+TKEhR2Rdp+sYFiwH/ljIndZeHBMpj/U5QBHEkI8vz03iNMQrhVfPtB9Rzp
a/gFr5GwGCEEGexUrb9SflVMY3a4L3AIsTILIy8/3WmYExvRL4cILMCvn6ehaJ94
wRuUz8M+IQ9RzjMH6S3ch0jlSlaFsxo7MJMSeUycdz1VrSrtjSD2yWHvz0rWTgX2
sOp8oE5WPk4OywaR2Iw1oTzYVdW9H2RKaG/DY+nUKseyiKXN24daOu9EA0OVLmSz
yG4r/EwRSzOCtG3uq3pRWpbV4AM8WqIvvmK8zEKbMBoG3I3jHcFmt/5RVQ3C4vxp
KI0Z3SevrtoDd88WemhyHXaA4OZcOV9WKrhjg39lID5Reznx78XhXoAjOft67ymC
ifKy5cgcQRn0RVcFxbY3mdv0bzrveQt7U5DboFBOoVVhat9z7kRgNDZl8HykFgwt
V81iWEtmzfLaIhZs6Aeoji+1wVME0135CV0127wM0qeZB1duUpV8SPw6HmD/4cwW
4XuXOgtNF0In2jvfchlCz3abjNcvrezYSQJCxj0HrRGk2ZPyDuuGmJr1JbmYBs96
swyvEtcaQ+T8NyGSBe4/hGyJjFWApef5JHSHTQUDPedLACx8Bxm2Nkr4G2ECH3IS
Gf1GN/w5N9jzdeFDWqBz1L1g7cLGXZY1fp1FgKtvXCeVoYmuerFYCnuoi0LlT+k3
zjcBxtu6DNPLG04JZhD10Et6g+qw5pkCJ5CK1S4OZkeRdo/aNHrx0v4zZabjDIGl
qdUl1wqVEvDft+ilpRuHovhtrXz54ezdjg8VrrNeqyV26nQuP4JmInvNIAs2QiDY
H7JX35o5RNUyBfF9kEnQkm5z34ZGRT6wlew8cPt30uZDszIybWb/Q+/nFQBhO9Ja
QIq8qrophPHTCmDa3+WzammM+BnyclKFtkEq0wljIZS2lMzxsXYuQg9gYPHsqzPR
QCa88TJ6RCwdyRu8QooAnKQl77ji7YcoD2qULinU4Mt1rmrdzA9cyBbDYjW0ViaK
mj2RGMRKT3eNlzrRhUZMMmDnmjnaMr1MXV2fGtvoeHcRi20JlX7PKnj6AOTBEjL2
rye8lDYjNffu4B8YnqtSlZnAWtQG6aw7KMqDGbwGAd8xZslEIcpHYM+jZcb9BLpN
XCJdAl5jtIUC1uF20RIJ71DlZMINPGNbfB7q5tKYDUSCjAW3LTIpcbgMSpTejkir
FQVU90xwBFQlcJU1UNdHFUnlSS124oH4Ws5VXyVHsJjkkZxoMslQe8o8it75uS4Y
aoTNaGYzSreKEDFxnhPp10wiNNPfJ9COfMFzirRqY8p2QACHM6JlLNI0egP22+NT
oaaQ0rgdNaU93GqUWnNtbNmbdiOH1vt6UooYZGkHlZlBZIEJopkM0rgwUAc/1UQu
NM2ky7QxiQp8xUz11PIUMk9ffvyWpwxoj4iPnv12McVhEwlduYh2rhnrmrGA7GBD
e2N/InoCP60NzC+o+WY2ufP8qzkIzzI0ec/CKe5thJtx2nlMD8/RSPP6kyQWLLNr
6Y6IXUnSa7/F2ss2E0UWZy5KlFOm2EMTzJjFQxRPgHxPCfR5zOH0DY5RUpQiwYc0
69pW9nc8U+5v7fZab7jg/6O5hTpmq4PYqPzk7y7wMHOepM/H+meLGhoxq3I6DX09
xv+KNwo+kmgFQ8ibJ0m210C0AL0SXprIOHNB6c9p1ilSQ7vt+XyKWQtbvPZjGeKe
ZY0m55PPe/m3V1VaM2VQz/M9lh/y8lFBaJ51+fT1USrImntxs6eiNiOhzNVvakAO
N2PdR08ZclLCzt7+z+P/PWDe1EZ1clPJCwZZf4fnIcNRyxDOzU8Kt+M/3eqaP/0f
uZtWe/yofCpsFb3hDQeM1Z2qJlS8EcfwD5jguYVFi2Mg8yf0tbwujBuH0jsf4EWl
J6q3LAqXxqjk7wIwCIsJBXVYBiNf0SRuAVDOdbUjkWvw1nuv3q4sCYo5+YcNpBU2
oB883bcTQH62U5bBiyRWgflV0ZBjrFouHQs6zvAZ13SZGZtQcXqjfGR6UwvU/Wxg
fgb+p1j/wsheoBy0/Jd4ETIw1Wdy0dj5dtX15Qh9OXHfjmkAQtlwNSYa58v55Y8e
j812IPtnOxYVDRpympmKidbt3BNZylzLb9JYcL5+ZOaSACSNraW9lccjj0AsSMDg
Ml8Z+I3Qko6bQqjNmNCLvNsMW7WMThQZEMwmzX++/EaQIXD+Toi0x6RSFWchqmHz
9QgDnZsUFFilomv0/DZoECX5oZwD18ikkoKLzPmpb7GOzy3OIhcj7MvKVi/mZmgD
OcW+FyL/10obQep208m3VlXTcU0KYT6x0jcR2mffMR5gVeLIGO1fb8rksMs3nTHq
Ey2WzY6YU0701NV5ydd2VzXPQBiiRjFrxdL0KKJuRM6DSSWchMU28pbDDXwmIoHu
3JI1iRwE0iwfx7blWn7EN0Sk9ouS2xWVf5y7nJWV4bJZvAlP5KsOl7Rg50H1AhCG
ZKP/H2Gn4A7PKs9HJQm+ycXaIs7CpXOlMwB0txylXE8p9N11tHPs6atK3+2D2ey2
D6BOp0/OKMdqdKnECpsX0GGLOpHWqf3S4iqVatcK7sIwrEIHKz/5OFK1hi/+Shg7
R5RIHqokc6vQP3Q0fiEKLwu23O3GHVPEqJSilDqumc3bds2hVmt1tZwb9QN4ZRfD
GSaKE0rIqQkmlrlyX7lOoxy1OfpO0KGGm/IQJMNW12K+4FYmNAxcwBM6eqCDmmnj
kQdIaeveaSTzMqcdwYHFf4xxNq3zuBNlAM0KlmI2llsyx9retLs5u9miNygGjVub
FGKR/Ot59BoVW9bBwdSoZmJo6WJUpdEEyZQLZbSjcRg5QYC5hcmlcBFV4grHxe0g
9FAfvEbVG7js6tB06EnClwWVRY+W4MIJXeUuvtJfvIjmwtaMba2vIeSFBOKAsgLp
q9YGlC0CwszhUR1mvPxjh0wWKSCPsxwu0XcGDWquobple94DL2F3SDB1GJRMkZPu
Kgl/nHCbLMFqxQd+fsMZ8QbR7B89NKjouXfX/juywTyVnl21afl0sNPPzw9mt9Xx
DrrOJSvyuCdOtjhn05zLymMYtNySpb9ggYowsr7KIRpX6mDEakymar5unOZGXFzx
B+lcIHTiAx3RLIksB4/eH4KFueKknZHGE1n2wYu+Elruxi/WbSKz9+A3FhK4dDAj
3R+OQJhixgUCfWCvsAd6+2LnWFe+1f99ZKSke0hieWeZZTyv3eRHQxDlNrGldSCN
GAbHvJrh7OP2o/B2ohYtxW7FoTosgjDmAbTjFD3T2xbIWOYAUFVePxtLUhLdFyuV
caUQF2KXaZUPx7U3soFX1rtNew43fffxVQyWXzs15o2KKgTnDlMZTRFYN6iuDQCh
JYbvqCrdwwqrkSrR+VxSiBkWGmqhVFmYT21y9XT4kArBqPLUjwUE8l4EJzgFWBzz
R3P5dAHaCopOJKviRDEbLwKWZ/ZnW1g2G3jh2HzRkoSJTnP73zJrJRYejYJfSMn8
nMCG3By+GpIqA4ej56qaW/U5cOMZreTaISHPZtmANfHOV2qPwRm4xw0w31tGF+WJ
4udQThJw92TzAG/4GNGQZ+15b3f8Ye1Ncuz9Sm1kUYX+fOOIq0usi8bQGmUuBKQI
/S6ds46Zvk7dkBsri4W64eNljI4U7aI1evmlING9XYhBVnpmRzfDK3zJm3dgIqZh
Rh0Ze8iq+DJqQPxao3/y78Rlp4x2kv/xNUS10EKbticlQtFkV5TwhxenGXXAKWhL
sZFXmBWywTFl/2jjx6yfyumBu4huxvDi79H6cUz+UTw4xWCycXYZDD9fknGeb/NU
1nQDxfPotphvtFATOMMlGPI/b5fUGGHbnjLb2b3rIcX3GI2gccnxZjOBRh37reXO
OqiQHcJXiKY3kZWVo64xT7t7qr4Yebf1hqSD2P2y95yOApaPyGYEx8vn1ODGgbM2
7Izvq7XgRGOpBrX+MHUSfOGdNeAkLGcm5T2b/jKChld4R/NPtnXBkNXxI+EXM/nY
QsEBahJZCf7EQ+rhLq/QB6Mcp7flQY8wJNtoS6nuayQenj7ueCLDTMck8x1PPADA
GYp4g87C2vdGTgazOyj8J1xGyJjNTwsTDdTaHtSPVvSmK2vuBKT2Sx8OseAk2blx
gVU+Se5F5/XfKuA+650yOoPuHnylRfNx+oVkeCWiVFSO4qwZMUiqapyfW7YqjQJo
CVKQTUwd2FbKWcSmB8VwJnr60DK+s8uwdOEwow9r0ATzI74niDKOdAOhTNe9fSwB
0/VmXlCyqSaGXQwJZUuuyGEnA2hfdn99ZALwF/LCpWnIf29KEXFtqxaSI2/Pjbhm
DhFVBil5l9yhvmthQ/Ir1vU7TTirASE4kbIV+qrElgHxxR/d8MJ7c5mAFuIB0tZb
8ft5gwV5uLSNA/hvDhITPMWt/i1tqZgeeyZ7SUIfO+XOt9+gNZXOvpe5vpQDgVpE
uhulaAWy7lAzDXC1t2RyT38yxAzzk7RqCBIzSNK90Avrmnvr081R33dsDxpr/4Ym
h7OAmYqM7HP/315JAlwG0esYkj+SrFqGmWLZ/nhgxMjw5IEDn1OOgT1igOhRGfzz
AcMFU9Pi87tZBj/V1z2Q8S1PkM03G1bNpl2ygUowCz8Jah5qsH2YToiiHDo4frqL
JhC7hq9z7O4hqeFS0frS39laJm1FVHSGbR8M8fNBllW0W7eRtmSPuuBEo4ZpCqZp
1DoNxJ5wzHVur4RXUTIuuzY7Avh4kXhmwymQULIFKnK9hb0fm6W2T4SnRts+ZTfg
fVq2YhFtfmIBao67tLHwmx+gt8Oqkhu0XqWb6dpfcXcP+rCAiMNNb/WeISeps6pl
CKstAV/6zn5ISK87+9dkk9VRZRylMTR3rqojp3Q6oGWFFNDAXRnzgExKHQ5Y1of/
0B8TvPcVz/L9dvoknuNZ2sw7ccC3clhj1yJRKRCGonrvJCk2lUaEzh/hlgqWIZ20
dcFVyLGmKSOBUulz7Ysb+WaWgcUPN3iovjMaBHeCrTn/DTmWmuZGfzC0+q1G3fLf
H66hiICPkHH3Pp3WsVPkhFPMgi9ddfi9GnPUOQgJkY85Z/PU0EkinYy8KgiqfHKf
fBD4KI+3C4gnev/fjuPADE6nc5M58/hc9bP+9rDbmgJOBVdAbmQ4MRLuR69/Wqa9
aNgU8Hdt9OYSult67zU6vlyZkuRvId/4UUDBs0ek8/a/eiQy9vxU6QxuafWHOJjC
UCe2z+yIweofAIKph1B53YMfrij1A6qWTsbtbVXnZBTp0d/hLWXJ5c0UPb8+KEth
d0ESMTHdSDJnQw2aT/+xms9lXb5jTI8ZsJdhiLutvReWqa7J99EKREpAGZ+koPwr
UojrHTlKeSMW/6OaH9f5QG5nUDxFWIwcEwFqlBpuHk8M0Ko133hbeqfh4SIvxbgL
OOVNR+hjL2v3b9256DO92KBLuUx+qQ/vMpc74Ui0Ticknr8a8HHhRfR7NJsBnbHl
yk/pARhtY7j5RgkaaYXLOpOaauMNMc5G7cyMEw+dsvzQT1DSv3l7OXfQL3jUUGze
aWWeaGbbuihYorPXQ3JXEabznxg2o7zTIrv2tZUkV0Dbu5bR/QmNio9kusnHcvAY
HgG9gp5BtEDy4JJExe6EP+YDKdsujBpvx/GleV9cfu1T2VdrudOjNaY7BMRt/tf3
CbvdfK5dVmstRjVYwlllFmEBIJWtuQwZvBUlIueCtgCQGaWME2x/LC3RKlORLMUY
SarWVHeLpvz+8qfcGWDq7Nv2/bqtv0+BmbZPVqzoTtShhKL6Uz02ntnmC4YA73iP
2YtfeCsXYcl0oUcMK0cX8J70tU9XPbVqqpVF4R1hkHG/VhUGoZn2p0Aqfzvo6tIt
tA/+5H0f2WEOw0Hiz5gmgpSCk79OsJ9XykD246DEzgtWpfFiV6bpB2Q0NNidTWBk
z5htoi1nFCbEZN/0kqGRXPeGShUKeJxP30En7k7DdsDvsg7Ls0Qa00Lvp5tmIumF
Hc+sFSjwqNBLkbVvWLoQicgQra47ZNOKpqvcyztiHi75Nz9nN5Zf0bnkd1kEHAGv
IWsPNjzFZVF47iHb8DHfBsd4s88WV4dary2gQMeDMEFw2k0pl7vXaRN39D7+mLqi
n0Tc0JqMXkWZx2GTCEdIhqT/Lx6rHyLkw5Qi2+90Coe+CDMOk0UuXgtwEjTdmRA8
jdzE86c27eDL4835AnAss0txvqU2bsD0aWrpitLSoaYdXlYxR83fnAGZl8EIvrSy
2O6ebaqWMH2ERSgVYYjD3WTuvTdLhA5Zj0vTk19r4UUSYYQy2FoBKpNreE38TFoM
orRMoCFglyuL/l5T7+O0+PKLv7MF1nN2kEkU3fJjwh2y4AkpNLuJ+L7LyQIYJOwe
9Mp1X9pVkdHoSeDiJqdaPwexsE5fOm1V03YYh9jRLf9HnyutU8vb8nWJBNIlHYcj
W2/AALJS8wVKziwD6Ijg/CqDrYiguZzvguhrEKMLzYdvwyOatCgzx3opJxJQQJbG
6C6TmhcXhpZZ6MuJEQ7nUTjZUhSVu9pfXwtqDK6jrNt0IrewmQPyR3jFBIJQxqG/
9nInbeyNL4m3/DUqm9ngq8p+TyU/BKk1J8jboERHNQm/aEsfNLTtOo6orUYPZLYc
gcUp2knU5dvHaDDOb+uI5645/hXZv34llJyv2qzW6B48Gnqv2EUqq4KQJ0ruzqTY
Db/UUZf7Ps0RXR0LB5E+2Tp6QXa1VjeHyyXJTQyx8SxrdH7NH/94uL4X1IzJ5Wwr
jzJJc0dMnOG2es35je4T6MouIjY8L5t/4iqaM5mvR4WJbYfv3DFXbA/NrAP7Ta2h
tj1rVAxjaGehHoKlO57lfvsYonwWH0tbJn89Im5rGtkNdeAPfgJue2wXL2SGdbCx
04ZJkryU5A3l3y9Ww7X0XLGpCPFwiCxZJh9yeVYPIg5/XKZs4Z1WOJhFIp45PiZV
NPe85YUw08YE/Forox0SJuJJjoxgxT8S59a7My3kf+ZRLppOJbuZRDo1ECBnQThU
Gx8L/PC8UI8nV0N3R3Q1VUo/9ATZ7oRbKW7TDRquQGL1j5lA3IPPCB9NLe7Tk5wk
adSH5MMSfn+oUNa/0qBsiDL3wVnHJwiyhMf3a784mWKlNZ/vsA4dvGnwGXF/9UfJ
ghBS60Ulo1B4hVx9wIFON8dwWNrFjnNTXOf7kxep0VQYJ3Lv8MlodsF3cLOVyUeC
msZQ2ZuCpEVFKlj7A7eDC3CW1B1yLMLbcDdPiPRtXwIZsxXkvV3Tk7pyitaUmJes
JNrgaMVoPKSyivYKMgKdK1sSV1qko01UC9574j4yWsXvgfzjgtvteUp3qQhaY5ea
m/FtIR8uncUZv1klnekUjUYo5KOPL0OXPA11dZ4eEIGI6cKEM0qkPtcaQUwja/Ax
fqZUr61zusDYmCKhPcEba76uswj7qS3t2AqrYRv3Jhs8kb628aP8NUx+O5B8bjHj
HWiBDgByfh8OO/Wt5uGe41yijeL7A/fYtFTeChKyjkfpn7aAiRH6ke/Fae60Pumb
E9dJAyuBst8IfPi1oY9RZ0P9Ng8RKoUhljeqrP1Cw87COZIEUlWyN6S8at6O6r/A
DZ7T0gEXAxkMk0T1MyzoNGiaozPtzZGygZxzbV3xo3U51+c4sOARRK7Xo80f1lTN
gNF+2KcHaQlbHJcuVu12nbCah2QTZBd1kC4CpTibdpNqEZABNYwhlazJezASxRTs
iE0vLRBFreZOJ7MOivU72Thei9Sk2enWATUhACSEXDvz/OY4DzfpinWeOY2hdlYU
Y3+OF4A1yFQbnOLDL4Do5jiyEDIyoSYdd3+rL3ibdl2zy3pkDz9kjSablLDkMq2d
z9QtPhIbhofnSZcan1YYcQ4oBffqOWMrSqmeiKEhlEN7tEKDhmJPYlGERoHl3q4l
Dpr9ysTNy9R4s9QReh+tDM4iG51DczBh+nxAEDnfjNiifTs/dwE+cDOevfM4hWwU
6ihLBX5mF2uR3CQzn5tGrC59gwV7HXvHRPxAZOn5JljCWsI0plk23cMJ+jeDHn3t
vcJl3UQVO5m8JSEi06b2fhrFA24NKoj62aNhsxNTlRPIPZsuniLdZ23muGOM6uWr
ci+TU6qtgTqTcxbUvhSyAmjKHX6k/bLqzpfm2PUwmX0+kz/utYUbhb1foVfUr6yb
svy5ENZJdLWb+PxdSsS6djrUfpCHYhNiDLfC6ZpBlP2ProEDLVIt3+lkfQ00s2Ot
t8WAgxnuGoBZfB6e1NO0+iE5zKdnGsQY0tilQMbahHVC8oWdH7HcPzgh9nL6mTtf
r96Ckt4lUw1E35hdwIdxXtg+I60lGASesbkGe4DV8OjC9RdKCBL8mCVfaYJk5+Jt
1EAif9x8prP5iFsPAqsRFWafB5EqBrqTHg+bQilKZDMyvCIs0KzE+OG3+zt+L0TQ
VLb0iONrTv5wyZHtjNcU5ens+BRrWpIWWXnYM/CUYWz2EzIe6QHshYwrz3oa3NB6
j57zu3G0FqhyBvsNjLydECsxNw4weWUKpY7+2YsAUtHIjbhtp5/bYJUW9+8OPdVd
fCUcaxMEYMdXoYWgHyCy9BFS3UyHzaoAJcVzA3VdoDYeG3Yl9i/8zec3YSGW3tvB
aDWIRwQDKbq1kIhBmoQjFh1A5HQWK0Cies4NsoeXKgxGj6UKN5nJVR6bgqjZrnF5
JvCNCBJN4OL8LJcexzOiRel4kUxTS8pw1AxTBIuk6E2fUDCskHluHsb74jtppnV5
e/+EEPckn6YghvXjv0WOS6sTiOrxOKUBoJFHBlDl/XD8ofk4/StnFxxGb1oO054n
H4ejjtS+jDgA9Xyok6o6EUe7ZuVfMNCbMi2viW3nlZk2OhC1cm2FhEenFMzxhPtW
OofrpsrRpdcRGgn1uG4STbx4bOjBlabDE2TF9i3oSorGs4IjhNOGnwKIGLRX1+d2
ceEPz7bOwd+QQ4tx8xY5YA8Wq0XWjj71DBJz/jFr0hmYD9MT+YcBy+xuNQcfNcKA
LNg3CiivWmRlPHaNdnq2R9MHeFc/U3yOw52f+dDn0hl7gTLDZN/zkR64XzR/lIno
15JFFcjueTeUPf0ie7CoXUunoe9/v7PS4MW1dd99wkNiCYiS8I/LkQ22uIaep8hv
f/MtD1Z4HMWic4OkI5fuwSmvIx5SWamQMafYjfur7ywZZjK7NS0w9NjT85jQPqcf
n3bzMwDpAsBjm5ABrqkOH/i3M4czpjYTugw68UUb5D1jo+tOyoJDpzHQi75wV5t2
3BilvrH1XurhZqZcJJfZa0QAmYvJGuiWkRStD0+abSVBwBOYQoMS3r2tJP+BuMu4
RrRxwUw4dw4j710yfJsc6YeViBR+23vxNIWlWa0srEUSFY1aEyg5NGThEuAPrhd3
ssvIC/7k6syyAAMQAyPfDwtJR04Wer9il+6h55INXdvkowXaeq86kSdwVYBqBxjh
1cOouSqO7p44si0Iw1JwS1uXWXc6svaPCSpFoMwll0qp25qrLZcf+AFVLS2H9RNj
kQsIptxjHWa98vMl24MOWJOrPLRWY4fgAJqgVJshpT89RIOTmfA40FVdQq/3ywli
v1/S3KNCK5ex3cUN4pD6AMnoNCEH0tpuhNpXKdnl0A6451osinNBD+3nGAqgcLSp
It2K//LpIUys2vs5I90cIeBhrckn3s6WYxLmDATRy/i9/bw72Z0hJVu9O0Sppenz
dUb7G0G7WawmrMuXf9nnozoFjU+oY+X3TJTVeh8bB0bF/UDau1PJ/FtRIWnrynlz
fJfgQzoJIwCQCzQ8aUqMcwlUngRreNuuDtnUV+FVtYs6VBNOdAzUiyvz7fukoJ+5
qrT3oBXR9k9pB9+H8WYZCJnd89Hp5Cq/L2hYnbmg6M8a0XnGCyZTp2wYTmvxk1CB
oLYx08oqO1ch9gLPHYwpmtRC6KbLIHuYf6gCMH0CCEp+A4cPWTq5ONKVpzILIEPB
1jPE2dD10tngfmFWlCD5oPmIjVBO5VeBoYJY6kSrUCibmeJ3us/2jwIj2Yqm9WQI
IxbT0eBB0itIgZxYdfgovJX8wJPlVEr3h+I1qeHGJPAVNOBulwntbkn+tuYF6+0E
wv70pO+p3ZzeZt1zAzzdBfWqZ9c/joN+OdOg+zq923sQsBQGJpeiDg9x9otjwkAs
01Qu2AN7gc85SodBMrpoQB+jF+G+h0cix9kbOgTKMPb6uhJDOR1nEc21nkvpHhqb
4TlWXM6rJZmWUSyoj5e6k40riAiI18oCvApkqgBbLdJACQB1duyyvEl4wU9AS1TS
NtQrqKHuXtFSSbvInVbkrFBsQi1JtYmhREjiCaju+kIetRreYnqfDjLR9LrW58gW
lMJ55E1dOLUTjXov8HA6uslw0upvjsVD6tprhqg2n8aqQPnq7ubTmMqytfmVfWzt
UuJGKXQcKGv/InAcqJQYta8vlozKE5dA79ejTF/2E4yfsAX5TIZh+UgYbgIAQs9c
l7zjciRPUooqQR3n/+/pADTPwT/Lj9InqMCe10XrO/Hg45xMclIQS474nc4/naCb
znttHvumGwuEZfKyQG1sTmeNkGwYclE9x60m2PiGP011gmIcR14NWFMbPTG5dVLR
HRQHmSXxEZdHArmFmIEWQnjK8PFsaQmjI0oiOQ/1gQ1TD6gYxPpkNoGLREQK5zV9
wBVyrBBVajiWNKqh98svL6JvG13rB5JPj/k6k2JV1rEkFxNPltDiKexK1O5VVGd0
0QPg4oK91pgGQZ5YSoOzgeg85MHSzCvz+6dZmywl6JcBnUJrQ8C6TcPOzOEWcQ7i
WdxwSV7f2SXC2+j6mCu4hYxAz+1vv2CrhUdmz+MbfTU2S//Yf1fTL5iF/JHw+tZD
HqmweIP0HVsV/0Whn28+uKkQXjIpQ+R+ISkKsRpv+Hsq2V7vf+Y7iaWKxCe0B9VG
e1+yT1bn6rqPZr1fmiA6AY9hDt50WYFUUHbn7v4iKl8gqRE/UFfL+UG2lqY5yOzv
r9ZyIxaNefekPzTjKjMU0JavCi6BgApVMW/VJWQ669+HCunxqjeOljDfT6itFdxU
3ahWY+9FmrWjK1KfMd+c6egwyDXvnMoNAUYswuUEt8CGhh997gjPITxeVxaSLhE4
rCBOQ+InVn+GMYytdE9lnqGR1oSuQUWYyEO6L4dfFe+wHLcEPb8sSOrBZaR/0Ghr
8VMew9rN/a2vJj5z4uNDQtzOM+Z91hSI0A4+nd6LywCoGMIpusCcIddzLYXhNp2d
czvjezUNh56imowsHGEn5bOBNl/zFl9Cv/bwvqcm2OqDa2i/BiZpnVr6T/6ANYae
YUFH8VmNeg661yb01hqh9yG2axEpAT5lnb6bLY2+j5gz+Ef4LMmX1Cq0D5XKhuKE
aWmNooDr/fXMEXXTL113l6CHVYZTY9THomHcrhV27a45kB972BdIppq3BdDqsmYE
5hE7aTxg5dwOCNOZEb7jlRa6r/UGT+j/HqGdzCBjACiKk84CUHv6U5GHatgISvR7
LAxLsulUUmG366BTFKHZ2b/KVmJivxX49WVxNbqu9k9J0F5OccXcZe7WtUHglT3g
ECyfP+CMgdlO+NwT6atZaLp2MiyKNENKjKh+9WdjCI2BROVtTJUH+3AfCkQq+H5R
lrBrBtSsBlUvxsrf3EmscVHvFV4RhZ6veKPFP7EMN9Z7nV6Vtem4cnyLOYVxwMzv
hDWOI+i0AjODrHdeklFGrdVwWjeELgM0gMyLMCdDaZs02VCXG+B3bZOHrP9foead
n31pyWcFMK13/TQs/ACWltMnodntmoF8V+aVPc357efyzxveVWF6lGqiBXZCC2Rq
elqgGMtIxb4het1aY6LJx4JkIJLT7tLRol3UMyVTinw0q7YdX2e7hcAKa2PPMjS+
3O20HiSVfjvpWPCxTn6QN3/wHwwXhchQsiKORnM3rBPhiQVBDrNe5+T7nVuX+QMJ
iXkTqcGKtUtGfzqiGCcnmx3Q1ykMc/ZEukyF5W/rZAWzejIUYRUtL0LTQzAHvF7T
h154/SgrEAStSWg6/2VkXd6mwiu6uIY6FpZCGkIfEN7fma8BotlgtFB8B8ryoFJ+
1pph/DhaUk8I8BEekj7cwVOgytAHBe4ym8GuRSYrSIGlm7sGVEiUMtuO+WrqqXBp
Ssxc9H9Alq0eaBVYK3ppjjpznukcviHKKmIj0UNuOfBsPbTDUfNNs+GPdFfpcUTk
E3rFC1K0xNP2up2bTZVmZntQdVy99xRuaaUnwGac1Pwh+YtDq/zqBzAGFAvODp4u
5FqMAE4sezj8wJKV0ygt7eJmorI2hYKhUy7d74QjUwAywt8UBT2VJJQxpIdK0TCd
jokErq+sFzakUou/vRFVWw8+SwSazOY5+SfFthFW5CDZii9pxQ2RO5krjNQ/GAlg
boFyuRSLgqzAlDVeYOmrJi+ZSA9wbFYOsLP6/rTdGrehnUrYOOr74BODrKIgWCoA
ocMR5DoNn+rKZ7fUlRyW0wXFIDy5Usl7PUhsNURDMGuUCzpCeknyg1gR7fEeyD1X
taC3gn+mzoueaISc5yCKuRRr/XCgaDH/mREZ6Lq6Qy5SR14yg8kxnySkJMkweOQi
HnLTbuHk4CZOBetDF+qjIT3m9a788nLif+QtWOOjGsi5/lOG5Fozu0iRRl0sDK+I
2U2vRdkKpOcIySlag9O6JAciEHCrdVGyAncgPyoKa00VGjoBfaCjp3b7vrJiJpGg
h0P/F5fdJcHrlURtaE9EGSbCpJ6s5Q8K5axQVb3DD6eeO6rF0YyKVfgdCh6tJmGM
ZXrdRTXPh76F+LzzHI9uylnipmCw78JEaTSgI2f3YFgcBfUEHvovnXQoKrRKB0im
ztpxxUy0fGKL2DlG3LCARbc8uiRE51tDiLrX3ddpEV5EHdWK6nkvDJKQvsEE30Vg
6J5LARBs8xSXG8qvpxl3E3Qy/iDQUYXwQpt/zdR7LGJ+tREiB1rTCJ1TS2+Xlk9k
5VPdGO0lhwGE2A7Rg3qyCtnQUfJklmNSwWG4C+qRDuP04rpJbVUuSS3WNfBjf0Ee
cmz0us4Ju8WgFUdyiRI6u1OEe3I+a7ybpI2iU7ZvyzoTujU5f3NpbIK7OQum0c1U
WV0kIuLf0AQXpHbr1PbHYAse3A5v4Mi8xgaKKPYVmjeUSgncQWmQR6857Qb1Xm0D
twK5d5o3OJhxv1X9ALcCOzpL1Z/nofzm63hA4aBO7WYaBysFbFNTmv9kxx5kWvSr
7NwFHodEI5nEjqHVkpwNoVsWCfNZm4Pp1RSFZRjF507VZiv2pFIh7Ftt2dROK3hx
qmfu+Tsj4LdiJvjhKDKnBLLguKTXc4QC2Glq8P9xkNKC4vi9GqIxZ6+IVvKAJmxV
W6I7skb+4zopuQv/eO7ngSicClHBnn128hZQl6bPtOYxGyfM8KR6ssFBHFjuKk/w
pRO45iJJGGZPeZMMI+hOTYwyIGmUpy5+xxnqH2CRiQXkUQm2xAcD24LTvBYb86es
TAx8VkTE0CgPyQXbas2HYrqlG/wnm/gnuiMfqgf6KHl4N78fL4qkYPLoMtvoB9vT
IanjoX3yvsxNpcMFllG/92KEbPNcczgni8R5vKKFQb+v1OWfcgSEkiLxBnFxE+pI
J2e418RS+6Mv6MVgl5hvADZw1VxVbectw4wuWqb/cdB9vXyhnlePr7gU4loPpuPc
rRxKW9Ci1Y1jPsY5awy8wlFw14fSnBXM3HR25G1pp7mpSMVNRe10F+CBAGLHAh/G
acTTCJqwxTvbnEX61KdUFCpLrBvt2NZYIL+UaVgDZJUlhzPCQi6VqzrT7wtghA+m
kmG/CnFFMe5ajN2fQWktRISZlLRwoQj2Pan05GKaTnOAVI8hKMuLITZOh/9y1YM7
Udsu3pUFz09NcrMFgh1ZjVMGcGDkxk5BBvIUn2nd6K97OnwZSB7O2wPhqx1nuR7H
3/axdkw+7qpex/j3ReQ+jgivj7Bfrj5g/QHEV5fzte9x7wZV+u4wiVGuUvjUFcWu
zkOUH/7RzDD6SDdRwXNrvfTknvOL1RTluqtjTWXEktqBDsV9Kl+ivZpopBM0YrD+
pvyJa4kVTZMEkPahrNWIKax84grr7DvqWG9W9bwrJ4m6BM5Dp0pZq7Db6JH/PP77
I/sVgLOp+THh4zVpZoR4TCMUJFLYS08CS8Tpyoh4hfd7Rtx4Lg4c9aktRjyDEV1c
X5qhoM9lGaXHtwgZYyDyncRAICUgOOdF64K+WiyjLYSPyOUM0KRexLOnJFWaYzc2
FITtzGM2ausBwSkB/DIKVda1DTjNdQpahdvozEuNI4qoJxk5FKzsjVP7n7dN4VAn
rvZeFjCR4zz+Uk7vorMBUcDM8mobHqPar/Sq6+AHHp9LZPk0wbkvU/ytHNNR6Y6b
o93J+7coRRhbZRxZTH8jv6WBaGq0FlD23pMxff9uJDL/2mGIAKNtNE0ZVgxBK78W
abiY5CjUo53KbA4yXu8jvGVqqKAmPvg/zXM5dDPXeVeu2k/pxIjuYA9Mm/N4j3dk
n1T/+JOWLsKaIhlbhFgpPJNu13YRpoDDMrJG050HrVcCt9euFZcjKom/uN3wmKo8
VCx1vdzTEZUFWU+2KjjgRIpecurM5Gs1PUsgY3IT1FR8iOY5tMTe7T3h+GwIvE9D
iklb1DmrqnhiIwfnO5w/HYkBTz01I0EROxWRkhdqAv6hmq7K7UwRpn4zbTa+fssf
5f6Hqw8q1NLdJlIDdOSUKWsf70QZSVKxqQZluWG4dwKV4XqWXuk/GSghXcu7r0v9
VwvjivelETQ4i2sUvOoQmu8q9IIPzmUPbczIdhmFJhSoOHdJig1CZJeyqijCR8xG
xohPoD1hGLqZAQ6or9BYjYGwl9GTG+qZJwbvnTVBIQVBte/r7M7ndKq1xy0QsvHJ
pF+13k0FBvevRvdFgK6XxJesD9f9QuaaDBD7cTkGwEvW1gAyBnj5vR+rxgxOz2wW
g5U2gnVUY3FVaeUpH0h+sTO/+xtTgHWbwJKFwqr7+SnEfeNHpFIV7pvMYtb2ROGN
tD7TvH3KdTX37o1FJGTJQC8+u5R+ViH5x9cltMlux99d/tB5D442ixHZdTAwz0eQ
BBmYuzO74MFLOEZJZbtkbe0OoysMiIxo+NHiE5r2UJwT56XhYRn6P7w90Uujy1tx
UJlYnwMN3Ik53IA597BYj5DriObOWZlLmbrUUq/a2hZ1hIXVvPawIigvd8VzBlYV
CPjxzo6dYiSJaR1gQ4GiltJ4vRQ+qS9YVtukmaLa+roMGj9VzcoE+WFY9APul7Fv
8WKpacn68rXqJaxP02jyiPz4UjK7FyNoNweriUk+RV56CvAbSi7dhFsZf2FOPed4
J+sWs5lBILnrBLIgCssfsWd0uPgEAf4aZpcsnFiWiFPRDckeoTz0Phk++08j7K50
0HhYDuw6WxsTtROCJ48ysERqyroy/RF2e2HfbacCQgiDmiJn5GeaNxNtTOH1M5F1
sCWdGQ4JRt02iNCP0tnIlAnHSa202r4mdtjEZwmPZLiXOaHkuiKQBlxWsMOc/Gtz
SKRmk64aa6w7OOX8bddAMNG6Wn7mzjTGdZWjyVa3j8gJ8vrybwBUXT76NF1hzfrJ
kB0/XgPm2kvvGe/22/Do+oE+x09PesadCofbL8iTlc+A4LLVSvyNqEa2OB1jRpWI
fkxe4xPRoFcWfzVXrpj81+6IQY3zw7vHNOw729elJZHjxq706k+cQD8AgJ9BshvR
xmsCVxWJR+d3tVAmm3Tj2828NSxCcr4sXL7ewXj1+/IOb8qVdj3i0M81YJSp9Bz+
CJb81R4X92m5lJVsZAZN0hLzkscngO0rmWiddZCpahyvxaxpPdWeaFDGLWxerfaI
BQb9ZtO0rhjyZirMHShbnSMYTUmVNVX5qLGOuOPjpTWeBR2IPLGV8p2I07bMzFGI
hxWID7OAlcPcDKNPJxbflVweSXMUEtkkLwHqUmoVwebvxUg6UUKvMXYxFfIyBxZH
TIwbL/6T+fKGpZXYk8aZMTYtALW4WE2lyDiLFkVVXQFrHwf3gm1WWpss971vs8Yf
qSG5UQXUy7+gMZJhPorCui7zF2vMcPraeTsAGhMy3OX8NFXYgsrR79zlW7YAGtWM
t6e+BIi7AmN6jB8FeEtnMjKQa0BmetB0DOEjdbBHjD1k2bXqm6Kp0cEyoOU83u6J
dymMVk7WUtC7+JhI+BQjtLCL2ZBzk5qfBH7fnXWTbkaUpDNZ3a1hqsk1AYoKV/DE
quyt4iY0AlzvegMWu2J83HPnht7wZvxDc1fUtah6gi7KZVQ1ZZNj/5F06dSx7a7g
tRMBNrEsE90emIgB1aQBLetdv4qV+idd0l5PyUtK+Y2v3uuHpUkAHHdgov/BZTNP
9A03AXM5ZNbU7syqDVCy7fUdtOao/yB3/Gp+QPPduoYD5nZkfbTzUpqoVOuSJMuL
M33Z9zE/RUzH82RaNmymdejM/7ZP3kd94Pl41R1qpyhXeM8Lw2U4y4jZA+NvbXq+
6NGByxXkwlHPBJ4LbSJt+WICg+O7JW3815I4DzeXS+pL5r/S/93EXJs1wJ/7LhC+
I3xi43ZUVcST02vNjRZSKtaKUUz3r/chN2mrLyUghbfCJUZ33xbB+j5GMVc0r1Z/
I/bYKUZl2JzTcb3zIWSI04IjaY/eGfnO8B/CbZpMJ0Hj+v8LRwjePG6leG6uxZrI
LF2BPaX302Ss99HJCIODj2RoWAgUjM0YUm2xV07dHnpGfggf1ThT7UW3ay7Y0uCS
QcvZwzo9jd3YBzdcDVlrp17/yfSlmwwVhGA0w7BeNFKgcu7pd8+toz+7sA5zNsUP
nJeKQJhjumTvAE+GcxAkNIzjwx902mB7LpYI3Cli8wuag3o3DVSOfb+fJ6kqWe31
8yI6+mv9impoogqmguoyMnBhYUDKtVB3M7w466lhy8NyUm6nwNR62xm7lnHlBwa2
3QxnZGFvrEwrhVt5wUdwA7fiLF2j5EtVrCvIc4/PuOIKu8ri+UrZkwdAMcXZ77SA
NKTG8taNtLe+WWZFI6krpFEhNB/rY580MN7+Cv4SV6EWPtLWq+q1cBsom6uFG2cM
pzkZqDcp005dAeVjYpyw3oX88xDahW44GIO4MuvLoYcQCBOcF5XCfZzYIGtOGree
wkvso7/AYKJSJX6FcgeIWQxLLmdGHH9PtDEA0cYNGgAQVcE3MwJc1LTC1YNQnYzA
NWklyZs9gEkQ7q87WhEDxHF7kbPg/0wRigF45km3QXdp6slSNc5A5mhvK88RegWU
aIdFZZzzZWhpB8qgROybv+Iq79hNTNf2AjCOYMDmD51nDvo87Hll80q69zLEm6Nb
fEMjt70gudwmvN/wto93jo+gql+I8d4G++W36dh87WIhfzPvqFntwXzLMlFSce1/
Z1umlgnAY2oyZSi81JtFhvlnyrm0LieVUa3JAfz8ExL2RDspJqxf1+fnNpX2hnII
oJsGReYCY9U2WW5IKeOcm/sjs9Jt9w08DwfV2qGm6isxb2MwkP15iGbYvuIMvdya
3j2UQEnKvt89cQiOareUEaQU2CKWSnb7/bRnYBiL5kWdTBuQJ+rp4qoN6FVHmydM
hfopWJlSKNdmeqU6KAFXkINGLRjDGlpkVq0K2vHYl52I0SfY+WkDGCaicAm3Ye0U
MfNeWROf6csO9gHb1Shm9qa6hTJHcXiRGTOaXAYXmeTnyxUlCYZ4gXb6t5mHBrRw
ASHLCtVE2MO0QBoAdrDU+cX/ZF8+vbJxW2sZf0mrYla+6LefqZ/QGtmW/0JNCcq3
TKj1wslzYc7I7DeZacvf64z6Fz+62/pS2rPvEH/ZqtbltNNeps8zGC2d1Rl0ohGH
MUACHui96LfR242WCSpYilRCiVZCjOLmz82gjOkuIMP0p+/NyGBGuvcAMQav5pCc
stj+U88j4cJ2gr/5bL0I8u0KS99n3gcEJe+7vbAzyzjxHWeguIydi8pVeVHQUsSi
sOp+pGQRU/7hINSkNSZ75IFvDcgEj6M8RX4aUJkGb4xO5KvxBOCcJAke0jGMqyx7
e8CA3kQa0A57vKF6nuGGi95gR3GLlNB77ZwJY1kgzbrS9hMumYEgk7p3vZKx5Qvy
lnpqza21eEwUGvg065AlvZ3CToU3nO5iAsD5NSCKYfBSQZkHklmO998Cl3gdbqNj
DiwVU4zy53AbLi4A9GQAhi6InRom8USNO7ZySvo8sGUbGkIZNljXI1E6oq9uREmn
bYvujxHRGQyM1ZAkZDepstyLOqTB6FLoPIM7VEDreV5wpqdRld2YIpeptEpwTR6a
U3YydjIRSVwkYt9TF0DflFE4pvmbRPMoMdjFUPj7dA19hgTeNqG1Jv4GhR9zQ9ri
wOTG+wcKTTsx6xTXYCEO5tYEvO/HveuWi01rYhQqNg9n33Wz6EfXn9PotAyC6qfT
TDzUQz4xbvMVtl6vIWzQbjp+AnCz9719JIDo8dB/2EETlP/wpVHORFcvB+7Wn98Q
tN7inSpH91Tk+1z9PuPxckY8POh0dzVsNWg+3VyGrdop1ifpSPQ/4K9zIJWDBhDt
KlZLRI0L6PNHh/7PHnJy7SLyf/xPRukXB8E5aWgAt242Dr8wgvwuXdwKF3RqZpeL
mlA43jryrF0fRNnGwlnhDxoSkchz+eVR0u0V+yWACGuQ2/aotJpHlSeNmgwtKfYL
d70lZnCQdXJGhdJ3TBSPeD+HUkHMZMr9k4gjwA4BI/lmaw0icrLewnjD8flBfjWz
C+HcSQMI3MMnToXnIJbO2wI4o2ICMXJb6gDI9hBk4uRVse5s/oWg1IMlvQ+A8wMV
tOxEKkWAoGZBnH6SC32qh7ajNpcZin/CcWSLtlyQPfg5u0OD7hJJFt1DO7/ap3/s
OsDMCV5oxLuKTD9KQa7AAi3ELizSEDK+RU/3U6ZWCy5EjaxuHCWRGXDNpxbMtYLC
XkqMaAWkjKqP2s2+bx2qYJj+6xoIL9lG6+AeWuRLIcQ2f6IHtuZWJnVR++pYWphC
36XLpsBc/a7Fe26og7Lr68kvGQ8dlTyOFc6O8/kYY0fE2hAuaSv9ipMe9jVN2uN7
nWDvnfAGyGKPloGQq1e9XR9JHBunMVbDq4s/PuDk8OtAytPuStn4ac+7/EVWIgG9
5i59i0XYSPya/xlO2R73rtci6U6BF/tCpHNr0bpB5VAD3kVAiK4HyiiLjZdm/DBB
HG04YpYyKyahOrRwLdG8rrqugE3GkjWSwWwezTNR+VrGU1q142tUQPv4iZj2DrDK
zWLBS6Jci2iD6dOYcjUFud4ye3rruWAd7r+rqZsZujhIzZnduqqWVA75AuklHWHj
Y6tI7c4INZNRLhU0cIRJRpfa9XXTQkzGpvANpqkfrOXCUGBU3/po+7wWZD1iYpp5
p7y8xt7OYPsYbbltuxcDhB2obzixvXFntj+b8UDoRkNb8UAuoZF/VU0eV2K4t3nO
bXzKMR/QtD2YktP73Dw5EpTCuCIpyIFtI9gF7Q1W64i1bOB0YIT+lqLOzPlt6kM6
3gIFh9hbSYHcPFqa62kSlteCgfC1Rx9+V+1p3NF1rt1wTQCMjnXmLv7jPZR+tcjd
SO8Gp+NkB1HceoC6JuwfSUAmDahs9TzuZP7+kr7XNiqeEk6pAr7iio2HMm8lOGkr
uNaNRAn+8I3TBbxn9SJRRCYwCimQp58DQV5DZwEM85Ef4laZ2L0wlXGhfJ7G8FpT
7MFLvIlRu0yR4aI8B/eO6YH+vaS4FWjUXubs3mnSTxYTb+XTVw2MtBalZF4g9jiP
cWH4F8/YHi6RH7OCQRtcCXvPACFeuZfWiWyeC7zm4VfMrOnESCO41m+PWFyCLtHR
IJpTl7WhSa7lrIo8LwU+ZPN8GydzqJutVqTowZ3pfuNfQOCjFEa6/XhAXAqn9u3O
FwnvwXSeImMmGOQXZFyXBuS/iWawW0FSCnSSErEqLBwu4NmYk7q/cqDNdKLJ/LJ1
UD0gPNGOPGLg5IWWE2UaZ6BItwnDqWPhDwdZJGv6rTXjtXK4pWsbGRwP54VLwSSv
NpFN0OasyttATrTLNGtQFbibJmekVIKJpRAl5mEiTOXigAcKLVx10q0hNpJvDCLv
2NeO34N8QubR2/I0Az47T0xCDdtDYNrFYo+Erf5o28PEd9c/axD/DBJi2FXRz5cN
nTKigATTmHr0ZRZubkVWDR/z4vNmJfLmbetmX3/xLF+XBZibbcT4OYbyrNlPXHeQ
QKHk1jAahWYGmI1mqvRqT4b27AWyxz+pH6ez4rUExT9e3cZ5EHFUx/kuNe+05ymI
XJy+L1x2D+EzOLI4ob5hD73EycZLeIBkmpp5N9mXLXe3NJcWJauWWfl0P77ZOqBX
gZvvzdtyDwjNCWqdNF4Bq+2XIUDzJrt257tmBxhsetCWcooOK9ePZhIFoROiY95U
R/w/nt0TEh2WTKppRHLdSQDkGVhDVuVRNHgbQlox7c3awEThenvDPHIV7JE4HFAy
wArnONsMPtuhwP/B7kfBVoe0qX4FHl4OJJaitinn0SkMpwOvGTz0TCTzisGOVgkf
o1tTd5gkQYkW8Ub01wFXAvl2n3Kd60BVwcgvixlrRZEFDVbICE8FtHnrzFE0TDkP
AkFhww+1wqF5ixNKc6eneYsKnJ4UeOHjRsn6k8JcE0vZ0csTVtRTZVXpNVNEU0tp
cOuooVICutgmAB5NLerKpJtQ4FcnO2JkyBF7XdQYQonGygFCMj1aCLXCK4qCR+xa
j5B4tOvtxNuNStUaJP0xbByI43jBnxtIjTnP10OlcLKjXIEvJYt86S4C8fls9v7l
ibTtHA6vEJ0qOa4rBuNpi+CF/NL1WaNPh0oPlcESg0Or3Yd27zGCdNIRcxWAqYzq
BWgj4FD0k5T3XNKluyYMik0ny/TEARgz17qZtTOGqxv8uOrNC5i2S/VR3o3rJNMM
0b75wnsbRDFRUer+k6R5aLNd660WZCFsUUaO1hKhw7zHC8aEqiMOSKbKI2XJimti
I1NxvgZVaKelCUTjNo25tAElygurSlmiom82IPEgUkmD+SJS5Ae8NxTY0b4BlV0W
GSorzydsjZ1kn9UjpiMY5X3CY7cMDP4NCQrU22TG5f2yOr7rob851uqPPw/PG2AP
RL+zQsZdi61Jha4Qc12agicD5RSdM3sgcJ1gyGjU9Uotdf8BoTG75YdRoRBVauUk
xlBU5TI9VAuI4ZlrPdpLX9dUn9imjw/daa3pmAwQLSIOHKI+nJ89O6NTPX7dpjJI
7uGBhDoN7t+bN2SOXKBFqctsBiD5K04YuV/xv5gRMdYKRKweAKRaCQgmmAaJRgt4
nmYIvZPC3ljth0hbUfMjPCZxPbViy0S8xLNJXt5VvSemGRlw0mGm8RVSLy3bE8UT
lxoI/ETgQHNWEiPF74C9NkRYIyAq9xs245lpErZIsomZJ3OwHaUs14LaGkay2HSa
vZFIL8TAd4Anf9J3kFgRbE/stFE90ngvtMBD9XQcaH9fRIHKnBSicgLfdu6gG5+n
5DdLeR9t02sOZVThKtDcZCRLLwKnobBHISoovXS/4w7sUA4HmVu5FkUUWA70VXiu
6fOvv1oHFgwHNxG5Vnv5gWpKH8XjeneBVYe2c77c8AUBcUZBu4OE2wIhzBJysmyf
yOQMyd5elspCkSBeTf7jctk+k4PJBhpwUXyDEIxpEQlzqWZohrcxumtCDrKJypap
zTMosrVmc1VtjEfixnharvwqWsIexZN4kWTN2Pm0ZXKwbtofpdHz+ApKrp1JL5ed
oX0N6P8nm6QCrz0c3JNMgDy2gfCLTxHT4Wpbd0FboMpXvhJds4aNMqvP8QQOPgmL
5Jja4vD1Del5MiVGI3UmKrMJP3wciW4emXsyLF28n3xYaUZzbtYO0Ec05zbGxG5N
/iycsKSB8Z6MevjLGDA/wt5glWS99VsrBgUUBLKAUkrVb2IYKGaBwQnrhsG8/j4d
Zo36Zb6PHYJPQ5guL5Qtbkv6Kn7S1YHg76NEsMcpUDZMtBSugGiqfj2UEZiLB94h
KiG37di9dZFtp/6PiQ/FOat5FpQAQ0SVgFhUcsVIxWzh7W0MOvw/MKza/Cn9o4s4
7aCyyZlHutT685nvBbyeIa3td+9gBGxjYDTyRz17SiS7eaSvI75fcBIh4iXqLz/4
9jh812fk+10nT0wE4pCJdGhDkifhER1SZKTJrDTHD/+ggkIThR5RiipOsfz9fwuq
WLlnxgZfOud98RKlMsEglP8//ytwesBBgSTut9Mxhb56hWXR1CB6xpO1SKGFVlUf
8+xxPM8rou9GHtSyHyyPs4R/RqK4CAfvpa63wVvM6zNrQ11VaJ501Q2B25H/XjYT
cknEDGJpy2/YMGuDOu9lib74vohPCSumNjcR2jKNoCcp2Itrk8AeRBoSdwAvPsLn
OV8Bgm5ie70Ttq1L0UOm+vykDqTsYCSN6ErOvfyFugBKdMbZeFm3rwKmIwRwTLca
GMxefckt/erc6SziqRLsX5IfRJIl4nishzTAKGkSotcrqE1LjnOM8MC2unw9cvYk
Ylo0hAZ0ufIUWHKurjXHxt/AtZzukY0n7VfMxBQz7Bxk93izDzK468Bz015JW81g
u9q8HjM6OD1JyHDMsQFT5zM271s0Ydbo3L5CwDgUsBZbzgGPCkWoD5/rO/kJcJAz
DU3YdoMy+PFGi2x5bhi3u+75HZS0+7t1KHTsuZqtq+PPd86fpPKCmQT297VfGEb3
Oxs+JzmyQ6LenF3DhJOjKa9CjPEZ9UUebjMNLcfWyklsmm7Bm3n8iDj/thfuS66Z
onox5WmYCXAa1LJCuLHh/rEwdljV+KRbUBKxL6eJoJdMfytsXqiv85usFygijd4d
GaaZ+36RaZfCKcRfd4yabUtG/Wnzt4lWd9BVHq4nggcYkxCCgGzXEJEq05/Y/8yY
mFdAyWnma6v9JFjG5VZtynxwb1Ld+stEU15rzu+0mnSV8HeGyvGs4C+5duxgOWVA
sQe86EGroRQfyBOAjUGig04pN8ODA90dNsXercxevsLaQE3fcmnTGuy6aBADqj7x
KuBcPNGsJ543EmmAHrirJ2yNHYv4j/qcOJWKvxFbWujFhk+hWuWTGue6ERPloou5
ihuqdkn6WmLQMterpbhLxQG/06ix1ycYaN4jV/tKr0LyYoJlw9ZOyKJFWuHwF7o6
SjgVVC2/+Gi8HgtIxqYj8MS93bcYZU7tbpOdehEaGIXoVUtZQ5qFYCQowoabTE4L
HIBBSSVk/ka15lPhP3xutm1/PakQSgZh7FyH4LNmDZepHXDnyoOJYlElb2e32tKq
A189JQJ1BcwUSrEbZELSzz3kBAomP2VAXuhRBx+3I67Dt2Crfk9WByqgekHsIB4A
kDa87f/F/HP8RF6GmKrdt3ALOLsoRsp9b1Yy/5+RS0lfed3pMiIvlBw4Fc2Ynj9o
maTNchm0dOh1OZ79f4CkOKm/TJD5kytFLo0C1v7gsMDkNioBS7yXsVgv4r18jHB6
aaEk1fTsUa19pciUKvLUgNgnq710tu0QNRFcKYjqYxQeZ984omliEph3PkMxsGIv
LsJEuNUCoL0gEjTP0qoxd4n5bWVoFkMvpexlMzKYZP5RiSxsJQXI0BOm92XE0OL0
2+Hv+nF6p/InhxVG7sgVep9UHAD3RAV68GvqzUQ3z14v7vwYMhJRuJl+Rmi0axxL
rBHSpOKj+1NYcwuB+frpQif/pbvk5dcK4Ux6eP7p2vGiLGFjS3Z1TgAjNWPDFInj
Y0W4hteG+Mx8p431vF7rvnvf+HJDzyiFrmfwcpJkJ5lWtOBEdrpk5Pomqv4Jv0eV
WkUNZrXyfqpdrgyxyshjPc6ib5B4pEEijGVgQKhG5xaJYZ8hMUY+kE/zoDgZvKJh
eyMvejeV9ELwaJg5eclzGGOAMbo9fJV2lLlVGuOaEXR0A/BSNDODxWEmX1iKLRWf
ZNRDt03FuWEwIglTyuMlmF6qOZvczuZRgMSLjex0GLuLCMry3axEAGiPWIRFsAs2
YX/myVfUw9a6nVIBAcuD57Ds3Ywr+2l9FNLChaTBj951CH9d7x+CRK0B8tYuJPQR
RoJUGkx9fN5G1IfvZiZblNI4jmZKkkPOkzachq0zMFEZyZYFapK5RQ7dY0dODulu
H6dh61Gg4DIyGp6QEFZaWWlAFvRtkstfvHCWB6FaGATYDJv6RGG7zlLa8DSeds0L
EBNFpvfItn+WV6a4wvFdTHC1bEMDiUXpI8g2E30XOYcx0HAq2xSQo++V9h2Rr6U2
hY7lpHbMESDIQGtFAVe8ytjQH9Ez8+6j8+UQBaehNTeM5BMY/h5Bg3EfVwi0rHA1
bwASslO+6uPAYc6rb+lNjpjKhcTicu+01UDTise4gccc/0TBRjyYbrjMBTgd6FS0
USe9mPzp+4jp50V1EdO4uePIwHeqSUelSGbN2g2E/kgbHnGVIIWLYhP/ZG8Dig9h
jGsTPufpRFr0b9ekb6tE+bJclp6H+qMyE/qf/+5ddqRr7CWIoy779DCtPTL3DT9o
BwFawqn4m7yJzEjGytaYJ2wE/pGaDG/pq+JkvH+flVX02xMLUSqjP6l2iKE0EvHc
77EO28Nz/hnK+wdvnrSQkPNaNu95Lr+YlgRp7tUrrDcebvFfa0opt6WmNyxpJz4w
Tc9a7pfh9RQfy1GWb23CP8+9S/3yBDAkrCM+/391CfuHb9X+cxdrdEDHUx+p2UDM
E4V4Q8F4hyBgbF0PqESDVvySppfNXzOISbDYJPwQP/H+4nPuhXEtPRiYMBdiL4NP
VJNPdHdbVjhaAzBM/NfDa6z2iCskTBlsYGaXCUS3vugaFPCFkAALIgg875qk44kn
TuJ4r80Vmhgqlbez/7ZZS4ryRbwGacGHY8GkGZ1PAJyX68/ALPnHqLlk5TKMYOqy
wsGcIQjcx3MmDsJAB6VU3z0+m7obPOB/FAfAWeCyjtr+3LBSGlC5A4r0oIeLgejq
EaTwjn1s7cBB9jfzN+3ZokMEC2bgE6/4U20nCAElnuiGGrmw5iaNVPxLmARJGXjF
cR3RegG6nthXPRdCo5s/7iEs7jdleQXZFi+DqvDuiyn6dTUla+tkOv6qC/ZOu2Nr
aip6xWxbS/0GGH6bVDSCH0w60EB6+Ca8m3TU81bcHkvyaRCzWN7Pf86jjwf0XEWD
KsAUM0CN25xpQX345lWG72r2GeRuyIIUbj7Q9IpnRMot4Cq+20c85B4eNe8jl6nA
RIh5fasA2PDqCQUrPwDIP1ENdfJyWohfhxtISpfdLx7IPYAHbYm04YrX/1tMQWVg
8mv5dx7DyY0uFJ2kAZwtsAd4imyzHSb29HvL/2PWPElHnuBRgr9HQD5hRKrCGISk
vM+X/U7vo7tpZNFSLEPboOArZ5JOyYzRMVhKTSHYu/BTJiB14D0F2iKcMy6BD76D
mY+JbsO0Hq3tq5aBSTYugHWfwBRbFkD80B4Tib04Gnxif4ZkfDortQKzG3SyfG7B
qoU3Ig2HV7LBuy0HoEZU7GSMs7lMtSzKQcKGy000lmGGJYIoAWoaw4iRBxF1TOhC
ASOdqYNEG2o8niiiOJBoQ6g5UoJsimaLxUinG/0N6ZsTePpz5w47bWRYOogjIl8f
aamEAjFjgkFDke7ynAVXDnDfLRBFFsGAHxkCiBCsE/CSWJO9uiEXeiXS/WFWMxHR
ehzBteYSKFYyUT8aa55zlOrdUy1YG2w0DrbkGS4KI02/0KRZpb3TQiPPrSyPgqYD
YhOOC6Tdkn/tcOrvHjxLT5+3ayFnjqfYNOi6TpqnKebugcbpLxRAqcLLHFGcqC6r
itYw6bFs+goe3t7aCjXpuAULmzmmw6nZN8jxJhpiXBwg1WIKFPjLTjAWbl9Yy+aC
RY1LiT5107yu6ZFTauiUzqktxSK3M4IBdHMxvWp+9CmmGO5pRTdHUkIAfwjRNo3s
137Fd67fiOyFHqciV2gG9WDQVAwhcv65UDtF+9dO8dShcPbD6BXppiXWuQuusAOD
74PMGGhrfBRjtEKgErYJuaQci6flPO1lybXLrROyigpncK3tQ/h8ot4gjOF3WcGT
tW6b9igidptP9oZAjMg5CMXszfhAGVJntLBbxd10CM1v+FJHu5UT2wpzLjXl94ss
wee+F+jUd6/Uba94bgjRxtgHBjrZakNzAjBTik5K5WRmjH7/5qsDesNMqZZ2UsVV
Ys8txrECaX3LhE5FAGiV56KJQog4bzqTCrJv9Q/6ohLVFbQgVY9JRZHLHmtUKsLJ
w1meqsxATUCcCbnCYGpLdZH8fbGMNTr98KMh+VdAzVDho6oPjCNWmReXLsqRed/o
Yu71hZb7T2WtgCy97mWcpEV8Xkm9W6+7sZFgzmlL+CJEqD5BBzluUmSW5cbtAn8a
jIlc1QeGj2fmqrTWhpgjapeLylFmoUvffBEUqDIe1GArmJLVHZXJzAqpi70omGm/
U60iHkkfKlKNRss10Zd76e/C02EsbjCpLQnuoAkeqeRV1XRRSfAqnbq8ts7Vk0ai
A3zPciFjDeq8G+vFP48il3hnx6YwdyDqpmM4AjbNig3Esl8K0xlll/31qiGdV6LA
rThgC4dpQ2xXK7fmbuVmoklOK+ZMPjy3HGkYpGzNqGUHURXqnIMECLyQI/3B1F42
lmEfhRRya9dEJEeUiyDJ0nrla/2TnbnbqcxtEgf86ngxOSOT7nnUkDQzxb+N3LjQ
5Y+7kBgL4VvUycHxEY5J6YVu9Ell2HgNRY/6s4ki0dkXqMtRYDUyi6UlT2dnjJ7q
ztA2H85tjyWsOhuBstAg9RMYTPXo0aelTrHiSYbinpqWBEdSYAfBRBZATAQAhCS0
tQgmMtFJWBFut2OiowdBV/TuB4dyWOHeRbr5MIzho+bQ6qUradH7CiSyJOaxL9dy
odrOd1TRI74oMWcFxSd9Bx7L+5MV9tkqB2V7exlxcQbpEb1M++z6XGw0vp2FXrIi
hVLg20AOwn6S486WZBcVio1VWBfq8ciyzAj0XnkA10B4Coobq3I3JYuQlQP62X9b
k5iot2yJPDDPUW8A76h6uBQLbo5QuVE60XQ60kPYL0/WD25K3ruUf2XgHF1kw8o3
Ieko21YVkIGGNZpMjnDhJmN7CgOKDg3Amot2ys91Sw1WOrGe2mxddHEaLaU5QFc7
pnHox0ypRnDEwXwwKJ6oPT9P6XSeE+WZsDr6adf20HDBpC4x+I8TpazXCZLebkR6
gWoRgXrHQ+QAP3cR/MiQSRaE3PjwWKrfGAoEC/T91EI9khlHY9OZH99osDyefgos
hTQocUDh8elrw9w+N9VgOwhTDuOAOd07v1GPDkctVZpdO7GaMxGej3Jw1yoxBYp8
tbHxSwkOVHdp8h4K3V5yfzyYCn0knqfb05GpHJ82wZv6BuqhBm9YsoE2AhBo90nk
mz0Ti3bP/ipD9VCrEwro4KrMdn5xfneI9ZclN7I2dxRieLB7kBezSLwtlpN6lgvq
HZpJ3Phcu0BoOFkehjd1zzCgtw1TCC4R6rDS3W9EeJQscfT4D4XFN6gm9v8fxrOv
W4D6PwyOwXxqiZ2we7Dqx/3xUL7JxtWqDslUbDwil6S9iFiJci31ygCMp82WpaJ8
N4LTONayzkl381/sHPTxM9hYNGWh7CXYx9MPJzt3eEHK7XG3S4hHkzp0BAdkU34J
yZNkd9SeEd87I7kDGPNLA7y9A76cJ3EygttgALVAFusU9AZI1/vk4BeOkuARfyLO
IokRtf00jy00xeKey3mjFs8hchVtnTx5kYrIKzQ91yZtJaiSHlM76pIK99Gu11sz
70fYsHzn/YUQAPJi4pMU1cLlngR9bjQssRMZhFS9oEypLkzqbF3vGvmExLACxXCM
P04JmfclnE06GD0OE27aDm+X2/aeEXnuj8hwe3XyW+LZdo9acBC8uis0gaFar9cT
X9T5GMGwowqIV3KtztMescYY4YFeg8rAlSKomuO4TurJn1A2DYPHD9c+8fqQTIZc
hdtCjuKirHiqukgY0dlUWj1YOL4McAjb+aLIE842Q1cA//xR8GYXCL7A0VuojctR
6/SAJ6UHP60MAPGcF67AwoQEwF7QeX6074Yn5Jc91fCYw5ofrOo++gVIutif0OY0
GE8xXNe9dMPt21awKqkPWkiJop8L2Rn9A9jugdYPCFb+eX+v1QO7NoiC7v+5q8ik
aLGyPRGA/x9uIWkisz5bYiL0w5fn16SQDHLbCOisF5qcEtmfCBn56WqmMY2up9OE
zG3QD2xl/mclqmL2nu9dINh7NY7eafPHHNkPnD1+16hBwd79/GoOe7vbGjoWYWV5
4rlvgxrwmLNI1yvrDAbstVimulpJUDDWIT5jXYO6ygHJnjnlQUKdzS5DROLw8uFp
B8fP+MENNbwbTKS571Np1huDvijMs96gaaalntMNq5/vyBlu2gYdZ3EPhG7h5B2S
Zfou4fWT03+ZuFCChVkgkKU/kNTvPjjciIOzJel4F5754DqReSOhy/NSDfiUNFK1
7vQ0LyVa1fuonmSAY7wypn67EtZLOs9dmT2QzHIKTFfljKjuEZbB7UM8Hi3MXw9F
b7EIit3/1KH7bhGdguulHNFanvRhH6DHjk1p+Hrk6GP1LXGWDkBXwnBxkigxsaUz
4YzKk1rMTnLwu3YIj6jBXAChTpLbYq8VT7GqqjVnOfgS5VZ6DmWhhng+x6ryjlB8
LrRihQKtTOBQYDuxFsBTumhYbETQSNWD3PJcU8nLFYlXX3XTqUbY1zaiIfujw8tB
QmheWDTbgyIywFCXQDJRFOPvwuNMMHklZr6+BMlxjX/+/srrIYh0t/2CCvHqcwEY
Nizv/pBHqKIAGudZd1iX6qb12+rIAIK673HuHF+4+9ccNG1d5CRBvCwIaNoREes2
Pls8O7o8Ypr7Akb//U7+uOR+pwYTPteitLOq83gtcZWSO6MmitKWz3V9uqpn6QYV
FQwV1ljiX2SZdGIItPXVdiACB05UlRY7DaGlwXtWDCiNu7DV65efZiLFe72GT9ak
vDjRrXhz+j0AG6IMwVnVWuKLO9pbnxOas8ChElJIdtYDYZSUyqnM9rx9+Es5YSUy
JQ9koiHTX3YnKXLopF2QS/hER1RZpNDzw070I5J5KPzBqH5ttTba3gfsruo2imG1
MESFZRYGKZ33hFAzvMu7WHLlwiKwJiSXE6jgb8RECzKuM7kzD3IExXqOdNVCyaZ1
xaGDT2sWtmVjpR0kkTfaRxAfXRUzCC7vfQXtJOGp+53ZB1o2qeCuppfw441k/Ka+
xhbFLvTpxiqeMu2sA5wvgr1+JnZwMpcG2fUyFqAnxxQWn+y4k/NccVoZRAGyomk0
NX1pMUEibfdZCw7MlARZ/OV0dLlju/q5oCN41GupaAz4AtCjsiHiK+uhivn0nGKP
2ODTbB34jwEAGjnq4OjvS15VAekC4hHyTVSE8DQs2EoE+Ye2sRNFa3hjZpIU2G7l
fd/AjXoQNOzSmuxgA9t+r88uJjGtURNtNvr8iiKdW5G9xJO32kJqxtdfDZCgdmRy
M+ZIub7Tt++9JBXvW751fXNG0Wi6daepVeGWtA8KZrxVWjex+JgLbEaM5v8Wgw+0
6SECp6ZsJnxtgu+PNJrrsSEcsIo0ZoEI6AWk87JNiOlgk3L0lgcBJONkTpuQxcTD
axLvBDOpr4+FzHMI5+Y8hlBHyE9acP+RSFxSSe8uXP/jytlb1xKbjsLlJWDDPJ8H
WpFxHJa2/t7pTJ7KXInRev71VLxnrG25AHZFq6KMQTu+jD7iKA/X592tJOtjd/DX
onIV8Cfv5Ob/hcDNd3FdxvVfFABn16VC5jqPOCaWDtKrLfUoij9VuX63JRYD9Do+
27bwn4n/CTdqep5t7QW8ikmmd0zoxLa1MTYWPuMrQPGME0RyipeQ6bkkfZV01IE/
hzoghHOtFUSk4+YLJnMvKi3x/WHn2rTtYjBA98U3X3HH+R13EhjCY1F/OE6kfmg9
pepmyjVtjACtWu04KVtP8RXrHt97iMmG4blQQEIje8RI1aFutsFwDqhnQAZNtRvj
6l6/VIj0m26aoIUrbVnas//2zlR6sqGcf9tItoccA6YxzSQM29VJrVvdjfeQHPbD
j+G/oVXWO4sdSFK2fLHK+och8p6jN4aDOPBrI0IDD1PZjLcOvtjBW16frHHIdmXU
km3i/1uVcyWRdUpOlsC82bnAF12R9ydPyB5dZOjI2ByoEsPf2kJMIth8YpF4tVJN
UriXnEhS6P4b90MlK0MA7DbfDUHwYrjm/owhyDAfFvOPTIJ8czyHj6xUVa45mE3R
lw2M4teH0akttul3pFqQ6tFKSNk0M5dIjzWZsppyOhBZ9RcQTZV6nkyY8JOLZk4Z
BQXKb9cDGij5hIaMwxR5Q2Nw/4ZRkbtfMm03KIhERhjduQerVVyW6zk9dpiuvnxD
rNXIiPg7PN38m71ObybyEKyJFaswiUWQ/+usHCI9xNIxHJegVvCxcopjaAvFiYkw
8xswzko6eG1MFfUo/Jr38/WkcAQjrspose0YmwtEBnQEPZ+UgMi4GUKcYPWPBvYm
KtETJhIsyPm98iOBlwC9eM8Ps6ILiFz2GK+nrQniNzlB87OGOgXumqk7hicriJGr
CYl4cQ9hVUnAQ/TGwecQnjgIcIsnNGd3AB5Gn/RNv0J2Y32HYbsLY/EkmAm2J/kF
h0TcXScTECMSSmC/7ucn+5BQzxEuoNDU51o+jzwStHZqoHxm0F+JDfRspk96WJQ2
NsFiwvWWq7ZPvlkysS+7veSsec/CTtww+lLAjmqgV/sXhcJnPhgBKi2OsYs1dOfo
dGTAt3zLc+Twv11/54tCpUcigpFxlg7HWjLgBNZ8wxEvptx/IdLz7XdBlngVdUJy
4AZ9m4s1z3pJ+gt4beKZkF0Kk1hnlLS0Pspx+VUGwDo1ThoYDQigV1dt/XrZRczf
dD4UQ3k7NjtipOVXMmJvjplZmiNy7R8BzCC3wLJsPLue0AAqsXqgWcM5ymZZhiaI
6lF3oaXUkcJFhDcBxMt4iVJIZ8MHLDLim76DZjUU/1MS1lh7bCraV0eG7Ws4Qe3w
LJoiaMkSQLyKtHILzM79xSPohCX0fele2O4teOctjKcKMc/mKKcg3PFJpH4hVx+V
UT3cHLt9oZVXXtFWzUdAjDDFi2xgnD94k93hcibSe61211TxYHN/vrXNsXuIVWAE
jo8gVBqPSnoXq0GCO61Fqv9OGLiWar8flkYFBh/tTvLYACjMkU4A89pMvoJoeRny
k8LEsKc25h+ciZ3XzaM1zaEi+USB5Kcmjy1Fhvfy2DcinTdSzZ5EC2/FHA0m0d3s
UOL6lmaAHXpXBShxN2hGW1Lqmq0QGIEJTw6GvEDfuOVw0wIRFKLGKWeGxbLxj93F
uUm/iHjzYaxsjL+ALuAzcJQJqhuCrAEDH33OoWz6Ey50pgkm37WPJlhmqV5JURtT
gvxH90KzZmkUL0J7iVYanz+SEiGrjDuOw3gKWofIjE9xDzD84GRN+6uFVaUTvd+N
T+AJDyqgG2Fbg+CSbVibR6e4I4W/c8LNBZlVbz9f7il7DfWeDtnCJBKOEqaEzvmz
HzXCFuYIdOVq/Yh5pMdE9j8w80yL7aLR+aPRE9A8z89jG2dGq5gMmZ95hTdcg2lW
n67EP0+54UW4D2dN+WJ8d9PCszOwhcX+X96CzJwFya+ol296vKEGHHUP4qANbaxS
KL54v74qYg8IxI6Ck3uNaeqU+h17oByrp+zaTDVXRLM1VmubYvRgv4SfgP1DqZ5z
3mEteS9wVC9i8j1MDnibYkIHeJhBoo4n1Gi+PqyX4EX6b7VK7nqArnnwsfFdX9Ug
kiyipRBbEoew7yzyn3e9zEY/2Wlo4VcZyuF/kMCCEg2miG7BhQKUVcqwrdbYctNN
+LDB+gDOhL3qvjJ0GzruLBmAvy8uqdMhtVnFuQhKJoW08XvnKKqn7OX0/wP8TuHW
NRzYbaw0hIBe7b8z7t+t8hrzh5zkAKkbnsSb77AHGZU6TZ0gQ9Z3W5ZHXaW5xRre
p7TMJK5FesBDwZZzWDGf7qQhYyFv6Tx6xDrnUQH6oSyTCjD5+OUfR7+qHV6xeXb3
H+FSgaf0Z4KcoWSIwW4p1jNNbUOA1jTigApVuxYGd1Y6ul1lEYVe0HP0cYVMhTCe
B4H4xonoqQ+qconnxoBTLgKlqJkPGFrUj79gKtOzHvyyYbtsNkGSIE3o0esa2WNU
KWc/l7aS5EYkxT+W0zAENBakATZeDW2yh0SKPKDq8F8avOtfvK1it5muLA+McI45
I3lxUhiiPm/kvP8KwrftTuNLOYuT3RGXn/RVkzvV/BjF5fOsNzxtn91tFR+1MeDz
sVO/oY53PTXW+zlZ1nFLSiBnV2pOWIa6FRF0kSOSq7+foUOxDOOXOQbqHd6x/bnf
vWhR9bapZ1jiSfiWKBmWtXc08ZaavpgRuLyvWxW3lE3yG87be2SxF9V8ch68e3BI
TTBZZglZbJXH42GvsXIURNxSVfANjRVARuBeXaweyxg8FILSpnh7OP+Y4cEu7YVf
wrQyz6wBjCZdYKeCTBb8Vwsft5bGGdQkAXSPrfmIxzvwCB0bNciK9Vjf3AV1mDTD
1Kv2YHf3c7IM4bOuUPAQWuW8KQyJYyOlgexQspLJdBnJZewLX9LNxf0WJvcPyDJY
OPwIC3GtbD9tCOFDW9H36MTg9v4WHoajtVgDwk2OYTXBFrk2W2J2Ty9P+g11InOn
woi5PiMWxs1z+A0gPHMqbMEWwjtSzimSIPmcKCJvzusRSS491jInYYkZ+OWpUwjT
dycSyKgRWayuWBlhsljHy8IA76S0Ki4cAOOJUntXW2Bzj8TQLo+LFDnBhkI8/iwK
Y5P1wCImBSaWtZA2zK97742NovCimxcZL8BNSa8RRi3eXb64SrUFc7kPLSEfWePO
S7Ydsp9iC1xhYhlcXK+B69qYgbfUTX/ps9VErjeytEC0TyYlLQzwRAv8/+l3EntY
k0hdLNEYmD+IM4Xx16gbKFI+mpJwUG2FgYVxjHk4MXJ5iUyoJuKMWsnkUDbWGYpN
LAcePgfnAwlsJCrBG9SVVGQA8PiuDO+dEDY2iXbYob+Ks6wD6u/JL6FJePv4LFbr
aKjvFCgsmjOl9/s8J3PHAv+Q63AUVGULmN8KX/sQbU2Ca0xhP9PFhhpHWNVnE6rB
u8CMqjPe6G4NDao8gjZUN/7zGl1VsAd1p2wiuQJeJ39vRjI+wyCzB99BmfPDzK0k
x7J2cA1SPYJfHkvp8M4X6/8BpNGgiMIYmkjgeyYHClkiPNpBYq+Ytxz/sN4Q9pur
DZxK3KA/rFhmqQcFc4hvu64AzqsbOGKCreOuUKQq/lRdr55t05IM3OsImtbmhyMY
QrP62SU9atEiqBbx1uj+ltzPtBBXsg7543ywImUTmhUclFv9L9Qv4+8zAdraP5gV
dEKWUZ0WoVOG4af0kpmGwgeM8bzcU81tf9LWyz17kk3pmqxgBu3R3HPnVHZ4QteQ
rgenXHjTep1QUBr5GvoKHR8/7zbN6slFY6EzpImtAtT6gxwNPBlxM9OfpZraLxoS
xatQ2AUS5l5UFZF9yK+zGMkoRaNQMUNgtqjrUhZKh5hqeBGOqszLxDjwR4pSQDSm
Sngrhaek2rqI7iu0xKxX7N3o73dCSkNYxK4XJPKBzPevCDrsTjofiQ74fcLwPdQF
59RojNgqW68Fn8EcHOcjaO2F3NGggbIaxdbbuuHcpvA2rOiVV09DOO0cO0y1JQ0o
vMllMdb0CeXi75ARhV7Y0Zj8YYztIGR6D3Cf2alYnfKPl4uW1ZMq83BCRNrjxAnV
AxS6JWDU6CAPRZqt736SkACV7Lu5jNAajrHYrS0wUnptPK56gIUEe/x4IrOzscqs
6e/TUBX6tpiBX9X0GwJWOPePZ6ATR+IRg4cLaHvUax3JJA3AduwwlYaQTN+ApJMN
wkx5WDdGh1WfXDfgk7ki/JG7BjZMGI09c3wts5Nb1y1bcAJ2IiP0kvEB1AzkYzRK
m+LRXXtRxjAa4hkB8/7pZOwf7SkSTlQmXweprwQClTMwI+nOuoG1KStc6Js7YCpb
uPBbC7egsnRlpjF6qEiqfjb2XyEXxnuuq6iXcq1+f6b8UPAyTiD2ZGmVfxF3O0Sp
1lGdaMvuuODXU8NyNNO/zA/I1AIo05tJ6WPsgSrc/Yu3U9C55iNXzQ4l9W0C6UjW
Gr2y21CFKPgax7AWRdrwXRaozNaG3J8Rx2Y4+Mf9j3ix2DnTeM8a8ejTtiK68aVY
s0nzJzNeKfMp0FZEl2GmTMb65299vwjxtDUNsvITS22epgHafJEQQlJBbaBSOnyF
a22xjLDDyN8nnK3sG8se/TB0ssrvkoZaFikPf+f1oOn+BsVFDhAJLgCm3LM1CCUt
b4Zg5D8QZwhiBGQuGF/FO3NJ1Q83FmQetmGUzPjjezZQc+yaKD0je1WL966SHhFp
hVXRlgKFKej+qnMDcp/vCDWpoOopsqmD90/0bM15zgvZTI3W7jHa7Yx6yRDLi0yo
L7CTKewFZNIzXrlvn9ATiioDkxYwdbf7cemBS76y/5y5ML+J5rNls/5IoMhr2ms5
Coamk7Rtss0Ja8Zf69ilqgdu41xj2IxqA8S29fyyiJgzJLOwQLETAYkY0ikc5FYI
ImGnHMwLbyVvBxNfDbXpI9tmbmRo88mmHI+AQSiBa9+ya1uYfs8G/Aq4P6oR8eba
6J9QY1y/Ytfar3m+2FZCIQJ9Y32txxJi5aayx3sdW4VscAcicmxxd2baL4/P+KKo
c98Co1sHcM4dzaCDsJxuqzGhsrUqp7Wnm/4FRNBxGFXhzjtBnakq5Zjrz/cwlhKc
dE/CqHQG25E7fuBMDdlTEzVcNesKmVoS6SonWPJkAHHplTGKB0BOQSMm/mxMKiWN
tMHC1mdkvMz55EgTYf2OSufy+B9Qq1KZ16a1cPHsVaTY+zI7Cbo3N9aAXNDJl8ly
JnXLAviSA4n+V17JWWJVo9DPMu1EDOyLNWo90uFPDO1ecdAgNf7ytl0Fxtyj9mxH
PAnOFrUxkGydRUlt+JxMYu93qlvcRSwTrxFPcewPKP/UCKXlmYIKcACQw97TNjaD
PO3PnV4le67KrBo1rb5CGPSFTDfX/beCskRGvSn1bUVk+nrsJC9NYGFWw385joKA
94OoKLzSJIF/xbNaXxny0Br6l3Pyx+urVo3NTBOT8APvCssfdcpvFKOjcH9L/zAX
aDjkfxuzOURtfBYhPwLmtbMoCeSfMZpzPGYHLeD3O7XYKiuBrYHwMRVhG6h8s6Hr
I3Yv2IEpnGNS2U5UMMRvdqrtp5AatCpQldqzHJwd4Ylm7itVE2a8Pt5GFganxjgc
WLrz9A7NU5cKa4Jg+JGG7QAhJbum3qmlsI0DqDcc7hWSqWDij1Y2YDRC1lw/BzQl
1kN6ENe/+vk5GMT+Zk7o/HWCGSObEc1FNgSyxmNY2Q+jyCj+rcOwZD/7YhJPyT0w
9/n/TSRNtoK44rQ8wgBrUHdzpEl0heFmYlIbEYlZqaA5CLksAlQTBS0S5+DtAJeC
PF6RkhgK+xkKNyWRiVqL2s0O/A8tHxtBGYaoUGoMwgwC1qYXRshpZREIarPe5kve
X2fsKga7Mzvh1onEPn6qw7+dQOUh+CiPZjaU/Biv8PdPfzGm26Ne56u7vThE2vBe
Yekrr1wqkOWjBq9Q0JtXyCr7z/zTrenHp61t0sObNgNdEz+U7bsh6G5UHDrAvW14
at3gqFNjV112Wyr9tIV3FEjYdy4r94tkike5xKTYqUmishhsHTVHBZryhlzQmfLr
F+EjOIqRjrZG94O1hAqWu3RTQd/oPlVgNmvvjlgCSsD9Avb/10ti1Ha8pzEfZVpu
E57C9SCt4K8QJjgaHLiV7NMBO/KBVjBDKPhwKVLpLocA1ZsmHLOCHzfA0CyXdtQe
1Czoe+BQE0PE4mtwYOsOP29xDYfRDhKP5+8oK9geRLAJ0mqz3swNM8uVgvqFauNq
qN8A2MfC96BV1XX8whvEF4MdbZK8W7q7oXnjekSSweiotp+8e+OdMGUOrETSPs2m
o9iEsgiqnCXDIkq5XESO2FtsBzt6B7koaII7sfzTBdm/vQYasssPPjOh1pQlJluj
vMfbydI35OV8dNC3AmVylDQnc0OK4ztAV+mOL2sPxr64ewxcci1bCZMB+0EjBEQy
mxDEjavfG7XrH5mqXC9zO4kH3x3+kzGzaGFOo7A/QzKffS4IFsOePkywFaxzbqND
6bklcaYL5i4ApexbPDw+oJL1MFkH+Z9It/VBaFAMSYxgGGExLXCYpNPqtypSsjf7
CU22alM9clPs4simhy0r44QfSEZSpIIaNCiU6RErmKzFJXZ7Yt6cALxqKvLTS32N
0cULroy/sJv0ZDZPGZboFc7QnjQJfH75HIYA7wriNP7mrMj22rnvrGxKNyzk9laS
mvzxJupNEzm5/pIMzHvdT7Ey7axK9dq2pHpobw45Y3a9yDn6nIQu/N8i09Fq3UHh
ZZs7IGVBWXOHY0uoNqLi03k7YflFcFJJZibJdnTnPfvzWvDTa0A70LSWcyv+ZUTT
UnJzx8WHFpuIlRaOSeatABgDfYW/OlnhcZZueqQpUKIki8vnel2IZ3eXb1EEtUgA
1rZZYamBfwpaJfAvhb6mOSqIB9J+NBqL+7LHUfbSJzlzKtpz+sSTaDovZcFFdZnX
lNVWEuqIOTi15G3Q7a/CESbiBZfxtFrTghf/zJkkYMdXvpmOazKgUJX5iv9vC2dr
FUvbgDsiTG+JhoFiYUyw4j7ZL59nGS0GgaTtDLPZ8Zwxw1Rk6o4l2HgF60JGOywW
PRVeRYGhczz53iJp5TqdX9sRhz1ClDzwACVr8/CYuBEyayEgRY2RgAxqG6qbb24B
iitUP9aHb50zQoUd8mcMbAj/ULtyxEtjp6VpiNffTr2v6CvE8LQlXcvvR2EKFLrf
9VyPBGPUpJbPzCu43xvIjbRUF2KlNcKZqw523BK7Uiszix1cVqCX+8mGwWoVaCpL
Fwi4FZthToYPnynlg3HtxsB2xOMv/1Hpr93PWnG9ybxbrDvpB3eDOxgTEvz9a2RW
SBM7sADfsA68zGOKKpPK+QzMyFew3n02NcUtLJB7CMKLFV5D1WMSxLQWWcYK0QMA
FkFN1xNu2FmTGy4RXYPU+ZZi11wwqFYUJCvEKUjoXCwYkAlD0wCXeqssbsar1UjZ
9B0WMjOCRdAQ/Ee6AhLvCr4OPXi/MhrBuuNMeHGNpZrtm8TYfgi0E1ETKC3vn03N
iq4p87naG+TOdeAb4saLtxxKF0+UPe/TRPxKVLG3kcX+xfOwd2S48jCQBHCsTW3/
YZgkmF7NWEZwoAzxrcl5ZolS7FQ26T/b9bTidgDSC0Kuwfcni+mMu384pLmJ1iBT
6ElU7DNv2fQQMHye90pwuwrMlLsWtdV57zo6avJlRMSTPgx0GC8lHsgpbSst0PeT
3M+yQ41vRBO6WCEveSz8Z8KVc825k65VfKmL5roDhjUAzUUGydU2dq0UxDEVo/Dk
i4JHvZ/FyJZPGG4VxhvBkscNt4zEdaup8lXDgmQbK5i6um4+TqHazG/GyJ7gh4zO
SzdZnqAc87Zw5GyjwbTGvXWo99qvmbrQENQQlfW3+U6Vx6hyrAvpXwEkXKu3GDzJ
Z8hlOvpx49fgm6EmfG/HIWX0M4rS+HACvpiWUJn+N4+4K8kmn6h8qMbVZd9pXkPm
/q9bkf91CDBaIVxYFiljk5AY4z7yUmWPdqEV3icH9SoW2zW6Yf7RG4AN3ebvEM4r
gsJCpoHbOlMlERvnznkbINAmDyi5TSBx8IYa2LczI5wMY5STZ8cGgsct2W61lEOd
XeDLMBcaMsnA6soSwNq83LrrH0Z5PmOgsCDAcqJgYJqnf5bm0bX8uoXnTsXqr5Au
UFfshL0uN+QT5uy9sV6rs7P7KWESxqpgb60P/v0Tncci89DI/44BJRWMFlnYMhFd
NnsA/tIoWfFeV6zt7fN3epO5CshFUuOny0lj4k0MQzepLPyJWclG5I8j2VOP+bJT
MOT8sNf9kaRGJ+EKZ6dRkccddpHcToVH06eY26khXS6Xw7163SWHaD8b18VBLEOI
jxyICB11gH3ZPXUDb9jlqOYpQewJkFRi+TVKfEl9DPYSiK7wrk5CqnCG9WBca1nv
32128jzACY2saD6054+DdN5fvofIjNkvti1pJQv7Cen5Pl8U7KULJ3zXMS6ery+W
txkm9L8wf8h9ZE1KiRad15dJQqmOaF+KSFB/P9asaRS0YKWKr//Z8wmSmifeDo80
2mcpejMjzyEXCgDDh/KgXiyMcPew5InAccnVOr/VqAWEZiwowfJFK58L7iahlBl2
iMKoqrbEOutHkAObv1/u9d8Tk/OAGL6unG6j03fvzJrJYfA62gRSkZ+t9UKwAa+K
XzwluHYP277O2zVlzbU6H2LJEMYioH7zUIzj3t1QaE2gBCD9iB4q8M9v7KB8h3CE
/zKiYxIMhipSdEd3kpV0AZWa2peqh3syulOdg/Dgtjsglxfm0zuYOyE5n6ywNtlW
e9rwrGGryNu6h5qUDBFyOw41u1nGEErVoBrncdvLag+DjZ8bth1pYqAw3i3Aky8Q
cohjhGcIVYptiuOl4IW9A2ksRovdVP9SxjYEkYqEUC/7LUXbjIswIb02SszG6H7F
ULferNR7BKgJGoX5rkNTbpT5I5w6htU79zML5U4QTcCvHs0h2QCKdMqEJu/LaBNJ
z55nH+C2maeaVGJxMc7QmXPyt9F8ljfwl5FD9fHZyailTJ8eLEmekZ4lgFOy78fL
xiTWld//5YpA5gfQvh+6zeYoK1wSxJg92zWUHtSvKAo4kxLdYpXM+O5B5oJQdVzc
0CwR5gQ4UkK3riN2Fmoj2aa4r0JSHMwlVvLZjDVqK2/7qVan7K9yfdzQeTNS5N/r
2OYqodUIpSDmJl/txejT+c1unKZIwzltvpvRYtZjJqzeu1dLQBEucLwOjQMBK2ZL
Yubg3ZdR304cIXwSGumSGEX3++eN5y6HVir3+uwdqJdLHjgq4sSjtwzIs6QBB2vK
SWe7R2Knf9GHQ27zwQf+a3qsw9eNt7R5UPq7iL16Q5Ibyh/Au+I5FaabPKrloqFx
DT1IVoYPTGmkWBpWEoyqCWjKTDvvBo2JvvDl80S6SPOHjmTuVJ4l9PHCN3SpWYoS
4sYQkmJKlwDwC2jllYRDtOSCeUYDMi471jNztpVkxH8Cb2awjfklrZk/B8GjGP6p
TzZOw3FOd6E4Xkls1cdNARmHO+OOj7pvw9bcZMYzRupK6WOgo6Qf4XYd95TOmRwX
S1jCavdKUHLH0V06z7kQ+BQYfcBnB6qpr8Idv/kVCFR20fXkTjn+wMyP3T3qQqNj
USbI5aPwanXRsCf7njADTyqI4zqFXtMOsH/RSQSwOW3/0a7hhsCInip3GPWpzdlw
TIIs+GDTqKW8Bw9pmrKmZcRkAzt+5zgvYEhMy/n/E9qo1KuUu98dSsnjNz7j8RNA
4FDFPm2iJYrFNYtATf50p/LzQcQAodbNGC/6y3Y5yw3KuJM8xxvWXYaHb5tQ10wU
fp1chq6rhVofdEPQKgmYlT1pSt74q3UWORQJZ0SAaD9B3Zt7KRCD6gJ8wicPRhRH
5V0IrS3EusVZg2iGhdQwFO1+0lHGFOoQleBDaK33MOwT/kxjv3OuAbxB6F9XuYHX
XOYILCMJa7SuqkcVbqDe/2DBq5Eqdb/jyKc5Lyoew/WE17pabsceukl/51sk8D+p
AfsGpdynlNMy0kiBqdpgvu7ZnDijMajPt9a/TYZ2a1Ew56l3Gpyb1xZ5iQ8pLvlN
K07FjkAcO3ZT3uz5sGHp8g9ZcYF9+qveW3Vw1GX8cw9lA91kZ5FTVc8e4uYSBzT+
2pwPm1aZKhngHAlDxTAbHBBbak9ywli9t0HOSVxTWyDcE0ELfPXmsGUr5AMzXq5f
+NMVSJFIPaIivKL6ShmGG3gHw/MoKKcNqokLVjcq9jx9PUTg1TgzcLP/tH4ufJdt
93NH2BxM7OoZKCEDUSYeJ6Gquw1J5jqv/6yRynZ0IYckKA+v5gktoK88P9a5Cf1V
wPZpmQq2SMUP1IMkruiXp1DBisqaEg9qcFKtJOhqGkE5MZKVuRWXLfKIRhUzl6Yt
UVg9S0IQr1bUjpASE5AMLGMIv1OwNIoWQf2vhJDDbOwLi5iNJvc0LVdVZkgCGQP4
pLo6TTIUQAKzobCUrNUVB5M3y+gOYWTrUPnaFKsBoDwm4LFR5FmCzYHvsHRvbNZq
T0bq7n9IdrP/h/nBnczgsNlQmfawqCk0DMviZ0RshwnLixVwJOyPpvQSw77S8wBi
jtOGmJZfiyQsUKfhZd5EHlTYG1KzQu9xgFxV5GDHvywAEzIKIyuhYhxNvQLRZFbF
AFToaaBCi4cuiE4JWGP7m4aVD26QuFgEPErIiDc2QJgUcT9UzrAzBjZhmDAI7oN3
bhmX+Bbpwx9KZBb9afagrBkVVPz0Oc9hLjhua7eq2x+Bc3HzwYx/T6YZyBMgW6W9
tSTIBsAtnLTwGqqf/ef8QVsLMlAQld4rFkHi0hblxAppC2GeE8kfN+agxmA78nzw
uKGYOnf6xXpJu/zV+buKBTJpaP6STGYixD2Ky2NFGYSv1v2wuwKyNCznJq7l77ex
bVvBi8bJT8Ss0ef40tw7l7BWtpuiNNavwAPqRKnuw1EincY4PP0gScFVq1IBvPWy
k2WkPYxR/Yehemd91IdWid5GX8Ont149RQqE5nw4rPyPxjzP+ANagmQrZfS3QAi0
uMGAO53Ch9yQhe2OExbXTr71Oi9LlWz6Q9BExRgc1TdCHmAOObHJqEPEVk5WW+G3
CulYDDeVYjFNT8/WE/snAg4HT9gE++iSVDsgxp44s5/dATVXReyPwPirrlJon7Cn
QJiarFIm7w1Rxq5414V6fvQ/ssO5dX7s4wESnX4jG/XuA1PyPBt6G0n9lrZh37NU
PFBZlHxGqTbrn/7nV6Cn4duxZKUvyYgqPyrRp80TLrKJgFkbX6S+uifhijSCEKGV
pSWmOnGr3cTv/8Yb+80HV8BB1qVbd8bUy0QgLaPyPzjdXqlzyN0Cdq3LHSYqY+/I
5IqgCvA72f6g2glvSc6WMWQ328qrRQR76Ce9IUDghQzoqEbWCswekg7vKB4lrrSW
XEOp3+clR8w2lLV+fQBIT8ged/o8+S+GHUv8Znm8tuiEfhWbcErUV9rDAbgL94NH
3XA4f4em8xcwGzbqZ2lHbbCfkdWENo9x6ogCQedDblQIlyrX5fYMSkTyQYODrE/4
hKjnzj+Xs3IxKdUaUvgZcPPoZ4bXcQUKextLNEaF8OBlT5ghJI7n6aRJr0Maj5ks
t1MSDwuggkbPcI2zF1b/wiSVbvRy1xMlPFIngaqQ3h9TgDQMKRHrVkJ57zBJIE8y
N2CbgrK8wcfskZGsNrAumC1rev8sYauDEb2aT1frJEJz2Jfw399jL8o0ODR48a4l
vG+ELEmOD8OHmAH6eYcuAnY+FB54hh/5oM4AO+uWAXFKd7vZqvoIG3YLh4Aq+dAn
p1IMkSh0wkYBmg/8omR8hht1cS7NrDvG5AlE4gr4vCn0k9Frj1R+0hopSsbSW6hS
dEgi6owb8mMqMBN2Gl2R/4YZY+JYh7XLLzK72nod7FMl2AIMulBVuBvr0RCiqm8E
UvF9YftwsXnf7a7UYuAJGDciZjvReDfNiF5u3HuI84eGIjA0iNWmPft64A9e7+3Q
t+7YOFdqk5BPbOpil1y9bfMM510qtWKtzq3FtpPAJP0GE4P3WhV0d//aoIKjrzVh
NUNjWJyY05QZwyA+mWq8z5AUEo7CumHnfgZvjCu7BUYxN0g7JTqqgh8ahy60+yex
QN4eWXjEH0GCH7YD9wcJ3hZlV6Rt7Uf0cMxUw9POdmWKV9DNstHc0r3Pu3uctLjR
/yRBeKZI7sZznsOeJMOZow1+rhF6zcvj3gc2iMHBUvBhzhGAiAQcAN46FFH5Uguq
BRRUtxt8+fRH3619PqU6X0AlShJ3al8eg01e+Qhl6hOn1ao0dCKes5nZ4zFpZlOi
mpQO+mX7FRQX81K2UpBBwGjwxljoPD4dX1iwp8g4EQFkkDRG57wDF/9xpLwVaNSg
aDyWpS+wCTaC4MkcfYQFznUvG3k9X5Iz9d+l6mVw7CiLbE8S2PrmNgiosuf9Ck2+
cXS7C7FkqTlXOy/Ans4bFnFMBdh69uZ0jHrXOj7+uNHp+BAzFuOGBxyLWcS7Unyh
NK0rLZ8pYSc+FKghqFPp2c4hM0FEBggVq+2ZwCDzltQxLzVRgQ2Wi2nIIUoekqv/
3KQVWnrLOHHe+tBFxgAs/sVnm+oxYvv3TSkfDdDK/MABjlTIBgcODnNtdhR1LH5o
lTivhd1WjlzUgFv/G8eH7A8QVSdBy+TOf+k2fLOw6ly0ZO+VxFzjLjQbrNv/4bsv
YeVvu2BrTe//Re/THHh0ze3edlQwEKZVNQVqsFwCubQJihF9p0xfVuapUVUOWi01
lVes+GFuFf76aqY1zbXI2AW3UCWeh1nhj3RWjLD9o78hEZh+wfcB+htWgrcAx/Fk
ktGZ+R/ipUfVfqwaWLAczVGi5fhsNUEsJ4VZnUmw5mvZETxvK+yvfCP1CqV+1IGN
xROzPtBVFLGi7Y98rPRH6VRzfqqer5jLNBOScluRLBFmLBhBmh7DzUg0j6ljh5Na
9uZMlhjSCf0oDWr36oo2+MBKnOQ85BbkcH+bIcAzX4u+zHmFJQKaX1sPaJfRzvpQ
34ywWjuqXpRKkopopz/1BYUDxTTCkzPvbsNWsTWxS1uALGeJ43MhrJVQAsUMjS3o
jD5i2M1Bc8X95oSMMjeJsyjm7JK8X86OOFtUzX8wP3O93mglFM5Kqm8nv1kti2IU
v2p+iH3U0t27d85yYmCDi2xWG3DS1JclklLCMjFZK7WkAikHOXxdLtVV4kD5OP6R
KxaFRn2ZKk5rJyEyxHDe+0v7eDe5DannyPJJ1nfHKAQgFsWzZ3S/mAbt7lyVwK9u
CtTWfzNqT/YwlujJM7msiwKgKl02Fx3TLFTdWpM1AEI6kIAnEDHyJ5x46d9C3np2
WRWFX6phvriL6WWt1zBxz7BYJMxLhTquWSauVfPgk5NZB894i8IBPtVPgGrNPHnv
TddmFC9FJNbgDlKlM1wh5or3wgERaAq030F4Li3jWOnWLsXB+UkVqOGYlWFkNo0C
iRLDTKWqrqRlvPAr1eh93MZVcxt0MkAl7UzGRJGde0ji5ikAo8ZQr2q975ssynXU
r7L3pySkdBXyp4jXNcF/ji6Gx3NT5mS3GvSivMeLTIzBC8QcKkMYUyXJlwwIgp+Y
CLIRv/+1KIptVK7ZfMpwA/mu3v2GcmhYDly2j5LdQ8XL+GtIgo0cCDAFyFLISV5O
Ud1/cmmlKFF60dNOakJIFaTw5eub8iKkUE9j08exLMcvHnntenlHNu1CONAccMaJ
sFuv7FnCB7S879R1HZK0BuhWfQhA3JvevZHkUcpGjddjTTBF3VKoI+XsHnRWhFVS
GpwCzH2uMLqyP8GIbOxTAqmwDkZtYkwDLOYqAHxYZTFNqvdG8CQWthKFjbZlVXUF
05TUuMAErq/+jU24WGb3Jn1P/CqieuEmYi3gINxCxsNdU0OTpPY85OpYn04q3xKG
oGIih9E3GR4b5jwZvFYLAhF9ypHm+UfcS5SbxO6J7iswPBUk5F0bsVdQjVXBimdm
cgFUBUhb7Bm+FWC6kvyE5ClQOeSs5n3Nh0uQaMuc3WXCghBSbtt//Cythxg4EBN1
ysxFVuLqxYiJK9+zdlZUFiM2F2FzXUoDbrL4aOKfslIVqQGjSnrSlKh+xrFqyI19
M12Nd1fEbHIOrhHWEdXCKbrhvci1ud9fQdGOYW0zrNWNc3rvkncRmjHx54ZGKbUp
/0rLh4gXhBSMdeq4T9Y6h8sRCtCxgxlFl3CBPrZuMHGgdFs5C9KR4b9P5/yeMn1e
eAKmdthdKTJ3hfElvoG4EKm/9HSvtTSw7EignQVNM79bzdpBtWqj+U4Zj8AcreOt
nUTFWXUY/Xrt34x/GRNfGrYBDU2vxOXbMdcM8ZzxOjMlOUv+2Yyott9GV0mNlNL1
O8GphcE3l6JrCiU9o7l/NCK4VEa9VA90Zquli5i0UFyojyiza/EBDulpNPO7ZHEY
qBkpja2O+5VaNeIJkwHp/PJFrRX2cBepGyx4JUmuS5waGRJ4m4awQjZcBL323Ifm
+kmP7X/z+VYSKvHaMvkyrbYdM7K6jWi/7AS6YMiS2anapZAgFyeV3gP0Rj1gsOJq
isCC4PsmVJ3wV+4PiWkvdOH9Wyjcoc+Jaz4dQtU8AGJBk6Sexug7Glq6Ug4VUcck
2mvvZiw7qBqbAOS1Gy63nv9IsZMsCnR3FYecjlAjHs7Dw0cwEdkP11uoUb7I8Eja
WjFRyBJ0bNrADXn7UYwzXDCIW/+ZC7JSaVo1gwVmkAPLBwbZrvFIGy/zGstobS9u
G5hnDQp0hkSdMePqcqn8yocaqp2aRbK+lVfviGbwmhTtkbV5Ta+kYLkhfKufgV4U
iZ6dSV74nJLc0Dv1PdmLBWo4+jUf75IlQ9G9vMtWJU0cI6h1LOCEpdr3cTl27OZR
LImvcoByNBXA1yf6Q4n8XSKiqdVF1N8TwSZWvggmhE2J7zobSlsbTZ7/ODfA1+dR
90kCkJsLasZdyxWAHKAej6YgK5aHdVqQRbyWqLOXxUfqxF5BGzzu4sft6Bl/JX56
3kcoAIF6CuZ05NPLVDeGuztUYtUV6kcNEpo0T90WFKwR9XEJAse0sk7QVKAVkayX
E9T4RURYwaYC28ZveiTnoBo/mAFSYZ37Yyvohd9rECYvqYNG4BysMNie1IoB3APT
YfKsfoP24tW0Z3WN4Hj4j8VFMYiADWN6SQ9pazgY8gaFMTVfeI/myK3EFrMGE8EE
zaHuhZ8m5IpmfIlGNk41cGRbmErig1gTRcS4aBJTQ+yCB8dCnI/B3CnwKTVgwhPc
+KDlWW1N1IUWBQrb3UaORy2Q7GXktXVdV7CZr7RkYkpGeH+d2QgZW3xMhtTsZbs3
vI5vslzbrzTGLE3V5llIgsXUeMtNLQrTsZ9gvK/q5O+UMirxwjh/iUJiKCYFVpo6
N320j8cY9Et24OmXKBgYa7RMIkjrgVrqI4kduLwPbQIs9EpAvAxitjOH5AgRdX3v
gOpev8i7SYaykMGEbNx2IVMDJj4jJ7p3oRxiCyqMX3+hzzXp8aWMepTkvvNlii9N
5RYWQev81dEXVOnmgeo6SnwC3CCySZb9qHia2ZcwKLBCFP9jPKVaGUtvUMFWXE2y
7JLVEdPSwux67Ajh26HlxX2qgnAHJu3FaM3v2cjHPghyC85QFFOuhyejdoIY8WHt
YgDJNg4Lhi4F0wU20nLA5mjKM935c/BMLwFnhWgpB18zMDBkjMC1eiLQC9nc8vR2
l0wiGa7KKw/dKMHwAf6mCsDMsPfYcxhK3JCZIS4akaB7tzO3XzkAuZPDhowrn4Kg
Co6PD3YRw6uOq9ASvbwgiOssT2uAIrkmFE5BeXOWhkAmA7gdXVhbmv1pOvxUk0Jx
k2PpnipBU8H22JFmrLaLevbDTcAoILquA3P8Jar0HXb5+vmMXhgt64rVTKcqFNsV
0C6ta/rZ5iYHCYz8CLKWGrDNvNF0o4KlLv35/ppLyt7c8CzxWhstEOcmaysBYzoR
+4qGZftONAhTJqQBLmb8D4tU0KE6ulKG8bwFT7Xs2RsZkSbP5DZKAfy2rCAM2/Kf
yWkGzi8qHGSzY6TA0gNy1C2iDrh4efXTnFSY4I8Vw8sg9zp7GodSWnO7bkPt4y3P
t/BU7Rxavr3xR8/55ih6OovLStbym80Ie5Fuvw0YcbFdsOrLE57aWwSYx3lxbdj7
Qs9EUYuiBVxSzbeXnICRqFLpTgzMDtc9HHkh1J5kIRNleA6oUGbovMxqnKB6QoGW
ONVf9I5Eq7cjNWyTq+KTVHX0LDuB2+cdTjjGSm9qCWxOciO+BYp8CH2efJVnOZCy
UpjkUWR+8lB1PFSjxoyGNCtg7LqHRdW6WWRzXp009VoKr0TlQ8v/VUbRDE8XHQOY
NEMGMUvD9zKQR0qAJCT7YG4YlSN/Aw15POCBmdcWcKGET5FOIDKamuokOYz8mEdH
doOeqaYpJO4Q94NeiyOG6CTVCT/ZfLmdnYIU5kO6GYTna4Rz37K/B7kd7GYqhefF
6peshdN8UBr8Y+MnmAF3Q74kdzQn4hp1qRFeBcE0IAVWmiR/CoOLVNHICA3RqPS1
XF6cUzMrfwNn9e9nCkiorol1DarIW9cqr16Y5yKEGJt7VKaX5IhVL4SHmz4MToGl
cainsozcGBazLACpw4WXmFGGyDEk8s1QzGjZodE4w+Ml0XowZ6EfhlTRwNRKsELM
ZqzgJ2xk6nhxMxaYVKQP/u9cRMuT8gDf6KtCNBF9YvqrG6qnUUatCXQ/pb85WOzr
hx04VvGhEqfWsBIAAWVWQaxT661kXhXix666Jao7fgchNfdz2YyKgRDKuK2kbiYN
DhBLSd2F6IwC/qvsjvwLaHcoTnsyXcoxWDJeC0eOScZta43fa4f0KMFoM6WOYNjN
0ib+Tsvhaf4/5qS41+cNNjIKqI47/bhSqMe876rukqLdGEEpP7OO712ik7UK3qvT
uzxS7QauKd/5WJWklJSqPimZ0AWn7NIKsCEUUwzsIOOA22EKveOHFtRfR/sJjqZM
A5O6ShpuatdIYC9l+k8PHcFBBa8RE4IY1lXfZ69xMoAI31oZYpzb2XMYwob51ul5
nK6wZwohDLOborhjuZpFt+wMWwezOAYQFBS8/SzK6/RFIBFr2TJM4For8YEVEPBK
ODw7jxUVigKJPJufqvo5X54xTBQjb5UhzmMpXDKA1Z/H6RaV4BPGODdX+mzsIUgE
MBQ+Acli6Ti7YdpSfxhUoPihBOoaJBJWMREafBz/YBWIqavsp5jt0Mz4ci85OQFF
mM2WizuQJ/46mtaKp/64p9dB3DbErNbX3ADaBz6flbu++W/TWxI8ThtRNCCNE3XD
CUGcUG1RfPEQThT28j25nPbhHdltzuzWQZe6y+LuNfoMSmQ3x34rlpvQ+0UYl3yh
9KvvG/GLGjso/EiYTwrRAQTYzUh5lpcP5S7dNqYg1s/cvlnCEJTrs6ts0V9znETG
L+ngm8lAoY3i5yC/73DwV52wDlwHfvMSdraE5TnzRWmkaRrAutcIRzDzYPOREzVG
ZNfkOBsB9LKZ7aJ2UkIbYjpkO9XboHv3i0bvPEM04/XYcpgUQq3xNGztqpOscCTU
J1VDMX9u0wf67m4BkCJMP3aF9rs2j26av3FJz7ZqzreQ9+Q00kZ42DI4Reqx1sri
a45leXHHucGQ2GB6y07m+f8SzOwN5JEJ5ui4rPu/cRyVDrvAOJ/Qnk47wfHC4eUv
VIyqZaxzLETmrDilv8ENFZ9VeRaruRb85WYnVqaR8+WY8u4gOzeINI5VvMntdh33
EwfapyQnjm1c9c4HqCa5giMdusc4kRtgsxF268AK6lpqo+YCvoAzwxsMMC0sQxcX
rCjzJL8Ls0Rg7JHKcAK2fxLeqKuEnJe1HAOau0ZvUhRW1f9raXrVbRgc7wav4PY7
8PTzWqdrFob21kHzLvZsL64wPiDQD7gaCifehsgZ5q71pfPb/1Sh63skar+7Nc1o
rXRwRa8sTsnThiZnW1uB+U+NLSn2n14/+lwyLtN1W8J0yRnaUV29bpqiIpVaYm3h
AEL22EdNBqbLbWCsKE0+GEX1QjdIWD8vBtuX99mP9oeOlJxOHhtRaW/HVfBVbH/+
TIPTfHE+hVfdZboFLXUjPVA22B9k/2yF+nraSEwZIvXkOYwllliAG5AFYuL8DYcY
bsUyFziqmad31VZbK4SnINeefCc+1NkMpJ54ejfOLQZMvU2gsQMYubOUQGU6eKgo
sxmaXRIee0tnFvutjRLAjKPYUTu6S8ouE2MRzFRR0o8oAspnBpCvR/4izlfX2GUG
OhkoKeNjzFBFV6VP7FmFGXvVY/qPWshniD10bgqQ2Bwgd3vTr85VH7iBxmB1TJeT
/GqiCsGctS6mSw7zpeI7TeaMfPMSuRu3CRf4BYN83PAP4uWl7UDyBkDXLTWIIvaE
Q9xw24LvpYS3Sl+ER9D5HpJCgwVFevzqHAs5Z/O9X9dFYTx1uNnntYNuxxmJvB52
yx5gnDcejylw+aA+b77GTd2djdvKlFHaepK1Jt1q1sgpzD5vEk8DynaXs1U8Lg/k
YXro7VlodFKTig+//Hy6tsOH7gDCp22rPORyeh0hPZRGzskX4lMOJf9oBi2LoHD6
/aA4iZuh+mij/GpNn0gasOtq4RnAVNoQygenD2QHRGv5K4Y3Dgi1WVIeS9OQ5zMt
1rYUThEc5U8UzSqKPBHT5jqCeHdCmiOlqomjx1mkWL5GqiwBF+/TWsA10ocP+/Qv
KYEoJvNBx3544PZNkF87NZXpI5M+tuelSP9SqHsawL3nABdHkApKhqOXYUXQgKaa
Zhuc8t3NdUTACwt9EccXHHaOHhcxu0c0kL+Rf99RSobmmWcBzg10KhNOkYMqdSSX
Qcu4BoS6og9vHSgL0rVV4u/U1/XEWWe+9lGp99t2jyHawB8q1NyOugK1Mj9GQXOd
p4IxIxQAI+d7/vUb0RzNZm56KzjRLXhEDbAAieESbQb2HXMfI0DgdmOnH2uUEHLK
x+Lpi/Ca1Zh73iSFcBTfgAxLKCdOc0nX6aYgSRiIxWY8W/d6L/tcqlRv8cjjmh3q
dc1hl4/ey4Kzl/nHX7sSwCT+2RIXfHXHX5+t72h+QFvLlX69fDjayyFU7oG98Y1H
gWOp5B+qY2tO/y94vQbEAi6i31eRBotOVRcp+/T+b9xr8Uj6wsm3czNAzPMfy+e8
GlNqVxcr0CQ8zRsC013FPUDgN5g7vUKCg1arKGrXFL4tZVPQCh+TO/a8akCeAy+P
mDIr3mWAUGeiqe5PfA9V06/bpbjnx1wboxOTzOFRYxk1uemVrqBZuG67aBIhP/9c
QMCtV96Zj9zh9pIqyLfJW0TO6fjfOpuAVupTbBAN5kxcPteP3tpS1o5tPLjRs1a7
7K7ApxHY37iJ8VLyZS9Q/X6F3EtslNDyYbMhh/0I/h2aFh7mHlIBMNcjEFwUO3LL
l0GASRu2MjahxHQvSADnW/IMkZwwkW24vT222Mxmic7uMHFi9SQGSNDi48aWKeEe
P6QO/8JOrixbUve/rvFvOiu4aGCDJaIsbDplbZ3t8HTFWuRqh4PzsIfpGNo2fMNn
V3TByY7PjtqpuQAOMkmplzUesP9sEdLx++yM2RydtZcTTD8B+wdTgwWxPI43hvIp
+42FyB1nVPT0TmGfiql1HdWCfDSzW80ECx/KpitjX5eTva90b2wtK82GHbysqLY+
kQ9fb+AmgpbIq6OMI+QnBadi2mKQzzRkHGylljn7co9wNHTr7h9/lpGQkAElMkFz
yfB4W8G+Z48sc44wx3DAI4hpgcKBBW52y6M7RCk5LSk+jThCHL3lU3ej6mbNfWhr
M5jcx5a147qIa3Va7sSPJViLjSCeTadwEfJ7F4BiV8HIze9a5SRFI0iKW8Xpb7zd
v5Yqs9Vfu4957Mgk8p9VuSEucbeBjKQDMMeKQYOvcTJ292xd7qafg5rnS5zBmFrG
Kv6CmhyvKp75rgWOy6JbojXDhWszJTL9UFvt/VyQgj0mDJLEc04B8FYIGWQ6aEQh
HbncgCeRrHWKgjMmfhod21pLSnDnn0wV1ePt3H/t7Frf3+u/cabo20sp1/oNy08m
rQ6V3dMN1Vl8z3bazTdasuFcOYpcXCKPBU1hlT0zLWPj+Ya/XB+MjdyaN3fw4G9r
KI1q0/yNeLeC8H9ceO8Rnk81sT0TiFscjyZ2BsioooctMDQtZUY+EA/QEdDDIJs9
+zu08cMh0HZyRh0ctEnvgpZ1LOTEJUAhU5aDnAhe/TL4hU/5DEk00i8EtmoyVB0I
8qdh0NaViFmgmrlgOlfxdxjN9VDfAjirVicJxYJTzkxqCqRBT66HIVTfjgZvlUcP
FZ1/arLd2DJg8kE4OkWsBq+nGGeJFPhXSUWBTSZd4lSBZbXTXBeFClzcTOwCqRly
zDgMGj71FwG34wfMdIPMs44f+UDS4Ozw6MdJnCkwQQETEZY+tGnLWChSovphK3OW
FJ7izsbCrdxyH2JoJa6LK3QcbsxIefHaABZHJ/kGXG7wN8r+kLQtXEa4lx5Zu19v
/yAE6cT4Wy4BuRsHYQkM1TCcYtR5PQc04c533g8nz1e9lz4S224H5S0+rVD146Zu
IacqGDHwePLmAacSZlpTfuKTPzhWf6CySxVNGlEIU0391sM0KojDGRyCyWP0A57q
0rPsdAnv09gXuksYzI2xIAdm/b5HWcYU4EdPyrQx9hDpkV63Zl1VO0I4uPpTCYTJ
w3RusmrDvBUASExQzjlwTiJWrUDxM26LOz2TJza+pU1Nwi+VvM7XLR9L9kBO38O8
8E6xS82BeY2ZYzxWhCCC7ZyGgwO8sxxHNMZhWMu77I8ILpoy2zQURTbD9IlMxT8i
NN0DNEJi650q6t/OHAzSwM8ln4zSUxpw3lllz6f+kglDSGObONP81thrft5gArSL
xus5h/LRAmahTNDHEhv4dGXrIvtpvODRtUcNCkS7ZQa2RmFMszau3Drm8H0Y7qYi
VvHPYAJ7YPRvSgS9yjA+HBCY7URwkVaC3/6L583CHH8eDjLQO+NOp8fx42rCrUV9
Lyo0buHYHi9zksmWnmt2irnrGG4RLpHVK3spnnjKHzUb/N7C7usY9vlotdOrKYta
xJ9fas2FFJBU6bNU6TDOYHTXtyt9Wt9ANAr/LyorT9GOAfYU+dR6098gX0LRJohr
7kgS8iuGBZ//uJ8gkhhLWru0XsOzBtisctrChmeLBs2LnGoq7rWQe83rYvh2W9mo
Oo33GorO9/evpXROCorL9af0WgZsHOTHuXbM4HmonAi+fdZOU45y11QXUUQ6LD9N
pngulEM3AqliVrmon/LL4Hpk8tBq3RzRS0fJPGaHX9D5MDi3G69bg4TFAFmisEXF
ofNzh5Ki1rmOX3sK1gBBKYrVZW4seqV9rhTmvoBUSZqFsFVz+MwftRQ8novkOnTX
e4CGDwY3aOprmQD25DqrZurlWW0IQVTf56uM3MHR3F+A//ASJg5AgbMbUACH3Dn5
ZhZAPVouMjkRRxBLxoMZ4kjWEeIKtYjzuvyN2i9UjDgonO2S6vgc/ezCLKoMwag/
NCOSf88yT8lojq8bxYCDCpkcxeiQ1N2vPLk2V5JOwnHjTSZJ1m8KpUZNXsN3MIys
Yroy5rohOzRBlSQ862QEJM2Gu06/DGi0dRGNXb/KC3aiamtet+BIOJINrRDXCilr
nZlzk8Iv3XjpUAtuq6dsV8ql+7GRHRoArBv37reFr7rXBZ0IxlgYhn0vFqLUILBA
hfFXkLkXcZM4H0lY29P/acEbTik0yctzLmx64vlzw1cMGTlDfQA0cVfo7z3y649G
+JVrLA0BmzooDccXpSJhTq7MgiKCJ3NSpGE8QuEUUjE/DXtoXdk4BoERZRt+Wkmf
QktujU+mwo0QrQIxErPENdpidoddoiycdmk1VM76Te3ABLcB2TQO2LRp9glTOzkl
X78+V0+aMrtKOaRG2vrZDekaT2W+WsMAKwZocYbusGyDc9inpK11h6ui4VRO1Srt
KT9bzmc4L9djYSjYqYDt0iLc6B7zYUn9jjbxAQ8O3rMlM1ABgGVmVLYYjzECNy6l
0wlTbsXl60QhJBJfukXj8q1YMaFRGV3/PK6sCbB7GzOhTNmshRKfNIboXbCy1yQS
i0eQ+FOAYTP1jg6TotWr6KJuYzwZyFF2t+P1SuWCuhOIE/fXH+WUZBlKot53zzIL
87tunvWB3oHu7VrAqJIslWSrCczt3trTme19crsZGdjt3X/8gysATHEIJS4zwowY
5+Vjch/NProEBs4PV/C6VHeVkec3Ni46gtbOM1V3vnCSH5qJseh/mde0BtiSKWR+
Dtfav0XrymgFppNHwDr0RMeSN/OBONHHXXLIAULLud03LwlcT246Yon6zBw7MUZ4
XrzC3RzDzbYuHX2b8+tIGZp4eWWEkT3z7wxYTcp1YE9pQOFPLYbyHb2rgvSmDvtO
/SVkVFUOP7mDpwlEY3U5SpHvrLbx8L+mfWFgcr4nCL58drdgeGX44o7JrgXmrFUA
IkW3B1ISnZROKkNR1zLrR1vY0M4p2AK9UM6lJP8z4Y0NBKCmmomP4++W9K9zweER
gsAX06YuEgBnFtclnP7m8SshwojDlHC6/NXO2jRKoZRGlNjZg9ZK9gS1AHnZM64/
HrUiGqVSUkYqdiFg7PRZOpIOPHifqUY8p+xO0VCRG3WQJOEcYLN/FqII2eCybH/T
ReoJdhDqKmxzHROZ3B7CiLud4BWsZ7yeD59tT0hnG+hcKkkeKCIzNsxrFKBxktl4
jgC/m0bCin5SWzlFuEDACKOzG2xK0YX+fWPC/hWZlOeGjmqglyeCM1I9oeM/wtt6
dwJ5u4WNytx7Hv8yBLx2qXONLIrNiWya7Frge6OwFO7atJ3Mzv4lWSfFY+NFnqOO
vikv1GbLBwkvttRkqkpI2BvR014t5PDQsSffrCs7dZgWM1wvQLtH9QBABaTM9wLs
ibxwGxnK8h3Z3Tcm8kmpAoF1x7ww7vst3BWq98d2IG2huw4/W+Pl6OH8Hajr0E2Y
sp+ewJb30+GcDWSO6dvFwrGLwGvyg2yHINobXs9ZQXLEXPHcdN/OqsccG6M3tmQv
13God3Sqcs/QCwyir+nYzfSSIAe/QYhoQPGKMZK0GEppa442+v8qwq/Tj6fXbpr2
V6XktwhtWe3v+y0WsyHVjrnv8LStisQA1/HGuNkQp9wwTgmnFyCTiL9AlCQT0no+
EM8x7MexRH+svxVh89ecOTnCZycXJS09oU7I+VqxjJaI6V33erph0FomixVxhWqq
dKfO3UBMXYIXTBcZ3/YbKDqHzFZqofLPqOtAcoEhUR1Yk297nze/QNUaQpk9diYW
43fEtmIJenjI5zvKW3wzlfTPEi34vRxNmwPJIDhIE/PWsY4HrPhUwG4Rb58HbnYJ
sa/7BOxTTAQlVv2CK1pwbzpUXx4my63jiGro88oCjthf68fI1WiPcBV46BZibNFJ
A2VimYqbzGIJbKnfI5Itb4wsJjCtevb5Q8OAcX3k+6PZzXNqryL9tcItgM09CMSC
rYBzSSp0AHraPNak41nwqdjomrP+X2Xm+Aipld4snmm2Le9DvLlfvLSTpkHrCVVY
fPVPlCV450uUHrzsDQ/R6HSyeLjsZyCwegc5+tggMQCyKL+VQg9iRPH9J6ObyOF2
VXn0Zlitjjb+RjhFcWThU3f6uNz7+rHRwzx4+x/1mHO1wgLYYT2lhUjmc9FTMvSU
DyFgmQAgXmiLwo+5LJZd6N9nkZm4Nwx2sui0o3Hyakto2yyAj0PlIVs+ZP4EE/fa
v+0raIjrz0UJiC5N78S4N4hGCTJXq7VN2Y09inw/MfAdap3FXGqtDYcwDTGjwcAq
6ZvPeiPD3mR6WhhrP+oy5DpIHU8Kq0gDJFbOEFkRGJ/U8CFte44+ciXbqGs+1a3P
ojjjououRIIBgUGpolT4toqwUtfjn//k9o1PPDApOcE+1wArsJIRutdh2UDq/zbl
cTxfSZnuzJISIS4N8pktnLtGFwzlpHou7BrKDk7wEanD9ZHMtPh/C28cXrCz4jCa
6YAxlV4U4s4laWX1vEqrXATqu+bzFDvjwqiVKc7BvNwIJbWfiB3DLT6arFLYN6PS
Pg3KrrxdjyA2Nez7+gcetIlbBPZFjOCcwu3VScJcAHdvTT2dHbmxgewQTR0DiNlZ
2XUgAbPop2EzTW5AowznpoP1ZHzfdUtoSFUMAqhSDNlYahpOtDpxqyxTL2si5t9x
lioykOl0GRduY9Gkk6ujjKnYs7aVjLdiwLsX9OxBt2x00239BpxNJdzl1A2Cyp7S
j++qdy82bAAlREIHyvx0+HC2rEilt4BjwF46tDXU7rKDiU2HAI671s7uZ44pyTZk
vreuopT/jjww6Ubr58nFEdvteH3SMjkzvLRfQMdDdsz/AfI7UpZq6rI3Zf4WFQ6f
+us9kufFRzNyS+EZVmulUKpboMXbbQhtd+BacDr1OWdHXr36r6qAj6TY6CBU0SZo
d/IxLPqGGq/e5EJI6GGBYzlh2oa/MAuIZ3EYEsG4T6HMRQnwGgkk82VxixcVy1za
4EWXbP4C5Hlv+lSzlnKHiXveGzHkoMZgvUzTdt6eUHGxXJu4adV55Sf3Ps09s7jo
3JFjB0SFFsDeFtycRIYJXi9OlxBEo6823MTlBdnxHmTskw47MkyL1WcIaVAgg6j2
mBauAODFJOfpkVR64Xuw5ju9CtZqNVryNOBPsdDBRnBQkK9jTbA4wFzR+oSg1top
Y+2oMTfPV/OaGzVRn0je/Oz7dMdacKW+K9wDuo4Qc8bZ419lSbDPxasL1n9d1rtV
GfuyzzwmmZ9vXotGRQY6yM8XHRRwDoJULADZLRfeYn5E7rLJYNO10JsMhfi+xjX6
Fo2tkfG8302sYTQrZv7aj/bHfYGHAe4F1GC+vDL+NNN0qhA/JzXo9G6c7kRaghIE
cqOERd/+ntrmApBc/Vxe+3ZbIGXsmpw6hC7Eepjo2uXWMeQ64hFWqftz4Q8HDxIP
eDDpiGTbiU2dz4l5EQJAGHzDCCnOy05Udj9S27/lZV/cFcH1vbZl/0iDipZinVSB
o+rMFjb03+d+9cCqR5Qh5ZQJlpQLA/qR/4sKi9mI7RND8cQtVcUAMvmHQljBICIV
GXeYjcaDzMundV5NvvjAZRCmOl/S5JPw7MnSLEwur2051Dfdp47/y2HOIWxbcEmm
gysLhtKXW6X6o2fB/Pl0wKUxil28ZHBt5NLGIw6yGAjZrQDDm6eyQElvdzODhyBD
rEOlwjYcs/bt+ZBVGJHO7eyj4xYHA1QABhZ9pNM84a/bjkrLAy0uWG7EWglUJNd7
r4CRNpFydkR2cig7s+YDiuJfY00efFyVytGqNSvi6Xadeq620lq/7rB1Meh5q3TD
n7GvBgc322ITaMnDtUszekLcWZtyuX7bLPiZByIkluteOdIJio5Oq54SYa0C862m
zPcsvYomhKvVh90vYFrIiXyAkLkgVYWcNKD0nISeFOkhakYoIag1LqwmDN2KhIv0
t8ulTpOuzu+aIHrs8AQHdOnUXVJvKHBgFbG0tYMfJp5K70p92VYEe4vhPQ5W1c1v
btL6tq7rc8zZXQpUVsmvGWd6B1kGFwV37HPu7zhKGDXH6cFrakVTuGo3v+WRqmDE
d65yiYCSVVoALibQ37XNySY6ayW5ufilVMDCaUXdpxoe0uSXQQ0GU9zSR2k6Tg5Z
Fuc5M98aW8SmQztmV7WY6Ha1aV4Z6W7sKGqQqHIbB6RjRqOs+FJDccEpyncgi+bH
ViZtLW1OEadW9iYmbx6EGl8NMYN+Vc9iNcWYU/A8biP7KoWkLpTPd+3dHJ4zv87v
as5aeMpJbDfRszKUMtaIWIN2ZQY6KR23w2bGq/6lErg3JlNM3pnqq2pXpDT352ZU
KYA7YH8+fwXvPy5YMOvk9S2pleuDOfvFXnZcTQFpMyZIDjNVotrwdAFyivGVGcTm
ugFBWwCDY1ytyAhnJ1oZbtlp09qoQG2uQjS49ijMIUH4fIwfftki7A33M8bKbxLz
LDiYw6vvJePOE/8cDVMdeduWjvw0iXauba3IJk7wDx+oKV7qW0THwrORaC7TV9W+
+npRv/dMrbFP7Z4sHjKGIYeqRPy4GLysM37UFQAirP5k/0ipm49MfsV5AY7ehZ+z
r5NWdKdQnSnC3TfxhLs4KEp8wdzqDjgjEz1FWPId60vpMJjcI9k08Oh22l0IGSPD
Dg8UD4/JR9p9cOUba/wdbE/B6kjkbbgEsXibT7+YnpME8UtAOGr/JLdD2XynMvcG
VTEDC2R3oKOwvS+JTbabMU+fXdmWT7nl81zyMxll4m4kaWQfAE6i2Ait1Ggt7QnM
9WNlzJk3S+qyIaeYt5dCCfReXCwOA6N1ojG0qoMrI0j3oVkvK7VqYubbU9LnAN08
1b28ujqr9yc4kXeTD95bp8RrwOsHB2tPjO3/+kRmSe1UV0xOVyiIRok5KtFNbV4s
n8F+Vi5annhefxulXQN2fSlJSkOlqnhds/W3pmiASToZxBkT0jePKOODEslVld+u
IDMyut/VjjFRB6pp9f86+ZFkdpbsSAAEUZD7KRFgzgFVt+SBGDDpN9bMA80ilYJ6
c437URotUFlbmYBrQbxabnR+FoXUoYJJLxetv73XwmT/A0FhbWU6joOLbESqlBZ6
LcfNiDX1LQwV+JweZqLrXBdCHPuigabVFIupVoPBYJO3GW4jdhBhY/rKKAkS+vdF
SaIZ2ZDe2LL8KJe8m3/VHfCBK1EsM9y4QfF2wmwvUjDN/LpNCrJnvt97STllCOpp
TfyH2ZVqKi58cTdt9E+oudDOOCsQilzXdyqqztkYL+ovledC42VyT+RzNv8eCV/N
v23ItAQYeB7DesZKVLXknhxgckcFf4X/Y7doX7boNxyGsbSMWWZGAcEmjQpCcon3
sy421cgwOy8tj8nyNnKidFSVe02WdeD/aMCqEARbv6mvQXhi0D0G4Vn2pvu0+06w
xvhzCdAFFZHOngXH2+pTEvoTT3rv422v1dV+n95xvpwk+d/1dwVeGrdllt+t03g6
5Bkp2DZdn2PZ1UdGCiXPGk0k3V1a3rtfxWBzLQ3GZ7p4gFTCrG4de14yJVk29Efd
NuWEMT54a71vISbOC7XJeQ4kn/90pAEbwbACrzb4mVmAsWJui2jaCzHJYw3Opspz
9ZRC8PuP/gOmo0ZF93ckjZ58Z4w6STxdlQz7qFiks2zW8lqf6t7xN625qsg1SR7X
iSxu+XLVs++wZIAqp+fDA4HLrQtP9VCDO4jB9hYwVpxE5YqYxTloD8qUtojvuxQ5
SgjYt+dFECxtOf2r0ZHnsMxv6O/q5mgivgAvyT3npG/OGlCD7I1nWq95sMomwtHP
KQV2HR/O0lprbks+8WtzgbR/Qjz/gPly6L8P+Q0BrkjBCv+IKu4lnIG56lBWHcVg
1M7BfVQHijJo99qAZnKOn4I9iuf6Piz2uYoXQ5EMUA0mCvI6f83sSYEY7RSsbQJb
lHG5PSoJIFjuNKFbXF9EseF1a6a9dzH5DH5oWqQsQCxL82k8uqG7ibLkc+fMKFr/
hyfSuWK009sskdwV6+n+3hZ7pOgFhoESuOa3UJ2dTDS0pKduCOgHbRXWhv7XwAFG
/x1gpRRqCco3n88hcCBA+eTsfPRwH2ODRLMpVuxGQf4WEjqiigckLltKguV5R8WN
7xlkkGzQrZJNodgjQlLiyiBLZWDsLPKG5IhFLDzWoSIIvR4KKfuRYtP5iobfPTFD
XQD4UvcMjjKWdDwTc/A5e6uHZEPnmBeuVOFGiLML3GhqPZk7ZdN3WKE+/Ryb7XoC
le3QHjrkZQPJRWgTXKTkhi5PCUBJmnsiHhu5epqtSI21Z5bqq582RLvZ0g18CGkI
dN1eo08LGBq8DR81r1LsIJmWFnPbxTGGXxhhr3j7ubdLTCEHTHx5FS5oDzScFijb
5evByopSWQawV9dask7Kv5JhgqfodgcRmXZZjNedMi+M++FCRn3f+MOZjncDR/Yl
VeAc2AtI9Y+iLRejSMr1/6uvRfvGe8qJ/kvaoeakHD7YawJYN5503RNhEEZEm+/9
kRst4YbbFEhUNHkMGOWOaCB4HgZzpOW1kJbU7IdVzN4soVsTAIWyf4u1JanHDSol
kxWTCDWAlWAlVDz0CC9kEa8tvX2JcgFvaxzfeZBDpv2ccZEkZTUjfSr9SYUyDM3c
+CxySet5XQymuunmAvRt7jnbUvXm1JfhxGBQQSbWxmjOLIcgxynHEp4Yg1CdH1n+
taG+aIpERxb3uekax3Z67FdG3VkEfvHLW5taYZ6L6nMVpbIuLi0nHQMwsjzqmdy0
l0T0mg0/SCzfNNkQXuA7AFzdBmJ2VI+iiIdhsHAcWd7REnkKucPr22HFl12yswr7
lbbQfzfc1fYIV8lNeb29aAW4b/KWmcOzPgN3nCbx3Te+Xp66uUWtU5Wh/axzq7qa
F7IumTZkwfxKgHvbb5XwS4zbaxKaFw8oYi2jRFYtepqMkfFRnRS4OWly4DBXngmV
jf5h/kgQ6VZm2ElPdel73HhS+GabGToEg7MSQthMsRxiN4/p0PKXUcma1yuRmM5C
R6E/pZZdvuvZK7w4FlEOQlxKI0Y/4/meGIxwAZDwF/ELF0iz2DspyM8Cmb7FBgPa
NiajcUWIkttI640mYZ111/zVALTKPNQVbYcv7xl5Fk2zWw5jU9DBZ6ID9QolApn0
XtHXIHWodWMUtDriBSxtvnIunDmivDB1UyejwSjjR5caOo5H2zlob4zMi+V22zeO
pxlmNm/5VnioiI95oRMQ4/yzYSoMqbcKtVA4PRdAbK73zqppIUSUrU/ZpCbYT1po
yIdv1Ap+1uwFcpval+w5Hyh2gmradSAVZ/BraXGYrpcPepxtG1kylW7EFp1TVum1
ZnZkeZ0H+JfzzwCY0oD24Xlc90gQUSqcL2fwA07LXeeKgVy1UnT8DvbM7Ms9dV+q
m32kT3iz4/xWR9gezM/OuwOnqXPCarU9FfCBL3CmGnRyN51akjgF41O3yhHzIDi3
5tRLwNvjo6Nnzje7UZFZFj+5jTbKev72WxBaCeLO3Q7arxbJ56Bl3eBoyg9HPF/4
FiMyowE8xftRfGZZ9ka1QJnXZkaQ32A5pgrVtmkzhZrYHIxIpVQIByUGpzT8F/IS
c0xc02eLUx/EWtLtCI8X/UkypMn3zi0Buq0uZvO4NOVVjfmAD5DkJKywgL2vOPh+
9+LycKGKhPiO+RQacwhs5gLqMrxwN+M7+THO50eo81tIN9vChQKU5XSeGeeKHKIb
o0uFyHzJ9M59FxMM1tdisaE//RM3zbyqYrNnEVrvffvjGCTNpX8k4l/LvP24Z0uN
1/7UIExboXuFtkt9OrWkPfXZFQJzB0VvlPB7mNMssYFCb14x5P3vrlhOWRpTXnXJ
cjCXOTEdOSx6Q57+JzAgaURmMcjfjfPlJLY34u25YWk4eKB1TjxQO2OEevSX30ge
P+YMTEwnGHfgLupyuZ0itNpcfx5TsMgC1fPmQt+gqSG+jRGGxZot5fwdTX/ie+bd
cFIPp4JdVNeM6MLlTtr4Lgsvd0cyFlk560dCzB1D9hk4oCIVSPyKquJOuOMNtWFW
7M8SEZCoBtiIgaw2A4RlpeWUV04Ahu22WhjVxC56r7XyfOAXZGOADrWIgLGnu+pS
geaLLgc9zC3LALD4wn9wP9Fkjto2X48K/pbLksOekey9TllrBKShvqgvNpI6K3Hf
/dQTiYXkf2kOLzAQOMETb/7rpIMhsJdPDjoVAKxJN/rmESUD7KoPHaPGjWIYlGrJ
bdkZQ43PUWWR1LnZrGrVl6JraqG04HBmwdr/ratgL85LMUixHtnCnMvCbIzuaTkk
lN//VEbUkpkSxGmCgsHoX4h6DtpJqlXESbNlRMPzG8ttAgFI/9L3diUQprWrx/4X
breAAuuU4dqvvBcOQ2DtM+qH6i11TzienjtczG2okT+R/MVnCmy+eS4HEUE5BaTx
h+rnFc7sYzWVyjGeRzrBXW0u6kOeew3oXTkRTruKDzOF9dSlEHZ+i+QLsI0H+xCA
Vn3VHQ75oviWGfEpromliRBcyZw9sgnszitnv2sEj0EgTzLX66KOU5G96qkEQ5rx
QkAYMfShdoJkv8zAq06DVdZ4I6DAhYZV0uTFyAwmJQ0NyOKAukUK8MMSD/TD76gQ
GbGq0Osz/o4JmUGpj9ljUndfRUkDrsmBopEWavoUUn018WsrqDmpQaJfzy+LLWIg
mODYVoE024xVDI431+BYPQsYUebPQx+KFM/UgHVrvp1tmRaksF5hlP2Ikl1eLpm+
Hqcb6UH4raSCjad9JsV+nNYNUnuPasiFidTQioTWSaiai7gMR7/4nNWU6OrzTpEv
Wt6JIB/LKaApQBbh2RfH4R6ly62+IHw3t/+9WO4wulqxFK/wPsPnhl483nKxStCF
I/XqRkTR5DLAsa70mn6BH6UbMxoVr5VBaUhIsG9HuHYtp7ox4b5AwDhVHMO7/lfk
+UyW93MLriZlIiTSF0Yv8A2PwOMc6TXQBtoK+jh+czUxczziJ2+vy7f54X0EBM+o
pHGv5kwWacnWFlXEugDWfIoGvLGGM8NBcwAWmPiFKah+q/OYESB9oQDXSfbQdtGC
TVTwRRXobbU+TmZ7en1Eq2qfcYUD61teSRfmz/KlUukA3loZP5i5jJUt6dvx0S9p
2sqTJIyYbESLodzxL6ZP3xKM9SN1N8TUoNHlNO3qjVG8MvK7TBcj37fG/u2haqXs
2cLqyTiJsHll1KSkLABRjdm9/RdEgCI7m+OVMA5kL48Dx31N3/Pb66ARHypAD2+9
2vLCUI4qXseVkfc4es9u6z3WQUKLQhXliyUHY7QRJ3rr2vOKMSKK0guAZUlxq6fN
3XKCvtKUEL4Bxs8DqHf4iotRGm2VtE0snuo/xlU8WdzSVIkVDu1407DKosEtTbWq
ZmUEHErzL9WW2i5fi76EvWlQhVo98PCNe7QpQTvgcvXvdr/uYehLKtCAPxGeGDAq
PcakQdfM8xLWCbl31wdunX05CdZiMeZ6Rpb4k00PM6DJQiaWXIdI5Y8YQ5a3EHWD
POP0WPZjtrk0QmMO7O/LIzbkT475R84/xfBCBR5IM/wWKwKbubmiKcDjlK5U4SXt
Ac/JvsfrJ0Kbin1xNG53QaUZz2iAs1XI3LFNzgw10iJ9OP9zscqCElKKWrPCmo+R
hSN/BtqCvZ4jko4399PO2If2tYU34BCpoluOkVNVeScAzoZAi6NMGct8xvydC7te
COL+aOLCslp3FakHFlXhb7wNXimKzvFZiqQ403LIpXKYOBYCCvUSD+kpf3yDuzpW
Z+jrYd+P6E+ac+c0lx6s3l5vPgRUN8ik+knbLPjxDbIlm2GTbFuXFUQRdYkSOqQV
fobstGAIjAvrRqA2RCK1sG0ZGjDqsV3qgooZ9GVkIuvCk8Z2z3pgRhWx+oKkOr6k
ENVrkNcMEtQgZZ+ssDa/kXoCo9ypYxaxuqbv4Kd0SHs2VYA5mz1m5qRSD7m5BBp0
674zB/6XmqJZsfao/ZGHYGTcNdkJbejYRTbiQC4KNVIzeX+yPT1gnFog5or5FxL6
V77q70li5uWuercAsOTR21EXojhc2RjdlaK6dcVOQpmh0QUh89p3iWayWw1/EPEw
h0+i3bHbY9Qt1Im1wmSMTq75gDHkW63f7PjeTwoScTITG13RN5O2wH5yTMAf3Kj3
AFQnG5vtK8wAzcacHPN1Z1zkVGBUracVebqtlxQ/OM99fATrrgdI+O5NVsNceYla
XrgWGt0wWJHY4Ry3DrwyH6a/mllbfU0VsbXl88rDlm+Y3BZvZ8/qsDipKOedyTwy
6o3P4Yiam2l+escWtCpsFWKE2LF+U6mzmMe792+SChcWXFghRW8DnNRjcaVnpgeK
nZCmFWvXUm1GuMDBMgu6BgOl2pacN0wXzGEWStI5C1onfDc6G2osnchIUhyUw+5r
g/OkDS1Ea9YPsFhouw2nPUySO5jwKUhzfdLHS/2JBkPNjTS1TQkx19bgLgc5QxQY
0ZjZ2OH26IC+DeaBpJ4joHflo+RJy/rWHnBYvmd4XZiwkN7pfVgSg9ulDulpjRPc
adXhpYws1OSxJGntCsyJZ46/FOAAef9OECeJanoTNVIgN3CdY8YvOKGI5+3DQDS1
NAKKWqn5iA25G9TY7jBWiAoiPMydJTWkbLHRnn7hsyJK+2yZh5Y9CbMEIEQzJW92
bu7dArAnGkjx1alZHzcav/vgtmBEFcdqMcN0YAi7h5XSGBUO9tIx9f9xvO3w4EEp
13N5MOU05GYZJwdMD1/ZrqPGKrpYz0Czl+x4cTvuCXDAyJm3dQgFYlVtkAp5GIhF
kmcnhxtJRXwleBQUR+VHN9WQS6A3LmEbLCLlREW6NPnLnXqXusaQ7YobmBT5AWX1
FNkGPyP1loq6hHPuvUBZm+jWzJI2VA9fWVebB1+KDjM++HepRGczSF7aDdej3MUs
winncask6RPp+d7/KMQmnTWlaSPlm4xHTqxYz9VyPXNycEhCkeojeScpt9RGt02x
2gKFDjvlsf5aA/0jqkybQtbZgEm4t3HWgcotcAlL7Zo09m8rO3z6xn31N3fRnR0z
Sx1ijwJQeMYCOTeRFoOi2Kmc5q7RcMYaaRYnyEVC48XXOVRpDnQaFldM5V2MZzwc
IQPhxzvMDz8blDiTGBq4IgLoeFx8xd5+bEr9QLEGdizHV7pXsVm9E+DHPXnw5/tV
6RkttSnpOwehfFgV3IfzZlxJS6Y59d5r7wlZhsi0l/yRoHZQl+i1GPtxFLJVmx/6
o34xz162FuYPEP2m/ruRb3+ZhoWadBlB/tMLYl7JG1+pwylUswUsO6WguT3FsLBw
17UcflD/dK0WnErg9Pio5j1F3F6dQwl7n0IJ/W4RjsANjEJrIE0sfo65Ky/HNd6k
pIhiL9ipQ8ZbRr0GI/Gd4ZwGzEaeYYzhPX/680gOG8NsTe5PR3yX1sAj3QHyToMO
pz76jPR5RV7c+M4x7GwK/GGeeCtr7nF0fX6Xw2Q73U92AsjbLSXm5EoZ+sboiFoA
9JAzgLNCa8CS3Sltmk2cto5293AofarRLXnUU+VqUj98b4VK20o2ikd8kl2gtmC0
0DqacvvNykcX87YWW0QYSqo5HjjtsU24zoObn+5fjmoDyTVltTooHnzev7YmmYVs
qH3v8oTzOcQtTCupNdynYw20FbPV7WwimHKxzZZmOGUmqIki/h/c/jHhu/snKArm
HekG2Ff29R4XsztZ0HZ6mzHzlja9ZAFvxPgHetf/EZOR4/1Rf2WC1XN17DyuYOzh
JOtbK7mI96NZ69QmAFh/3EBCwa1mvbVJ7Gj8JplLqrc7DIaPT/JQ7okNWd1E8SkD
GtYMzm1yoQj2aGtwyQhsJskCDeyaYT+r0aW+qn5AvLtBr0NaC3Nmf8ZCzcQu1prN
dx9ErvHwT43ZUSMzuWa6zzQef9eR8JP+UqBzfxug0q4sMoCQZpIXAwQS1DLyEub1
EdMFmD7fx94W8OdeOnHqXtEptp7Ufx1I6/mTCSEnQ3ShS3zk1V5ncN++XDsC0Shg
MtkrVROTLnAeQUNu9Pgta9OwMivR5BbAJc8x6/mNcxEQqWwVlzYHypHkwMSfSurz
7603DKnEZ81OipsM7TI0Qkf9UNSgo4AGZDqRcoH5/Nn+LzpQ0PHtdhER60alsatO
0LfWPlH2csbadRVZ42d3qQpshyaB77tAw/gFHekJ/x3a+8JChgClbXIJeP9RBeZA
wFuunqssRcFRJORMTM96wxyKdgO/HYcF/NsQt/UrKU+QYo6rnKlhkIZCJNgBTknW
8AGfNkKnxXuFj+Ti/MNSJgFtxPmg/tDH4RWIV+2wg2G0Nl2yziHtqOqoYXJ+C9Zw
C7u6Y5g+XlHMsMuAOfFTU2L3xa2zU3X9Rninclb7a3ts/vjeL6/oWMGMqoVebyfc
NbqWIE5xBSsJnY2NYyeyGPnJhaIxEwuIvovQnA//6miDa3ugWUEvORvxar4WsQ1Q
dw840GooktnxoEiy77pLVa9vGPAFTsbztg5ffmL1Yg0hgMESIrtXO/yeZFsoimK4
hW7IBq8tCxAUOHIMar1ELewZmzKwdea11FLWwpZOwxhmZGrXLAWETHgBVJ6hYs1b
pJVRRNTGOILfkSW+LYMJtEfwvVNg7M43bmYutlB+o4oVqAhON0gEh7zKApzccA+7
s0AxwDLbc8Rap3HP3drdaCA9YYu0JXomzYpJFE1rVc/1pINX5nBpLLBTtBQk0TH4
tzeSH4ubzb7DWC5CNbpYlvUuzUhN5jdaH76LHPGminaFGPARRvBr6YuR/eRhpk83
QmjuwaO/My9vgjg4vorgztld4+ogHeHaYToJn27Ln1tGX3bQqe7ERZ9X1eZ9kQcq
ANjktBnk9eEB1PfEv+AVxW7CMtUOBDOEFCPv8M4CczMWvOX71muWjjcy/z9bCtr8
mWgTuQwfzKbZZ1OkXA1va5unEbPC6Mvf2//CGUNBR80AJDNtBCu3z0dKwhGZXSEv
Lu1D26bQDTEhXLGMO4BBmObnI/KiapGYMC7RIuZ6WR0EJm4mboEOQL/D3gT2IJLs
2UICBSi7FRyoQE3yYFwAU+8tb09c6wRv/DFjg5TWmKOeUpPDojpfnGjgTxyJ/Wbk
dM7koaYSh/Jsk59ktpXd8E0RFqX2KVBqlJ90gY9pgXJT+ipFbU3o2T1MEdBGpKdI
OnfQ9SAszzCKaB7Cu0Dd5VxzgCJgmn++0E5u7Nn+GENdXLgZcj8A/p9fwSYIMNaE
NMmUL0nHDriT11ejeoT9OXI+Qy9nJjkygbyIqCZav/F9AbtxBTwa58RaPwmJ+H7J
dafjFkbOiu9+VgNWXTQg1IRGKsMIE2b0giXrqvXBWP3h96loSPVCRGMB19mN4kxy
lKJGtcyey9bhyOn6sVBKnw7iPxm7GFjbkgYwZ8RAx0B0FBXRu/XJ39aCZs6ugUbr
NHBsu2z+cEd3ixzrA9mZE6zpSRWB7/AG6xyZpdXMAEHRePLD0fozW9beDIERWAuQ
oqEzdVLhs9nEpj3j03uzGWZsIs0KWLLSTf0dsgz62l8a6NcAthoG4OFTW4edIEdn
N8OomRHgspZdxwUGQH01KhzlwMj0cc6ykw2cJIL4RPmar3yV3zN2M1HBbDm/7lJo
n7Ts8wScnlj0qvgIw9TTqAMt4Pm4xgQMrXMQ3Y8dHsq0B/e+X+4/fHxF/dX269gQ
EcRczCCY/axKB3AMuR5LImIvTjvx5vb/q8XH9dik11xWALThXejFVtDdK6mFL00G
ivAmX3ymrh8Jii1b2XcaE36R7SOpBIZQqUpRfB4IukgTge7G9y+khK77sbVnZu5w
CUbPAL9EGc8Y4vEBamom0QaKsKjP2BtZzn0JvjSrs9PtCb+o7LqHmSgq4xE/BvAc
18LueMARSHxUEnbvyy0MwUwSUwg1fz4GKiDjIGFt1HzZvyL9pA3s5e6nsWOVTJGJ
jLVcSO6JqrvAU0DOLF32PWFk9SDcVo4rN78JphmpgRQ0rK8xEHRyvlWTIf/yaxzc
eJv0xj4s/94yqAg6zJ6bvycj96gGyLqIIM3HgUEb9dypUjGzY3EfsgHJxj5qokmf
MQBLFn2vll9TRIPflNVwBWHCbvOY84y0pJZpmy+AbLVwbSLIe7lkuQdxnbItrwsN
qoo1yvmU9zIq10TPZmbmN0gr6ER3i0Pto0QYlNyaZ+6TRU67Y+CYczm9b6Pm1krx
eN2aHC4MDHmPte4i1R08OCvYvNCIOxv29RxB/SwAQaTtXHyYHYnkYUWrwRhn5dnv
JH5rjup0yK1PDxzXbLTz9uuCbFkohfWP6jlAcYZ61HlSfOzKtXp25338gcVbHILy
UQyU8s9lk3TVV/t2ghDFyNHL+nI/1O1Zl/29ZO/miE/0NzEGGDb2Sh9Q9qWd9T8y
Bt2qgNpjYPn8v5cuhApqZMdZjQjf/gkOOSPoCs+x3ZGyi1xU5++mGNfp/uVM9WII
JOmaWGO50lbFR6wmN59hiSGdkeMhq26PWKvPmwYk+fgt1+V+CqmE1aTzseVl/kAA
/FERyk8yuYBKCrJKjcHZF1iqdE+m4kQiQdku/JcQjogZwNgxAQNVxET/SkCfn+oW
g0Jg7yhdtBpgUuup57BiFG4gDl1oHIOM5NKRQQyLUM2/uT6NxSHenryo2aT24cA/
bGuG4JuLH5Hb8yTSRyJQ5pjfUqrA/5AQZ1Z/PMPaahayRgtx82gmcina7WbsTtQj
vlXlbwUX9EjR7DuzzCK0UYwvL+bs+uSMscp0NUdfHlJWtCI5JboyBg2Zx7AE3thp
DwHokDEHGAK6nkVRDlgMl6QF0VpEx2VgW3LH0Ls6vGoQBNQuGjC2bGNSsupxPQFz
gRj3ImlSTb/ez7yoevjMFgeNuDJxwVXt2glzGeU9UEUHGDRN2feyxZ9ZF/7FpMJl
SvUvDk5rsX0hChuBTRX8pxRF6bFwGmN6yZOTb7iE6mwsMrMBQn1wmJ8OwU9w5cZR
7VCH1Vo6he1WXj8ksWiwJZK0XuRi3QTRj2PVuFsved4WETBo6+7sg4vKnx5eE0/l
/XRBLjuI6fUMxqZu2iiXZv4Bg0WCvdd4pVD43lC01ZIpwrkqciFX/WRT3mzVvdZ4
XDfqNf8JFwd0j6XJpYpLMXdlJqNhrlsEBsjOszd0v5TQ889fFrfuweGC+AR6zLQ3
Xo2O6CX2Gefh7Z5OdDSMI6HI4vyNQO+HH5Ubq0BQfjMP036LWHuOL1snjVSlFDZA
bM3bSsmy8naUHAyyW4WpKb1vm/A6JpQX6rOxOrWaYmnPBk34fG1QcZjDR82vjmcg
e0vnUYjTAwO1QE3jTIUCN/x2WG7bnMwWUH6pZSw6hFlM9hosmHyMLznrkJPNQU9V
BpGyZH+p5EUAB+lf6DdTwF1c6jBljX9On39uYTLIxMKMV9iiCN/pt1ZezCjOpXT9
34/BqMIgwsOuQXeiPEeZFKMauMr0Y+XjSXOJwj7TcA8YLRO49Imn1O/q2bj5YLTL
aNsxMidTpC9JGi6Uma99ND/WnHpyx6xDQTEEm1xqRaKdk5yZ8UmeTHkZj2ty0bER
5UYVbDUGvnXkd5xDr/1ikLZAwxrk9KLYrEleYgA+rvrSHueccnB5zG/mkJ0JF7xm
fQVmKF9E6InR7y0wUhauztCrMAP4l25uamy5Y47WhHpqsMC7Z0WOwBrqDoeJE32o
9yEdXCwjm0w/cbIYp31ZBf51m+W9dIOjxO0spsrXNjjdzEDf0j/C4NqUgsQcvwnY
OVLyiD1ToRG6uPpUDq+T9lrXHSIkT62ugOTcmIdZSecA8TrsdOFig7SHz9n8EWt7
C2DiTvGoPZEXMAhJ2FQfANi+QlrGt3b9ycEsdkZZylusfdMCEzOc5XLj9fUgWmgj
+4riSQ+9XVBzrPy1KXvLFixYtUNq/izNmIyZ4UuLjmgdxLfovvyWgYYGO/M+hyHs
sPY7AsvEO4oOK49gp26NfCwJiPuT9fCngfGjfyMLAWUdCtzU9flUR8YINZjbHpu1
v5T+wdrxHeDxBeVIZcsX3MwIK97IXCwqEnMyCshJzNUUl/Zt7MlQXjLEu/yDdY3n
4XauxR4NCeNre+BKaLcQUGf2zyTLQ7LMMjITGjqEbwpgE/d9xrPirwVJemmWRJEO
Exij7cB51sjiVAcEp+Rqea0Bi65l1B/9pmsYcp8G+IlxsYen6poQcC2d9/9AIKzO
3DtVJL2Uz4jyshG7gGhWhPlG35rXYphEO8vLIWIFo5qf7P0hzvvMWHgfSPI+rlyu
VU6j2GFqGkd62Z0dFLE0ORUQL4QF5TC4oTGlp3pY7BmrUMbqW36okgo9K4E+8k81
H+8YhnFTccYFwGODOx4fR4+CqtDrSOZfng05KzSRvEdfXn3yFduWoHsG90zSkCfp
TZB7QQXAu2oGrj7STf8tYYVvnNUmlgNWiE0JyvP/UhxWTHfDmG4S7d//rHAFBwef
8JM0q9Z2EelkvelepSh99OUcHfdyeYzzS2c+vns8Et6n3neseEzkUAONSGtoZBKP
sEtIhVyRP+Z7VNm2JK5ugfd8rPKJpzRQpk0K3IA8YTB7k36RCTBcTrqxs/Te1ZjX
PoxkcQGejW0wuSLzzGfbHSBw1nykE5G6g7HhPgabPR6xNlaKPrrO1siDGpS62x0Z
QE21dz6HzrIzqXCcxzJm26KavrPk0fM7wWT+dFEWW0w6Fq5wUzEQ2uYUcGnBF1Bm
KBu2QefEvPG7E7JJpwwH2I12XQ8Frkj9pXoImBO8vGj3XISTUikE8L+4/6Ex8OAt
r+gXB8kI2DwLDT4S6xIRh/tVBTGR2hoaA3cJezSOaoXgetvSE6Bx+WtWIpjNYRzJ
0O2Mdl6cthVzdCmH88qh23EE4wlvUe0Jm5gOBWFu/Q307v3C/klN5uQoYjAiRXnD
4M54YAXq4ar6SoLsGcDVmXechtkAh0M3k1TfqFb9ixVpSAkSy4q3YN7AaHGs3qQ+
jceV+Lpjyhvjhz3TQhSEVgCl2cQNPuvJLcR8h2YHU2tDgBSF7Vg1RzD2d2SWx56p
1xEwDQr01nFYceYnfYwy84RHMgCX1FtxwyrO6l1GGet8CpKzqR+NkHVbV0P02quK
7odG5aUPEesaRQEWhdQRGQrR6AFix71kWnHD+XlQJpiw2e4IMNRCCln/NeuubF96
lyNdxKX4zqNDDwN5+sSYPxbiXVUvFUN4guXYyH+mdkXnwPgARjKmYu7LEDIH10XL
b2WPhoSjNOyNDP8yeV0vgo1catA02GxmPKxDYHmsB6VH2rKgTMukqVFk/4eU6Iws
ACzWlRgTdu1oG4JzXMPQfMrLr5gzCxqxuLJ0NnjO0yFq8+GkjKzym2nrODPSBEwo
k3OK7V8MTAeTZsM3qGqkfoDBBzgzdfr+tsg/JxSSfFkWrNpQjNA0DP14o/VIs0po
G9VUoCM1RlWnJqMcI57I25fs1BqJPpFR8hQbJSOwv227LRnGfGhRwFtTH6SU9JCB
sjlS0T6IiCiNeBdDitExxirogwNjDn1mcTNlaNSJol7M2iWPy/nOv1A5CRf2y2GL
xB9pUv+T/0v4b6Uf8EUcQWFZt06RHLj3Qu/KNdeLqBNmeKxDJ7B8UXk4NzI15ta6
EKuKS0a9LzL4FN10MLWKDMQD9r2wiqVfzKWUOOW0nacZFEBrEXjuQYCic+gdNNcm
SaTSz2hk1Prl5C6MyL8f/0MN1aOBCOz013fW+V0U6i+PPGKU7cpeVkJOgTlsa2mi
NL8De+hL4rIGddQuqrKKZRd/aFfk5CgUnSDVsoZTp19VNoUyZH8KVB4osjVNZhDn
LR1Y0NOZT+RX/PPX0TeDlb9m2HluKAHWaaiRRaqgxr9v+pljZjRRs5/1fUuCW/eI
hcg+54ozoifHv81vBqynHzyqF5qWKsQ+xq8VGzdYlCCq95UYuZOeCMJx/NqOuUqI
IjUiRkGgO7vyBH3GS+2BLwd38H+aubIC+tnrRuHDJt8bY1Z3e6NvgeRcRyj4ngH8
KB5jN+XwxIlWIKuLFnnRZDPAKXFUi316luzLiWX7MqPs2bzb4IK8p4USbqeFerNl
iUiI/QauXloGzXVQhWX7MkQIiKaKrmOFFMpMS4Pu48YN+DeE/ugoJknEriBXKkou
YlbSTVoABivH0wXRWHCZ0kaiI90+9yT9l4DUz6pOeM8/pQfLKirlMSovbhDJvWV/
PZhb6wjps3gs799Brfql7FsDgOYCyIxRu1Ih+pxqF33PbvY1DyvssB6HYJHJLzsX
eU/UCXfpJo7tyaVXNOvFWasco2A3AdUHPhNkg6uYnCEXKZShKfuS9rWmgj6Phgrg
jpYxBMB3KtrPGJ6x2hF6YyJbysfgqluyfpa7skpWHJXvwxC0mFI8u84FldZ2yD2m
or4qT3PwUsYdFhbl8lo/rD3TBPcO0M2R63kISzXQ/v0AobWAy10x8AD7KCQ2nvIS
vuhzDxEWe2INWzejX7QC4o5ZU1z0ImQned16iI7fh7RzE4lRC4C4A0jf27xWDjcW
TjT368pnTHrA0D2mY58k+11qnyjAbQOqtmaj1rTOCmCR0O0RWd+jOyg+odmiuhRt
9hiKAirjh+P5dxdO0kKqUzgcbb9ZxQJjCPcMx3eA0r6lb3OYuixuK9iWhZ7KqDDL
xLLcSpKQz2dVVU2XpUkXw/4e+kaDIWIjQH9Msc4lwG0Ols0cV2mhUDDtHzFzX10R
sxNk9ALOyq9LiMpUNuuOEDoASU9/+ocs4Yrew877ro2KOoUzS2eRziZrP2xmm/x4
7ubbTOJdMnbypAwZmF+UCeOvoTVQhA87I1g3tqWbIyzR6oHK/RpVVGvl0J+VSXeB
On7I/HGdRqIULRRZ6120t4WMxS1ttjUNIGHRQ1ngTNMoxg3ysZnV7awlQ4OtO4oK
YSnxauJlXBBq6ewx9cwMnd4IdsbpUjHw6UcH176qR3lfaW2iKUvF+nfz81mqaZWH
Bfrl4QF9wXVN6IGE34jBdNLfnGJAcsoPljWfGsUz+P0YE2ldnp/4FOB0yt38LAxm
E8Tr3j0J2++SC5dwnRs97xckG5wNBaoo4Cm/GlTpdlJvkJ8r5fgUC72katXI7H7+
RXJpBe7oj66FRKK11b/cr7p2OedsSn999oVh+MexvjjDyOYcZMAGXxe2guhEb2EP
0tCBc0NQgaNlEKrGDL70yV5iUodHUxOxRlAVzeS47TD0rXiBLUnnl5H6a6N/6Xgb
w60s1xxUfhSlQKd/qtpK1PYlP7tqX4Fp5RwnjjiReb55iMV2s85UiaI874DNOhGh
5bbKXNt2w0OuVtw1selL4UNEagKR5CkE4cDK95doUo7nv2/AeIxsR7JvK6+Qoepi
W/Dwy9wAm5+M+0SeYsHzyEsrsPR2DOCBXUq9xmB0hm11H/skPUGmlSaE7kYVr/aB
g56wXPHkxyjZvhz4G1ofl3phA9EuRsweqjbLvWYfd8OfizduUvWIx1/jAgPkOoBe
MJAK6Tny/IRgHBI8ogF4HFeYze35b9Z2aIrZu3Z2W5saW9IAvZ2JV6ZZCnOgJXEi
xRmoQ1VJP1rSF9ciFPBY1rQktYaesYvukHTp6Jb9lgUSks4Fd/KiCzB/tWH7OM69
j5nN5Oy8F3EMaT/tLZJ5UzPnERpCulezHhcE5QSq8iVkZgT4hwI1eIf0+EmKQo7N
iMrRra4dRQP5Kl7jVyJiaRE2ovSG0i0SB2kPJqT2Jl9tdVX3BOHLDR6E9MuHE/er
ENRaftV2R2R71PfvM22jCYRttatz2R/POgGbrj6zwQWxvSzExT9Jk+1p4M9bYXo7
akzX2TBa1cw9KBWC3tmUrz7wukL8mGtb0mwM6Uh5eyWRzlElcyXy8AwrPI/ct3rD
ufzkLZDHrhpi/OZroxA+WTQ/nL+9Oe5lVIrXuMmNHy9M6gEl8naT7YbRLGWZm3DM
EVOMlnNiqG5MnVcRnh0WyCMyuQCOsYJ21KpiUpFUwcM/vYKGXuERgd2e+k4s/tqh
/GBhL/UEiN9TK5PU3yTa7V9ewsZBEGhk89U6wWgSZKvSwqfdqgQ/yer8Ow7X+IvU
86eQK3H1Mond1dK1u+7q2Eap27EVNWW2P2mWb8hwRNdlDo84gsusgjvGnc4EVd6J
ZKtOx+vzXHlFdVheEwyr5Qlf4wX6GcJkfp7yjBCOiVEHjZCRo6wHQ7m39+Tgrh4f
48jY1GtM/QaJAuxyTAAbl0QtTnCqdkwmBVTAqyavkrWscnKSlhTI8L1lWZWYDltC
SR2/cndGtpNjlvZhX9e0+YqiR7MQ5gIyCWt7oreFLtTTmTJm8ONvA6cKQBW0RsCo
l8tknpRqIKrrUdp0MZGiAe15RB15hGSZOVnJpm5t+dHCcU3eUi5OzY8Wpy1mt8Le
jvdezoILfiOPsZEnODhdvJGOLTbjedU2DIMaQzBFEZFeDmb7J2+FqEDNmqz3qif1
gimrCh87CSiCsqwtoAAcDoQ84DhLorekJXy5ZrxgYg117YDfbCjT3PozT6mHIPxR
ZIfFaiujj7cyZMwwNDALICC9WTupwojxt/iamNjT+jhe7/0t+Of0qxoVDIxT6jwR
AUFwO48AD++46GgefsGGOyEIDMOVBQg6QNktvPioDOWHWzbEE7PycTLWqQHz2rsN
k4u5sVHoZ0RWL6vPmBRy0DTfGeZ19UZFF7x4lCtsREzNHfyqFORcImEaw+/GWx/j
717NNp7M4uCupNaYlMhHP5FqcRNEX0YmND6xJrMJevhJY9jnTOc2A1ER2Kd3goMU
DCXb1+Z8/AZLLwwM9qJzqWLYj4qWlGTce+BZT3JOzRtHVH6uHlSl4LgnRaI2I84P
qoB9I9eXfBJVtzQsPNyMf/sK9TqcAy17bMsCCJNIwnPIIMAR4+YndsABr4r3XVKH
ybkiT2JoLuoYT/LEXqEFRkt6HrNgRtAd7NEhhtVvtznhsUoVzDeTKWOxiHUzdfLx
48fGt2ULnBZp3DWOtGH0NW+zDg/NHlC7fsmbp2p6YPQEQwQl9Y6nwZbMfdFE68Ba
VzLXMUrBFx6KrJrQY7UPlwuYwhIVYM4vpAIM57nxkB6DYZz4d9mbv/qUGywOfXLx
byJ5g29KZnS9JAQ/rlTXSsjx/zhqnInk/vzHNHqGWeWT+r20LqtchG9oKGgg+8RT
9AAE8HijCZYiikeRP0/cWL+noHYiSVKrCA8kCDPxCsv4w0cd+/uiKWZ18O1oUji7
Gqe2HhbT5GIWh5vXGr6t/HNN9M67pRIfQLvp3/zi4Y3KWkxksCW0/0b7y8XJWzQI
D5wq0LoD2BiUyYphymhf7Pu7hDLgKvXi0Ip7t7f8fDdAJ353SJV4xp6zswly7f5L
7urWQOsJLU2r0K6oz42ovvU4rydHz8G9HA00/6ICqEwZtm3eI6jb12wjzIJEVlOS
GMmDYwvqRJYtWTVLFTnniWPYyzV5qYsm028xa0Z5pA9PSebmUhCecin+/p/A1DuT
Ygjj2zArvtEd8PkVLT9QxWfUIeafB/Kt0H7pf7NcVkvF3KjEhnqN3oCodTiPXogy
Oylb5ZotflHPaMDln3Z5h6qOg/F2eG4RE88iE0BGk1ZomZN65QFX5ND1T8UxLP+e
4YpW0X0TixK3HksLiP11sW2azH1QXgClTnnjKHtVnNkD3cWqLOg5rq2iKg+dUmrD
iC/fRy/QZ9uRSC949YmvRyxyRc8KLh/1srHOWEQyz5XIa97QaWKuvsfDruB70GkE
V3NZV8+muUbSSffYG+DBQhVy7ganPtozZVus1JWEW0QqZmYJ8GHWMATJV6HEOAl/
H4qbvhXSN7mXOA+VUzWdSStoxj2lo5hDG4ktdwqNBgQr3nGy2X8VdA2mVnjFXhty
rH85WUQ60eeLdFi/2lmLFsM+HzoUlSk9Xuu0egKkwpeocf6kUACHKn62eV37R5tN
P+7L4ZwsNQoT0xVQM9GiIGeMgCnG+2PLMks+kth1lnjm6jyDB1xB6nFpg7YQ9wjP
R8LtoT1AK7s+n7fUiWsiv2500RagU+7GOUVA/BnRRyg0wiCE0CkntRLzj6U5lwXd
GPs56NL1e2ZTJBNQMBQ6ntH0feZ20cz/fmOPFUmOU1l318V3VCi1/iwjccLZeky4
sIAVf4bTiCCTcQphZT1/H8yPKznKFTn3Aqv4FM8QBPagvb6iJPrpBmF3/K6Ovbua
pDDHcHz1iWaqIRIv+JuXZfqsh4XAhtcLKgyJJaqiu+HJGtjslvrDkR+dYRUyw0Pa
AZBprSbYa7vG5lF8odlAjKOze4E86EVqtsL0pUBxp4kyC6WcEH+JAmNQRvvpuXGf
mcl0FMRq7RpxYWQWqCyFTQBbLQR/NR0kqrdisK4Y3M5EcXcz3LHHs3s7OgGNdU8I
QbE6ZcjrBa9n16OwTWBrFUckBqDt3WoRroOQuRnLzS+AGyJWrB/CaL+RJIxCHfCO
gvu29HT8MqAGD/tgPuEgRFt1NxJS+xAubCzEiKS7fp0ux6Mt+2Tgde1YP0iduAou
nIOJpUcJ+IhQqiqgcg/3mLQqQXZmz6kP4G2g1tvw1rJg8ETZkvE0m4xdcB+t6ieB
a0znEpF+6rcGHaLDoO4YX8ouxoVYbnGQKFvAfvQ70gg/1L7mmfNhAy+laEPPKV0S
G5+SxvgNjagAlIIbDlxqnYBEEruYr8dBCzjUT+cGSM3dAnwZVOpIyERD61kDvB4P
uSHZdqKjqaYRvg9Ryj/68x68S6OnCQKUczPUWgeRLZclCiESQcViQ3cNamau0FtM
i6JopF+eGJL9cY255llUmdXrtz6kFa5vquF9WlwbhyA1IdekdP+Iq3Z0sEvNZ5Mc
yP7eAWtiERc8k9drLQ5mdESM/lWXktKV33LMGCexdtX9jJmSVlx6mNnZ4VmaYePA
Ygoo/NCtIPO9EvMfXvNc7ZIiGunnGdkFge07M3MeTYsSuUZv6zI86HI6Bg0klkFa
FOA2IH+2GTx2FSJLoAGJZG7TPiafOMj39m+ENRasYXdgR/DYYYayqXbtNopRId6x
4c3SPyE/ncfvKByvDX2bDIPYAkMYKw+qpkweYIvqkzoz5luu7zvsFiD/p2rFlaOQ
5GlkYN5ZMCifVDFIqoq4wvPFlAK/ttYIqRj9qqWkAGL77QTm/3ZkW74ptotB1G41
1BpcwzjkNOAQFbiuVI/sINpT2xuRDhkcgD35tm6yHNU030rpwhCu67DiKQpcYG34
WvjYN1b3ZJk12K6N2yUfwsJmXY1kwNphtLEyCNKyVCI1GXrtNrBxoKSu9NIsfKBR
OfoHodwz0/n2zsApzUdYK0Re2ngXvaF2xb6CbHm56e68onaPH1MAvxUVT6w/HoFt
x46dZnE6QQRyiaqZBMTxFP+qUXPp50zSjlrkM2MMxsVLX+9iQ1TyvfVhQdJ8hTaa
ZKpNlpPQLOBitW63UYhhUAgKwXlMKNPGHlImXorTCnA5s95zTG1wMq8fy2zM/e9/
I3g51EOcEcnHrEY8/gYE5KFLTxoT3LA6FbaftvdCrWuYH9pehE2BlgZ+wSLMm3i0
fRgpKnn/c0mrqK2XEhjkkWGE+ngOB1byCZ919qaKHViiLCfzogEzMCC8xDZnBpgd
SSBghMPu7OV5BLS5V1Iy5hMcZ2nbaddZ6VSQ0d21NW2zYBvFr2zqSt0Y8KjBCCVg
8WgErVpvFdSNE6PGeW6fO9ghhCtj6C4GRA97FMFTibiZ+nGwCJibGde629IE8Itv
/vQ1hkKUhJgxEi0EP3XYNnYlE+FBA1DeMxaE5MMsy3a2+53YvhwYx73SICkcB0cR
GY7wHkiIQSTb4wflo8nrxgWIHc2RPCcihLwf4sYQcJJ2c5hcbx2ei7PZQ7i1KnaJ
7LZmket302NYLxN8ibOhENjHloR9llO+c6NAt49OpMFAjOFCPLayvjvBbCsIs4LT
BZAwlitq3B6ZDmp5PitM4Jj0FTQnqb2QUug+Z3ih8rOr10Qhr3Vjxhji4gD4ZVtI
28KiYXtAUIs4FaePdl51qRKokn7VsstGwXVk5bU2uvpgGRtdgGNABDgaQYg42QHH
AGIv3ti50k3EebMzmUHkIMiWbjPOPXenaP4btSGzphTIsZmfVhmIVjcXI4WmxvfK
/E8+QpXuRP4pZwhDQ86PvHz+3YTlw7sdCfWFNmoBGNitrAPEsYHB0NceJI/VTVDp
wi2lO7UQI1vTf7byhGAr4kYfiLQd2edMx41amZQ3+zYi+wLW+wnVRAxaPqbpBWtp
rAPhy1Aqfc1XTvq0XYgvzS6NU8U2F+ZgThxmZ5S9kZStj5LTU6vNXi4+HePrAeI4
BbQmi0s8h20jpp0mJIqLiTwYa/HbucrcsoEEY2V9ivkRisG2p/SCNy20ASmjOHKb
PsY/fd3pL+DwA3nMVgcsENh6I6r58XhlrwwtR/YvRox3qQxzky/jB3R/TdZ7+dok
siYVjh2Iffx/seZdVkbAINEZ+NtWdSx2pnDnUZ65blsUaDkntxjBkVw/nGsMgz2Z
+jTm/Hy7WBI0PYbTb5c2sJiLRabyo5gtHWIt3GxtZqCcuUNJAgemtLSHwF22iFGc
1hoNUCz6CD/yt+UB7PRVxGVQSGqCYfPhCp4zk6eaVcxZxhwpvJD35vH3hP/qVGPp
G/OPles2LD56/+a75/4Hx3nGfOwie+9wkizK8LJ/FAGNbLm0o6SSYec3RrlN4xZy
38yl0sAyYD3kq/kGVsAjRnN+HaBiovIwOTs1jwRT+xdOeXpTTvx+LJO2Q4J/XJxQ
toyJqbC5jTWzc8IOh4EliN0y8eQgT09td1dNgjM7YqItD7T8ducAwDEPbVftkReP
LXgLrIlOqRsnbv0bkR30ygYpr2sVOg5qadPKuA4ILljkqKerrNCuj1AvtgvvIO+o
yuRYxpM1WMoBaUllqRR6plAYK2BAEq1IndZQvOLCqWy0xzsdR1bgHheSVcNaB27C
5jl/uGmtGW9OxLf9nHHNA1vpbOPscFQcFNmhZYbl6sYGghVGCuWDioCqRjgVLsas
cws/as2zIf4eTW3+uiPSr43O/eaZPRaYifcmX05WEWuKrFamHXRJQ0Hu6g8ZJavm
E/s5NWnA4GR0J8CGa06OTPJYuT18y2zoDKlrwNCsEoX59TncwjPNjFMY747H6ZjR
Q7y7I8OhJjaYn4OT8zwVxTJmwFGiiItLSLuOTvF8x09yi5Y/FvSiaGmKNwdZCGuh
5graAok1wfPSBT4mQiZU0mE5tSMT2Oc62bk0mp88BlYvw81tq/QDuCKWDOSsIe9I
zNeQrHLzMs2FsN4CC1MxSdZ2jeZsq6m3HBbrJOn39cqwrwKm3F+jsS6KQ5ZoSNgm
2tPGTZ9CJ9EQoVYOF3Ramqs7YfiM2bLJcxeGdZV0AVQh1qDyWoNIeAFcM8JEH+8x
vxhPQmSOjPGt5HBfFXIsA9IcdXyHfDYdOwLXj19YA8essbhqe/RUrh82D7ANv0qb
Cu9OyavRyuUQYVtJu73NwFeUNm6GcpaUmvT/+QkIkuzd4NpB1PtoQOi7YGZ+MAdi
yGb0GVQHq7P/t6cOgCOwUT4L7nlgxf+ctjeqSeCd/4hgL/0m5SFLATBWeGlcrQkH
frbBuei4dWANLNkIC41zTqBkcNY3IkjHmGltcBM1gjwQ4pJBjN2nxYeGf/c2FCGl
YRWmnoKpclCnejTYNcX0XucX+tmJiNpObPvB9oGCqEJoJwXdwDFvu9w+41T5zMOs
LFRLwzDSoKHin9aUuOzORJMa8qV5AUUrvRi1hAvmLzXD7zAlZVuX7SdKsKXgckX3
AFAUu8JZvTxkrHAXGEesUE531USdURLaJu/i8zdV1iIUaZzex+pQ5cP+vmHRFBb0
6pemSpIOzY2r9Th8yZUx8gpduW3S1o7T2U40Jb6CzYL8U3vXU2E+PpJEDEpY7no5
a5jGg0gpuawX8DO7DsMAfzWW8dm6w49B19c3LYa2fu+Fj9CPPA6j0UxQcVgwA8vu
zdTvcRaXBq5l8K4HhG/+dsrnyg9QVvs4yVhVR0zGBCfARxtvY7LUqwFgWzXmucbr
OCUx4ekXnqmXRMvpmA7suHNxK4RVOp3+ovO436hdvCrteJLc2oQdOtuZ45Mp18Kl
VYEGsF2ILPwpg6P7XBQS0ySP0zyrbw6FgJlidPe1Fit3XXjUhbi54Kw41exjx9vI
XkoUigH3WxF7BP7oFqwTAHnRNuivooIk6EOM1McBWQRvLn9H61qGh82jQrxkNMqb
HAJEwzcFMtU31D/nK0PXkvs1xqbP8+LQgBNtiB7MSG2f6m0Urd/y80MDhX0EhqJL
YKvY8juMLmiRkEZ1UdMtgNqfFku1KdJZ79lHL/xX0VLunnrZ5CUChEHX4vbGFfeM
o5RwyUS4nBImOWDbqNjdsr9zFco1yI5k13vIFGVOuY/7fIzxcCd+QPrLFXLSeFnJ
4CR+Vf1VXznWwJxMqmEy99CqtrMhkI/BmfUV72yGBtGHi90uZnGL8ee+7zTB/w1n
UC3EaKVoVZ/ifbVDK7fmjCgC4wWt0KYBsnq1Qhbs8P1Vhdlx+hNUn6WMW0CVYHss
77tGW6sgsOCTd/z0si9RqpRZF1Wrf74V7x0qSADScWKHVjbG2/s8n6APYYWrJUtw
3yIeihISxusJ9CUnfzeHoTg1cOF6r3+GuSQt3w+GkELx3ssgq7dptVayrQGJUS5w
RqiG2/7/AFBShlkIg4ElfgTBOc3frqjpeUKagTCf+NCeJ68KYtg4WVJKamZt9hSJ
d8qZ9fEsicXi7qe3B4yFdRvc0ildC8tSsabRjkFkez1hFUhXPZ62vXoRdk2TD4BZ
OhMWalEv5ekQk7gZKhJJfShypvQmnDVl/Rzas2ILwwZf8TPMjwQZ/IdDAS63fgPc
09kzaBQ7V5Z56W+fampyfbHv1bnq3Mrd4ptWmjKS4XSUBhMhTNoszGERidd+7zol
hbMAZ/UZPZNfqd5fvp51fm3RUKmzIsRY9c+3T9b8tu444WONA0fTnDhwdzWYmtJF
pmAtiRK5bDd6tcnQ4XOG8j4mHJnmMstBMsPEwGjOzOa3o6RsGDRlyjutFJK0ZtKp
pWCwOEy+5yOv9NI5aNDRLnn6cQhTC4BkxY6mXT7j0/1DpATFfTxsTB04d6s4z07Y
auwdO+3yzbjpe/4HiEQjP+L9jQ+Ve4+r/Yhn9CzuyoCHbG0xXZJrE8wnDw4NfDkD
F2q3nomypbQrLRRtZPMA2IV4adzRjhZt7sT/nILfYF/iAjaq4V/uwqHHhsjaGgi4
apM7iuu81pFo8/zEOCnJMMCN3UpMH9eMbmGCNeOPyfvzyO6GGi5prLSLd58eQ9zt
w3eQF8i9i182NEg6/cxqzjHyYdgu5oXtKsrFiuf/Jqep8yxdzLoAkTbm4vwDvx5j
7wLiEMBiAwPsGNsq7mEXtdEjyzslFUrQh4v9jO2iByQLCei2nr2cag7j3xe2PrgK
1j+X4mI/mUIZ4DydUjIupb2Gh3JCnuz6XvCHDD8joa61iQni/jpWOr+QBc2dYhrm
8I6/iafk61T3jZP39kyb74ZXtAKpCXjMv5LyjJPDckyIoSUh92n80KL+o3KLHjm+
EPiJ23bWef/GOm4IWorm1qM7Fh9RDrYKXjYpO8vw0bv4UdZnRg7oUWKuqtcbuvbH
Y9A2BNttXbx8Dxj+40wEYpm2OSeheKXaaqpTL3ePPrNVbu1TYcIPKfFfaqys9yfM
W9LzRNpEmdHfOPMOYqdH39m9EkijsnWOEjmYFy3kPS6Nm4qo3v0qDipJKrmxu3g9
4HVrBihIGR0jE4sucoPDgU13PZRUkfVItTd3AJDjLjrt+qkETnQpywEbk7LyZgSZ
KSZ9xtQtG3u8LL3Ue1JPSFHZn3R+PHXFFyUkum707NQtaUJmX4PNelYhay477mvR
uaqoRrcVM+bWUKsDR0M4DjzAPhQ1Nw/3n2D193jJ+4WZp38rSQzhTaAaZ2pD2sXz
Q/glUaUJcU3F77Md+uHLk78nl68+nQ4Z3pUcpbsFj1amKYwM/KUdLjMPx+DDsNly
RruBz5tNcA6df4jch/kIV8tQ/tOVMTuUD9H5ClaThK/7hpunA8eCIZOdhJe8oV4p
6+aD3hRlfnYmxNjGMk127co2R2hPEVYx8IkIJ/HYKmIwqCYHAYRVCDOFvKqlfrrV
kRfzpugLcaNUZBgQwCbEmi0UgzyPbMNQR+1cu186i+rdEBE2MXAnapTQ8IkED1qD
xHhenln7B2BrHQddiiqJHx19G9dGsxLLeygJN48xTxReNSrWgGfkuXuPS8TK7i1k
NfrLpo6ENqtd5M9DZrL7q1+GUkaV5wfi0ue1AyzW3OlvsN+MmQBUvai8mizBfdnr
kMAtQCp6iRsfYwR9FbusD9ZCd/WSDmZcRQ3oBb/D+Jj0DG7C+dwQ6gQRpi3fQLEb
HgaGOOXMl/c3R7iawSl1CDKBPr6UOh0nkkdp0/gSDas6fb9pJqsx4TQ3rekJ6A2i
YOEKnP4rVezAyYuHDrF5G5caMicEQ+d/644/0HOSvhyF6DJ4Dq0vk31j31dnVvK7
d2NIgNdtPwqUyy/A8SF0vmwvufZWoQRK4A6OSWE4YkZxuyGxi34Tk57GgD9XktjZ
TO0CeCNlrHqDsLC2ozZbLn2hsMcXqcNJ/i8rET803/R+k7MBBR0P/RaKvYZyPlFa
g+Ben1Q+fDL1ZdnMHc3NtNCwRT94GXDIgkHw7lgufkiaHyI5LWzLVHvv/ct10Taz
szpdhLK3tw6j85vMBcM4vfSdt0Cwl2/DVzJVYpCjNXaYnLRPSb+EqJFn2hB2abwF
I1A7aGCn8Wyqzygr0Tk7ZaluqGOl6nX9qZo/XX3ah0DmHoemCC8d4yVo7X4sc7i1
9snbvG/l4hkCrb3Oe6z7z36ARBldmZIxhkqxdSyvw8VlXB4+T32ZN+Ogl5cF2Rto
YxTIOyF5tPVI83bCt4YvQ6O60ZhZH4YNf0yG0cJfccHGDks9bYZzLnxZuonj8Kh3
PZ/6f6duyToIQn9xg6CrBm8GtKx9P4jOFE9Eu/Lei3VrnmDli+Cl9m37GrF63NQD
84wEXpviGyoUQDtt3nxiTmB0KnVUlzu9ugW2UXvXL8SUFY/sS1P9IqjTs1R4TOTr
UPXkRvAcU+eAFDKhff3OA+N5VIM93dVlenFjFKfu4jCaF7lmKCdorG9s/prUn8Dh
mfrIUNqjrwmaQyMegByq/7GK9WpibCfUAWzI1VgryRAu4cmds3WDxgZeXBrdJw7T
l6WDckK+xykUkYaEX6KqflIfJsmVxzasgRRqM/6USl2LxqljZePYcHjsefkTK9us
AW/iys8Ac4Pp0b7espEfdDcUe/kouQf5Kqa9RqCjlp463WL718Rz72Vd93i1ZGEW
Afk4uPXDgWzzIaxdWxCKjuoaamVrvN0OcSNXCk9xC3o4/e4gGCWF25CahYUOfv3s
503xkXHBkfGRNTOBUdA1JA/QBZI7tLoRNpX4navCxWiDMwN3L+3c7xLUHkGp/yhW
ecPFE/HrMqIMLvZ+aOC56tVMnTU3DPrxwBsYIMvGZueJV7ho0hozAaM3zKtlTvEc
GI/tB0u818zDm9qocY0S8jU4vxqT7G7FWfzn8NEhyKGSF1Gn0fSAlbOZTXYRYPBo
E6mdXVMGQe7nQFn5T/4Wf6V6aI9Mws7NEW3YdCeBW7eBQBTf3dwE1rWcjkliIgAi
SF8QH5BvzOPeMt04/0uWHfjJ+A+SJFen5e1yRy9X8LNuU96oKKcabd51UCN7w+er
PP45mI/1wjLfr5XbrFK2lDzHeHz8AEcEmkTaESMxHc8EbybnB9IB/+XA8fgF2a7c
UAHX9cZt260XRUv2h2v8bc5Z28WfWvZjl/hX0CaarWB2cpHlwWUMerEV0BCvvnG8
X9ht37kvvUJ2etaltC5sl34BtX2UV15kyv9+S2JcdwbUDwy9eawe3Tejzayv+x4y
aOfw+QR8MD5qhNwzXHqa4Jwy6qZqM4vcdbPkdpYbOsoksUx64FDQ6dICoFMicVrQ
IjrBz4nXvP1gZff0ZQrvx+bFd+b49p6eGzFMAJ0egdcXFZ+P+9LJit6R4ngUmA7a
o99LDjJgK/OrtH6HX6oztWjAlS4M7p2XbSteufJvTff92j29adLuH05147f++z25
OcjNBKhdav0NGELY2SNRWzDaxTHuY/oVbxBpk+HvFFo/5r0C7uKksZmX9oQGQJVy
xp68HZbMosugPKtxXvAx3Q==
//pragma protect end_data_block
//pragma protect digest_block
LNrMFu6TuxoeZj4SuACoUZryulI=
//pragma protect end_digest_block
//pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
liFRn2+8vlNZqFtgK2fBy5LTSvtpzxXBB4UKjpDp1mmn+SJBcLTtoD4daMAwHn4P
E/9ZuUnmGoDT5dcY6XAsr67nv3QAcfhzPJsUQ3XkW35Hde9qQC6ALOG7rp6s2k59
1eCqwcX0TI4oMi4mW0Hf15Qy5zZxC0YrHMSq5N6dL/4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7568)
7MYZxeLZkEhKnAy4e+g6CzYsq6hZ9L8KmIPnZMVz8sMWYy/pLEtfTM1JY8MlMFvi
3xfJ/Hoqj39KbroIJ1V/9Uui00DIHKNp00UMBk+aELz5lTlGzk4LczXcv5XXQdCe
7UoJfgEHhnikjtJ+sUJZvn3LiBhSGv/MZzHTNINRO257VawzkTRnj51DwGWJ1APl
OkZ2TW1OZRCOPdLqtsakf30XoeGaY03j1jQEzHhzWJfe1R2Qyh5DulKaTTK+dH0y
jYM+OvXFRyz3+iyKTXk8uZRmmUB0z9JlTyHAlAbTyMEoKaWWE40LwtfAxHJZ1Oe0
kLqD17vWLWDLV9h6nSMqVCZCvr+tw069cmuhAuA3h87xBfumnCQdN/r4NDwjWPem
Iri6tLWferqKrXB4JXyqEJKEIIHw7DFeOFM8G4wKZcacOZecNlcMQjtKd56h8E9C
phcVex2Oj8UavX5K7FmC2sUKpoTDRy+vEE8IOIoAX8ZYfiwTJ51Nskspp/sa7iO9
FkMqqNh5f8bZ5jBx/uBWeY6HZ2Lz2xC4zXQ3EbaZhCa4Pr/5wbCiFw+pHZx1M+3T
Y+Yac1nsOPN6iXjH+6FlAEciKuWg0/6icI1yMLUvfe189e/jwgG3rF61WaFY8XBx
NEJLSiyCSOGz7QLW/LE76ouBwTg540zZR6/fHu/+gfpDIVdsI8pI0DMydF8bF5CE
O4z9GhOTSpqOlPTcjxGsLmi1kySEH4d7bSmAkU95NEL0/oiODCtau03s+8xFmRkd
Rnz5gIX18Z4lkcDeJA4jqqIIAyE16u6Lyxz5G/0UkPyYlIAp2K5Ngo8Wkdk1aKIe
PqSpaJgCA7/ClNGM/MytBbatjzEmZZIx0GT3tp41uPuzrsOjLCFeZS1jVriBgUdv
lsKEvEK/pSxlAjrEEF4LW0n8K3VPGVLHCr7lZrAHmXCieu771SJOAGvqvw0LEf/R
79pAlZsflQdv48GbLDAefbk0lFs7vi1kiWObzNVNIr6u2WifM+rYdmCuQIyAKf84
3pFJN1p+qZefD9t18bGJMnXy3Jf1WzWajJOeCuZeBwCNp6gLuUtWtukXH29AMeua
6/VvpbMO26Lx30eSExoCkn4jH59RrLC85k6yr59KPd44++srrbMa0vTsqzlf7DBv
JBg8tyoPC8tE7NOhJRME+Z4SyS9PMGlz2hw9xHsBo7jEOS61DyS2Xhaa5yl2brvd
itjYjUfWFu/ihDhxmHGToXrTHd8Ku1Ux7sSWTyOVDLnPBfpHLYitVluWXgo/POuC
92zYXCB4Zym5UG7QA8PkuD6IMhCZhFLTz1jBVbUlm0FGwUJdeszYmA+VSxzgzvXO
N5yA+FDyIqaHbWS1Y97XlNK0MtBzdREArr2rCbb0u/Om7dxUeCnoFFQjgStktA2U
lTFW9MwgChOkVEkFzB74VBJa/v0qY/DgQi2mdoHWeK5FZNPc9Vgc5LzcTZ4vGzRj
W5LbUOsNilqxWUsqVNcXVCnjnO6xkuutJ/r8+aaJDUiSwnaXIGAibbIJri7N1L2v
SfcPww9Qzv2In2hudhWX7vj3REu7mI8iT/8gAJs45nCeFCT/JWx5pEKzEMsc/pNG
Fu6SoT0ntODqjRElW6PSHnRw6/3iVCVujdvNlWhzuviQsh8AJdfMja7RjhfjAIjH
89QPn4RmXhylvCMohDSA9BxiqBCBgSmEOtnKbPT1g0iNx0RfdSvSkeWIKdHKCfuz
PuKLSf8zxoxmSzRKYBeA++zzZ7mQa2jfEQLdIUsDBPJKoG5KcRmUkOs55XmIiY9O
0MWKoeb08ZNIpRTgC+UbAYHfqRsGGKoYC+Dy9FlFYO0K2Vj4Vyz8XDZ8ZOTMs1bC
G+ao4URDE0cD68A2LNrifz0h+Wiba/HkJO3qjA4O22plmdwm0Rm/5wcQ9Ea8lRco
aAexBWcBPGcoOkO+qI9kv2RvsoAbkZAuqoPiNwqozGnxdiQUebqJt/E7WKCQ/FB1
QwyS+WFl2Uc7GmVCuztcTUBCzDJ0+FcYzOSUxE+fCgncYVhI3iYVh5VDcHrhr2Lq
/CUY0/vAjGkew27Nc1pKs3ldjkhAqzYw7kOF2la3l636bEw3cTfVUDh7TLVZ6u2t
2ZFoTPOtMwAeqk6k8oKVwiQqJS9J01Jk+sLG4p630CC6a3+gc+XLzajmAqucF2vm
QXnMxUQ5B1/ydL4l88zdJVjTMuuOp3fOyo16E7uwo85x04PFZ68ofWX6fm222zZC
bY84F4qJHPTILwTGKfJCIAA/mJ/NHQTLTo7rNjkdMZuN7Dt3eJINgs402idHhWVH
+BnjBM/NnJftkw+yOZTmMhdfyyh+F/0WUtE4uFUQrZd2soJy827zLFWw5KHoWRuv
ERM3Hy+LuROWofj3elqJz/WohaFYJrmutJ01kcG23wASXq384jLnnOql6C3SwULZ
spSMLEu9+MuEWP+WXrZPBMfAiCEybDS5ZYKwufh192hbkAjUiJOZEtzszLsp7Mgl
X9+oDRanJhTx0EkUiN4kBbAtlQHW4Tihx0rv8WC3T4zvpSKUC2pa/4TKVr+j6ghF
F7UQ/5JBi6WqLwrB3OeZrxSGTOTF65x552IJ77RGgAO7+/yJ4M2BTBiM0a6jw9s2
z40oJvCyvQuLoMkaYle6TbslL/lgrFE8a/If202H+InbwlBI/H2uoi531b8Lltgx
99CuRwa063GqFxq9ht7+RA4VBv1qiXw8/59f9j6+ig/+cr4+7hgOnrTORaKBFgFh
LUQxEl8HF9Y4b6fX8TdGrvYROXd1iW7p+3op6rWPe3jpRfcNYVqsBGgNqWKD+p4D
l5VdljrZO6Js6zDXYqdtL2OmiCQbZ+pqo4WpB5QvPDOh2T+hc7hsSq6+3/XtVHbZ
Vpu4cAnVSS7M6lrZkOhRUmhV0Oj5886p0VPuCaM+nLoqJ+eqp1Q1O1logv8PsGM4
A3WeWiXv6UluJNiCud4mSoz/Q8kCMgghHJypTbXxUomwI2xLj2M2g4J9UvXPQu+C
w0A4ejTs2smTZj16Z4E4eBEu/+uEBMe0y22EOrxpCehbRlzK0xDQQLUhjERg3NKN
8elC7gYsLL7Fg3W6Lgh87QFdFj306Bz/0IXWYVCr6vhKC/fvyK+qNb7XUxJkerd1
yhTkU7uJeJxiSVxLv9PmUtJSb/m/NzO8XlX8m6osNB2eQDIId/ZI973PTf/3qL7o
Q1vIQ6lSq1zGC7UdAFxqqogA7vpH3GWeYhWzzkTrImTkTDWxQzd9DT5b9yOpakq5
dF/ycavWW4/VESBD4cQY3NOOrT43L34lTVEyW3hN/3lXTHgE3LiZb9s/N5HSuNfD
RHtUUlw9eE2TWdlkNAhJc3TTYQcQ7SBuBsLHApIgKzVsg4xpCAItWKlvH714vj6S
o3TXt5RWYP1upLgVuv/Zh7n7GdLbBSz84EUa8D2uyKDeTvasq2GAJTiRr8Eywk/G
Oj2+BBdr/sR4I8F8VV0eHYMIgDBsl87nQfn1T3OAVsIydMKzUKB5w09qIZh3neKK
8x8+bzoWMcPa2nKi7bRTtgL2xqaKsAZzSox3X5yJoJQOgdrIKLIiImjYI/qEXXsb
ky3jUlFRnWfhW61GLXs6H9wE6Jp1t8Y49Dt56G/eL7dw63/4ZpvUG6NHTPzAFgvo
oXNmzx7SQmdRrBTWVRnMB0IaMzAtsNRz3vACk0OrmrqP33/laoR3WvA4vi6A/xj8
8anEuonrDFZY0POJGETp0KiO8UqJ0JDf7tUYup+a/whoLqd/dQ8c3jNIyyMH3cMI
vy4Bpqfg9VEOfawT5HhZmCDcayJSsbi2an9F95o18Gl6sQtlLJosXcag6uK1ATa6
BKXePz8z3pv4Wt3qliowsG84XXXV89m1ky6YtOTl1HiuaPLyaiOFncn9cYSWS/Ig
Jxil0MxSjybffNNuM/GexcEOQpuNkNlwyfpEqpjnwMPh/zQnS07chIENYaYk6G4D
MlC3sSRQyUP87XoJsTl1MuvDVwvMbaTwUlbM+q24Xi5PXZROXumevfgTBPcSmiW4
XHlBNC/8g2QSOPlpKK+QwihGANvFUSOiXdZCwur/i0tU7TZ7+KTuAZ5BM4lZYA9v
nkqrJmeqEo7rzP7jeVn0N22pQ3gnKucVNtRFjeEqVs2a9PS/kR211raOu44lp1VZ
3XMjAxLyNCvJ8/be+SwdvhVwWdPxF8r7vh19MGtRdT3hD8bxPyi9Ip3+M8xCNwIG
gzrNcuvxADBz0SCJ+dOhn4Y5abiFwM6/SPXzXmOATlGuzuVjMovxNLFC/9iUdZJA
mt+4TBnnJ0hmxvjT57lT6LqqFN6rRdDDTqTTQWZm+EbQdkrCwR31axqOBSX0dasV
SDn4gSPTa3Bt+dYFrsGZlDWvLYE1MbrNyeQ4Zk5VbHwQCuYYNTMYB52EaKEYnUoa
GWIalOYvBzMbBv0bqvjUo2rp9RQLNDZ72gVmViePy7ZhEtXSP8GtagEsiMzaU8Pn
OriDC+FEoGwHJSl3QDCZuG03rTuSpXGLD8a0Jq135OVi1lyTYddXaFm2fNkFULz1
O2ni60Fmgr+CXJFYyTxZWbQm3s68U96FWnAUN7PFGLhzLbtPvEYggxzAlDiyuv6r
2StywL2YfEoIxymEev2JkoyWOU+PRbWu4RUx203kUlvbIlUsNs0qfKakoTyL0GIN
C/lILPvGy8/dEZ8OBbHWtfmT2566MqsjztvBHiBl8dFv3f9iG9HnkWUrn63cl1/B
pZnHR+4BU8sPl5h3nvguOWgi70vgGtXGYwZhtRw8/ysESpGwQWvUqQTSnni7qSCg
LH5ODtO5Vhucyzs9gYt4I/6cRKdu//R3r1OkjiTu0gry9eiuBWYWNZmdOX6dnR0b
NZRn4GBEi9kqFjOjom9S455qGTfAu/0doBfRSHMiJntvUabE1y/hV2nXBStt35HV
5Ub/7tpY0lX8fZseem6qB9SSOEcTyvYYRxRaEv4y6g4InEsXS0oHjEWFPc7uT19q
Nm1EhHl988orXNt+BWQDjmmuSrJAP3VXaRNvYS8wAP/5biPtK7nz82W6iYpUY4Og
dK2v+47Q9SNWH9tGBbcpDNZJ+wJw+Fy1e5V0eKIvZNO1f2874eqSxsHj08UVLFq8
WBlOQvpJ0dS01v3zVmiJ1AryTWjkrg721zSZXXan/bl0lTs89NE+UL1b1h70coBv
F1R2j7qCCretb5VknVPQ1YCAAwuT7v4unPrCqpPdEKYoBcFR9GmpGKYj7VLPaNfg
r/b3+DEVQguFr9eeu/ztb9zgUdwyhDynQ8o0CpNmB4e7vjiEkm2ruoG1ULpRnFu6
9KtCllBnzxX5jY3K4EdtCZUNEQlvPU7+CDQMsqT0Lh1BDI/qR4QNf1alYXtHMkce
j/kCw5yZpKQ1Cd1GTuSzQzxz60xgvTV4OYK4KX+01aKO83Wtl4LQ1//Mf4vmMgso
qKp7MnRDwoXJBf+pJnZCpEDcegv/lCItDWNaJ/9lrZgCISBRhsj2/jSgbju9uqHV
duT9UeTBGTrtuk7CB8YFlVc2ajlCl25fPV2aqsRRBdhz2LG1oTQ2/5ebfPN/WN3Z
ZbypVuo1xPB4FFr2rBTJpXgiXruk5kR4t8NnpUj/ELL0uFd9KYV2WeMLNKHeBTF2
wspch/sbRNgPQFxsOjmd0j0E/RXPgEt3Fux/t/lfTvs/OXE3p3mgtrPPRmFVnd6X
heMt2SYCv5zHdzZbttbbKm0iyQBnJEHbRxp2A9EMQt08GxKRbSu953eiFN7342Ci
2+T3UlgfdnI0kAHYf39N4pRh0A+OUoRwNKDQzzP73hz5CsOfxqsumJY7aI031Gxq
IOZ1ZB6hY+7ihJ3mpda8O9wgMd0Cu7u0j6dbFP/NiyKrSIjpCN7Qt0pWGOLAKOCZ
NmvV9gimy76mI3TfXe1OFjAg9Hw4X7vfeUFZlRJUtPDcn3kn2DpECscvVoaV/7SG
r5qLSjRav5Ko6Fxcm3y7tN/D4l0RmBdQRndeoArXMBJfGDY81TDIIjMMqtL2cB5z
umQTNGTdr8cyfvOVUHA7Krmf9NSzVBVxu4J5TD1ij70UgChxYXyjzaVi/CztMCo/
ENSJ/Nz1L9YNwPQYIqoQR1bqdEkjmCGBgPhcokMSJGqD7PcMeKn8MpnEpd1O0G5I
NZSxUSTFFAqFOMYzvAoeHSYPRzQvPjYl0GXEXMa9rp2dhmq3Ne9hiK/nhSqSO4jf
2vELF+ByYzUdxkQwmlyeAKpDNXjklU51DDUAWtzPlMqk5i9dALFYLDg/XLXOggOD
K1tK5Hr1N/nlJgGWjao4XVJ6K9Ky2NouQfEUvqIFGzHh+YwgHe93PB/AvwqCYJGR
tu95PNyFDuA8ay07Y6pJehBEHQqTjcUgllzw+eQ0aDPSMb3A+cZM+etMl3mbbFIy
Bcilrsv+uQsA1mWcbDhAOv+N9SSEVy0ugn2vC3y3hFqCijAJoiNk+x0YY9OiGOZv
tSGj3Jmg7KRN7FmAtB+0CU1l4+5CdkKDZLq86z6Jl10H4aLaawxcOX0K8T9plKaj
voaVoWAwU9hDZOD4jGmeqDKU2MTwzT2/UPv3Yi1odLcEJzoA2YV3pjizcooeK/nj
7AoInxImryArtUkAiWLLGAFkIUv051Wli6D7UBxO7yQ0o15AImhewe6pRvQRsf/9
aPP8lUjrZ6tmbmjpw3/qB4emkY7S7NBwW685uH4gzGbQ/BhKKcLeKzCJ5GT4ov7f
CO5f+aLFzCnaW8YvGDUnKpRk7APpyQp2flznbJ92uVuzcXWwUK2wHT+f2Sx5iVFj
eYuGw1CsI9R1o51OiMsW/mUznSrQOGxMea319COGdrl2Kb7GSk95BMDvFKVt91d5
NsrKokQ2JxAer+iEv/bNyPeDcAswHA4dnLkPMtSZ5YccysJLmalrsvioxlYG2rgd
zkr7R3rf4ztoDyCyz7chyGAxkxPCUtXT78ZeJ6FtRaNtSU42Q0EOZVqlfM1ujUrH
0q+P4UP0BhRqANClbAlluXrUcTX6X4mHdDIjbeEI6mooEqjC78frfUmvIZzgITY8
Q5pAImUsHE5Z0lQDHHNSaG3mP7jpmkY3oDAjGlTNF84WXX44CQY93MPcvrct7kMT
Dy4Wg7somo4zFWcIO2086iRNpovp9BBc4uHizL52J7InBwRRifqdw4+sumNbkhs4
CN9Ex4WYft+KzxZbAp0ATbP8DFrRNLW48u1pBuclzMp47x9QI7zdKw0D6WeINfKm
DLTjE+6axhTsarzBRKsH6G6WXYjxWkFHUdjdFkgOzKC7gXAmjtLuBi16Zs4FPpoh
vOxujrLAJZyU25+pvXolRspMp7Wl6z+eTmCjodm1VIpkJH2sA1nKHQKke7V1mMGS
jbuTZbMfRElhsCRC3X80a+J/RpgdOWg28VDM42Rd2FOSmMqitbTO1jbR/s5slLVW
ThCp4/NArt4C4XokqR18kv8eaasDHHXmwhX4MxCYqmirRGHdcsjOK3yn39OvbB1e
QrYqMPfqwUU7cMhTeqURzHS9OnMWsCQP7ZwkHuuFiSw90JB8pBoLecbzXUWhOti2
MqHq/FiuMO90BjW5oubMcbmt83vX62mlQQRSZYlM3Ajc+Cw/THpujjsSnyr24pzn
uTy93fRthIdcrNKOGq6r6KYo9dBC+IrmWJvm+NEfFJgYzCJX1VZXtDTjSHo99xVf
hxHCoqK7Xi4yBrD9tVJiHIqbAjuZi470caNOYUQar7IarhQLouDRjIjuCj+da0fR
eU64F4xJ1tA0ijkSY1dQHbrYVbaryKw5dwIKqlXJXu2VtoIztr6dKtDOn1mpHjfz
9uYUcKv90vfmW+2rnrteg6ucfs4rS17zit/3IEdxDArXhAMgzeYlkaRnEc3L0iZ1
r7HNwUZu9l3sTClhMqaRGV1F0GxIr91oRW2SfV2/O8T8+haUBWBHnwP2QfoAKGhM
sIY4et2ik2HNveTsEvDKx3gRHlIiVGuIDDfJadch40AtQ9N7zPpa1ZN0svLTm69p
AJVwAc4RA/mUoYB4F5SnBlxYk7PGXzJXfgNxD0w8RXs6R0tIhlMo7jow1SUZEqX8
iyzA7IscVRjiL5lNry3vmF3HvfxKwa6hZFxm0Yv91yRqk37BdHzhpl65G3f/fOBe
/apz/L3P2YqccBZdikM6Aul2iLm6Z2ZdVCx0Rlms2IOHkF1lh/S1wa5lI7yGnR5x
jDuNKb8lBwcLyH6s+G3HDPqY4GQcPWDOrTMde08xJ1OfzbJBG9e0S6lx57ETtAZh
PJvVfr9oAvt1CiCPvlsZQWyyeo72B0FiiGqVWn9Z0m6g/r0/AfkO0QAD1fTsYa0s
5wW1WF3GmKg7i9blErrpalivAZ7A9FGFqwvp9JjLhCv5JUMC0vDfWzk4EE8dgp2V
kaVaCdNVEP9+Aowujcpvk6jCvanu2/KTrKqj2/2k1sfbAbyaRXik3OJNzPP165h0
yuIlGeVLwlpQYZka7AClARdhCZLe104GHunkE4cSoiUhPxl1jhryd28U0PSXRQ7f
rxw8/Ni8jUVjaoG4SnOzfGy1FyP3loqHzZirrtTc9vWCQMJS63U9WBW0ZEGBXbRr
5DTfkNdr4UA28tZfuUh/h+UbzdmheIr8sSOEgUcxeU+nDI735jJSxNA/3saEodge
tl1nCJHZIpxNgTaPyOjRu0C5eelPYTx/NqfJ/rKL3FlcY55ThoJ68RlKtcd5mhON
Nn4Fq3FgbLrzqOElCWiZU/IcTjNwhaXqDElLBXxXBlZHApiIvDO5cYz6eZ0NQdTa
CzCaBbj2TJQoQM55Z5PqzI8V0IlwC1CO/p9dh4F6QpZDg4Ow6NFD8xbDVVNWDWuZ
stCM4jDWgyBaMDLf9QllmsvCuGnzF4SjhxEzkUEL70yU0mNi+fd2PzRATZwvBiKF
MPkEBjZPvaZxLi+3OMGubaO43KkBedAZz13j2zsJ5RK+B0Ro2AeESkHIAQ8+ey3L
y+bDNU+bJPd4vU+b6WPTqI4KQhFz9KIdVI2BnqdMCLoyfMMXMHlU5USq6MoYMpvP
lCL0BSW66ZI3bM02nXmDCNBApnYYqFv3QwTI275BvetYanz6pUy5hZvC5MH1EGhx
naMxgCjzkC21skolANxqB2ajgOxEyenEe0P0umWKxx4ruXlQrw2HF1+8ho3hz0rq
6PifRL7K6q4L0Cj8qrAtrjvgepND4KBWQ3ICQR4k/zaOsG832BUmhkuKkytK+03o
tYJBwiJrsgsE3dFnJY3R5B5KF2EKdA+xq5pA1poHeH1pqXWD+8IkCj2/dUUerwnS
DZDmBXK//8VSL1L0t3lfJ7uT0QECM9q7RMrJRoxmFSEkjeiRVEF1klEYQf+21aP+
7fioKlniKi86CLEtTdJP/eZbbmKWBazvo7f47g7oYYYfrr6N6EXH4WsmBemLPcqA
f75rJ207PntU1sYcGMr154e7xpbRAnVAMlTmWvZjoCblGlRUixOX6qStgO0SvpMV
FiTcjaQPB9jXzWjAj2xHnfHS6eV6pEAWhc3TAFbhNV8tPlpD+eQC4iBTruum2PQ5
9pb0wBKvAfPLnTiJ1tMNkWwdkE2N1kOMt9ob39DkKQB48ctfMV64W/sXYfCYrlT7
wwEWt3WhF0BNwm7cKC0VPlMMjZk+FkxlOMnrqy97BKyt54RAOQN+/5pq7+qoOgmH
rYo0cmpCWzXny808/eyqKgvBQOyfF8Gre1RbwRq0pGvy0ZjTC08vj2pvyNNPsbXb
preytZplTRJzrROJH7uurjsvgxOl2vvg7HHN6ckAeMLTGxqjrA3p5cdNo79Qr/Xn
ekCbxWRqXPnpobY9aZTrSN2eW3R3JW1REA/eN4nAygmjduNtLDzfWdtcwcVQvD6M
H/Kp8QNPiyUzSJTJ4liQnDRucs7bbguR3OJyg/1kY35xSO3QWaxEwav5aJTlGvZH
9EXSfyaYiklUQ4hlsZjE6zJKkIlki6fwvlKvAiKbicETMiZA4xiuQQ81+zj++cyw
li6Oz3RERwZitdItMMH/ZhCp9HzucFVKXhUADeI5oHrwFqMFaS76PPjHiurrGTcc
I6pO9jGt0xn3fonN9PfGEC6JDcm5DOMs+XTA3mEVRug=
`pragma protect end_protected

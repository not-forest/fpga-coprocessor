// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
QA4P5qYVBAaYAtZhkw5bQhWyiTBh3aXdmiunVDheV2otZcnHLl+KKN84CTfXQJki
euvwPAPVN2tnOv0pu3ZfT2PNRW7t/QiB8qs7Ni+fnE7sHi8SCZ8yz1JL7mKo06qT
FRqOCxwjJzcF1IqtZOCo3yldCozByXpl1y3yE7x4cIo=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 7568 )
`pragma protect data_block
EyCFmbqGqnZrARxEM6FleUeEavqziwXjc66Fej3MzwJ6z5itmrdG7oVs9PknsHhR
pK5KQOaovI5pUoHAIy5GZX9krLnLY/BoPzJMB90fZKTq6b34nSAfUK4U9vBngJv1
ZHPEYdKdVYkESE67aLr9ERIde/RfcykMiLyec5rqhCqezn8KgmEDGJXv7Oq7gT14
FFSYnQYAXewsLTu+PpNWUEw8zTAmyn3rG3ZVzlXgThOQ4sMy6U9xnQ98262IR77y
WPtQrwyN8bhtUWMZf/Um2uVqXQwJCt1+hJQzr54SbQ7IjBLobFISeZ+jZKKC2yTL
4lEp03C88pXZMchunoKlxTgJqga9gmXg6jUAGkuA2VcqWE6CyDfAD7Ypnp+Pu2vH
O4nP709OB278NLdikHxAHN4HffNeG+86FFZl1Uinfj5607rxcghWBVt6ne55UnMC
FCpkqVFLnx+Ljq3c34+EQvsZFsvafxGGpFU9nXedwY2cu03jH2wwuCWyVmiSQ+UG
aVYuOCLHjmzhJIUiGF5Gx2JPDn5qXLhG7ADcOVVsaPFmw22DoMSxll+pIho0sV3v
qq06pY4Y5j59cpeZGuMNkGaiCkWavTHU+0TXFXww7aYsW1h/AGZTu0IG7ihBJ3tG
G+uKhkKEpVdIz3K9Iqdvfz4rSis+9y5alKqZvrX0whLiYJvjG94bOW5YKe88IqjY
LNtPGe4+BBXSShsEDgp4K2z7PK0FZW52FkgJi+NOFdjG+3uX6/1DVRWeoHxO5qHt
d1jVHJilNYR4x2knzkQnCP+qX1ak/GKEdibXjYU0x0C0hFwSNKn452INunmBEru3
dnSCie8h9qUbMl3g40CKLMg9XNztoWSzwo/lW17OXLo3XtBqy3R+4/Fzq9+mlkg5
LszJQxwef03eLgLnoFcNqED/XQ9FABbQG3JIdV84ptN4o8Bf2pI/SHE1+CgAURpe
RrqFBIyoScTydpPifjmBBIDy+C34t61OSssPUAyjp6HZDsBMjq4pmtZ0lhI6Fa67
br+gM0bBup50Y400wKwkSCFCt46dpSuhl1P9IXfuuKnBr7uDorBNV2xhxWpXEWDf
hJtZvRLZiOSkYL8prQHu+BkvAlrO5SRMEIlTo5j5yM+HW1E9AwKsllcPdnaKInC6
uumnNxgW/VNyng8wVE5kIPPgsOeKjf1bTu9j+VojX0mfmh/xOkRr+gyilDFgwJF8
dRR1cB+8/nZvjIggkHhmWgTdBsI7hVFA5C7P6PbAtHK68fYF5qwh6PrMQX8FM722
cJVRkCdWZLQYkVBQkQy8PsJLmlxrWvSRrzDGjxOa2NMo4ioNzO1zjt3jC66kqJ7k
k98RY1NyUtnlZRLwOD+cTsLSGYlAf8DoAFX5N9s0wS6DoSc4rUYmL1TB4v3dZkT7
9iJ6qFb5mTKkm7H35jNIjZOVPZ6ZMJl9mJy310xBNbZKUysP+a8lg0197irdWDll
xk0i++n+4gBeR9tYJ1XBiNe+Buw8/N3+I+/Yr6v8G6LgbqIJwmf0JXmzLFyim8BT
dCaM/AcLg0ZIx1+2iqnWY0puLgE7i3fdXChg2CgEWxgz3ph0WV6Z/bvi2Ji5+DdS
CGi8X74KlHw5aYGlvL57eouiDyDG0jqbkLgsyFegnTdJLgKbHZY53swk9InQEuJL
WLzJ0rjvGgwIpG1aRDYggxmCpuE7HSqX03SXeOht6DseuABqCHs3t1iK3pQ3XZl9
7ilf9lJLLTo7r+AzTGFV65vloqOnI2xCJVDPN/PG6rRM0m8wXE3puQJFKXMoKKv1
pV3V8I7cvFeazk/mwT6ihaFX/5h65kKbDJwuuIulClFA13a7A+r5y8YlLj/2zzsX
IJxXBqf0DCsAt5n4ZRoYilHxp0MYKyjgcCb0l035JyTsqJb3JdGDmALeqpjoNxvb
zpaMlyARmouMv9eiYnCS6W7RvXFMwk6dpbYlET3QNq5D/krvZJcsFM1N+ogTRXL5
GSx7axNwJrikOsG+BmMi9olfVl5/iuyuE97qpl9SQxl8ddh3IVjzg7UYZHApFBl8
TqJJDGsiALkChxZSpB9C03dWLpsaHPDX5pBw7KqwRryJMWUrFck6+vkD5cOGERnx
tQi3o9XeMTSJlASGf7aaCbHjJn+jZQeZfKQQWoYDIz1sWS+kegUAxSpvNjrkPxo/
wObvABDy9t7B4cPU4xy8H4yCYJeDwD1lyTQSXNX3gXHQzGzETmjozWC+afNCaa4r
RuKQIcQrElTeTLAOqN9+2n9odGKRyrFKTPj9txnF6oCDzYSbh3+qLYGV3BOJzZX1
N6LoP+/2QRxOauP87/0aWF952X3CS29aJhhKNJIwM71tFcdxBCo0JFp1/hXc82oc
+it7/8zLV3SI41C9ywbWwNdU1Fel8+ehpgv4fJO9hZgmhKvnYjT18n/3ekml+kyb
26q/5BdXb7Pcq5VvTNxvq2fwySn/ot+CXIXBC/S3emrA9DgSE9hg4gVH/askfOaA
S822vDeCTUbdmTzzltTvRGzz4xDsy/JIhe1nI5PwO6TxBX+tovyYJBWg1V49e0d9
TV3i28W4A9SEYsGw9kHtiyFs8L7TzjSkV/ZA7xFONhqlQo16rrckTHz6u7pfohai
hAdQ//31CvlKJtwKB+eKNXXi0V/yvNZdOrpxFc3SPkj9W7NF0eqK43+TEoJX76ye
fHz/BZsgPvdPgT1xeBghhQb2NJTg7GTN9zkJ/DlVRvCZduQ6qyNjUCLC1K9hgZSO
NSUEkYeDPNG1VaSPm/kr46u9JVeTW3Gagjk2t4i0slp1wDQyN6F7HT+D+tUx3aSJ
cArsGnpEKUJJFeES7Zaw5nZYpW8A/7/eiw7fxl+4uc1bFnecMyX0Ic/XV+Iihg95
XtQH95fJNdddoDcKztOard9tVnew+EXG6gYFj8TrF+LNo8TwiHJSJW4xoRBD+St3
ByPd81iORTJpYaizLyp3mfqL+9YcT3AvTNOx6WnOJdHuSwpSV7FsdftO2Ezh7Fe7
vroBt9ZzayOkHXHXXGHauBciR/BAwJHGrdVFnFI56SKBYl8jlmfjbtGugZMdzO2H
Bjsmh0LEh35dytCATgEzp5JHl3eneLDdu9laq+sy6aiMwGRA5+aRHz3xyZLe/pDH
5zj4aOnIvPaB0dE/dFTk7n8WPbaI7WyvdQOz3BymGDehfACkfhB8lxz3y2H0hlX1
ncHbYKfA/4VyftPCNgt27KaJRsSRXkyOtH0hhZpr8XLmrMPPRNiG8ceHbEjKWtSJ
khYAxY9ZaHUX/AlrXznAS4BkOzNGRxdr5rDPCPKCY8/U+f6ww91AL7K1CDdJMJCk
2l3BNMrh2int1/7/it4x4hJpnlTJ9xJJjNPYsWWU2+A94NgQMsgYKPi0zHfjlrji
ooTTOJVtSU/xSNQ72w6TOwNah1KkU0lmCYuJ+Lyw8VTNIHxmenmABSsvpw8rAKGG
z7i+hazuKngvhEkN1mcr+zW9WZA6qA0nyyQ9+LCvoASGHN+l0nNtvTERht3u06+z
6h3hwuT1NRhEG8gOW1ssg7W2as2xIy91hTRLiJU5xt4USEZg8Vm5ZALSPUCvyaPi
+/7VKyEf6Ut09kYFceoXhhsPwN+Esk3aJfKdzIL1cuwyKWeXFQIBkFidZ5Xts79G
mTp76vQwC0t5ld96St3m0HQxXdl6NNOALyT2FIpSxF65cpXMd2/vdj+0OplCBVvL
TPEIjevGhlsL/wNPPPm08RwLMUDmvW7xCmf6a+gFWPv/vvX2BJ0R9QMMWfwJiyUY
enE2mK7WNw+GMXCzPuZh1Ztsm++RPgLpx1UnpuGn5vxdz3aFtrsQwhfa65cSGDdS
d0POL4jJnJLRAfmGP0Q0WuNJzcnHNYjXlpjgZC2c9KEU/CGKECKc98rLjdl6D/k9
3xQiXDrtxcguOGsOxP+xrXQg9nA5vjLTtOjA8GC6OGKxq+gXjXD4intUA/DowKEd
M14kjci7huz3IFrmFxcDAmWKyddVZH/2EzglrElQccSn9TRaGOmae9uRFWD5mZWj
7liLqTwvHFe3Fv52bMbK9vjF8m3t/dlU6CrsRBnSUmLZ1yOTyCCtHFSdyM3QZwa7
dXk714f2QMQPz/WCqgaXi5LJvOS9YJBUmKdEn7qFP+nXQ+FePzXbO7eo6xkEbQbw
42u09ZkZWsvOc/Ip1l/EHFe9pPlDj7FZk83zB/ESonRa6WMffesyFGaNP/Dz0sCC
N4kVSXhnERBNYHjgOA2rst5OWe+2yd5lxXy9O+/EkIqG1TMCwmSAvZG748pq/EqS
cKPtFX0ZRNKqJ9Qo37DmdVD60AfySkuCnziLheSxw3gI4NwhMctbzZ2QPNH4bGN2
tRuNLzxudLtHMCNq42lvJhcPPjLu99MQy+SLHcoFdbXKMxfn8PZ2x3SE6Dmo3jB2
iyHfLPc3sJ9O1O62iyubQytod0c2BrLFdtqZuRsXxhiJXgjsLPE01WGDcKXfTM/H
bFYs4U2s/jqXS/fT1o6dGyoi6BiJowOGhVQbSOvu4+IBYguKHjrh7jPTxnee4yAl
FIrx4zI/zZ7SNdqaWeoBGRyZbMnhDarPbXvT038X7GTSKm8wVBwyQt+niio+k/KW
rSkw90Im8uBxfQbe0EI4bS9cqLQiLCkUpb5oH7ZUCQljHot5MDSkHrMiR/29M0Xh
jvRJoruFn3l+OTzUQTWD425KpiMZBFRCQex8sJSzjhup0dpBkN9T1xeI8wXHl7n0
WXTY5rQvLiVFJBpMKWqDgw60B1bDBhIme7v/KSiq3e3TDR/fpl5uLIZAb8yPAVyS
4l1o+mPg/GjveH/92yLTju47fNOolgAb7Vb96eaUGVvQO7xAlIi00Lsc2enKIPB0
RzBfykb1xrCNmAjBvOu36YdsQIDN7nz3gJkmbn0vwkXMW+Of1cCcpwT68SyApc1R
AyUlsPCF7HGdGkmyVwm8ft0o1l2gPHJRk+ik1AAW/exzzqDRE3cPQDX0AS1xK/Ty
AvJy5opwoDVqWz2l1su8COgK5ikSytLRdD079rTpGJ5w0sI7MwW9ChsQ9PxIuYno
keo4j56KiP7RtxY3id9WvuiEk+yVmYJtcf+eoJtfwadmt/QhwdBXFxF0gssoISCJ
uZYKYsbDjPlSTS+1iiQBqoBoiM8K275IyRCBAyGkCfP/gwlfU1xnd65RJ1HPzjHP
Txof83soRLmL7G/HVzkEUFJ2CzE+Xvx0ueIYeEpZfrWe+BbzvZ8cHD1j9evXDsu1
89yXo8ExB/AxRRR3sBmyFy6OrNqjSAqxB5aqr+EflkexsflGnh6y/vRyhDBoxOqb
WnXkkaaVTesb3Sr/JtcBZrz5pZamDGGvdgmW8Z0bUPFHuhm7OG5TLdHSfxk5Z06J
VXEQYKYiqz5dmOySNGv+Xupfl78Gui+k/jb1Jpm1z5KVoFSfCk1au8WOBTp6emk8
Zjm9byhcaUbCNWGg+9UGtQ7JqpPO67jK1hbgVn/afT264u6UO/OO5pJkS8qD1rww
OnDVhCHj4AptjEo2J7iZCaQnHuoUEZcsVoJ5NX0pJeoJ8KAsOZMMdPu/fAO4Rc42
tANhRpUv7ZtOdyl+uT8uX7NgTmYeULahOr8kvrdvR2BUWsYZwuu5MYG8XXZWaFGT
zQN+RHDou8BaMht1RPPyMC9Cv5VegjvOpRC8uC3Gg/I6JNeXpk1PaGecNTxkVZ8b
NakEvFwqEqdpBCF1L1iTQaEcvYtTdQLkdwwZBuBtpfvxk7SfDnOLH+BbedgmxnVx
PqlRzA2jPPunPzSMXMrScwFQtYSXQauh4yb146X3VSnuXuCV2Y53iTFfzFj/BIhX
B48nuBHuceExYWZ9YMMSMwu2607gO2A3WUg1jS8E9obp0g1OmDhoF7zQcDRfgTtX
7wGfhQ4kXskGZhKPVC/RTbtoCR6IEE6k4igcHw7qgOWomwv1MloDWLXog1w1BQ4m
5tFe7b1vhxsE2+xkZBCgPq65h4IBWYH7+QZDV/vSzQ9x5qu5xoUz+Vf63Kso1hPy
UgeSbPKB6L+qpmv7cgbDCq6jNOpiP1zNa8stmZ5FiXLLbG8ShvF8eXYWoX7FbvR+
KibDbaRBIxu57XIf5aXkibqApNm2gDH/S54Vj5b1TrDPWi+qv0zJrbAfe21zFwdt
qGMFtkk9PNfJ1G3Oy4LE1q5brreAH/hnFLRSvaUtW4i06cvWtu0xy5iEqEu97LN6
aPmwc7Dm9WIN+JR07ZsPrpUOcfY7c/CmYZsetNAlF5/uZ9/2iuEhAWdY01lK6b0K
2905hpVNAwabrS35C11r6ISHFlXBc0WSSfKsJxXXzWGspCKET+6kNs3Ow82fVbSI
4YDo+BCu61gRbO1OlsIzXZ2mDiKLcXUAS7cNoexxkegiAWAS4fDYSb2E3wiLSLBj
a1lZWT4WY2DsOQBPFcfKBQIPqGp5pSCeVmfUksRR0p2zkbg72EUgJ1DxLGO2ueDn
OEZohd0YlcOasxmBWtrCJxZmSq2QqzBleWuMeEFoSERUjHG0Xlf3+6a4ROlF7Ozm
/d0fU0iOAEV+ULxVje/pJoqIuIWI26Xfonm6QgNudzbws9JP2K6NBC+JPvxDZPmJ
y3R/ZRaJ4KzFBZ8KwO+cFWXDKyPSxv9yVoCew6csuPyVwNd/43eburUBUYV5sQYI
XBB7/PPeenpzekELFlJSD3FSu2bjBUlX5zw5JOEc8c8XxufOCaDkZ9vjZ9bLqFFO
dBmTRcIs36i2ju7Lf30IN9wkxcVglh+UCnxSiHucS16o6OqSsUZa2bsO6uJekTwr
Msx9IN2pwYG+qWd9uFi/l4MoAbU6sMFINR/9pz9aDF4CT4tkvucW0XziQ0ja1Gu4
XwdGQmJnbI9JPQyk+8KJgV9nNRZFoqAhDUIsK/hrVbk8i5Ng2T86PWWJbIyrnxwf
0VdUFzDrkhbzyEBcdZQ2sshoIKiZY3k9K34kYgZHR50pn1GFdyeGPTawhiqOB7zX
9148VOZ6E/NUpNoaUTo4y7mcXiRpmHDgdd6as6HkA2EloAg6VPQn6qKQR8ZCBbeX
JJZi7Ehnm3vyANQX+qGRYYDmqXOAdNZ+/oKn8U+LYWN6g5ghW3ydJ5lexMxq6wKt
cyDGNLo81YNR0CYG/WNB8HNIvbmcFf6Q2WFzSW7G8FM0uf5Xh0z1+nffhWef87/Q
ffdhEgThcb1fbjS6/guKrOZ+4LTvthh8IOP5OZdnmVMB2woudnP6ax3C6VlVtse0
9wK1lM5RT+Vru5y5UFtcgQTtHFNaAR8CFstiAPQ+gA7T3+vn5QjLxgZQV2qcQUhp
tV1L0zt6CUDwSUishhkfzC+m7iuIOb0F1tDH3hQujHkEO9KRi3GIx/tOAO1Uglpn
sBe8Q4UQh/NuTwlVHb2FDV7hMGS90cJgSMfjnbHaS8pAB49XoG/smcv8zshJ1sRM
f3nNV7tcIVCxbyvyxI3LrqVwY6d03FVqEKTs0gbR6rODY6EszpYUpc5vOyvlB5EP
ZrSsWtG1JMF3SPuag4p+QcEhTJdeZCWc7dv2ylk4oQQjpMO3Rn1VPGHLDViOabaX
WDOBjXut5WGWr2OnSRthS/M4DclkqT5l9A/1OhiiTr014loZXa3/bc3tphtj8/7U
v8YNuaSgV9ui+6Fgcqg7LBSiEBHcolmC3I3F4ELIz8Oih26VUVk8NJj/AY7W/uYu
oOk2Yq9REAzO9HcNVXMDOeS210RrxsyT4c4JwX7u87LwZNAnzo2Zs0JFy5AcfO/w
EdbV+GiBiu9V7ZC3PKQrxmBTj6ZgqWzvz+8pL8eaRpXfFhE/SDVmYkvKQCCZjAxJ
O26i34TMJ5zKkKkO+i/OJDBHVxlASDUp6VCvXUbJGCAQ0DnfXmS9cniDugx2tpIN
stsX1AvNRoCN74oV82ELbCQG/Izs/mBCyEzr7+eeHGHpyVndSdXlHe58PQ7w1fXP
xV5GAm6RFkMU0xwBP4Ssk83jneNNnKJfm3mLhtkeeUtKOqQ+9ZhFnk1us+hwiMHf
KQ/S34B259jXmrBlWAlf3eL9ZzlqbyRQFRRLggKUATcA3LXLcBlXpMdK9zrLeyvo
qdKo6egIiSFYq/1jJYFKBY/MKXkqldIvJ4QuAhomNTrJ+dbw5XBJqyuATKcmHRzf
/jU6ORkhA/Qq0EgzeCsxjnrnSE2iEbfdsWnW8661+w96Bz6XFk6OGGAgagRIMUzZ
hSz+e7YXhua8iOQ8fp3c4CCUpzg5pCQAmTkXsfhbuf1U8YLidjzLlG1grLK4Tzma
138Voy0LhR98kROOcf7FBTodDZUDYghk2pSu/zHN8dFoGXE7ywfYO7ZuWbRo4dzY
xtArIcYDpIafvuejf5DIulrHAJnZCyUcp/chTYjiz8x9lf5v4fSgv54zAy5GFI6B
EtnaOg28aUQDHgBw1rOo8MZijmUCnB9T2N006k/KNfR1m6+w76CNREPMn/2GTzME
NXVqSyHq7FzT1I4kGg6T96+tN0ypgI51MpxvTtWNoRNlfB5I+EGL1A981DSnRKEV
x63eRA8NMra9HTsLOTdq9WVJG2p3j0dm9PCsIQyvOmAV5QkBAHljkLRYQ9JYpKMG
BAN8qWcUy4LiTnseEw1n2cX0Dm62yRYqtphBhF0/faE7q3KsPT6yd0Qu7U29PTHI
TacSnCDWsTjnkOkDVQFH7/URoIvPH8XAut/92UvbVi+/jzCeQJ8Vx1HdWHoHz6De
na9QMTxTUQibC2/3AKmDFgjIIz05A7n3zU46ENsfdKRunW2/8m+qjTzPuZveq7Yi
Of6uVilyd6XIn+c4Fd6vyXYBGpDeRD8vYdSZiTt2ckVIQRZmkTNLuNJAx2kfrdIU
/yW+nfK3/mHsQ5YCdCVT6WeB+mFUODD+Pj55X4gh+FpTBf8/B4BIE+iCkPp1JLVC
K/gMY3nSgyJDw0eaQL8Vr873RGnOrp5CKXgd7bfKUJr2qHVur4cGOLSQ3T5Y7Eah
H6qy1vA5WDCr2tynV2nL+PH5YmPo0SpAaR0AqTe2xsC12xK5i5IU7apEDToVniBV
DMJw0AI+048sM10Tb+so7jCbL65ahCzZ75lQTQbZduWBAiWQckpcyFSLbyD2tC4v
7/w1v5y2RyZx2b7802ZCvnDc6G/WLxJwygSDxmwf8p2GhoG5/BRt/HQGoT0hvbfe
6SKi96YyIsFNRzLGSIHcamB0j83uKKY8guTlVAjovtRkZCf047Fy7BjhOhzbhYTf
JWxN1vhGVPIgr0DsaZ9Pt1JrO86c31JM/A+cgPzIpyfbFcP6nrvOK3YsBWwJwaC6
FvN612lFqCJOhElipaBuZcQ+Ah2QFwFKeXJ22MtL0f7MhdugBUAVtvsayTq7mI7l
kEe8i9qn92CNsIggzf5WwBPI5WTaG34/LC3cO44KIVv7UyRgsddK25/dUoUtWCcW
Fl+laPpryxz08fi3MkcG6suCxNYNJHrNcjhfsKA8xHzvZ2xyuzrSKpDSIy3rMJE6
ZXrSF45NxuNlt+cM2+42zMjZcaawRCXmd8xTLqz0DQOvzKGw8/ghOOZVCwSDpI0/
j2QU4QyvjmLJcsO1POb7XlvwKCFGgfZv7s/31b9rxMOzWfEofaxTyRef4fE3aOMV
0xWF7BFl1eRq8ICKIP4GN3OIeINv5PTA2hZtTcVZJWIQx67Vn8BdBIsf/1GVw1jY
6jIUehzmMMb/s+KxW4JQxwoMDqbSN5viVU0rOMaKHqkQ/Y9GFY5cAAbXJ4vDbNk9
edyrzn15r2hnOaTCHGS2NaRJlHWj8v9uKp3lCFR+Za4GOtpQgzp5CN4IVXb9qXDV
FD8/1YOU7o6Pb0fX17JCx+3JIWASFxh/E9B3F9nTLtUo90acXUI09vd+TIrSd+df
f2DkCmLpzX1zCAGUDdN3VeMs+IBZRoQVnlQqMu2f1pojC9ddx6036UM7nVUoyPel
sQfg6Yq/Vu/ebxAMTNNFiTm3hV6eoyCiJUPoJ6VtiEUY9gfuy7+J95b+BYOIV0wn
Nipdu4rzJ6vh3MkQNwNNJN24Z3t47Cf6NjjViloNBZJUzFjOzi/KgO7hhB4yK78H
t5LdXxkShUYmQHrmKPhm22J6yWIN0cTsGvlL3IqnswQ=

`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
YWXGwYe9sCunY2JYC/pfrKGGbJZSmDLs8cWcRVtYJV2t8eZoaxSiVoXjLLh9NYsNfrMP1D5EYT84
ZyCSi3fE4rKeEG3eSkyA2K0znEfbvzxz1H7eWYTp5ka62wWh3AFWq7/3w9ui6v/xQdUscpjWN0Aw
ERMbEGjcXvyHf3XYHeIiP/EasmUOULiL3zXTEFHOwl3Ot3iS/QzDfWiZKMutrT/17XGhB17bMyXD
Uk13WPyoUgVAVS5TGo4QTxu72ZKZ11AT5gkt0U0QEsBM6JTft+sRAXLi6FnNhQFcW/rCOTTGMfpW
/sOSggckQEG2a5wDiYJB7WEJB5WnWc9Cz45mGg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5440)
Xou27K/OoUHgPwqYTvyMndC2W/bHHXCZly9FDByCplTq/rWzm7V6qF+8av3ymWtF1suooBXfmY9s
+xUStzE4NbmaQguo50qWpOddtMG21gG9G2rQHPlH8PWYulE+zCzu0IK6154QfxuktJfuVSQZQOTY
u8g/TRyE7nFEzfnh9/rAI9igioa+FdhhQTXAxVtFO+b06BYxQs3a5XVQdl8dhqSWQ4BtZW0xeb7s
PLdpbDgLbauot+ZFr2LcQhe6ukje4VzhccAcChzeoxZBb/GTx7/lHpm4NEz0nOwjY2gQ8wqi4/gK
E5FXAld+7k0hxwz0h/L4aanwWAyeq40FAXq+R9CjK+80kNkGUXWIDgCcU2empTegxrmdgZkReisq
9QoPT58kcUbMsj+OiuQvRk29kOUtx1ZnWds99hx0ifzbr1SlkgH+91OQ8oTlFYPNdlhryMvvdTaU
qcuNOMGLFNuHcr4OONzQLuf+hOUXoxZ04hP4KGYgz2HaJPOcAyjAks4og41gHLvY8+1LIqVdnfPV
nt7Fkqx/iG6IeP1KVlVXTCR3nlpXPcFAubQN3+WgqJZJup+bTmlQGGKOQeTEx1P1jxqUPm13+25F
ECZUNclDYbKxX7lsb0dFF5vS0bHJ9mYDHWrXDheYKMiVobAK0Pa/N+rwcOF1HQlFL8zh9s3TkZjp
IERQCcEclzisI+NtBv218FJnMrtrbYiuDTRSoIloo+K+vgd/qOTjwtm1qo14NEA58d91KkmcN6ba
zt2x7Fo86EochWdf1XvN7ym/7BdwYI1jNaB4O6PVY9qVH36SOb5W9Tn523ZL2qbYlFteeJO+XUHc
2F3go0+kQ9Mi7qjUyOEtNzgyZ48EMT5acgk2BSh9mykTH2qahXkO1mAD0SFTqWJ5PVWZtKGipkgn
EMdTr1mfDFypvT3atFs9PudBZXzgiOYiGXSmZs7c2Rk8XHvjQ3pNBQnkrq9NaD+5MbIRvATG1xKP
gQVZ/K8W+zaTtmZjzIe2zz+K5jL0OVFxo94hcYSDF71R04ihUAGzVJBFiA1whfEnP+An1N1PcxoV
Z/7wHJR0X7x0K2UOw95Woo4yFdHWwXGotjiseT+w0IQ1eTncebtI6Ms4AUoeQ6A1QV5dw8isQumm
cUEamIxa3xpcb6s1Qb4VPcLUnp3x9QfjMrN+xb+kb5tjTcNw+gm0p71nHa4Ofnslxa1KTxsglFwA
sK+aeb9EDgLGTpRpazbkFit6Ziz1tLsUFpbhzed5xrzGQfbsWR8x/QcUrK/DsD3Mjyce3Ta8MabP
fzxmY3CZWSbP0MxiUiSA/LryWIH17AatiiorgITnJJTsBbPICOyVw9H+zm/3G6ZFAz8bUW2UOGMX
YOGT7+w0YzuXz68qs7M6LVppVQm3KT0HdNI04IJ4AHipOJpcskVNSwiqwErVVMjhX2kMqedXvqJZ
ttMmBYoCUiDc9U1Be2kiWh+BEv/ub4PU0NRnPEGBiHmViZnsp5ZvXlZBxHOawHGkiWZTjlqppudx
5ZsPu4uBkbJM+9mzIaJ+NCmYJlHRCDjkfzzANzmAp4peaaZFDn9+5kkkgNPglpTrgb2DEd67wcIj
idXZmY6s39IY9KKuPC2wB1votSqrjnUDB0lIHwEqWBpq4CcYgN1W2JXoT8yCAcBWSaoDZV4v1XA9
Cq1ZGJU3aNwu0NYUE7EqGcKckZ2EkozPONEGy5k5am/86INg4CfjF/zLoKoUtnPVHF5OwFyjENYW
Iw19dhhYAj2t9IAjHKZzEhJgG2V8DR5u8uHWbctLlCDC7/1MsMXwVh2vgZa3727yDyyTAPdOQ/Eq
8hOKaWYmOVfrD8PWqzgin/apBeK8iXWbeTsRD693bjm53FByq94a/Dw0owAFzxcTj4RWeEKD9TDg
T4gs5NHLfhcO6dlAAaNXPrFb3wCkqX3TUBS+ZpkUGSe4guhnnMK9TAOmRJinLN5S5c/XhEy9L1nV
E7CXI4ONVW/q0phCJN9mMxtwTyu9MmG6M9dg0L49ygHem1rLAmUzEDyuw10sjQsdXGayELk88ZR3
l+LrgYf2gBRRDI9l+qDJNL2Sc3ZkyFvWqcSKGwRONj3AtMG+CWZzx3ceyjf2YZ/1zP9cXyapKOSI
EJ3CEuNUWuL7ZF8A8RnuHIEmHw8jWesBhgxOudgNINFw6fx7ruIttpwJgQovlqk43C17+BEfKdoJ
iPYD9Fno/MGdlTW1R5n2JLujM6CwO0gDLHt08XUcrXx9EdiRGGYiBDSTM/Y8iSzUsySRvPU1+Yjc
1S1gkFmNGB1d6M5W0kGYkaPhDcUzdlCt+0HVVZTi2JQ5Y4PoVTlipWWGRiY8yEHB8w/Hs9fQDN/F
zEmrNomUQIkmW3xx1a9idMsWDLgIzBCiXwQnwgnsnGFSDrZydupad3uq6BAgJ5vvbawKo8yabjxf
tOVAn7/3Ktt7So0x0yCwL7H7o+1/l7Vt3j7iNH0riDzmsXZxMTgEcVnh7O9AOpbZ1QPWsFDSVsdD
oE7RYwVg1G3F8lY8hgkeik86a1GOfnC0QMGoHjgz488DKFmmTi5rFl0gy3UODmi0JnUd7L0bb61z
1054mfoDVJ0+j3kx2vc5Owo1U2MVDFiGqwPt84xaPEHUd1NaJFpGq91udtrCigfIOHmLxLzy0Hld
n3uKy0X8uEDHixIWCJ1IqeAhIZGzgNp8gKnxAPasG+nnS9NF4HWoCuTulEUcerXy+2jsTuTkBDb8
uEWkhQO4C1SHz03nPuTjQUU70VG6B+boQ7fgfRzPCMWHyaKgTosi8BkWcTZd0T44lf2ocpJuEKiE
H+052O0fzESrJ+4Ivl5JqmD7Wr5Ng76KzoAwCgjklUYarLUZdO+POkj+FBv2a80SjV4cj8Ap6CvA
uGNlKqeHn+LywvM8h7P83AXYJk1FhACX6R4SoaOhkk4U608RFpqUUJSzxA/wDjT1Dw3F2OuiTy/s
bDLLiN2iD2hjwqSLrBp6789rAmniQ+VP9yI40t3k0JAiKur/7e2Xf1DJDlNoD/fEA9d2Y0I8wvv2
IzQa8w9M9gmSluZ9BsW0Q2PUbDpV8gvpRSRzRo/90D8LkGOaTHpqAtDNyHhfiMJweDG0s8hEugVT
zE1IVxBUMo0A7Y6lX5AsFFsBKFCDD7v1w+Pqm7+19mbZ4tWF+hcyhI/HHX6WT5g5IuaWDzX74yez
yv17JFyPk6OnD5ZKQeKdPN32bz/ra7Wez3mvwEFe2ae6LqXDbYfw0n8FAIocR9l3aoU6WNYAeOaX
Gcov/XlrFY/Z+0qz0rCwkNln/VPt0FAcQMhpJabg9A5Z1Y1QZvTfP/GM/JL0IlihHRehQtcv9vG/
LIl5/ZcyfhII2NrI4tiU5l4A2+mMJHWF3mfP/NLwZBiK1xfgb6HyptkPARyS/oYYLkGmuAaBC8Hy
9vPCrX0OLa20m2cK3V6g26/VAU9fnS4MZugz3AgsczvUuCtHk+/gIu2BH2PNVy0XgBJ0UlJ7PbUx
QNJgEKEMD67TbsIUOY2BhVIQVPllJ1MbJxGaEIKt9RBMDdCW/rtsxX7xw5eamKhW+h/2as+60bkZ
7SLTxnQ3Kcpq/6JzVAu8XLYbhwxxo1IRv4d3cHKxqBGC3deTs3j/3QLhyFI3vGyvUivoh8MEpmju
p5oum+A7XWZsLt7Qrpinse9m/T4mRpdHRze6Du3qiuE2pyBgoSIZAA43O740XuFtH+aX2btz1aeW
gtKEj6/2A6iPUsp6eAjJUsCAtc/3N71Sqk7XSzEhIsskDFsM+Gu4WqzwYd6mp0Nd1WxLIUGNEI79
IMw79d775zy9+z0j+K3BDd/v5JLCFc2t3FgvH8O6ZRTfFA+kWZDGmY2+MlwuEaAgZk1arcN4nxAv
VUf9M595+GuVoYgtcrruXi+8djqMCncAEXoASaX5yQ159KmFd1Mauy46ZBa0lvXNAnWm8aaPutdv
ZjX1lEJKUD+6DmOVX48Looko025dyILVZcUqya8qQQf3cimONyywhIW+USo1GAhLE7lchLXxybXz
P9zUOqi/DrTH/9vcViba039b/uBcYa0ghdfPTOMkSwQTUMLsw2r3zEJNjim7FGAOuw/aANI8z3sq
/O8l43SdV994trVtKgXm7s9NdzwOkka9ceyg3zR0SW+I4qiQrB4Frckn0S4xdhAioMGmKN+TFRCh
pYZB3w9he+S2kaya12s/yYx6itoOlweY7ltYQznn1OuNL3jwkix0AhMwzZPh3yRuprAgXNhl/j49
MjP5d4X24sOK8uf5DUDQMg5wlVazjRn11XCpP9b6RnF0yNtHgJaq29IwZanQakYT9scwLFpOtxt/
rDfH0l7Wiy6z8mlLTpuUflyam4pO4jGDRJkYJdXPFbUaVsESWczCvgNd3qJhs4TsttIqHpc6z3Nm
BeqzovZgXoIbUZHqGsFMp7jMJ/sFsHxiQi4+n+4mvS0FThENzTfRLV9F65iF+Qb1Hmer2x0G3btQ
yKQGsgX5H3jaW0BIXPjFhVYs7h6W9uay5dOY6J0k+UEl9FRsT62DhfdMwjsREvbGr9+wISWpzFgP
Q9Ph+OYHkGHzN1IFh1AwL5F+Q5Kuwxa2Ut074n0QYAohmLJZUBp39UHdak56MMAeg1RQ5KxXzscU
cvCPlLg7XUKBgvwXb7xrR0ATmSLg8ulP8jiaJgTQYoD9A0Sax04IxhfswW9aOvRWf4jdHoc0+Q4z
XPheIAVDGagY8ASdMFgvrol0kxZupgV4NHaT7MQLrTHXYBL+qhCg1ixRjlJKtQoU+GItq1tbjkQk
lScw8QWBjvSfzK3llY+IY2FAJOGdPNvv/o8TrqQy/YBAJ5zdYcNtOe3Ua2AQvffytNTRpR6+XzTa
r8UiFk4381FwbpoMhplCwMB7E3ufrlu5/KuZSqkIVyi2TECwZ0xisIunclATiicjNaBHYl/bmdnM
+PeDVE+/cO5ebVR87doLR0LaMDWBLuO4xIGNQ/m7+LS2zRsmdDcKT7R6vR5M42enfII8u7zjBksy
p3ghJDsXypIJAvY09MZJ6m3pOb7wCqRbcqyCa1xv66H/AtKGHthkHe1p+sFAlfEiz+KokkfkdpyX
W3I7Ff57kQ8a77wvXZPt3IICa0OM8NLUCVDCD17PTsp1bis7CbtMq1dhh4OiMs06RsMhlPTbm6Uc
XrLhs4ePga1Vl/eqjkKKuoVVgLhU39bhgHZRRPSRB8VsH142GJS5slAr0ZXHfrs4IzCt1Ozv3hxf
/bkZIEzS9vNlEecQj3423HiqgJ6GvXevg7FnIr/h8NcYYTYhy2d7BiOhXTIaChE5mdvUavRr6TiE
5pV/mtOaEsc7QYfC7xVPf73r/wV+kJNZIMT9+3hfQldfyvlzWpxLMiIEFnaHbdCHl85RaBrqt6lf
SJ3aaxyeRBu5MJg6NtPRWWrAmNG7+b0x+VxSTGw+/sPQMoya+XemT+jCC6IevXXBZOtfFjeaCxz7
jX37652uQGpqvQpF5i0c+17MCkObN/Jm0gOpbmKH106qqbEnUNUsmty5WSMC5f8OuyE1pGJCzwjw
8RrDuRrHgJyG9g1Vbybtudpnxx2X+OwAJ/nbdjBusilFbuGTZ7AO7H/3mp04epae142wPWfSYErp
yKwzqGUf+rdUeYcSzJgiuiqSEzMxhVCRI6q6SBEi6CjCzlod/JwmzpaBnJjw6+vhQ14138dWBIc7
pCD50r1IKniLhHujEMicn48bUR7m5Q5jGoMEBhhb+PBNAhb9ebyCw/qBGFOdAiUyQTOPfIyKjgBv
8lhWrVu03R82Mo/mESTc+xC6fkBFIecjaTE2NsfZkRMa2v91pOD1mJnpF0wRYN/Yn0FQoPFcy+wg
P8kapHHe82ZDzueAZQlzX4ZoLv0ZSjMtD2umH+ro80RispFPxDFgFUCtBNp9/sCbFlkOxMh5etmL
9JQJwPq96J548XVzHydxMQm19ANLt1McoWRIG4JfohsNZkJlcv2YHYNowMbNXwJGFDNFqIoyaNsC
gs/ZnYo5W53aR88rD/38UGZ/FiHB2Nsk3sU5XQ1vO0vL1tvVKdXy5Mf1Jp1Z2pF3x83PFXV6IQxA
zucFW3jXbfEGUm51zocnlZW23NdNd8UGLXICIB5O3Q2V9iRCVsXeG2YfErFCQzzVQV/5FGfskU76
IbW4/hZs4FCCFScrfYQR27m5TBcpNtEUyk9f4XKmuee+768GogFNRcBoO8IsBF02ozgtVEtKu5Kx
guPLWqnbO/dPubO/mTbESXA33qtCzLeVQCR5C0CxsbQVuMZzfePdsUokCmANPBY0Fr5Wuqd+Yba9
A95j9dGAgjCcUVa0iCvoY6W54RJg3CpC8ImMJHx728KyPNGoh2HfBAHTXNSdIdDuqbX+5m8mRo0g
sB1E7v2ZSas8EkXKJJxPf9myWY6nB7OPDyAMvfJAflkQwGPzQobccUz2CPb8rZ0UvGZ0qIb+AlLM
8fOlO18FoiXFiB0yaR5Lw0a2shSJIbOG+shlNp15nleAo6vquO92r5n0gfJW0wjiPkwkIJMBK1ZF
+9U0hzBB2oZ6v01QwzT92Gp7QE9Xbs6aq8Wdpank947StMjY2yCXnBQNhLOlpvJswlkz3Zt/AhX8
0gSr5Rjdt+GeVcoUIkJ3ikDGX7CTs3qyvtOvGJdP7RA3enMSUtUldxecRicp6045iWixqWG6QU69
hS35quhVd0BotpJN14MD4rtZsVmB4GqETL4xuK7hZNduoFHuBau3cBM+j5mcfp5oWwQalA5kIVOX
hX7uZywyFudPqLiLfXxhKTri8EtG61Nd3K4I8F3hylqV1K+eRnRS6EsThA34Fg3U6cuJyT5m29gB
QUCUzlfutV09HGh2nzC5ep1SPy80k11LJDjduSPy20b5xPRoBks/Qb+y62d7AbnaejH7u/gI0byY
f+/INOxIvOqbxcTLSvVQ8ihg97ViWJdQXV6PRFsPv/mVspgFGW/g6l6viGG0JiVBvT8ZoOXzOGYo
6HK/jNnSizIAhlF/EmrrcSi5fPDmDaMhPhUFqtnyVRnGngZEg4qIBUB0brP6ApyHlyBKDtvOtdPG
xQ2V6dETr/cs2c0MZv+rCemtUCqIn6nnjdCYvmfkK4A0zyGO3DizyvvitdHDGaTl/bA3Vvm2YZ9a
oi+5ewq7ohfKkw7tT7KYsXv9ooCHw/+orP8eBAdF3HvZpl4dx5UJbFsMTavL5peS7UDLxg9B3ouc
JPv/58pZJvM1AAqINSIrONttgCzzgXEfxg==
`pragma protect end_protected

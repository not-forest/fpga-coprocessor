// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
RzCHVXk80EVTzR9PIgW+UNBgDwmc/WouCvY+bgocq6u/cJBFSaVS3fHIZkNOAigA
rVNMgXAwOaScZzXKrubc+5eq+pwXz0P7RhT71DJtIFanSnQ0q5mAJbfnP4wGQhcJ
/YESJbs3sq3cXS6wQlwkI4Oi5oUmDODJ7W5IX7u8gkbtFVJewDhO9M0Jj2cN5fWC
UMCWyV+EFkDi8R3PezevqhATM2z4+OG3J/vcXhn32fb7emMpE9wg1M0RMUSWrkWF
1PQGkJsIwCLqCu8b9pSgvbs6yDJoj9iK522C69vsT48pxzzh/mci5Sx/b+dtVwLy
zKbZTqVFkEPvO1l33zpvxQ==
//pragma protect end_key_block
//pragma protect digest_block
PlMlA5bWPVKEVPcsNsJl2/Bsw34=
//pragma protect end_digest_block
//pragma protect data_block
FiXsmmDKGvpVJntQOgG8S+tGPIGMcZHvKfvq9yw6ei77PvvsGwGPFeemJQYy41op
CZH66uNbimzQoF11YZybkeuNPc7DJlfkLdJLrghcHvOyuw/LUdabeFBbNf1nhQs6
d3Vlmtxwo6AYK2opdWBYslWHX7HmWoAT0GhObGMGahAknegjYoQ8IrwqufyQiOXa
9MoEM11JClk8EXmeUv8iv2vjYVNx+HbwQvcj9yBCXrOVMlp3do8J4vdgldWx1nDm
wL/JqnZOU1K47d1yh01gqDcsp0Ka4PaQE6RSkUloZnJMM+QpRvDjh0wrnKRb7/wj
GwXOiE8AB1LtdCxpMxekt4jPR84nQvtpXqn/kNMUoqZcU4E9B2aEVRA34rLb6c9/
pfHX0C5LE8Ei7yrdSmGgUJz4AGMFwFVFG2fZrVQFvH3R3nGuDca7cCTDWSiD4GUT
t8dUbhXRckfQOb/PbwUBfA65Bl0+ytTK1xN+Ezpxw4XkELA63FDuS4leM8Mlun7H
iEaRzqpNAEiEdHheridYOOWqx7tKrSkKcY/vKV2ThlKVc0jdqBK2cRu3URfgm1sT
KSCwYtjLth2QMq3ENvtvElT8xcgpVtd4QvkmIhGujwtWRDVmts8owwBLPhNqPjcC
TJubvbg8zSGQPQGreeQrMsGd0xKeQMXfAigO+jsAl2BKYp/YKQX17PHYZ6VBnSua
mIeEO0JUpqcKaYt9sHJ0F11Ek0F5Muik2Y4DWyB5VKj05hkEM6r3Iro1t/GAe7Dr
f1Ai2fUnx35eTwrz5jWhz7Iz1tCUwbyaUYX5u1cLx4SwVPKy/5myWEMp5no3SZdK
Myurt7JpjG4cvBQfs4Epd+BSPwQkbBKG6cZnhIww/6GiGcMQwOThQVgcIE875lMr
BMsewPBOCOuFpP4lSZil9N1/HMrV/SJyQe6EPFlF1RxlA05uqOmV7qd609q0GwWV
eF0hI6TxZBQBqheI09GJo+rj2yzj6VKbaYL0yX4wlnS1DfIHkavoJ58FzSsifzgl
yjpFUqaYBoLxkTKBfbtOHlWTxeke4xclDZp7JP60TsMwkUD8whrEOmFn92uxxTss
TOI0QZ/6BOwihEuhdN8F6m5YwuxH2Ru6lcQVCMQQfI+7DMqSHh3Y5pbTsH2OgMwu
tipPL/TopKbjpGzbIZzCzwWJAkJp4HEdFEamLgbZCb0z5VS5p7vJGfVZFV03BlTK
YtoM+FLOAJCapbVVbt8VmBj7PT5sh3S+NK43BLDEGPO0OYXMyvlQylDO9ciqD2gK
sI5tft9YAF+X20tfK/pRt2itZXfuBiinNnJWAsApriBoCHNNzd5kXZEBtbDn/H9O
HaOrNDYE/9EdUqgGhL4Bj0FtPsf3O9dBuW5uzSoRymGWDnxgoHBK7BDBAHbQfbmv
sWPMD8XGFWS5A9HOz5cofR3SuN7nOeCsBTBZbSci+OD1LGtu4Hvm6td4VDMwN0Ez
dwnl33U3dCURiCLFDFdrXfjNLwfRn5q6NTaFa7TTVagRVPYQ8rHLZfVG2Gl+BVVe
VrafowV8cLE8Y2opSTbdG/DxBJkYP4BCtqz3+RsLk37L/A3/YLb3tMbsd3sY2iMh
FsIp6SHZs6QmKUwuiy/B6xMdo4o2sBqe8WrQU5pZRcBo4j/kGtmPW+HQvwzhCg9I
deMEfgPCWKfHrOhcDfu3B4Tj8Rsxg6uvn9xbXGAzBsZLZ3cHtbCumgwmxDCDzoZu
LeQSTEsWoVo0aLkDb51z2qEk0F1TcQ9SfGpwX3CES8pWcq71/+58/YzGzo+P3D1N
7N/CAnf0XKYIItsmXeYa9lTxD0wWQ2w6f08nvWxTIPrMzdyBy2LJ1sraXCPFYVxP
qBcZM6qzUABOy1M+aUAvQVXUrB068Ez/1yt5DZ2IdtC83iNrxTXmA9NYitID9q4E
epib6A3sImlCAXSJkfClRnVic/MFwwc7zrMTgRGWmOiCanGQrmEFzViIymF1zt9E
1wQQUB/5TOTT0rbMJqFjoEpku796+YRGrpGUeHCYBQyB8NO+CtCndGt8r8JMdxrq
qM4fYBnodwMtaGUmn03OUnfJaPxAXeRJm0CFfr2fj7QW1/UACy3U4ZesONJDAt4/
KrqFCZ0tOyK+Po6SRHEvRWm+zvvNuSHsk8+ULrpVbKLxhx5amBzORtFXYYs8klGL
/B5KROW998ZTO2Wj+WOH2FiqoCZOWOqhyseuSL3vbmb1agw64UYhG07QHgLE/jWw
GwNqeWyd8XjwiWeEjLqt5zeuDw+X3pGMv4bs89QPZvhqSgKpGuD6j5UQzYhmlBDY
3fBXFWwO54EKTC4INnb2GVWOZFRak/yPiAD5dOxY4RrxFi1yJQ/G5I3tX6jyvyqN
jE94xXy/fUwjirQDbGtz55+VXA1YSlid0AwJvgKnhh9yNuh19PlDibVgDV1CQe5Z
Khohh8fYi4NVKzcflOBPxkIMQLBwX9YaqnY0B/a+uYKbeh5fMpB5ImwigNiZRC6M
JlkvGPGr1d9cLV6bIJVvczW3k/BVPYxyzoUfi7ru90XEV4XwPg69djVv7TDMqDvN
QHsP4WlNwD+0Xp7vbESttAaW3E+2DgE4iiusuh6VPv5DTXBcWZNqFHLhCIBWAdtF
vrPwJRIPpHM/s/wGAfG1JP2RIN59wUPaOksHkSiM+8xK6bU9KC/RYabTVNSjHTgo
MYjlVbHBgaM8kR6bZVvIfkklrAL95Zup+QpqquU0a7Tkgdcn7s++LmSiLRK4mmf+
rvrl6RaYw3iXj9L0hpneJQqSGqkyZleot3RFLmJ6Cr9UW3u+k8k6EeaZEuhH8RQY
4kZxwVuMJnpocqiwBFy+Ob0RteVn939Wa+nNBntYApqrnBXQc8kSWiDi8IHXbyov
YziTE5jvfhfQiNmE9tyf33ii8+Q+j+oztrKexbBEGSoKsXJipHWX+PnoKhOYED/J
+UIMb2pyKuVK+Ul+DMw5M03T01iNZxU8rBFJ0PEJKTxvvym1roLlhYO8ENDX383b
MclHvQNIKnPZa/nFKx3zUeIkj6YJTn0VPa14rRk0TFJDHMmLucYnhKrtsc+eAza7
ilxvt6gBhiqqOp8SO2UdmECOvWse3I6FMrAAIYvSY/bV4m5AXs6xrkk05qbkuvEh
xTTx/Vi3LTjVU3fTA28H34D+8l7uNq8XIJQo3PAvxYC65EG6qPHbOn2zxp3LS5rR
GKuvNPRS8Pe71rTTktIJNkO/6jhUvuxCcR5IuvTGqposnWUbZJEVDLetpaKTYSts
VO7Wj6ai/qPS6F5zv3jZhfw7UpGNjlHikoh6KdouO0Swj90IlF/5aO7pxCsF3gG4
FNxM+WEYu2fjTcyd14jSiBzNfRRVUFPQmip6eg1P+sCQIioQgQWXvcvj0iQpnuwy
ZW2FuYy0vajDk/BxK9L9fKYEDuC4X8XEvsHeiqyZKbsGA1jp0/k5zAREmW1r34n3
uHeJQ2i+mIESV/OORWCnAVfW87dUFvb9rFNUQ9b6v06L8ChxhUMPUgi+fB64tP7/
8hP5MD2Pe2Dd/SI4jSJMk1/T1OOooA0r7FeSkXMIJRF+7HzY2tjeWiZ5JONsvVHv
37iybYooN8nyqKeUFF9kaM75y5JHQvv/E9BAYc5Gy26zrIeJWcvNUBIRTR8dqrZr
N0s9KpCjWjMLa+9cfTLrpxK/n5I5zve+19+MQjrF2YWeBrAlkWOq/KBj0kflG/1g
gfuJQXT/fthN1VNBG+ohzZpUjgZ9aoyXANv8C+oikuPeQVdlZyiu8z/n0yEQzaqu
ncCJFx1HsmyGpsuc224ZMApKp5MvoNFWa4VGDNzrDTmJGmHTok7PwROrM3HFNu/D
CSiW69668sP4RN/X5teVX6PV2uEc9xDO8S06M5hMaeYTjxkNdRFdo75mu8sYlW3j
ExYfxeCiXGfvuuZ1Hz2djpzw9P3YqxzgYPwWM2ZoXRJNXt1o0CnODKWFsLQ10mX7
4npjwvgmJRT86mHMv4zIcBUC3MVpis0veQdKm8SoxBf69WFRHpjOzlZKoPp11rDx
Dae5/b1gzRRfSjD54BUb5Q0wD4VQWbmLIthBrsxiQGbDgiFC3zrhB4Rez1P2/qSg
nJhY8GnwK7x8wZlWZHqxxar2A3bvRd9JYxLzAwtzcytuDysDHrJV/he1ulW9Vu5b
5dviTq+sxE5kILeh8C992/cwQ/g74yjjVEzyKKI2SGu6GBEL27umh+o+Q7imQQeB
et8WEfwrgyPX+MERitXig4z1faGKZXl0dhomyPvEEhmp7CrjnihO68eMRWxQzscj
RLBn0hsvKcAlBbw6GLX2o6qItp96d1k8Ekuvn+dm3uabb1fsNCCWIXAlGfA64eGb
Uqgy9wQvPLovHzoJQH5xv/NnHzWI49YMnJEfQm3XOMBnXh9TfG663C+Hh2AbpbTH
YdOzuF816TyOdjIKeN/b+HhlmL8ceQf5IX9N3cAJ4ipJbubNGqj64GIqbN6vXHE/
od0EJxzlPQuzMYscDI4KIP5t7L7NjAQ/6LwpCzMaC/1AV9YFwo/F0V8DZ8ae4L77
LzWqhRweTYU61Es0DjP+e2gLepOKoRHb4MXbsljxWBIj7MkRiJs8YZkYDqDKNqWy
KXDqmUEa+Ywwf4KG+kKw3gyfyLvmLrEDTIziPHnWlCl9yDQYmP7NjxsIHi9PPCh3
L2BZgRzLiW/z4zIZ4kJv55sdEmKLF6EM3VYUAv48fMLcX6bqtoAhfgkVB4jMK98z
X2zjghUB2NoqsmttSS98A39UE1OuQZlm7KuK4+hRr7DrvouMB39v75ESQna8pnTt
67L1Kbye35gwGNICSqrdFTRJxOuH+faVbNoLJcgn9uy2H65cfsEkwosfypwyY88Q
b5FCdIXiQ2HgJDDj1jREAXn29x1NPd7hTAQCDrwTvv5RI0zI8gnJ2iAETo55OYv/
ElBoXW1k7n5mgmUxRbAlSGHgj8UyQxwlvKUHcGox564eri3ckpBv8ZveYE3h8inE
uGaZVqYzK0+F57Q/FFajFsNN+O4OBhMOpekECckpBdL6fOglmLEHDZIp2YWLSWVK
VDwXm2GM6rVn4BY9g0AJex0uhFHqUpVIKd4OKrgzADscKelrCi3mmJvWF7FM0Uuo
6LzkU/tq0sGL9E3xx0cbeOSOFTGxEQaHbBMEjwBFiRiUB9gc/Nbk9hRs4zFmAh2m
pkJRe3bbfeYnoSvdrJqYcle+ouVbrlvCL2IjE6c5AE5AafW30jNVm3oxDcbOKrAo
Hctmf+OQC/GnOEBLa2zCJ1X5shpiwI/vMSEq99JGbApCGtDv5RfWP+IZjy7FZgea
wQqtAPFSk5MCwoWtM3D8ctSEmXH8X5psJvvl1trhvHUbPVbH07b9q/Ysp1eryq+V
q2PCCODRaSjxBTH1R+NyYQ/swRF7QV594DUK4Vuv5FxHRY2hmlxHKJM0oSOqeZnw
D5YSuyTdHY5k5MhxCZyTNZp68u2oNbHJfKf7AnDXwEb7GtT5/i7ICF2FgzEeqyDo
qpFkA161or7rvGcADkbJIvK2y8gqFwmIKIz1obSGKZFqEj12J4oLIYwE7SL+Q77p
co3JhhVab55JxfvvI+wstySLCxR628ygNSquHB95IEkiqAObIfU9C+DYynZwJmx3
xleNSi7IlryZLQRLIXGp5v1XQ87qSpGECZc8uLa7estYlbeOXREBEZawheEnPLqS
wju0VyrXUGF7ZnGs/waXALm73QNS4TYZqx+Bhty8eJ4CCayGkIvYIPtsHMtLShtl
L4mJUIQOQPV2rRxf+8hCj6uvAb38pUFgwuuwzvJ+rHPVfm0Ih5rG7XDzHOlVY+Ir
yXJOnAzzP6OEt4HIQv4pZRba0pJS7pLHm61/YkAu7WvMjrNQk7Imhr5/uklKhlvV
moUk9FY/13WdzVOrBE55UUvX5ka9Vb9DSprkBgbZlTeHJyHKP9iwDp1p8ceuWxLA
FFTikzo9BlIPswJRIZ4mQb1r1vJCcLnPCh+Iru2b3fW03BAcdDwDQvb1XbUec08c
LXJ6Gy1T+StPY46MR0T8ezaLmCk3We9ciieOg2AwPtHhUc3c3u5wrBw5vEH4gTmH
Ms8A8a+vXtE1B9Bbwa6BzdLWggcmNqhkTF1+saMQMqAPVkA5egaj8oh7/4PwmUY+
cuOe05nOIDABgBcpu2aCAaNFgewM6EIIzusSILVmQq0GX3hscu1+gCEgbSk6WKye
zon/MKqn1THPpbFFDyUyWJqP9qUgEfnvNE4PpkOq0bt26fC4dvwXGS1cGQdbqWOy
x9soCLLXqgUJvGk+SBvV7HHb+3qyLmTZaoqZWJVTwFxt8Zr++mW1Kzwtc0LtqZ6M
5jv6o/lClLR/Kf5UkQ4pWOA2N1hmkm6vDRoU7U1/zyzo9ZqVuN1BR4cUJEIRCBk/
OkY+aSKAcEcIGVkNTf1bN8YWrGzFuGIspgtyFZ9Og7w/rs0BgLrZW5Bt+x0WDDg6
Isnx4BuymyAeLDd9VofPzdjRoDpeX2D18LyViRUDAU+4kT5xxw5Y3SzvNtMCJZR+
yVG2l/QKIrD0ifjX+CT1A5oUKM3FsLRqnK+dFBR6MecA2IxeO39eNU4gls5H7bbH
PFKgg8iMAhgJgYgX7VnpOLK7nmie8Sz1nQL5Z1lQ3TMtCg0/t+eoTSB2dgONsxRu
RdYEVRk0oHg5FnL8K0CapMluF29vpgTJxRpHgDu2W667SjBphmVMXemzxKBFqcpV
tauGh7FBza7CyXLf4eCE9DZATp7c5tzzk1Uty4RXPUkOSet0V5zRZkGupQNjUFme
72whrGtJa8jmhr/wmo5T3V492R5/iZXA3Y7DRThxGJeTbinG1mY50cuqZw+JrTbI
EVD+4kJCNPQnbFiG7VGIer3zKk9f9WtroW/22z4zDgo4Pd4Yc0Y4DjgXw2hlJlui
tjif2yjmewjZjEOCqIz4nURoILHRoGywZ+jpPd17LZX8xWuFJHXwvkD9ltwYjKtT
4HkILT8Uw8ixCAZpn2digYCPzJQ/7MtOEtCxXSb02uCoZo/Lqkbq6zmHK3LwtXbD
idJNxIu8YR52VT4cLmsBfUZIse/Nj8rLgSOBUa/ep2h8MN0O+YQtA1/D2EAoOI6n
4WvcSLPJzxASyyjNPaVWY4o5wutlzqp3WKst2CqNMhNQF1Tp0A2I7oFeLYyIEF1N
9+I/ZYY/XAHGGx943zsEiSw5vLkixetvYJ0FhAPzJU5buoDHZVuxtUYAoYgROwN2
tzhn+E5OHA+3G6FffhZURlMmZCtQTk3Sqz0XedOxnyBptmvNwyTC+mRnnIFfzuz8
YjlT8JiULHCdj1oT1wGZ7Xwwu4g0RDgdzUx5gbFm38KGLqncc420BpDM/GB7odYp
E9qoeON+oIiDUiLchkvJRqnQqJd5UopmYvPXFuIv9ZMCVuI3WF7xovUu1iRLf87l
aR1gw85MbgeF28vd8a2UAj5WbSEIjGWBe9aHWgEwjX1cEyqN+uOArSrnE0YQ/pK1
lO2HuW4Dtw23stph+jB+VE31YpW/e6eRRpNYizjGQdXZb8Q2y8KCGzWH2Nxg7kwA
AreY+ynSaFfNEFJRZ6huFnOKDHX8cqxDhG4U/dS/HGB37R1HnfacBFuB/o5P1qPW
xfzgq/HR6m1/66WXnbT5pKcdDsB5d7rAE3EQElKepv0fr9G9/Pc5O5hEl+eI+iNo
aLQFw25qSO5D6AB55WSSe8H7s86oNuoh7S4IolCH5pGab+FVv5eel11kpzFfkDaW
xtyjUa6a0i37MhCsakoIN5e/xEIzoZsn/Mp4RDTwLG0eaOog+a4YS3q76t43qrtC
pq8I4YjUYynQTsqTK1OdVTPBKf/HWvXA4PlQIf9sTqwyMYj7LRCBj/taoQ91Hoew
qXgjZlwToE6ShbB1zGl8b3/y++WhugVB8FyPy5x7n+rt64tD+MK5yWaTarvOPmJT
2WMtUinEWsoP9GabrcISsC0kJwPxvsb2xtkSjf3FgplJVK5tAFD8Lo1Gx+zOgYS7
NJ1EzJW2UoviPKRQCWhhu4lOpa5UEEudie+clSULIZkd2K2aej2WINVsZaJncmNN
j/9JUZAS+LIYUWTC5IkjWY5jMeRzWZhvtkVVpaSeqB9bLynb5OX8eCK3BKjeNPQB
4ZSnm68SZIxFUpA2TzS6phGuc+dSKaaDuONcVyeCUzn7USJK9mowxmgpntei4C80
JurWCOfejnN2bVxplgkZV4/TdXBw89G6z7aZJfwrc3RhoYB+aX9cNMCMVM/f9FaL
jgs7wFcFndPZeFnIizh3DYiGezHsmCZlKeGPogBwMupIj0dS0raEKiJqv+Qvs9UF
cpSMPnJ+vSA3nkCoSb3b8bGJ/bpu9LA3eLthnHA7bWGYFDbbSHysyzvmXyB+jfVd
e+QD+kFYr65cjlUKVvllB29XqcNUxEjab3dgsZZCi8b6FSD5tvfHP2BiQNbd681s
qW0ZrlqTy3z49wVPxsOCTpjQ2IaxrJ2tEA8zALue/eSTlrWSsb2zU70C+OQ/zhFs
nbHUxVbHJ9T1ucvbsj+uUrfi6++oTkyBmI0Qkbs3Qfd/j/sxo3I6t/hWndRXso9W
V+5k7g4VBI8Tn3sf1KXGtqhi8R+/Zsdt2Tc6JywIUyF1jqZJPMUkbgTvygtc1zPJ
NRPMVsOf1Q9IKJVT4nsUFdGQm22TBwmow4HhJzqF+fdI9esnlP5qTGP5rGBYDq0G
zGVPllD3lJ8cu9F7pxb8BVGP2s9MMW4WJXueDuwAF5sUpAnEJCETJjL8+gf/EKFt
8kMP0PAkPPUvO74GHNikQr3KS9NBDacUF1O/tUmpRaKqlzSEsvg1qhtC0g1pvQr0
7VvnMxLcEq5mCxoSYG9rsxD2k4YDA/J63f9Jh/pfqoqxISX4ZgWxwjI/vxLnKTOt
K2AQpL8e7t+P4smXwxhehr7KpIxVjr7KnLamiUrwCLfHa5fpk/1NsYJTyJ1ooPe6
atRLBmDqb8riflPHq3AvToW+sHegfd5S+S4+dFcTSIH1Ej3Ljysgll594D8QsvQM
kp0l5VKdFsARKhvMUofw3hFubjcPus0kMKEITOFYKpvDQz29D8p0S/Iy/nltGFnK
uWBwD3KL6W05TSe/qUYkEKpfzaOW7/UMUVNNft8LcgZQIL8l1p4nDL03kA8ivwPc
kjBZ48P2lvM5X7pjHhcAXzmxrQK6rd6W1mylB0fGkIQUagjpfqZ+yDl2YAaaSGfX
igvKVEQXPiGRX+44YKB3m/jEUEtnZdoAsxK7tmwwpekZZfEj5LBsXvHKYmCbEvSi
0d4hQ+/i5lTDK5OSOw7QzXn1DtAcbgcubkQwZMmdpfuS05HcmOyHfTwPfWYT3fUW
YWifPoSyaSCMTonZ0YzwmayuEtJ8bYJ4XDWOvmtF4YJP1TYm6aO5Rs1s02vrxExl
g8vHyeIAD/Z6s4aZcHud8qVDtySdw1CnZ58MwFP9bfqWclTa9WH2HpOF5JzZtrPn
cYjSaJqr+U/bXiJXLByfUxGNjgOdpWHQSWdQaRfiWEsUgzkzqwyQo2fTeZ87+2e+
fjZv5aLCBj7IDyzV/cHAv/JmfYX1xb/uJEJBfCx8wAkq/vyJQoaPD/xv7h9hv4t4
9Y/mOfkEhm/pYChnmm3aI8zGrccs89NgqanG5ecsKURdiOuu3YvALhUAYgQgalhn
TRHoFp/2nktMBaYfdDt6fLdlj3J7jldroCZT3SbVl2vzYnwsV5bLOUYbTY3VpQAU
VMx6dgQeAsrqvDqpxMGMRlOjZ/qHBSRZQRm41Ckp7j7KJxi7NtD64S8ZUsp/im1P
7x6BzLikfvWexWHKYQk6Fje/oMxz5v/7oMDP4Qs4zX/hj78vWBN1osiUII4aXP/2
Jzk8EekDPbPEGnP1MEOAQOVMpNXtrtcAipFmF2/llBZONlv+hgVkfqnbXpfuKuty
+ifHXLivkax2/0/ceomeMyzbGJuLcD7H6ZhSGfTe62Na6uFnbbwY1rfL1aBd74WC
XClmr/SQx7pnaVAAEgFu3xSiWstNm4CQoMIAVdWIdoTaeTBT0hi8galgGb83ZoT8
xAgC7HVxrJABDuk6jzBkSxsUDT+7de6fZHznlw79ylBgAImStGBkeGiYA0Pu1pH6
+g+VE79HyrU2B3HpNRPQz1F9k2ZGz0V9a2QUJSOdLvd6k64/nozOHPNRt8BoLdqq
TNa9nGK3yL3fxy2x5znts2R33wYYnNpFR+tTPvGOz3RMmm3+To6JNR9zMnHwbyf1
PGJ312eV2TGgI3jVMRcZAdKTCDDgdkd0sqWQ0F1gp0DK7m4fGGT4uDz12TCFBag9
bb++SyW/ftxXbQIgUp8iqa/DiWAhd5lqy0tlDxskQaXj7xA+dqAcDlXQt99DheVe
4qedSEOqrZWBvTLYc2uawtZHGQmeLPKx2UHMl5Yj4czltvIrt45kRh5EW+/rS1WM
633uX2NPJQ6DEE8MJl4/3wh6H8fs9GNU/8uPd27xtsjdEKWj6g4XfaRMs5DDyyQH
aAuz078vn4huHY8cpRJD/hLufMoISBM0JEMJZFH/RaK4f9CbhhB658JxMQHM8LXH
/2MUfIBNIeRExLkpOo+MG9lAu0l2PXL6avhJVPUC7Ka4DK+R3sZ522iz4XVIG0QL
QY4/FVqvz/oRpR6YcnaUIT6MRs1JduHyVdkFoS08yLdD3r0Lp2j45I37ZRSoWop+
W7CKZUYyWfU2gkQvzwUotgXbIzI3CzXHkckfxrQXuSTGgpHSCjF+g1/XcsdEiqY1
+x2NjWKR4rYQf5hZb7rN09CAi1fwU695kvAMsFUwcz68CxHWx8aQeeHXi05+89UT
ZuCO9y3QOgk35JnRA25fUFu77o8ib0g0KFIvJx5gtg3MBBny8oMINmwQy1bnhPeJ
x+UbRi1JigC7/CwIqi0RuSmkRadJ8GwnUor40zahlK3VuPhpResMuYruhh2Haupx
Dh1tA/MEc53HHzV1wgKg/EhLkgsBF7WLFZeo4sdjevGMPduaZrJuUP8iwp0Et8qi
XBqq9/og6qRKIeSGZtx1GG8MIAc97zouJd4XaFehyb4PTdg3ARPOmctHPrhrpeWw
He5pDiop/AFSpkoTlBAcBThVp/PksixBbrCP3eCzXR4BteH7kvyqBA8yfvcLaxVq
oYriC3+WP5k06dAlHRizszu/FmoHNKDJdhWVKDt545iCGeN0FdeGAfgn2LqR69jf
Vvi9NxjGQEUgQ7pY4WBiBmzGqfpDDijzQX4gH6hinNBIYYU6TKBbRxsp503aVmK3
P9zexDFueFbWJLKckFEuZb5s94AC+MsIIpcFZIXdH1nBkelox12Xkv6aZnqc1CHi
zTe48LX6+yZRcyS1SLJEYi8idX9Ch149/INETjXyOdC3Vddjarj0F28S49pUWzPR
LR599FHWtdsXtZ6QmLy9CdQYQVj9d3e0gPxrFuOhc6l3kssa50GptEzEpWmOOU1C
pf+YvR68esFllRpLsP8BUzwLmYxvLgS+NrJUZDZw9npQd92b4o/dkZdf0o4siTAL
0M92CaNQdOCCWPMcIXMx3la/c9L5kIwdGqxtbgNkkP76BeFqnMJoK4IMgK/Nb+mG
w/uDjKl5VUx6LIk0IYZAHzInvOtU2YvwCk5G0FKBG+RSNQu9hVloPakYsIKuzy5h
7dLolan/44UylnoSe2A63OV1F46UnokcDnTOQ6/R+Klc4ICmIqadbZHES7i3mpA+
r45OJZ9xzZF9O6nrth8M2R3sMl+glNwo9ojW/O/xQBzxIAKHtauV+x5xGVWpFDmC
iHjlbKcLohQNDYIFV6zIotQSoajQXv3kGd/lE8hX0anOW+wXbJ1oR4s/ZjCi6h8+
jd1JRYF6j35os2hPP9391aFWzFL+Ye0A0C1Bx9COdMHWYR76eKwJZKxcTcF1c0zT
STRTq3pYOtHMdOdryv6KuWNcvoX95Fh83K0BB6eXejf2ki19J1Edmzo602Of55SD
vDJaMNocpBFwl/p3VSnFGJtObxu3GVaqf6aQdiezjzgexpUbh7cnn0tddDvIUT6T
teVzPRgvzr2NKVCtFBwiMtlDB6MFZRm6tjs8H0TufNSk8si5jVA4S8DkPpn+QF/T
xbM/fdiaXsHxzDju2PqYAw3aAmuHcpov8+gftfuHqHU5Wxe96ovR/rAzvGjzv6tV
YDEuDnBoyzgi9OvGpAvaEkRJ4wvTOlDFUM1fXdxnGybJNnI8cRu+4bXPTl5wtrDn
T+UNThaKGof1oTUutlXBe/h21qwoski1Mr3PJBwKCSqEtyPMTea6FstSiedfe/LO
4qIVxjsp7+8XWpeRcZtfa1m/TYJD1+lpADdykDccxFUuBmF+wKMBe39moi3i2Qz4
pdDUceSmjukiEpwJr9omvxD9j5HblQQMZeKaAkxWAf+AZr3ms9UX7CjyKkgOX6V+
2j5w3uqJsx+cbgk3Dh9rXY6mHpcMiowGN/lAaiEK0pOm3tDg4wn3FkbIXLzmGYMC
T9y6xNxjc2HO0nZ/QZ4CLHa9rVBaMtNro+EDSxfNXl5qJZSQqAAOBADKRb9D4/ha
kd5tPiwsHw1PWR9RyM5k7JzlHZoyT+y7wZWqhIZTfmqlgNmf9/XJ11wNvaxz0GKf
7RkfpoG5JSgtcaGKI/Xa2hyWfJuVhtw3I1gBf2VgvfuBWxr/O2qnzmCr8/21iC5e
UkpGGzTg3ekZUrI8Kz/NnVu4dhGODF2+gi1Y14kbXHknTaG8IWVBWuWupgDAvSIx
QgrZivnIT/cKhCGPcbQ7wdD3q+0toXQaBC/9fRLAgTSNjrP3DNEas11lCWrS9+Yh
fwS6WktXdIu6HFEfmIzgYJX3RB50P2sGLYMUxcTfevddI5olWYSz6ueL/8Rjf5h5
+L8oy7Du4Yc5IxTj0FrZn6yos11TSZ2eDAXAjUwsYDmU6hXYFHPZNNnalRTjARuR
PIdbEBcHoPPXG1WcbuksOlIejopE5O0LMkfitwtN2IBxVr4INb3N2i0FaakVlxFN
ijZXzhPluIZqYLPSqnrUiGslmTBz6Z6hmNhozp27d0a4jyRwmSjOF2dh38LGc5ML
nVTgDfE/ITV7nvEIQB4X4rw1D9/p5PNCGXkp0l9hlRlPAcsWIMN6i+DtRcpfwOz6
/z2WRT7q3S45FSb1wI4h5wVe8Mu2kZelPHPnhUJTRJvkIBRyH4+0sH83icZxBrMx
IaTWHjnVYsSNUfgJ4GudQKhh8f1fXg6doiaHtbEFUgxYqH7532V1gOTVDADhEoBB
P56ZbwbTpeLVD2fxVgygHEG4/5PNaAW015vPBL7GCSxWYzht9Sr6jHQKSzb5/c10
1FhXi0gMEBZ33fAmERJZVoafqL6qXccM3m/NnMfB977tT4vl0h0yq3Y6VKB/gbPL
w+xVNpY84t7gwMH/lEevkxR9tBlXChlzqIGE2o7goCghK7RKmLO/KHk++WIeOUzd
e3l1pTnDdPmMoBJzV95Rr5wChrWMKo9WENnJdTpCUYTiQBkJ3RwTfO/qeJ7yk950
8phJot/VCeSig7/YKgLweldS7v5FrjB2RNkMCPMgz65xjjfhQMz7WpZA+nq+Yt1/
lUE56ragTBFolCujS2PLAKXsnFbU6+YUfOpN8872MraTU0tHLGr4pzB7h9he85yx
Zqb0EpvrjrGGjHMxnxuqSUkeFVisdS4O9SH+U6XLCjGbn6HqPwdMdT6mL3aZqZb/
5LGrbeS0Gsx8W89inl0SuErCamOnubXs2caW+AYh/x70Pe1coy+nMsCAzSajpjZF
qsEPjN+KqA+st9EjV6i+lI4HV8zj5gMoxpNBYDY8Be2Q2FMrQ5JAlBIWxcKbM9AD
4dj1cZihnzVBxmakdXnrJhbBNpdj3zVHOH5G76da1Si1a1yqy3VnzU9TGLYHkCeN
DO/GoILy+rWnKe1qGAJ9NsFE2T0/Az5NbhvkmVrpol4ZHu3/qqI4T9LGgBZzHczv
BtJ/pohaURBFqkCtsUygURfMDlaHODE5XHTzXqL1QoF+ukgEqdX6beOmzLIBrlZ3
6LaoEHeyLoxVoEYvQCp6DrbWe5xCTbZuyCLaHj60DDbd3CMiPhmle30DiO+7T25f
H5J52e9nNhz09lywQRii8qrhj90cKGdSZHjjP3Agh86ByOHBfogA5/oQcAoMipAr
c4jxvpE8P/+vN7g9W3zVmHKCRlKztS9AtEjBkEDMoQJSZ8iWyF5jnnbW+5cjdzcq
wt8IQVwEbPtY+ZSFfeu5hz0gyKt11sqC86d/AnuXPRLp0Jr68klWdC8InkxQXQHn
lfIRUikQbDb68jkK6A9oiv94xjxZgZa/qH/7ZSfH3ZfIdqdARlkTrYqcwz9F3CtO
lE1xbIolWAZVwuSM9Xe0qzWfJjufeNeu4mz+H7vbuJAdYCQuKkOA8o/6rBnFACs5
1XC3zl7GWy94YODy0fNkUCinw3D+RwfRDjtXPf8X4Bu+8sS4267Ic1jKEv6sKvNS
SDcOfkYCOhi1LqygyhZrsXXkcsI5/AvTC3Gc/E/aGNZtD5n/+8yc6ufvoEmBWIvg
1htNNSbKshdmfkbsCtyG9J2N1Glfg4FA/CTJPIeQRnkCNOwRRV94iygwv9tM7GhE
1piyyzAmbgx5rFpWkIjPDawqItw5mTdF8ByKri2CiUGju6qaIvqu7Ec0Y9cOjphF
4DB2QcsJJgdDWHL3aRHzVrJdFhxYPTI81KeQkdkc1/Fx6RfumjWArI23KTfsyaEn
WvuK+n08oNUV8uYyrbqY2lpE8NBXG08H7f+ekemOj6Zo8ryd+L4SMVK+534B5NEx
YD077WibIiSymQLIELVvleF/CS8nZCrKbz671OjiHwuOTLqVJJJ/s+9U1Gbfv5kH
DxYVflkl7UNH8G7hK9aWwF9J2vE5iyPE6FzWbgG6Hc8QHFrGZ9Hmh2J5xiuZb901
/GiKwMn/wNc8zQXcIIGvqh6weNOaOLas790Hsv5Xqx8wxv4+3mKxwKSV5ucFsAZb
f3ZiKhbOXy7SPF8YbLHMPaRWYL3VnuSdu8LVQHm96xoZNjvgwl4hoHVW4T1tcHOO
TPxFzlDU0+to5Xw+PZJCt8Rkry5F7KAWODJfJpYoSKx3y8u2v4A7X90oXM3vYKdt
EmD8u2MhvwZwTcT8IfG71djWz1MsqoyoCG3xuyymmSbKwtIsJipwMfRs1MHVg1sN
6Lz6Um28/3bxtLXnPTTWvkXSIio8fUTTMp9Q9PASX5mtsjJS8mTTqeWvdRbdYGV3
WqiG5QhrJbbGILoLZP1oGiTaf1Iflg0QHYp7mg0niB7yYzlSQI7KLdG0oUQ0lpJy
0vTJB1zlvmI2UiMmEr/krgyNNGNVqYCBn0MbxsM4RwKf8UyVRcs+34KIMkiFJ72T
QNoHUvV8PmCnP4BQYao8bqhokcqwG8y/uScI6Go+O2/oNYXQvWjg6SZ+K4MydonJ
+R2IZqoUBRStk7WQFjSo8EMrdhO8/twpecfjVxd323bod0HXYtLcqg8iOx9izdDs
Xw6w/OFu8I9VmEiGY6KXStiXtt4LDZXA2t+zKcSSyzb0WFSVEADkA7MFb9GyFaN4
mr+tNXuHBudPOPMvU4+n6QYE2Vkf+p+3T7gv2U3moPD2+fjHVwzjkJYqdQl71hQ2
5u6fL+D1hUiGV9G0+ZiLgvqcedxVTRciKWnY9xzGGi3T57X0G1hLWPbTUk/4dZY4
GPG36a/Yz+YiVQXLXajRBI94HlqIJyVfVI2VQ2XRAAopJ2vS8BSrCqthp/CxBWIn
uMm6QXvYD9sJq8y0N5ltukVwrnbOGtcbZ/hlmwkUt5jPd2sdbBz1DhOlxCpK/03e
wwhm0zLf4EiLKNC/W8t9Dx+R8S/1lySvtdchaE1u5Ynrb11te65f62nNC8Ttxk+k
4in1Zjo1S2yB2sDgO2n59aGhXAGpUKpm+NQ7RGdVGk3ekJHqSeLCJeCLffss35r4
6Uuvp+SGHpHMItpRk3kgJg9S5qYXxJZGes/GsmcvmINmKcyrUO6gyQwOVyhFgm2G
XhvRMQIxKvd1tmX0cvwHxdr0siSZp/HsptRi50nnADOJdfUgNIprWGNZ8/Sd4LYS
lOusRj1nt4Aq54pmqWa2KwEMzCx52raaMsow5J1dWffOGpMUaAkmrJ7ZVn2DuOgY
zZHrvTFJTAS+q1Isd36El6ieD56MTyiOVfyl1Hw+KqHpwaTpUW/NwiUSutInej2L
BHMF3PMsJALIS56D/PuCGdf8aA3jztpymHHfcP3IBfVq8IB3Gidp+0VwLiusRfIr
LUadNnn0AEa6kOu4ZDK2ZlEer7muOB8qfnFzHFiMU1HyU0eJrwl3aVQkIt2FUS+H
vG6DjZz0nTxnOZnK19J+vMI7SpCKoTjuM3tVrA0lyPQMN3R7eFlaTFehdk9dLhkc
DJtLYA2AgLYv1yF0chpPPvZX1xIWUPUAR/4FI3ORPERGDP0McMgNqGWLtVsQlr+1
e6n51ZKWEHySrPS5yPr9pN3cPJj2lbvIaDz+FXbXguHxhRQJF0hdjEwZhNkTwrVu
Y9g0P4fqAmLmlGXDbxdTdegC2MUcdS1XB5phtsst2J4HTgRxLQOCtHXf260VQz3k
OVwXQfK7n+a1n1kC7NB2u1PLmfvot1SWEEa/ILzFNk5IojyE3Ju5FmyvAcxQkznq
B5R5nk4PUtgmJE61vhlCjJylSVbAhwRn9EurWICQ5mh4tryaFFR+39Cpgz1E+00/
TyhKdW35hfhhgCxH0n5epTTr0lJN115AAmGH4AwFJ5HX922OSdGRmivItkDXkE+S
TG0o78HiAJrtHtjfGfh5AQ7nOVA1abuTBQg3lWXbnpj0+OqZ8yXPbxm3bkw2oG7v
64KTP0SSNs18rw87A0J6Mviv6Xw2i1OQQVLQk9uheFPm+t3XchO8e1oRCIMJTtlC
PRAl7q3+YPVeXLLGooVYGelVghUAy1g+GS+z/ZMZ3FPrqjzDoToRQlg2J4WN2vO0
TeRNoUCEaDH6xE6hXalbqx9464Yj/CmBEnMM586Ylfik7ocnIMzCK6tN/y04YqmU
APGZylEQ8DCUkMo5qFA6gOleF/A/+Cnp5NssQTMVircHRdPLjjkBs9EACGtNbsZa
6M3QRDWr2vTy5esTssuHMaG9CFMrkylSne6bISqVuSHjmP68oNzLso7vpkWe/3KW
1pgzigt1IRibCm7UZoEcecLPBsAlEXyZcLIsN3dnC6ocoC/HiRF/bqqKwVhy0lDx
M+XqYiJxTudH0qMAx7loqq2826WkPAry+8TlwsAaReWel2ipjrhg5CrKjzvZEDHE
hHGS8iWozc4vXkD1oMOVLPaDkqDS5D7+2jgWJx4jR/o+soSuIDX+xyjTogZKxVrd
RrmP/YQTVMOOZA1bHMtd9kHl1qrPYd7puTtOikGCue6eOPP3mVEk+xL9rxa90mu1
adbZxG8p4a3zJcGIYrNVquGmYch3OhTzRFXcijqGeHmZVGLiRfD8SAhTyVorEpaA
OIuPzDGQ3TbbwZIJ46sM2Nprf5g1V/FhxSnaqTMnHlXJJpgJcE+2c2aTU9EvnlWN
05RLKDOPIsNC7BMqA/o7p2u2vkgkGyHQR21ZxIQh7/Teg+fe3ZTdH5pExiV6o8j4
NNah4OLU+PDqhr1Ld4NwHlBH5eu1s0qoRdZzEQERj+MOyOqSSLnGMCsL/wgGr4Ml
7nDZ7CYMSd5voOXNPlFZHz2QhoZ8CEaZg+OHaAa81o4WDBuO2Oth0mbV4iHeNEwn
qUz30zFKWj5IniljC4x6TnelC403Qmu+d5iXNgtw7D+TuEdoGVb3Fr5+O7hqQufV
gNiFB6t2ZvSSjTaxmavkUKjvDo0N2YZRxOs9fGPwmb9I/N2CnKv5K2YA7GpAQraW
qmET9H1f0lN5C73T39V9f4PNrDFV+G2Q0dWeqbw+Ylefdx3uBvGpUyFckTg/4QF7
vUD7/t2UNQ7sfN2P1j7w0SuPUrIlbk2yEObyVQAU2yS9AHFtOoRblSY7gxy47xPp
eOqqb3PmJqdMcrNETNzbIWiHNlbAnVqAZTzpESACPiSz6RkMN+QKBBM7cpAM1Hae
j+d2FZVFUWB1ahbnxUp2IbMsFdGZuqHtYS7yg3dPzmq5uRc/Y0OVWUBisdn40+mZ
sj+YgmfwCC2OeqE71jlBCmdSGbLwZ7vJEBz0nA+p2HljFjFgh62QlZJldJSV7O99
p+iKfuFWxoFmTz2JanE3mAAGRZJGCaKOZd5p4nVKa6y7/xX8XFB9y1HypizHDGOX
22DBmGEwVRyY6+3N9v8rxn4Jvda92NJ6jn1nTMeOaLoL/1F9Fr2wapjSDwNxMmFQ
2k4FVMKNzGcrmlwzrpvTnFoXL0oR9uN+3ld2YojkxFeLSjaEfhoMNiTyphofGywS
iRWrfNpYvimrNFu1VNAiWo2v591XfhUxvArXy1YUudG05cv3WTdUwTCZ9Y9tWVGm
T7YnRQnogpOaLBGRoP5LnYyEs8QogmO/pwoYwGf98AwD6u6UFSBWxlANTkfCuXaO
Avygn0WxbjcHfNIl6g+XNmm8eSP24NVHGdyGr8jKgmk+2CYz0auOBAGhqG/4RXce
EqZuVMgRhiX8EdPcrFHQXvWiHPgnW1ohc6K/+9EMpMQJ/svVVG3xDotHgLD1A/85
k8snbt68emUAXPUFmqDi5RkYrX+y3UFI9Js9vD9/c/cuPxSw4WQSjhbL5RnnJ96z
yye05T5S9rZcqx21co4INxTBHt8HtJGHhI+X4q7lvZgXyQkwR4ckcHz4LB3aEHI0
Fwli0D3qEbZTB/gLY8AjB/AdEXAKAhB5iHn8bQruAxgA+eiZilRHoGW5zVOU7bfT
/34un1d9Tnp15lsfzjLqUCENCCgf59ytJEFlmRuDVTUl0mV4jj/HZDQo+CxCOTHG
jtODY6RuLW4qOWYy6UeR0F64IaLNQ5EYCchDdxh0uRQl+iBizy5M8XQXLUa0obCS
xCuL+Q6mT82FVlRMtRNpGXylki8OM3jxyzYHFCM5HjR65ozuqjUW+AueClGNJfNw
zmOAOtvzY5LNFBDkHdh90s9Oy9JBuVwsFOWna2C9ZZs1dUXfMn1Xn5x3gtT0zvMQ
jfTwlbeLs0tWjEw9GaBvdxBElJ8gnNptnVh+3ARimgVKtkEuSRkjIjWPJMiKOIUR
jAEIb9LVztdrga1pRAWimEZw8sEV5HG+8D4TS8xr1ngKSxLVBlT/AVKDFGlAcx5X
vzwqMppCc8js49rjvk+6g2B56XpTIpVUeg+U4kACdKK9JOp6zr54r7q6CnxnJEnA
csubK7AuSl9gorA85trbjRsy0oJA1xpRngm3/vqygu7DgNhqUOabyhAZHKZkBpZY
F9+aVWFivgT5WRmud4KQdthooQ67+RDhd7P/w2R1Al4sSD2Y/7zasyykQ3wVdtgz
tqa7qGid+0xQMzemLpYUI73S1OmTIa4YeYiYE55pxx0VefFSfuhI5eEe3i1EaiPE
Y/IbgrftbYlga4UfYVskZT/JvIuIdemVxWPm6+A0L6eWfz2qCm30JetGvqsmj9qy
ba7Ydhh62q6y+TRecigKvlAMB14mH9Q1RP649jY3Wjk5J4Pk5ph8y/8BpxCeNbGu
qX73Gfrim2mvTdR4ciYV1oHNkvjn8rEx6KzbvoCPQExBFwIYmCbpAp1VGodgf+Wp
1tmJeVXSsjckwPjV8W1nPPI5QJLVdwKlqLGuKUSSvjHd3XfbpzybqiKXAuNHDjEM
Wkm0Mo60THd2sf3MOb1A41mMYWTjKlggUmF67V2b6j0s/WQ0sNTtmFfRptx7aPPA
n4Ep0y6TBJuB/u5McDmZIb0Ea9UQGyD+SQ7aflXCEEuVpU7G8UDRzn95Xh0S9/rw
pAqdQh5y0eILcCbmR3b63CZxDFk06Qss6Y6wgXLV40X3rRi0CtwmbSK+L24gUnJO
hp/PprzoB43eXUGRqOFE7UDnFPT3Ex5ruSminDJmeOdlMrw8aCSnNVl26qTRI8gX
lK50KjT7diWjhiSGz5MRJ4MRDTI/YLy+ymosYOPkfBnH3RTv6n7BvBQ0mMTlFfy4
2tsZys9bATMm8OrikHxs697psdf9Tq1p3rRNVyaIn0pNGxFVt+qfBcmyhGjxys47
x7UuwiRciIG3lwpxn/EMJs43XpzCdy60MFjrAs156kG2jNwvrH6OvOGCixhyH2cR
3qj11uLKHzLZrXCSbk+FO1cbge9iI4pT7HhF98TdqbPPNXhu+OW14g5aYrmcOFyE
g7ppf85tfCEAD3ZmTV3xw9DwgfoIPkM1sDfyicuIpo7vcTrLzg3X9XuQdqnBnl3K
syQkQVXPgcQfGczKs5Oqy012Xd/ruB+hflBlznXcFpoca8AbcW3rVV4bOFlAdE5J
Xfyv64kOpd5Vv8bmgTUmfY7Zq+zfq/Wbt/I4sDdiT/UWlZ3VJXxP4r/P8tVr7q6e
Auu3EMYRgjHqzk606rvEoVEBfmoJopVbxji6Lu6GYrOlADqiuRIpPtmLadVw27G1
8OjPFSpfc2X2GI8S9LTRViyB3bxn2JEAsbyGJKDIDB/ClKilRarR0dX3L7jXyWPc
xfmgAb1FS1gOz/J2ECzJmlkOWAVqNxMpFrY+JBUriFCXmpmmJVNvgaT+haJg1GPv
coUROaIcydyg8/Z+44MKpFv/fs79p9Onl0eXfzZqYNjopTqjBLG0LklFcA8H6yRs
79oDRQ2L3UCcAmPdiCeCx2kUGELSC/hG2Ej1VR59JNVmo8PAfuLkESxbv5184O65
ZfHDfNBACH3SSMw2Sj/9jCAhqAoxJWeyDFjgW9CKxK9jS8Stv+yLggH6mhuYFufY
hk1EQnx3B/9sb3P04itIUdoLsLCYvu48ttilUdZdI0HWfkPB5l3nnaoAQQWHFNNN
uNBD88Qyc3S+gjrbqxRT7DCZ4mrrjSJILhJSYtm8yz0Na/qGYovyh9WpD3R8shbW
8Wz+Bx7epHFvCFJsKhCP01lS+M46v32rIwunoBuhLs2bYqQBtL+aYWjmrKW70INP
KQB0rDnfI4s8CBOSP2JS6IOjLa5csYFuOtTv0o3Xju5R3CmOj+bEpakEhSZQ12h5
W8LBeM3VmdOplsRnum8VgJdwhB6AUYsbOHkb+xcQ2mJZnVtgc4GUPi5c49V1/J2I
C1bxbCeMPhF2mwfzFFOixmt8Z8l7dJV7ZbEW46vTVHVQkrqfM7fUgCq4cAGG7skj
5F5AA8+PLb4r3BoXtzI62TX0g+qyqaNlamuECMoxfqswXrgtRD/PwoYEP83+VCJn
vAd9KeqMM06DUrQWs9qxF0BB8IUVNyuuI4LnPqJZa477HJcb71/Jh37VKvWOkceZ
NYJsQuFZWh54Mp4gqOwL4jucfOUGQiupPBigMst/1ZE4MyBBU+PHbx4U11YjVWvB
F9z3mVsxPirZ4n2e1MyTdjah4Q2C+FUJwfBzEcC92+DTW8tw0+3H0a39NvFXS3e/
ebI/ganc0P5OqGiq6fNaoC/dJcrJtuqiN0sw/UeVP+DgpY5upSrmRcAJpc5kc6yE
TscM4CQ3mwFLYZfeuICo/m55H/d4FKeKOHvroOWF+z6esSWW5sQKTFPphGMQFJsM
+US68gzEfBNejh5keXt/5M0sGcJvYISyZUEmStZOfBmsIFHT8EZYgt+S3aw+fbsm
fIPXcX/5I+kHbVMxLybSU3iK1AR2EjAMgcswxWqQoYHtGWJxqo73RiI9YA4Aqryr
UiFlVLNCa/nc6GBljhCS7XYbGfCjRYS9DNp20VuTJwa1lgJ9vPcaIkz5y+sKqSBs
hChYix7LMeEAIHVpW9qYxrUoo155YdxIun4V4NLaE8t//huxg/R83z49ozMZKKCV
m+ZGGBk2fJSx9O2QaDZnX8coMCn6WpxnzortNNL+j0AhSRnRzYykv6cvPP8CkDHU
h4KpWKCT6PZS23jiqK5+bRBTSNKP+ercdccECl+LFBGu6g+gQKQLN3wTrF4vIyLP
XRO4IS/aYU4teZaMfC5mmd2F3i0ATPQ/WIHvWAsDkzKzexneFunUGLkwJzQhNE0S
wm8Fg8uhyjEKnScD1sXuug8/hGbdi066EgG8FeMCYULboTYUgGNvi5EaqJROet9K
qxwQW9fkpGkVgpqbJ5XZtNG5GJ78IcQoY5rn0DEaUkmMpf/jw9RlvZS9JrFJm8K2
vmshkkedzlxvYWdQChSn07WeGztcY6ec5bwlzjo1976SZUq4r2Wfunmz/+IIYQuo
kwxuLBCtEsUNJQGFN3gN+xqMqp4N5bOKyxqqsC+bYyl/GKXBwN6r4vmCYvzIMaUD
2EShZvFlxSusO9ddTphS8bZ//Z+HGxlW8jIUjIzE4NaKvxnHnIwbAklrn+PlrYKT
UQn6zLBGJMb0hnZQGtATISfxRT+mXwtg8FO02Lc3ku71KFZS6vlNoD1dJvMHtfhB
jl7yWm7NdB1XQPUM8+OQRxQLsTUttz8Xe1Gv6NUPgQ+kjKVzA4/syjHtW10cvo1x
Wf+Ne4UAK7CdolIg0dlfHzulgdXK1cMJ1r6val55wTEeIWXbHM/N+q0HFtASUPun
XVW9J2Wk0rtGf2g4uqnIS4VFk00Dj2cIge8h6pflEPrr0IFkz0cP72sMBhiB9lxl
Dl5vsxcvj27shKAGCh912Lp76NrZtrf3xt9xVCt+Uu4RSgc4V1qc+P3y6hnJ5Fcw
cqoFBZN4BqoYxQ6cngdDvUU/eFlK+1ESmc3TZ6zsGSRbEJaRrWdq0VkwTVy26TXJ
QIN5e+qRp/qsPVbHXMcQyzoGXiFrDTtT+YBh+W5KoAFkIfhu325JnhRwXRcTwXDk
FjWdOe2vB/U35zRkNhxBwXHkNcMAvSc4QeLntIdhCazv4ji4QifaMXh1q5FBgmKE
49P63tW4RsOO+avIPwYudl2Oz2SyAKjrCOadvv6N3CywIKRbYBBuGpUk2W91MOYh
X/Q8GQUyuUmORy+JGp/3D86WLBpkwFHvkYabsKON+L/QXgAnJ8d33ZucQXStmZov
fhfGmkgHkq8GQnkMY/NQoGsUr0KkCSOOWZ3gRCKymYG24Ht1o0Pg541FKcUwpivc
3vClgcFKDNgscGKfQkZNUGAqf5CCYgxETaKhO+uD8zd7dDweztonQHwKQJRbu8Xk
aKIDoenaaIs/rPZvLhHjKFRP5hCq4kP1LbWO3ju5TkRAkBmI+HCerUO2EJaa0oK9
pnhqjFvNmL1zNnKmR4amolCAL3m1KNo5wnDm0xD9RWVrdFsXRzsYtLlgetqN0GV6
cC+ZbxnVkTXKM1x9fyBlP774XCBZ9scK4vf1GjRgDXVq3/BLmO0q7YsVNlwoJCcN
5J5C2UcV546+DTZDW1olY/P//6KseQvw7U8Mb0x+6O3beDHHRgvPS2NPRbzg/ZCv
X3mEZGohEfGpYBN8oOXgVN301RlK+5ibat51fEJ2hMotEUfcBgHS1eE9VoJG8yYb
LwUlu/w74uI0KkBXMZZbu29nv96L0AhEnSskGV0pWoPDEpF8w1kjH0FLb03E0gm7
YUu8EUwejTNJ/buLsjN10GSRM1XbIgUxAYTVfdAHpRclKZBiYPyt+NubGpfB5vBB
Ito2KoyM+O5HAk63Si44Gga7ryS1hBXE1KPsQ4H73U/nuYr5MqLwuD7mTS63xAI2
gGt542vI0iByaVCCNh24Jlmq57Lz6Sy2jNDfpnpVJQl0pEp2RuP9TDkBzP8YMIvU
WzWdkc8b6k1spXj91/BLHiWQZEBe4ls9uXWwJWwD7DiSVa+2ncj2MUun4pCgxAWT
0tNqkklx6/vASttve8wTINz3py4w44F/7C+aWe0GHi5bPO6dGwbZwE0yQKcFOPe4
xznfb2EaHQy350dSgEI4wmxAuKclcy3VOE4KzOe+ftKWPvFBPCb7by4HJsKXgPhP
sNdHIztDw+T/0A7ABNTCPr9i+VAMz2Ja08nduLL3RBZo2k81Vlfuy9m8Q2jIsowo
i+Kj9MV7wX1C4SNQ1RGeG3GXnIpcRYeW5WHbd70xxxqIAkWm59MS1k6GcTAWes2i
DOSVj75ZFjgm+wWRyXvncdpWHPpXQJ7A9BQIFjWFXk0TDpFQb0oEB4kfIqFQK5sC
VQNJXRZVHHdq7cqEvhRiYbmy5TYp9LqMGG9TpvuSABxbz8vW6Ng2ow65UJLDd20P
NuI9IRHdUm8hFOjf0ZNoVKrfHN7V1f66DluLiKLPobMrEhd2fprdkfYivtK14ckU
qc3O8sK25ZOnGA7SU5YhFZHYxsmEiCCpXXMd4yd+SAjjsr+w0QWTiL5P9byqHgSR
gGNkMzPYUCGye9zVDdM2CCHW6vLs132FJ1HhrEbBrTdo6hybVjRurp9mrOgchaJy
2ua6xMKLXh4t6MK7FTj2v/QzWaa6vLQII9sE0/Me9FHNVSyAWH5EJZLv+rVjEeB6
GUUMQJ07El/BQd5ZPeIWA/OXjQrp1S9B3WUY7KE+KKqCcWW6kB7An27W6C5Oc8mI
C/lUdamq+KJYbzumfUYW7apFVr9JLs2jF7L2pCAPqGcBlL2eg4GljYmeQAteyM+1
JS35f3RGOKWtuXjG8S7WVdWDglUC6m1bN0YARcXt8iIJIBK63ddbxoPVJlMmLro4
7kxoU4EB9vh+EIQpQtoBlj6VqbfHoesYI1OQ9zeyDfTBG8lJp5IRSnNQMTK/C1mE
rRtD4d0RZPSqVRglR7VkMvUeh1xECKes81OBDm0PqkHHdcNYPZNCDbSiHJ5lXoG0
8CDucmY0z0UjIUtBwBqSCmHkh8pkH+wECwnZqL1ZIQWpumfUO+dOFVqxgFZ+ePgx
6na5hVNCuEClDozdMy1gU9hPUbmMv9RjL6mFXYBEzNo1pjTmDOZolrygzZ5OS8SG
HUOzVABEWnmlkvt1ZmCDzRuYdgjRvJlerMHs+3P2bhLz3NZMtiEuze+Xi/c4CHz9
krMY5YMMe59s5nV5PoZL4oHncssRQhYF8Jex5aiUsDABkOlT5VO7kaXtuJY3t70o
bQ66v2FGGfFAQ8Cu4gnrlzxgn+iIYoy4Ui0UCPQrBWeDpPFNf2pD8v2ZQW1fdVcR
FUb5oXNs0arDYCNiZ4BHikxfu+thxvU3SQn4cs4b7OolStV3I8/wScGmifSgwmgt
0vMu4bTUmh7xMLV9Ohvtn0y5NgbHY5uUDVe0blwcyBHVQ7ubkemE0EKFrIZMNooM
yTnDRQKYp+nAWvB4g6VU2binPR/+k3jcB1QTf3iSsNg1N7uwkhRDdNXyYt/2IguS
Onta/yhzhgkLijejob/1KD6RLN81GnrC7WiqxvTtqa01pFBd4s1LkQPogE/JqEzg
00iwcbxIjJjtac8QcufN0jHeFQlfiTSGOR79++r11Q1YjYcEkUyQZXh1p5pUCvck
qsLa9S3bYBt6BuCUA19t6f1XUMPGlcI6cNzmn3sj0FPdtZxnhP4qJOAwIxnG3Eb4
7FT4/LsBWxhMnZC4MlZGs7lBPXpooUpxydX3r7zsvmtKy8s9HxGxw2U+C9MBMfZn
3dxKvll8NOKvhs3YXTZ8FQCHVupsuUKKVV3TKW7tJTGhn8qn9WxEQLbPdwNWrMd8
ZcJJ8FiT09DCvsVZuqhzXSs4F0fxpORoh/8MXepzSZ1xjpviLi/qBxMHElJ6sx8A
s4m9jsPD0ZFjkozZG1FA6O4ZHar2c//IRKPC+Gmfnds5dJeifaihfwb37x2CCb3J
8j8T+jWH0E65ge9osQ68ntuyV6vcKQhXuENPS0iox2mBguAW4xtH1LRl170cuvJ+
C7r5dgaiHojvwHPQckluXYRiedANpVXSF/8Wq0EKCSHYar3bfMLvxuOLPYnUuX77
9GnEi043QN/Pmie+bKnnZe0viDvPT1CmilMHoZCV4RfzZlt+2TNZgvdHqaA0/Bch
X8QzYFh//tz0tE7NdYfZydnuOP3CVt+h4Zf7SGdp8XlmfbuCLlOeb2Pgc83zmOBD
/kqPx4iORgQIJIXOD0cz2wXncrJI6BhUtu1X9E1ZLqdYkHJxFFaOHIpMxkQTnYlB
8svFE9k0RPVhKeN2appDXDreAlWfjXOLlmwmOqj8QmfkC6eSIlGuzJclbMzAR1uL
HJuf+cE97KsRtp7e2oyXIU6nT5nTQrtsdq9WxPNvvVwO9uH8Mvkl5WNkx1KzxfCE
vRph/7vOFO43F20LdZC8d052OQ/Kg8l5o9e+ppyy5tkXrme8kRPgqNBBU/FthEFE
XSZ10uF8UYUggTbJFbQUoEgI9W7dDMPS1Oi3XiUPM11sEK9kh8cCTPsjW2LQaYPh
gLidS4RCM8A8k6hX9vhl2T/XYbjEAUf7ros8Fjmh/P3KQxBOa4dwYEvaf6mAdhyw
br0XdXAhN1qyRrNWoMgDOafIFYG+fPxfDG6USzQDhVFe+L45/w5z6DgvTjei9rO9
w5VktGwd8p6kGwdBkbrLEjLGgi2SX8P6lhTsqe2yVCIjlUD48Yxnf09ZvfTg8WG7
d5mvunjLLkroG1JqjSwo3VFG3HHq3+TJ4QVgMZWARpNgGOHBnP8Zk5l0K1pqI3xR
emxdcLzrU4kcONiGZid17E0Jg5OjQQGxvjQUSoDbUN66TQSrz1CCj3qknsmW4iWe
hxiyS7xuKQ7HHRpWVEkZ23nH98WJkHfO1bRrgOamqlGv1mX+m2WAAskqBGHFORHw
R5KNlzdL3uKpyGej/YRU9ox9b0hmVBDL1+t9xePNLTdgDxVLacF/AssCb9vOFykx
b9tVSZYUDDGtVEZnp1z4AXmDTFpmCpGcL68/w8psU3+gc6kxJVrUEBBjudnDw9zI
fr6ITVn5zquFP0JFN7D8OugdWO+Ku0iYP2SAUOsgwFCV3nnkh4FsjNwvcaioJKw4
SLrUbNQa8QxsWSTO6ZyJilNmXXxz5tO21LDJ7RBuVlmRPJlvrNa7Eu/tQcUlT7/o
aHIPV2Qb41QUzBR47QGKvLYjjTJghdM1skco/8HPRsHLS8ecyYM2m7gWzm9Rhsgf
vWknKKrZkn8ras5Y41yTZTwW0Z6whOPLGVbdawattJfSNjZJfAuZcWqGThLEuJZx
fP/h6LNOOqX4XiAvdVo7ii6/4a1QA3pTfGALlFNnG0CAhdfo9mS2dDsIwtWLSFoa
HgBa4EdmBKNV2HnaoXOcG2wzspu8zM0cB3PWWzPYVR/nNPz0G38/uExXQhM2R351
zf3brEqsiK26H+lDy9PjNIC/RdYR8F2zcF08yfWqYZOBpxLDax7NZ16TqMUojW6c
yMyVvPXeY5OPew32dvPc8veiMtNbwaA9SBJ4eFU5uI8JUoCIXhU5obr56bD1x1Dg
7u0ZoT0aoVTMf4BO+PPy+x3T6aTPyATjqELGG4wYxCetzR0v25+JnsF2ohU+ZkBq
3SqW3IJPV6Wm6xRdznrx6bTnKr4E8Rr2vBaX9lUisDvM13FXhlr4RE5Tlz/iQ0m1
mVXrqN5on1vs+dTB08MRVmfv2Y7pL/VUNpFv1wXpuNolGtS1NZWStlD4cL460wKZ
sPSf3d19uxkjtGN8dHcc0qICs2FO1OQLX5LGZYnBjnjtFTVbEiLpIU1UJmMDdgGg
zW9fA6WUHD+d4/3oZF/ODIkT0NLvP4MkmUEPyzO29ubJlNZGHXNjY1Sj2j4mjvyJ
eA2SY2/ZPjofVSefEv0qCYpcEojsgRdgnFjD7M7M/kReopHp1uthj8p7yGcN4AoN
Uablc6KqpGn00XgtZdjIw/fezGnE2LAk98IiqrfTz1PYXS6SYgDpS1yPSBR0RoVs
F+HJuZzNR1YwVeIeC+Ge/AhUxvpLQxL3x89YaiHpD8gGXs2xeKIT5+EPaKiGtGcV
+DzlQQnh9/xMg5LOI0OapuRt18/X0z+nL9wNiiaY9fOrORtKc3MQ0WBIb3v40jsu
40h72hVsRx610AyUz6k+ATSYlVsZtbegNkTMqJiibIxhsa/EPZ9wUWQ4QSkUhHNc
phoAb3yHb3S2vb0dW0k4trXt/lokBWcKS5g/ctvMGyuP9hVEf+jfg3v50TOi7NUE
8bw8PcvOV3VcvRbruAXKAJQEno/uGSpQWWS7iH3+ZuYB3+E45hmPiLBzmwej/vrF
ZO52w9DwNozrlh6J/mhFux9mLHAq+5u72XN4bWHqFHwac4RheDnLUXA4PwPxFw/O
t5wvS2PnbPJBbHGLkiDOj+uGRQQYIG+WNfmESsyHLUEPxML4SkOa4Y+/qGZ9hJY0
C45dHPaTDVUyMSb+PjJoE90ZwISTKDhdCCAzyYDXyxsCBBOjPKce2YpQZMBmsC9x
shTh1LZ3khs+gDfDDXhdHDG1NeYcuXP0Dec2vSkKO5azD4URFsBMrA4rJ1M0HySz
bYUGvssPf78464BxJ31SwyV7inRRLdlCEYayuQNiCiIPD5BEbfSXYXe7OuTfqMiP
ntZLdxJD5A6g5iPiqTYHxtMpnegfZCRF/pASl5lCL+q3bJ5Wob1ZEaSC20LxbOgy
p/Ate0TmRFu2vebrSutgHx4rF0lRLdVRiNU/VO/DMBpIAEJdRhK5WqLU6FVI8Zh8
tU3+lgyyVqxomxD3nJtPWUAYyqlyl5JtNz5XMDJRpeDbEFwGvkkx6L/52rMoULBI
WeZEv6GJ7bOqhEgnf5l0+dXmoDTXUawDZ27QxiBVkVBSaVGExSBP4XlRqHOUeXyX
Am4Gcp5zK33Gw3P4l8EzwbZTTFTr7Jdf+1UBvNDtwxxebWRCX44u97RNYG/ghcHU
D+OsCMnhwkFjiEdCFO70P6mc6BGpT1RZV4mKVKPMUB49hIuyT1NpZv4Ie3+REfxm
lvPR47NF3tuw7H1+2EXuSxcOlM3X3+t/w+iI0O5CosrfPfTRaPKy5+bgcf+kp9Dn
Aj+9DRumXdx1GaY+AoTOYqz9pHc+3SpK4kfelrsR8YE4vPz5u60RBhjGzqZlUOH7
4j4fsKcKAoCEKf9uhA/iryg7GA/Tf8Rx1T6zO3GazCjv977oSjhEgZEP54Jl61Iq
+xN6cqecaczB4/3fkCUz+Je+W392JasMErrMwaZ6KWFdNvlhdo2xzXwNbQhOJ3qU
wj4+gmx0wBNNZEYUswdj7GvdqJOKY3+kD6PK2bzMlEjoEzZzpqGWH7qZhOZ7a5b4
Hu2dTlRNfkbVCZPfVjFZZeWpwVbel6ghHWfUO+vISCpkEB50by4aD+oAtFBefXmP
qmwvJURLQbwcZB5/0Ao+CjINNvM8KOLUdaiVVfHF+q4E2ZqbNijwKM7myx5nTCp9
muNTDN6HHwfN0avNN5HBQtFG34WDES+CgjtGDs1pPliArw7U/Mp5fbagtlHhqom9
Ao8swdtSh9mC53MTOS5q3TL/Yu6mcZdbGnbgZPUT9mzG3T7P167DiscAC9yc2t0j
lFaK0o49/IWJzJCGNz7xWQPD7Vo0TeK2kUFSIYqC3P5BKhsGi+/wG2Mz5p8UwZGp
fCDnbtta3Q2Ss6oadHKz+DznOzS57ywaOaY2Y695/Rl2Qh3CKww3iKUlgGBdC/Jr
QMosq2EXslBeC3nLscSC5bTvaIlIHcQzcIHtjkKAI7MCqpoyTri93agVPMVtDrWv
am7Bv2cfz69gnSwRJP+m2G79shvPtd8iIs6HcT7vRLtUkfGK4a/LA0yy4gaebNyJ
T4Vs9H1VTRWnkre2cK6k5V7MAq3VvCIN0F8jMNjfdYZSMZ6t+LlgKp4dIk6CIjRz
BrWZ4oxFbv4mE8vfe8F1fJvMrFkm9K2mCcEw7oHzHOX+OpSDh4mrK7poSqbU8scb
fdG0i2B/GcNHwpgvhOh1n5hfwW0o4jU6YRh5xhjtbBftjvcrw3aysQd4DlduBwjk
vSPfch9T+szZOrdp/sX7FkWtatV5TJmC/1qceRBVIeoq+3cwzLBZOZ19yG7TA0qY
gT5740GXPFW0tnS9OXmycuDkHxhjcYkVzpw02GIUIlEVjYV+ZGnGL689cTmbuwTI
4JxrHDgFmd4yOBZNUjuwBLmiTNEy+fMGUJXX+u/meZGHalX9z1v13zJOWgcB4Wh7
qBHpaqmHbaRplv5OJ3OjKxLlCeVm0tqvHIUofdk11Zo8V35qjW7DL/ZgssqSCeuB
6y79Tr7W1T9f9t4Qq8Ip8LS3eebxNZZd1lLajLvSSmnXoIjqelUFAENyFreplXv2
SMEArTxHMtZGl+8hsUOmHSIj9X/dI+WryWnH8267P+0Ch4OC2TBaJ9MhOYCd3sON
x320ZdDb9xFnv9HobIsPVcIe4ocM2bSvSlVi8L02C4ygCcbz4qkdIbA0yL+6NaJM
wdiYJ38h7Et2NxV071cmacwAODtHC5ynfE5hK22eeL6CrD8TcNLiQsagC3LTGF3a
RAUv6GBgYP931RjHcf48sSpnoHksXqiz7EuOtnQcN6fZRb4PUaqHuE7pgx2KDfp7
9E1Syh1pd7XoU30ZNTf4XdV98EVInYEv9iZo/RuOC0tjQyE/0HD0qBxtoUgXWXMs
jG1vEcNNL9t/pIfI9eE7gG2MEk416A0iLnGiLc4XpHINOXNGxgB6SZIU+2x76iUQ
lvN5mx6i+u5Ch9GU/XVr7o20SjVMoUi+Uq9mEcOcZh3/AlE6zpIbhGmIcGw1rH3V
ngXMsx9hby0sVQiTJET+Q6QxVXShRJLwyVtQbCW42Zfkctz/yL+YyrT1/Pc4dKqh
275mDxqpAa1QeiX8k2Uk8FzNF8ufBpoj4id97UZJt+bJPpQk8LXNtNa1TA1r3/fW
bYcBKdxsh826N0TzTf+bD/AaVpVf5B+LMkLAQBEvm/cxejubM55ElHShRXo4M8Il
KEhlwwOztuY32gmZ6Z99LmLLsYd2ghssx9gke6npv1JU/9NCVi5KbWNVtYxedFAn
QVzWJjieBjFoNEqsOft9GDbTQQMBPJUgtZSeZR7rgksG/k5uihWtrG/k5FL33XH7
ixL/VDMqyUY7RNdTAC7S/hVtTJwr2t4+Fb4DWmgLfHpYFVy37G2p+pp3aS/8TRTn
I857Vqi0euCpjZwSRnmi2aDM++oTFGWQr7hAaVC1V/vkVEUuy0pFvdIpNFJbcbST
AWPCGKm6HXYWEAlQncWGDIZ+6dsbivYTFJ/h8TQy3bclk0UweP8OhmvNa7AeCBK2
r1MRlAjFARdJ1qXOtUcM4GiqOtCzE5CD9ppflwhpPHO5Z+4RiiyqrMBwJBIk5cd9
zwAtAtYvYheMb3AO2NUuuu4OZV9Io12hObHu1rRrWpWFXhIo34MwFadMcKr3ZIdF
Urs0+ZW9ttwP7HdXD0P1+JFSgBfRm/SyeFlxuOtLbT2Xw91d4oV1Fa32+0lFATvk
IKIuc8LhLJ1ybbZBPykxbqBbR5m/cLapk8WkJzLhkplpTfWlWCeSme8yEZSVL3AU
YkmLJNFT6iMLwDmjOgmF2WWhyVjPI2ADr3nJFolmXxIYT+oKCGzTPDPp3zcN+ZX/
pO0f+zDhBwkzswOJh+A69aUNHZuVlt5hJhvR0hVqXqTSdKCv6Ev8jLL4t0CInWnr
dr5zz/50P+KB4PAjYzDvf3ThnllEyIRBm96uG0gP8b7ZYsPSBfEmsNcYsOJBvyG1
5fNfz9wR5E3SNElC758RF/R5sAfIT3LrYR0a0rGKxbZJUs2l6ZPVJ43AnUV3lLrI
RC8RCELeS0N+G30S2Km4iEV0iIQzkAEXBSXmnvSJPhoYHpfb7xjfqDx2LgcRkuHV
Q1kik0IyIPcQtHLFGGEpxgY0lrpWE6PdZuGe80FKxa4Zx7wwwZLI+hrNlLUAd8t+
/TKsw4oGPwbOlskMEY873E1n0ZWBUgVdwUcwXBV0I0alue5Qz5/+/xh9bZZHSelY
WHISDUAHKEHqlCcIyEQIuDsOMs86aDYGmoytOFkF/O358zJ3pxNBeZNtSmTpRmWC
K+0qnFYSDvyycYkrNQb6qqvNFILmqHHeE2wfca7fFypme3C2wsaYeRNnGRYLDwBb
XOHc1QTAQ4cpwG1JaoX3rtDEXxZ5rGol8XpDEBcCgE/eZnUcgnXlEjnLMx/iGjVv
C72BbZDKgHbG7CmPB/HRLEoAGQ8RxRTkfsA0kMYBV4sLvFBKhEKtOcvPXO4UyFsV
OT6Wu/2HRzajWxXtkj4aNCaCjY/NaAYWBEdQIDIEduu/z8IiUY7Y849zSWlhkIg2
FMG9HuwLXhwJjE+GsHKv7IFv8Spd/NhFKvaBfsgFFy4WmY1gzKw33JB+eNnfPQlL
MRxHC6r8+WPs+65t9rPSnFU6prIX/nRgyQp3/kcHlUXh7SFcOfipxE3eobcETCXy
YGDxbuuux+Ax4J1MZXFz3ODeTKDsxnHdi6TdtwA3zW14Lb7hfMRPKDoQe+meKVN7
TLNYDkcW7RGMj+oVx0+al28YTDU6KM+SydeXrKfMEjK94IySsi6/jJvaVX7jJqHt
vwfBseQzS/5CtG4LKUUxDF66/gvKHpzR5AT+bLSC1BCuCzQ+kkrTM6G0PYEaESCI
HD9ol+ipQVH26dhl8hEN28zQF3x5v3GQWaAnX764rCNy9sD/DgDgWqhDKqI1RDnX
sU9LIm1l0h0O2Id0zsFhOYqs5WkjvYgvi5UZ/ndJFagSRtFC8J8MkwW/2UI1VBuY
qAqV/L4yVyLVb91Hqq3or8r3mAvTocsUvGwWZAC9PcgHaybIToU8og3xgA4xjaUl
ZMhgRrIsJ1Ab7Z/deTxcamDk4zUv6Ob/uafya49sV1SvkGOHiMEXkekY+gLBsP1d
j8jNXnG0ZXTIX1JHmSOdadEUdYxTBsu578JGa51GZKdUEq7uGJRGwizcz8QSWCNi
ZVEzabPaSG8PNgI6ACdkP2U4HNPyOjqj/Lzhd8+2n5pQ4KLPeG+hF1jeQ9mBEKfc
Y1x0I5ebmk3PKL2e3BLd3h39KYfOUd03buvqq3j2ZND1r9PmwJPojM2IxXNzwFKc
DwdL8fWFzxTIjHi5N551gAm21oD8ux2a6ylZpuT9gK+HUrezl73yirZ2GM3sjyBG
TGfvUVZJxqHmG1LY2DrBF43ujxvHx0GA/2J7OddOc4NDFjyf62RLPZuGFT5Cd2t9
h2MDZB/wJlHYEFvp/0SuXOyf6m7cnK8F46JfiBC/yF8+5HEy5CxkBGxQF4jVB4al
SK1chdi/f4iyLdq9N53Gek6C2M+KQcV4+iCui76ReVC3MFvxnXBbnCwkDWu3V4SJ
qZCuuNlYrUuyaHRWyL6yoOnPQVcUKZqDb2PWq6DadNZAH5dx1cGhDTf/wtFAs5wx
5XQa6cGqZbsFt3dWNTR+t1FRyRwHg4mlVqC31t5gNO9Wrm6r0S+vMpiCiKlD6aWK
xNXBBUmAkGfr6OSaM8hJo1h+fi6u7NAYnykxmSR7e7L/dDEwOd+1VMPfsVOoumIX
eOI1iH0Dr1SCZOWHQ/6blUbo1ri/EgaxiO6qTRJdofK2lY1ZICQfPggAoGx5Nx6S
T0NqBeAKeQAGGVto3B6fDxq44GLGXUSmeOC5fS7MoiLS4FlrOXODtlHhMdBaKYRI
zy96gT8jYVUEc6Bd9sTrujm7uZ9Csg4+/u0mgDVbQ7JVVDf9PY897FsgT60vv2vi
vbEhW/6e52TR7B1BrFg6jVaLjmzyUI0hU++5bS8CRK9b8s6wUWB5VpS41x+7MIwK
Fg4qmymD4kS5q1gCn4yMd0MseWWYeMWIt7WSyGli2XLTHXlyqkNgjmd5L/ayUMvN
k6shGqL44xDyktl8RsUZ5Ig7T3n4a2I9KBZO+YmJDRPxGrHEmc0GY6GeQp697W64
ZX8yQ2vaLZ7rFpyRF5GI1St+K1Y39gLUd7401H9DMZq4BdHCSX3MGkh18tUMeXA1
8pXCysNLjDuKzOBPqkS4w1/5Lktf+ebumn5OuJu7/xxJCZpqmUwr497K+AXknsmm
YOxkZld8f1LhxQRiABldYcsTxRKjNmpHMLo4xqHBUegNtxCJBnHhLVUQgMYi9bgr
b3l/YqY+TK0FaixLWeGHd0YzIedkpCJCMpfVH4WyLLge0vqHDKfb2Z9qluyZ/P1j
4Y5rHp5IN9B3ThrhQAXuzr/J3nB7LixGb4MrVslAkKeScKuUECbqufxYRygyMO1U
69byNPAb99fYyp9D8c25mXZap+JcLJ1wON3mAOga/ZBniaabEuCP0HXAiHxz1jPZ
0MYcquyNld75J3bvBgpFM1awmNjhY21A4Jle/5F7onjJ0wQdHMHsDCVsKaUBhXyG
lpN0AIxDaAQxtxQxmfVRm+3wjKJ+ENcu6SIHWTL1r9EfpZbEyWrlJccPPWzuzXMa
OYbPAjU7bBLTJXSJCugEODhQFb2jTFB8q9G6w6p0lQ4EBMqNufa0h5wzpmiMp64T
UoIqLamIzlAuIvtFpzCCAujKt+8Pf8sy27tmiBh9rK8gQv7o20GP8H4ETTJL3+ek
M2yYbOEnxXaBU9OpK26yDnNu0eGEGJQphjS2PLSxKt7CkqDqxNWsvdJMXWHvrom1
nQ/dadr3FwDbuDXrJWYiQk7+qLZ24jD4qoArPsORhXPbGb1lwAkj/Togm+rekonF
g6kpy+jMc4EOeIO8tb/bajE3CuIM2eIWHEVclXP8ZVkeCv6YGfOSoe6fc/xYpBBW
b0WZY0WJPoiVuxqv/3LZmbqG1GDA2Ut5uO6gGneXoe044/veRMpqn0WOn6+NP0v+
Jef1VBbNS4RRo+gbjrdNBy1BEjRBwQ3ezp90D+FdIkNROjRewdnN/808mVLJ7MSq
ysRxeAYohRB0FgdvQGXnUgpgsZ1PhheSVLw15F7YJEXKbE/8KqzLeTMmPEKnQiys
9RWJrFPN+pKyw49IrjFUlDIytGYBMXsy6U4jqFgs16Kx3CSYyjgbCrQplQ8nJSPr
S5euqDExM4+Z1gefjnp/pLcZ6Yc53lQyZwE4r+3rjhyarfTgnbkrKiRDy3h6yhVQ
DMmVmKHmFugMm+hDY4PX0AHW5dzn3xtYstUjnVep7g0/BxEETRjg1W1iYT5imtiX
2/abgxBlB6FdVdUHlhkQKrgxl1rKQPJalqq3l+H8DFENsclELZ0W0GZly46/6N4Y
OZ+HptqWbZet0TIVOiF8tqoDqzxi66L58PrxU5ezAZS/LzqqK/6zFy4SZ9xYNpuX
2srwY3poXSXAKvylvDsrziS7UWzTn0LL4YDsM4sORUuWz4WvQEhu4W1VaP+pjKF+
bcmsVCsJQONLfghnuMMknXl/XAX5gpYoe2EnSBAlRWL5pAGBL7A2rI5KWacIa89d
RvjWgLaYSewHZyJ8fDs7zo2ENgAX5XOnOgm2gvtI+NzqN37K6cA8n4d5gL53FfAQ
AqLdh0Bf1UBh0dqKj+o28787CLRaXzud6ppSl9+i+n9KArftk5fWwB/W4lBvYPKF
9Jva9RSS7hxPuC7tFoyppHtPHMhiBEYMmF7SRl7A5KLwhmxtpAfKr4Qys0q+nOoy
nUx7gurk6WUGscXT9vWa+nbHk2qrz+RgUmkWDbLaQVyPyGvPpmDyAapuLjo60y8N
QtdMMvOPiA+ZkE9q2IhPJI2rn4OsLcO3nvDqSL7DCJXIyBskahNFgXmfr+P7w3mi
+REatHA9SyToBnfqr6sJ8/Pt4bPqBmzQCO2yN7ruuaoahJmWao3KLhKb+CYs2ZSE
KChVTonuG1gYEWqdjUgychAX7rRqVxh2Ek+LiHfu2soDzLGJ9/rBziXMClszwNMO
UumsAWwdgK1G5OkafCBAmkpsqCxaY4XfYgwch52GRyqRSyjcjTGgcb2zQ6sUjw5c
UBvrVxCijFJXNg8KMlJwg9M7dcuuW1G1c31bdlOA8djdgEgKjYSduaSaW2Hu/h9F
3pG0HKNqmodH+O1NjhzoVc7GCMBpvXN4GGSqTrRLnpFAy8oR044KYwSorM7YcwG6
CSBpM90tVFfC1M7Gvb3Uh3kdruZ/1tQk+PFcuNKnwLdb8C2Ndc3sfX+W+OttxtOg
4InEIRVI3eHGbgLc8gakZid5vq8MAqHE2oYQ/8psW4sW0LUd8OEp0wgg0hAE4dGj
VEe9pUMfzbRQKTrxWXdL1ZtSCi9guQ/ybF68QkylmY2SceXI2uKNo9jPTFFQkvNn
t/QSQWWw/6J2DoZlEy2mT9lhLKbTOfrhpUvMx4cW6fuQdP7MhVnQP4AucntEFaBe
MiqjOm8HRC8wXjFLWZkEtoMlvsi2JNMutKl1f1cmIQ3FK96uyiYbRuZjLbz+b9aC
ZHfHqymusBG0eUs7SwashvZngkuvTKv2V/pSo7aFVarL87f+xTpPSoK4TVU2U8SW
+zsRANl3rc9Dn3wybPimJYUjsl6JCKxORM6mizPE0WvlKdeMPuu0XlH0GULmacSZ
2QJ6732v7ZqacXExVolTsXnFFWP0JKM7BsLnQaWuHuymACqh0hauHkkHgzgk8gNU
2urbXxpwLYxGrsTGzhVJxfqQTa2788M4B0iHILAPySKF+DWJoU4NRaOaRK/Vwcvp
nHGHg60byeuAIwCi9mxvGZticbrEBWLQO0RXA23WGBiW1rtNYFp7ap5Mz1fJqZ1j
myP2/gJKDd7k2q7/kgKBeFVBpKomVNfEmBL9jZvTl66UCvy41XApdYd68SN4ExTX
Rjz/uSdjcKniK+jRUnly338kEtU4dlNqBW1q9yOm2NmlGS3LrnWJfCcjjlm4AKXW
0jugIXTjhhT5CmNhnkAMfnOz0KZb1lRlYoCFdh9si6rTiaYjNIYzVlzg90PFpBLr
QDNUWDfHOQjHkU6KRpgYzZ9uHBJyKuVb3SLtRlpBVepbmfE8tr/Qof56eTI2F3lf
v29pb0zplwQv9nBXuV2CihZMQ4mw95Z31ymvLaZvYm8M5bhllV07noR3h/bPnXBR
PpsjE8/kheeNjsjjXNIDc/q37g0VMrNKQYqytL3G01BjSBe14M3n7JMo6w6nEIMf
Fk4l4slBPiFh6l8Im7RrjjlUmHysWgWv1dQFbQiA6i6kIQJ/GTZrWcnBfLdKOKYh
+579HecTU0HdvELmaXedigvOFidHTpYrszl7wBiSqurTronVhAa0eoZ6vOwuPRtw
DRXbHviHmLfVttDrWAvwl4+BdDkFdU7We0s4lHwfFnjOGBcsHOg3/MKSCG6tF044
tPXrZj61IM5tL2t4RdCjYEcS5s9F17l7Ge8mY85+xGRZX9OmBiYED3v2zzTmvdj+
USQcvzAbq3H909QkLPPZhabYeWg7Ua5aRdTu9HoKM+Jp+JhNcTdBKe1+Optuzk3H
HhiFrpcFLAjOq0H8FFNJ7N+2Y82tlqWPvt9pvHj1foT5YDIcpYXFBrBsvPKlmHzO
ZC4V1/2alVGt0P1dO9vcZ1RlQvqOZEUAi73zaxQMH/2jZPjl0WDKhg9jp8it67T/
VdUvTFQre7u7enTpRgxDR7JWvgfucDXuZCgkDUssU3HDQJm6NI+IwuUdYgGiqL99
oBcAfr1d7zqVJkzib1PyTGAcyuiSOI5KSZL9+le8JqxkI66tcGNJPj/gGmIZOSNO
QPnQxjnTW2SXesLeVnAGjkxgQRw41h04C1qtJ0CapssSaavaOtchgAtcIuxmLF//
mCfCKXcelKJ/UDXZX2OSf98YnJDRkxW+ruDlRjNDQS0laxasz7trRS/UUO6YnZNn
+Lmzk6OGIVw5iWaBAcrzBYp6C0TYYnyEg2G3s/Gct0ljFDb9g9Lw4AnUqSEkpAgu
5RyyAeQBbonP8CDTUeO95CHtqbxAT9/ucHCNEOLXdMfJ481zzlOG3b/35tHPAjsA
8g2Ai19jXZfMizDsMuSbUcj9HXczPLcNoucEeoNkIMf2J2a4W9dyNAwLo1UEcsyH
mvwSs76AR6Mdv5LZds/Rj1Xx0u3DR3euTUOcpq9/Ibb0sjFgcYsxUXCE/zH2DfCC
4orOgRfHAROV2jjLynLE8ijW1ulD8Zw1DXdoslGV2AdAIhuw/8Omuo4U0GhxmT+m
iJwRennXMbAqPUPa2YqpxRzcgmgHpjQYmavmpTrnob9XNID7esHfdG7D6Xo88yE9
MuwrK7D3yp+A2F1FSPENryGzAWFQx1hwfKxUoSvYAdkZ5XO3FD4GNrCNwcNuY4bN
EwLRWB0mu75AchNrf6fn27ABwRoEz0rTtUQuWJtDli9y5woc3konzneUbqt3Yufx
f0TShCen1bZqe+2AGamJDkacGeVEWlQgO/oV2V8woSBsa/OrMNIeIst4hEMqkLom
oXkbZb4kJf8wiK6NZ5CngKEGDsXZqOvlqQ3OT5C8p2FX7CSXFGhthRIqwAdtTVS3
8ggPgL9AEBPP3WL7U3Si0sM1TVb5ByCvMImkk61eS8ZDhuhNz8FsDLpwBkOldvDH
mYjnMmkAQpFkIQf28PZbMTSrZOrJAsnDOCEHczZZiQGnUgqWhmMPF534nq/9r4n4
Aqp4Y6YMX2g/BkPU/FVHb+NYEDBfSIHGkBWbsINgxzPbfXZZmvW2r/1EWHkqOOH1
QRnP0pNse0suLVJO4oG+mvqqQYnb1HxPMDlDxySks2Q8DQqcZ0LXfgRuLtmzrvyr
cJ629JOBdTjGaqStV6LMDhF0eyEuky4YYXEhKYkS6v942kSmPa6FmEachJdTNw5i
p8GEmDPVqmIpG4Yr7e6R5rl/NQqhscqToXRON2y8zenYRJsy49wQK7tIQgCvSA3h
9AWXQyTgBsrHA02ERTZ0ixu2aCDJRH+9olInEqnu0aEibn9KpF4H/xbHSeIRRtY5
C+5fNIwryuTvBl9V3c49c5W49qDgYWSmqhStj3wTbHN5TGJVAmaMx3d2vg4c0WY6
voW9THvsodEtfzKYbSwCuW1fgR+XPCQHDkfbj+7rs4gtv9HkQkmcHErU3PSZCo4f
Mj3Y3QVVmI3MJH5oR+N6Lo9fu0lBCCkFjRxs2AfHVlOihbr75+oKrG7oakjO95wi
NzeWSVyVL7bToGxRNeOZP7aY7XnIlF5CTAD5p7ZTrB/Nnu/vj1JvA3ZP0U1yWjad
xPdbJVaoV4GL9muvePmOy1HNnIfHAeNjY8d0X+zcRQEJCSXCSwqOGwAfYvRl5W8U
3Ut+XDRhBe30cbMLSZjg1URfqGo6BqNPmmYSvc+ZSYQjUYPWK35jQYfPLSkHCQMD
9p0iZj9GSweHHxfP/iGgJaxAgzJEDbmb5JhnN7tdi2kicMkgI8hhPnU6lElMeSy6
/gAx1sQ3oOrN90FuZihFHRVf+bH5fZ28dmLRRVl8AuZcI9lEXyftFB8u5NF0u04E
8YIakmMy+ImFnvTm2bUXYAiNmj8ghgBvJ+uTcHB/QRdpUMq0cQiiwi8TxbnteD2Q
R/5Yq1g1yH6TFWICCAuXk77zKEOQvncSGgz0hxwN8OKfl+ilpn2JtYsvLbG7nxIo
B2Wv5vlbK2+ToFA6K0jMm4eDlYGVj/07Mjqy44NgN/nWxBoLQtof7EizkrM79ygj
BpSApAuQ6jHT/Kq9b7WiUXmZQf99wXgbpW0sb9YukZ1AIgQSt+20MPIDdeZv28Q4
1BLr6ynfzebMXyScPF2+5mdNcnWVRVjo78skLJcNoTkpMH5oaugA56ujQ2FzOLbG
tVBJStsHrWmtbel4PdWQClK1qqC+MT3Qg9lzGhoBX8qMAhdwE7bHcKDEA2Hf99SK
kf41JaBu3lc3wLCc5rHpLnyyanAnPxZfJ2LcI4bEY/5Sut5j014FwmNj3aOb5dOU
FR8uZ5gsbiFe3G0Mg1L8USRdcv9uY4KJWNVweb5Jjeb/vsEfLHB3aaUUfZQqBoaC
dAO6gDJuSlTlaDWyIivELQmtI92FhL1g7LhhMzHwnnS1/W7UBhN3UQd5GUtpT5PP
8pZ020r1tiL7XpY7BlYReh5eErfm4rk7SpbWFwtjMv5G1wu2UrGE1umH3CznHcas
hNGDI6+XGOfYvG8IKadsRmvRLB61GvZ6orF/6Z5yHQVN/+6103Uh4vIbf83zWlNF
8iVyHF2ygP2n5RAb9rYP+JcKLdOTANhE0siXP1rXxq1D528vQIW6nvaDQ/C5ELwU
cqvjphaFjJKmFpr4pmXskgS2C8L6943jcur6jL8kN3BTsnBTBtRdiGjKCIx/jvZd
kDUfDdd9y76FNS46s1XwPpoihXgk+pJ4SWY53U23X75mucHA7PpfA2o2Tq1zGg2X
GVO4Y6qeOtxBQ3fxcxHjG0wBOrr+l/gm+tOTquTeDsHti/LYjFWdRjm5J/CRXtMs
1ep01D1fOFU00waAmymMyxxxxlXEiQp60Sn8dNCxVn1ylxx5uVtGcCjaMqbymOce
yUqQpEDd4SqdD2eVGQ7SdSeuiHrEguxchtctqHOz/l82+2OTLk0HEi0pQiCnNJbh
96ik/jui7/97efRS1jdWK7NyJ+De3aPInWRsyGWsJVtRfMsc84VmAKNjCmHCBA0g
4qGwFURnmhJ+1h9UPmQF8kwlzqY9Tt+wK3Jb1PwOutnKWZSKb9ITECVKM61rJsYO
F/wf5Lt6C/OXoGYrM4JssBeLLiqHdYRujAjGN0RjeHc7AdDB8Qpme6vtqYG8b/i4
FoRcmjgjhAd73DDM6Ta2+0+iuxJ1hPLIycRJUnPvQV1nvTzJaCdr4PgV3n8sK6yS
ZrUvNKCKsUEUC85czgVG0Uops3Ry2nLLm7mM/imPfkzYhc6HX01ryLKKlVfJ8aHN
i0egeD7O7g+1dlPh+SQMe4W+BXq2smNIZQXhWXDxz2FCF6SvLewpTShwoPoo5u/l
62Ayb5gz54UdQYsZP6XiZT2hRhl6VRfYfhwgHoHNtz75y6OmKOR8p5O9oNauB1dQ
S/ukxbO3jDQNeJ6JIpOKDBC07Cj/L4kcaB8rXlWtPcnqbC+uZTJQ6yltw/0NmMBV
NGJ+Kx0s+mbmUh/D8zK9bDDlx9U2/2mcI4Tt2io8sFFDQgmoAdcuQ84t9GZln5um
7zcQindr6+E4T+odT5bMlZ4BndwzKQY97+aR/+zQgl+zOn10d9wk85h/GkoAdCzb
DXN6iQdVuNlPAyOTla3jKb/Vzqu41eOmAx5qNbyK8Tc6//ZaqufsKtr2qbfeb//p
PkLRnTHP5/mSLgcpa2ZK5sedxn4txZC/ZM2hyutd1oB3EH9mflqQqbg2Hq5Urfh7
l+TJMzSLFldnpLCs7A9YNT/2ca2WpwHh6sUcEyk5foswbkXfHMQIMLQcjvDXf1Lf
ClpuBhXnJlMbGFqmQ26dtpobpm46VUjgx/iNM0p9gvdjN6I7moAtES3XI0QqhRg0
dsV6L8kJt56ojmQNAGamgKsw26ghQwfFChSP5pCzfI8YVo9H6BfN7pq91YBBsUBd
dy9QsLtU2I5Y2MMqdpATVR0zYc2vmk6W8tM1bi+8LdE2fo63AZFUkMr8ICdFjho0
XtSu0X4/Pbimlu6CorhQdkF0z+yTwnsSoQqjATRxbmAyLIrE08q4lgVs/U+ebWAN
N3tQiTcDcbUVBc8iRCLS0eLI5/pHApmUpo3AbOicS9Gsyh6L5XtAJrrrnFYL6n2u
PfgLh2RS770oB1dLEKkIyKGFQ3OErcHGMmwtWP7fTrChcJ5XWvOx+7eIGd4N+NaL
bgBygdxjOSU+AHymZunqLo3ILjM5yWe7CkC+1yGxb2WfKBJ2nQQgZs+a5PwywfLZ
AecZljc6KUcEPLwgiayLLBTXaw7GJfGGoRdrUEjk1ty/c95ll9R1BKF+dZq9pSDs
tWhc7VTl3ckJgon/JpceUsuboCEEQkrhKlKi2QJ9qaWOIznMvAWDZ2B6S+KfEU/I
Nhyb0BY/y4uf6opXruW9MYQna0uLZcvmJkSN6Job0pkENrT/lroTQmJce6v3AXvZ
ywrt+2fJjqVOWISf5bO3HgL2vOG9tJkALv4CGPCRhm6YTFaVHCE5MpXR0Ks8RCnI
J/xvL+0JdjgASEBsjj7oZqfZ5MKSMQaaF63Lam3Kc6rJ3SFG0L4umjEGKrdZV3J0
xrSaASNn7G3/Fg5Khg2y713jMySFq7n92Ak1iESpq7VQABJTEsKpUr/VMLGhLz0c
GYHL/60lnL0sYSL70mAnidX/3Mp4lI4pqjDsX+3/zLJda4aiLz6FhWbprYxMSgXQ
FQWvtGmIJPfnQSvs9A9Yo5fyYFhuBwmw6t0oyVqbIpZhfRzHy332VFFNdC0Lz5aZ
7t4XtFL/8d6pONWAxTA9BGBChC8TNjo6SJPzQlmY5b71KH68EagJWQnsmLoxkqqy
we3Xp+k9B6PZovuQtpppG/1ncXZtsAXKz9Bsla/rLdojzHk8UDsTzrj/+1YmJJ+Y
5/8d/CrjQCkzmCdNfeyUofK4cmzlF6plaw+nnVe//KgK8HQqEk3mCSIUgsbkhY/Y
KRpFWDNZBQGH+j1DBEJTv6/uAjgqbng/wdkmI2qaAYulz36YzppjNigYXBBR2xHE
nhLI2p0aj1BxKyDEr+OjXiR9/g7Vx9bpSPXQdUQoJgKMgEv0a+4PNnAUKBibupln
YI4IETPSDwYdF1f8eRsBU4zPFw4G6+KY4QvuR9MuwvAFVu6Q4OjNXO1L8ILipUZJ
hfKgYY+UAjDqbjDn1R4RyZDv9V6ZBKtYU+WI5r5BT5JyXOUi6Nh2hXwlcuPyO/6B
1fvxYV4MNleA7RD5NzyRATkrjKBDHqj9pFheEyTo2wVI0tiiFzjfwz40kdBKE/EL
t2b1FsqBl30lQNpIbvTELygHTCsJnTHKSLDJrVmU6F8ioly1uYV9KOHvQJMNiBrI
GTd6Mv5TKl+E8P010XHxmHTP6uPVYNDhiBu3Ujt5WudNR6Jdu8bY2RVnC8EB+cVm
Mfud7wUtgals3tijR/SgewA7Em3TQ8g7HeljSYnLS0rnI5LI9mQQXA/ARuGxhOKk
wx+iW2o8EAQnP0xFAZmerLOtdYP1M49G76kDR/Qg+lY4S66xITRfBTcG46Nar0vA
EbTuM8vian5eKTmmHw7K7I6IaR8DoEPV7zDd++/fRk+ST18PcRPMR7WSyOIdIymb
SK1eza5LGLlj1QjrNBZvuZKJcJsM4PPR/1tEQQ9FB6QH8fo+ASiijmG6/WONiW9E
PMRIk5EtqWOGyGt21Jag9VDFNEvOiWsky7QBLW5vcmfV8xZ77Yei705JvW3yaGv3
LWdrTnp1ySaU+RlGoOXQb8qhQzcrm2rvMoECsKZQRDS1seXN1qE8WX8NSJJeOzcD
Z8sWFzMji5N3Nkt30SB0Hf8640/iRYf1ZhUvluxa/FDvq6saGe2kescES4svQsA7
FmZahyXxIV8Nfmb0L/Jzynm/JVXcUFXvvt9zgFomgRjaDAFDlxMXHKxnbLfBJn6B
uqzJgICyyzFew9GnmzsviCaro9Yq1bxMN8xFDNUObr7P/JgLyAHKCIRBmXUoT9aq
ViysH8cDJwQXu81LFR7VY7FfaxkAuXrLZsjwMsRdqEPCF3AKauo1L7QUEb2ViB3e
wkVJPqTexGXJFvsfI/P9DKkfWn0EymM2A96gTiQVDyhHypyVP8rmwV92sJHWjkQg
SzAX5QtEqLxn4z1I27npr+Gfu8id2mWQytHcW2U0XT8P2zzmqeh6PV9lV7sWHeec
CWXc8LwF1Bo7YuZ5Ai51OOIUQagBPRaXYV/rSf5C1XP6ph3zSu/ZMQsG/n9u0XrH
XUZfd5Ys61iKJ2gD4MsHSIMxLoPIAg5RTbFs8Ftj4bZ4T/WmgYXOtokMrFfNgFry
ZXKsiC/35EDQ3jyfabnGztt6oiKyBWCKENLenA/V5L/HcszEuZT7OjMNHuf7VrLL
Pln1YQG8mrFZbRzBzOUIJtBiqshToVnH3+JIjnTTvpTTvKuqf+0QHTK7CF/fq10b
dr1m91zI2K2hSR2q868Rtw/Wn/FCKfYZle8b2HcE47UJ5wolQgmi052VyT0N3JhK
W4S+vCxfCRLFue7vueTQ5uojEgFN5Wk2FrgFJGqRalKlmsH3n4fjJRgnUXWsHwRq
P54k0ulC96YhQttAX63gRU3TmgsLOaU7cgPlfmn8MmqHrNIPJ5jPV1agmaHm1gIr
gSQEUz/KEWp5ynPrs4esX+lJE5FjsOLxQ7TDPgaQ+1w4GoL8UEiZ0U1+kX/zc4ER
FoKUE1XKcW9nu6X7vcL2bI2kMWHUb0kGnSBv3t98yH1ZlgNDGFCUmD/Upnsd1dF/
c5l9JIWjIsC/oHxsyWjkqO43B8Jozpv6dIwCs5nCpwe4sjzw2fIZurY7rGPLPl9c
/M8Nnar9tRELcaD8dYyNJ9g8kVR961VMTzx7gt9nkKM65mv/22BPPvnW90+hOz7V
oFP4Cm6R/peJqzBzATmSGsVEjChAaUmYEAFbrrS27eNOEqqQLOSrwQH+k/rwpOUD
/B+FQKtqPkpiiHl4ZWN4fcU+un+5JxLrIRTcR7kAi538+euRBLf/Z0xt9ShQ9FC4
fSVHAktWfl+GQl2QwdiRsKYebMRuhWX9FgwjgqbNW2AMWZbGVS9fMQuQI5h/vLfY
CNvMO9hzJOOOs1b4725JJziuhNidi79TWxrDZvaimrSKcxVJuUwb1Al4br+rSzXo
nQpiXJoZdsWg2Z7PVdpUzzHknLdk/4XjUm9ySWlzbn2bOxb6Pr0n8SF+E8zRAyJm
+fS8rMKLDzz1AhitB5ItbFwBACKk5cH5BBTkLuT0v655CmvBekt6EkyqXC0tJhaB
1sT6igkuAmgZ9dsYrxPFN9gj+UTp/sv6jDcy2Ke/OBQFweG5Ot1+/tyjDE/FcQrm
k6UqTjnR3NGtRjMl9ZY3zl3R0C2mkfJp8nj/Ml39kI4FjPdcLmICPJOhE5nTAXVW
rUjkP/hAuduRo2McdDPtUQTCrNGETGbJGhAh2NXxKqPOsUyuhZ751rmIVjEMxrqT
VqV5/L2lLuH+hvjhX9GwpZnC8Z2gDnUgbMku+XSyQi4ROu72EQWidE3pZBkmwj6r
S7mtSpTX0VR73PJZ3ujor2m6Flsbh5P54J9M9POez2vEAVyfvIKg0W+ZHTQLyOV8
4UPyxixiarJh7TZ1WL/gXykV566E96QnLFtAPuiLZWAe4ueTo8kMdwegq5rtBHs8
1Hnh+6Q3hDkowg2dDeBAl2V2ZFs1P/xgrJ5finPvZOuNCFUJSbYdw5HGc0Ca6+i9
6RjlPo9k3QB2vpSmAUEKYUWVUobrP5IKaprxakSgaSTlEOeg9OxM8JtnRmXDZkvk
9MqJ1dYWrUn+F8cS+cDbZ1eqtiRaXJbGikiO1Tfa8VzgjjkXMDCsQ9o7o9qLTGkv
cTutAQn5rOwfkuG0tVHtceD493zGwzsmrhAuAviW8pQ2ewbIyAqjbjYqhyDeTzM1
/pVHX/RNtn9CAzS6cjIqyDFSImjtCRJQMEsjD4klhhkgqzmNYtKuMOfyfNWO7XxK
nwWLbp69jhgI9ifFUuJi7zOHrjc6T32XaeAPtxYt6xseuwUdDfwjnpz92AbrrIaR
Ohc4vBCIfS79gIQQ4KgcoxsxuKHkcrBqdhareTxPYtYe3n7L+XQhVILu/5qASqRu
BRdZIqnPra+fPIIoaO7s6Vdmik9y620ArqzDo4XkTh2hIuegQCwh/eesjdECrTPs
I8/u96zQ7zif834UKLoTNuNP1VD0XoXr0qYvrvFsy//YHmjkD80ElAVCBjFQEjjU
rpEnChqmcAj8xpWWSJN1+G9cgnX/lUfG49jzKNH/XDYCsVt++LxdeoeFngOcYqNu
VEEXsP8cDbNtEjhbyfpUX82D1iMAOwDOFlZ6FlrngJ72QKtQqV80tHLZK5UaXMGo
YSdSqKJ6XH7nLH4xEp+tv0bp0EJ+vw8opO/7oOvd6/efKu4PDSkkIxnRzyDW02hr
omzZw0rkOhgRGhtQOr05tIntlxcjk+GcyTQ0gypRH1iet1tbmfpKYVpYoPL65Rst
CkbfQqiBbC4Ft7A20ammwcayDoQcARWFt6QbVyz/hhqF+MwO/gmNas163gWjRwWL
0XZ2hMXjzi7eAk/nIbBKN2skaGvaIXmL/y/kHNNPp2ZvrkzW0ox+uxudBzD7jncg
5dpq9dQR+z0rd0zI6BJ6zYeMAekHi+i/X0Eyjzy6jfmYyEKphmMUucCQJ/IVOknS
i3eP3HCX3X/NxeLZC6Hs1VObcbutA42XjGSWrG+uRSecNy6G6bsMla4Aw0SZbSoc
eUvXtgHg7m3o4KySxUng//7RAVbKSXeC3CuXzW2wj5OQQNMFcbh/XEP4qHB2D8up
l8JVf55qO2JZoCg6hShryFAHs2SJVOp/du4JkdI7zFgxBO4lUoB5NqRukgWV4lXc
qlVQHVkZ5/+/OADzxBvFBfX4xrzdVgjBiJrKI/l+WBCZwZeDHr5oL+e7yPu+/Ysb
5lr8oYieShzSre+zieOOjDo23Knz22P9wVAK1XbOKltfOHB/IzXw2VcYNjN/72vm
bEbxivQ0BSHz4W6Q+V+ZWUsmWekxBhHnqEv3PRmlnbEIaeyg9p0bWNClcL4a1z21
teC0se8BBYBKBLElIlS47/TbrqNQKCr2dq52s6OwU9VHlE/uRFrXvcVkd0p6YOlM
2Z0V/R5twDcOvvi47biOwwnE18NHkyWL46sWN5GO2YQCIe1VTswYTAI43kB0jFds
E3GT8Vajq1oPo9Noa0Weua9sPm77f/TQ3p1L2rk0fnTeoWA/TkO3z83WOgxfDNz2
M8DFuPQz6qDA8SaESOG3K3fOTim3mdqn4vTyfflYUFAijth7xlCbouPd5b52HKhm
sphVx6WSwDGzXluuF/7+MY3BGC4Qx5n1+XhH5tso/X5qjYKF36vzsYuWVocABOz/
C5bBfjbeQbYwi6Cs4wYt6/GK8KnIHb3+r+8Cmsp8ZAvsoVZaPIlidvktR7jCmy25
O/jVMJ5LUdXasPyYnSDWbpt/xKmS2mHiU2vde2j/3RgU0KQnOy+zyKquh+hsxlQq
KEIrUF+aZBfKz7xOUaDdPMTNJiVggkWIM5BmmxKuL/sSxWkTmjQT/PUOFgHjijit
uwwRn83HnGJ/JchjF+mDEhyBjMvw8RJFMWGvXkbloJo3qYiVR4MTqAH7UlpcU6hE
E2OeyGU2kzdVRtwo/6kNrdVNxUgZOxJUCSJduxdAkLrl0cfscGDrd9u6U0glI6Pk
Zjdo/IkUUgrgZk/gItalXQ8fcUb1luAVMho55YubTYrEqJm1JsPC4Qk6ep6YiRKc
MUOj7khy2ywpurn2ZfSwPh6y5mShhKBRtlURmiSJqUhSVsAz0U7INyazJ2g9O9Fj
cbpLj4MqLkUcKPMfZNerJWMlWmAkUpFWFgPdeiL/msnHHjGE8vrzXNP5Jo5NsFZp
Z7X+TxTZaOaJ+t2urwWacZ01+hacHsnks7g2butRXc3VFeJ1T9Dh5yU4B8QSqJX/
SIoHwixM/nL5Fhr9rpOxFWoq4q18/3D3vMHYIPlHjLddbIT7kfzSHdM9jDfUe+MP
+pVoIt5FI3pkenFXs5Xz98rdFZDyAcKCmFuGHP/U2zKC1AXGZXyEiQ/gDWp3O+uN
bps8PwcjjrllzM4GieL7Xz8ZxPe9IlZDgAeT9PQ21WsV5QlhxOfPlI1BrzC40AQc
AK2aa0eCZPe+UdHNO+p3zqnZZIEjTD7VNCp5y8fmxf9SblGTzKH3qXJdldIaQ1UV
lXiEidk9hhcrGbjFyP4d3vwzn4T2JCFX3duG5p0rQ8FNpsUkP6JaiofGKdsd4eE0
jZzukzptVkmaufTCGkdxcQeWZhbl6SAly8MPaM1fMz7PZZEGtO6LKrCIpQAf3c7x
cc2DdlFr9LoHidErlA1bXIn79clY3AqUB4hwIEv/3XL1L2IL1Gj9HTbRrGSJj4QB
w+DkHWvY+yhzXTXpsVfoPlmjXRAb38zyvvmcPdY9UhQCxvvwEzsqH2gViyuTTlIj
NkmiM3/W0/+I0ybGflVGFA2+RYJxr1nxzbf4Bj5RwnNNEQ9ZHU2udzgqvWjTla76
DnH32e4d35BqGmsmKHO9Bk8OOBpUVvFssbp33QRDFkoeLEJZJjyTXRxFiSAt3Wcv
Z4NyXAKjOxvzluS5B0El5btqlUR9R3ZA0qUcDjuoqH+LruR8FWnu1/CpeSBwm4A2
boILHY9VSup2YlL4S8eYJcgoLw5Fnl+RWFwDfkBAp/j0eamIQTexDhhIXYtShEyv
YyUDR1LddEW6EkmTyckOTHRymqZtLwLrwSFmcBEf7aoJw3xEhvkLOIp6Veuasc+G
VVPdjxJC2WZVfN3LB4g9zos2tP2xdv9C1O3z3xRo/YczK/Gs4ZG8yQCzUFrIoSCa
PDw7qgJbskAzZMc3dNGraw5g10imvLxEM/ejlm2VBlvVKftp3bE/jA9kn2aIAKBu
qtlyhV8lEj/s+Cl0IqM98MwQyY3MRY/GnsGwshqzflVXdVlfyq11K9RAhlEsoAE6
NIdJfqC0WTL1aXeAmmXPNYVVBrMqAqZuxJyboFx9kSiWhHFlQ51AL94zXzwLJ9xc
h1jpsInA1XUE25HurTDjVfIVjhX7ED58WlfruKdWNw8zWP7hiLYcQ8RXsMn17VC6
G2PCBr2eBFEVEUMYspVBknP1mZwiGtA8D7bv6JmpL/nYtMiig3TlS20M+f0F6ZMp
lFOzk4HP8e6hjDBf7NovlWYQ/beG9rLqGFkjLAIKDLig26YZa21ugr92xepnNod8
BLg7kT7PH2ksJLPbmRSgOv6N0GZkkk5Vj7osZhVRUS0mzzGgC8n4KhrUlswsxDzX
RBTuap5tGOfOOufXkmKX5L1r4Z1Requ9b2mxYkhpz+UubACtMb9PxAMWEsG6e2Xy
CYVUiQIt4eL+MUwYtBFvkB/Z0w1lOesgTh1z3vHeMUJ1UVm/0p7xhhT49yenCERf
5fx3belCx1CFVy7SNjn8oF096bBRT6lucqI99aM1uBjYF1OFCdYa7+FjXR2LLhI5
WQLdVqMYYFT0i+/wJ5mFx9beLeqipKIIQVBzG7knHn90ywqxNQ4fmMABIuz5jlG6
gasentyoHsLZdO+met8XWFGUAMv0kJVmJIZuASh3DE5YBhLVqj05xRTFyf56LftN
xGBIkUTJcU7zhB94oa0rztkEAlWIpF5JU9+seXl7EjGjIR0w3A080vnrXVWeUioN
cSJnznyO4Ai+GLeJJByYrRsngMOk2bS5oaQJIUUKUyH4nnINNXdk2ow5MwphKVCO
xZGaUY7lMl4iWcjgNkUHraB4R6I4lNeI/dNknWF/x5qfMip7NcTxtxVDNeO/jkx4
upLLcGWrBVFjyhDQJhd0skVoSOI7Q4OvOlY+RQOKx/lEv6AHWeFGBVHjJ7SOqpVs
HG5SpImB4uBlvrrtxL1qtCq7p4FTbgZSMRWnRofoqheDw+A9CvSuF5B2ub5luwdf
LJ6TXfWRj6XVwOvQfoNE1XwNt6j3Oe4RmXiDpf9rM6zvS1UHNtVT+NLIudIlrLq6
snH+eNQVt2hPE88hR9uIHkoE/J+wasM/z7AxK70m+iuweiSSpyqu8Zp/EA5b8j8F
//pragma protect end_data_block
//pragma protect digest_block
DqFLdqV1eSsEbsA2TEI5uJas7WM=
//pragma protect end_digest_block
//pragma protect end_protected

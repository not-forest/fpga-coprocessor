`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ayUXcEUyn2Hbq65+XccvYWHrFiE7ukwox4S2yPaHdzcmTboRXAmr8O1HWU8NxFbX
VhHO6sRa2nlCvDcc07qYl6BpebZzXRgmcPb7Yl2r/AjPmcUw1nQLq49IMSiH2fsr
BFQTvZdfiP6qJFDfLV8qa9RbMe5xwQ/URXKp6vWWzVA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 36816)
nRcrYeNTe7L4hJczCXBPkf0m06SpqrkiIgCIEdox0Ve/dxV0MkPSqv4x1D9JFFWc
PE2yaXedN7g+92gHehK5l5dSkqfUXSVdVkWeTqE/frf2VxlkCi3PzxUVhMSPX/lB
avg/AbDoJcbCnyJIfBKa6G/K0wDW3lgoFflJXh0ouiesrnqpgYtIBqaAJiC/vqO6
vZ4tCMD3l/f7RTtx613NCueKxB8xWt6WwW6rVQnYgAohUcyQ1Oww205i+lKlyCaP
BHp3ow88GbAmzj625ksqr1Utl2wDZNPWGDfEk9+TaSIVTb1y52u867dttJJbzKjq
3pfkpy6ppFFumqCWQkY8ghMU4W9C2/Jp8bg5/dac6oBRFcyPXlICb+GTJ+XBhxsr
nYKgRmCRs95+fZ0a2JfBL1ZpdcXNr9PiZswOfKxSKTpEFeXr8iINflRWW8tPQTcm
HRQOMBcCSBSni86hsapNVkmJ8frjR+XDUyqC5ePMRB15M4Kyqz+oVHGhzbZXot9W
cAY8fFo7pftbQH4kAV93k6KxSXWhXJ9ukUeGpOA/4CP9l7PB2E5RFN496juJY+RQ
PgLWxjAhvhKG5LFERFg63FedURx9f0OVz1UFP5KozaIXiO/PcpwGfssi8qt1MNez
8YAD9g4M3BjW94n+NEcyjmtTY8H9oDuK/uF3s5s934hWpnta+MPd9u+YdHsy3tky
vSQDw57Eknq4mrmT6OlF9XOeDJe36vnGPMs8sOXNrkWY85mUYQMIeYtNZeDdLm9F
2OFAAnmfrSehZoBKNWVZa2UMqiBOAvJIjXJ9jG451NWN99b4j9UDHlPEAptnYYeW
XQAZKA8OTQ3Z+4h+l6mJvbhbS1AKsYbbh8gt/+v93DVD+56fAfgUARtH6AyzBbl2
GkAqgr/LbL4DvkoO69IRmF3JVffdujiSnARiOht1kPim4Uavtd6tAdfTwWX24N5l
xcGkEi//26kd3B4/OtiewuhgdacGLNBmQc1kOta7gWpO398LS9fAXgqFaNJmX7gK
Wp7gQQiooagnNJag7F4N+20lMMmUCSuUK8SjHHsnLQuhOvDQK3UUEM9d54zUbtdO
lu4hdj1xTEDBPmc9sVVA/vAKfbxMinKUFt/zARZS03IWsXm31/aO25lDyNEquEDV
7axPaUq0NzJ4K8bNlWDHD0C46x1E+5PSBRZdA6aj8OvhnU8ZK+WjNZtXeTAECB7G
AzOwZB5jsrPLgp+2b7bgdNq2gGBT3zXkqn+KyOny4tRxC/w9d5WfG2kt9XVfVG4C
mzCOQrHOhnyP4EVFLdU4gYban8FbtyKrxCAk++Uk+eZf2jcOyn/4xtCr9I0Elymo
9gepci6YJqgglTo3fzyw7vWtdKTy/tBpkNwnJmHmMclx9GCLrlidwuweRLwJrOZV
rs54U0qfADVdn4MWaItTljgucOxNTBWs25d+of4FbeaIwrPv5CGXYqs43psU3UOI
Qtso7YJlqNMSmNvb+JuPGFRdH23AaIGCXlAfx9RWvqkAXQ+araRaCOoVATbYKm99
CGOc7g0ZECRzkRfzziXtABVcHCFbttQT0mSWLvEZL77PnYuBVAy9HAFP/FtBcxxh
5ajA+dzAQVaeguaTxsQCI079LwSsZtf1D6VQdiuU6w0YHGTzec3mpRdqoejm4dT9
HKJ4fLZnET2QmkvXrkrrYsCEC7lIVBLfNUf/S8jImMAkDhaAUrxd6imv8D9xWXZf
JSgXSISn0Nk0hPQ4B0izDYJ1nRcKyfRPUQtZBA0YqE3QWlRuQJ3BoJlQRVH2hDRg
LsggsNBcMm6ivksfLDMtDBfUbDNnDmWs7hgK+qHoXyXXwz/3NuCKVDcfPnv7L0jG
sAn+SMFhOvC6K7CyXi/tI+jyIstfgzs4tYDIiV7DwLJxCFpgvk5Tfi8s4XR+CudX
oMef9f8cPKAGOOkdv/Ht3vaLgdyCgype/dlTi69NDPqNf4ST1oPQ3dNOdYzvjhqV
wpEChwqHx23zCxUQEEutJhiAMUsuRnZRA6rrvFS2k02HIXcl2slRCpv7PDLQzDkj
SUojX9SY8UPL2/fGXDYzLfxBXxoH/Cl3zm0ixsE9+p7gaa+8VhvTuaqR1hXhCalx
6yIaFkzXFHwFIdZAN7ANZEsdX7xXp/y4zuT5byaap8O4MmQ5tZWssJKkL3tjil+g
MOW7vg0sgcleTN2xZDb7/KKVWnL3Sj0pS1USLwkXqu7ZWKALSWnOmm2jZAx/34gq
rreoIxJAGsPYORGAjAtlfYjkl8A//hGx8dHDPuDRyyShQv8REBlQjZ2UjktdEJWP
73UqFtPuMQBbza9ULu3GlDkQcj+yNRGQgc+3JLkciLSMC4Z2EMxxLx0w8wISIF4z
40yw1oRit0sKtbCs2fh0RnOBPA98UpIXf0SwwmL3R4pOgKVqj98YFinYbGghM1PH
q04aCS1ZtlIBtpJHrGTkz1Z2RFPMCrXGCfg8lxMvNsQGHQLjdBdQ57q6hVtgjVQf
rSgVGXHbL8nZy2Xdw8c1FtgSzs5thqyy5hLx0QVocOLNtWMEqhxNH0gYDPirP1HG
C3A+j13/Fy97KnRVLXirF9m78XTokiB1DJb9pseVPtcTPSZN4E1HUAYXXkHErbiL
0i8ZSLn2pAMQj2FiJInziIEjymO3E4zF55ybDPvdnrRNT2qmyvukXFfiog2PrtOd
yJu3Qu0ni6El+T2HU9DSaYpvEmsbI7Twh/3kXq/MzxiP4M0/B0P6aDi3+oNpa6D6
VlArRMLmA/1P8wtrMjnX4nPbqCn4aJys164+asNX86LSwP7MiA2p0z/3VBAOQlo6
PHDXr7RL+xrU+6dbZqpSiCbLmH7i6wcXELd/qo/QYj8t1pu4l4Epl24QFsrFQZwM
q/mqezF2H2k61iXPMd36t3GEvZfSE/zVD0WW2bder7pxFEjSnB7j1Wm9kP20pY1B
iyYGW/w6dRaS9E7OQ5HA59j8XQMGKCMGwRDZaJlcsTqEh9dkByVqNhmpjaE/8Vri
gfL2/M6CNNjordu+DK6dNtYQMkR2MFR18cNWqWhVn2kJa8JqzzIfTfT1hGZVFgpC
+UwrEQ9hJ22VgiimU59WC2YsbiOLWq7xchXBucxT5bnGp8un2DWkacaH4X1fLaM3
qGk72GZIDw8gauWoasLzcm266gihzv0vOm7BY0+VE9/Ct9R1HVenaLBoqs7oPErO
fAm1UQ7HXPAfLPPpzMTxWDMbMxfgx4WYvaK1RWnLLd1TGSjD4xcFvcnWCMwxPl1E
lYA3HvGyhImz/N95ORbF+bf38mRbXcCAu6KHIyncO2wWNk2iitwDhovDNEYFEUas
tlLXlB9d1Td5vDbtfhEiFizMOwkzNB3Sqe7ynxGgI+4OsmksQU1yM9MYkX2G+GuM
d/zqrUEQ+wIOx1UnhzdRY2rQIEwBbk7L3ZfXYrwUbl0J+fv10lrDKBtI4dL5dztE
LfFNKUFo9taWSgQ2YfEhy//Xw31d7X3Cm4Km8+PoFnwBshmxa5iJoIging1K40A9
Hp12DZKIdQ2vP7AxhCVZzguI2JFj8wXSS6VKCAqQ/rZ9yPHzRh0zYZQOHx/Eswat
e/lUQwU1E6iovYg8oaJfiFrhFapbBd3Eqh9p/t0rZywdtzHp/7v1rFeGbn2EkOv2
DPaAxYrDUkdDzVOMBYxBx639BvXzJt0PO19Vd/pFuwivS6hO+oZvKV3YKikqolh+
TEJI+9HpCTFaHWZQXAgVJ9kChsbWorlzKcB4z5GLkVxImRlMTl+dQyktpvlbgfkS
xomqEEADTj5ZNHYWFlfPu5yMtvexiAB1KfODUoXIy0jsIsAm90FN9TPYzjblejND
8kIWfrVofYXS3x9p3pN98tyog48M5wgpCLw6Hw8JitMJIQ1+zzWnj67jTIrCkLEM
/SUZxBdMhJzz+SEzIFZb1+xLbrHLKzLylHTh0SLSA6e0i7M4YK30Pz/n2bzucsBv
fVxhYSQEGfqttnI1qn0q3I4vsb+qTfXoVaB5AGiOlNFnt1PqCtvTMd22SS61G4V2
aI8TdAq5G+2UFfYgCkISWEpUVZUA84pVc9QKoOaLJz//u8jPLiY2/+HrhkAbV/Jb
YcLBpJUSrZSZs8Qcp5pJ8ZjdHmaOoQ/zM2QiuPjOOfQvF1RQ41zH92yY8ixjGXGG
A4OaLqa8pR0Su4NPWfzx6+/Swgcdznho+eSELRbRjWxVNLKPgF20VFF6VI6Avo9e
TfEZLlzouUvkELj+fslO5UY5WRdNug/Jt914XoMhodP4yP8X83yV+QsYn/frUWUd
DZ13IH8dL0Iqf6Mg4roMnRrXAFmtSwax5mOQ5eyntG88quaQTff+baGj/qxv8OAT
rlKoHNAenW+rBCx3Bcdr2oYz9hYvG1KfSdTnzsBy8bKUhksYnT/pQK9xGwGRURxT
5MBKYOQl3xnLObpLG71gmQRPjfgCUkSHpSvZAc8jIpuegtHTVpSzNkZAAY/YX5P0
XsmPT/7drUZnbmDKoa+BmjT18D9RAY5pMXyHKoUyPlXf/l1Q7/+gjnDkdraSGsnh
vysfjoGZJlnaayq0xNOj86jzFNHHvnyQuvAxQQ5qa0CzjKqnB0TfzTYaseAQ0UFr
yyyrROOpiksOUrtS7d2mCTRuXIJ+8OjFBa03sLpjn1nj5F+P0XBKQ2d6tEfc1Bp6
5e/X/sRbwT9HeUtkcKWt+rQoXjRB1eVRAgATZa5PjkngUqWcxvL2jl3GsjQeTfxi
uhh87pvqcdAXz9KB2ExbsjqKyAhLzFqdShoPRA7IhNeX2TJEWJ1tvQW6N63N5zN1
poUR4/X0HOyDY4LZE5CDnhjuEXGBu3Hqi2HqCBdQ1TrvMF98DM4lgDyt6oX3Zm/Z
RVzMr4svc8+mrjVqSJI8dPI2yKNthsVlioiGMeQl5dZTIMAxRj4EZkcs3OKqvqZs
QjmuuL1eD+MeoggJsyok5cC8xcUAZgOim4I2ZWXPksN1qbFfOi+UQEbTeW8SkzVh
+SFH0PN9zkrYwAZUyK35YHwuvqW0D3h7VayluhLXQ4e8zzXjTsj9D6EZ8S30u27s
iv1hAE68u7kQtpZxEAXs1HDB7DQfaFccr/WMX5MXFzpTL58BSb3MZhWJ5jliF43h
uwNsvLUd+TsNZoubUihjoIR9zZiwqVLAu1HrutKOKx5RO8wSfvY9mK3bRd6H6zy8
8YvcuxtLXcV08TSqBWYr+u/QVTHtnhlqgqzT8olBSKCWbqdOWUh1imynH9FOP0TF
l/OOFZ5mPtxdU82ioc7AdTQPnesv0OJp3k4DiYo/CVbORnBbMiFTWy9hR18HGDBg
4zSY+xXnfXyzNYO5/yIJ3yFVNtXm+EzmwpznO/3X+vWzQYxPUd4CGnFMD6a7emOp
5qKWYwMnVQ7KNrA99/Y7avoMJbrWwQ9pLNAti+1V/ILYZuSY37mvUBEnHsE8T5TK
g1aV0ORd+Jhd5UaSnqALQMpzwffAxJ+ZPjniBw7NyqSLA59W2ewIU48UwJig/M9F
SEdIQ8dfWsqAaXZh0o/Q09HTekTzs1toVQfuGGIZzx9enB0T+PM/ennBeJlf+BKw
m2qCVpXmM1P9JtQW1IAunyRMkBqyMSTyomwDmjbmnRRSQrWMW5G2DdEWPG2EK2vP
h5Zdfy0Aalg9DBjVego4pqKk+lQYw4WLwu/jjf4dma9tQB/v5sEBRna9meRYbrD2
4LgMGz5hrfIXlho8oJbINAxETq9yJSlNDVDEMPUEbeDIu1jFH6xxKh0CacyPg+9S
c2MitE3darhBjzPnKELhXZ+o6wWnnqzwm3xYdFOlH5Q/jX7o/ZDK3k72lZuiVezy
1Tsf+4OtR5VKwmB8cflf1N6u9rWPSuQ0w9pSKyy99/jjjAgs1UnWtkclPC547eqF
RAB7qSujEkuhDcG6jY7TIkQXCFsuve5FMZnYyITBwm4zWWZs2lTovyb1x10jufw0
k/nQ5QB27Ylmp54dggD1Kl9hunfQuhPULFH2GDvtLIaKSYwWSzgkimHfysuxWF7T
4Mb5HW6Az/ViAu6Lm0C1nV2kz85EkjtRZYosDxn5VzfGFJplLB3+JOzi+azS8MmE
hReWh2HUXX3Poje9JdMSUsx/BOVdFdoz6Y6HNoARRCzJUXja2T1i3GyNqE8hl6c/
aWpgfWeTpN9AGulm3fJor/IIKgYpWsfjIFZyJFXo5hRR6uRfXU4a0axxaqDV4ekt
fxOGQTZuYvQnz8r9Ifa4rU891TkFFyHjoMmJk4+rZkC9Pg7ahvOg9P9ZAsQXj2kL
sgxCNbh/U2PcfLhEvpOTxO8ZJMUStPmjL8vFVvXRrRb6STJsYDDkIvEYoUKdQlcU
+P5k6wFK1VG4z5P1ec6iRcuySlhUJrA6qoMJ3YElk6HlRjn9ENegvuVf1DTuYTLH
xp+sQyGdMAkc2PcmSZNdNpTcRh2c3Vtu/u0QCxR7EmD47rjtXB9aMMAivVKI+uXU
dn3qF9ri6MlH/WUSTJmV1XsbJeI4X00t9QbUPwqz50XLC3NVBt2nJd9Tb72YzxLR
GI0D/AY1a4+uQe4syK+WfAdy9LgpeV4RTbl1aB32RKaAk+hW37tRfmsGdkATx0+z
owkf8uxRJFMWQ0FwDQtGBXu/0NAsOEzDROvoKPZbBmuQaQ9b8FWV2MCXzkf8uGki
KtSmJgep+2WaOZM54VVYWfjpvJenPgo5RGugSIfvZEDOankoiaek+Q5ZANvVITlP
5VCRAw0OMB+QFAxaY+8b6tJNKRI9vf5FetkgUwklO6gLQrojWNao7eafVdqf14sM
Q0W4rDaqgCzxywcA5dSuWw7rohr7UfkbhKAZ+NfIhjIdIXVUdqGSLoBZKskvmd3Y
g+dp7ThLnFNWtZLzN+I9Ess8eqm5cnqj/3zlqCtNFcgvSMbEHqcLVd/avs4lQge8
nKS111+E/OkORBgEvF/KIdvsEq6/nVo0UCtruuAXUMC4P4QAljOKg2V6Ph1bVCFa
0a10sC/DnVxIv5mZB6sb97pTuCDjshaXB6oZfjj3TnQZZ59buwm88Oby42HTOZPy
y+VGCMBFMMoqZjGbmU0tn9SDt2k1pavOSoaS1O7jk5Z63X1ZTBAyJVujx6DDDQlU
CXpifvhxOZFlNmk1+hHBT02QEu3D/b0o0V2DQJKDhDGis1Z9QDSW4DI4GU9KEcrP
pFghlio+n3cH7TNFtfOlN6zFO63DD2nygbkcPXgyyS6yZ4CIb2YcNgIS20A03Mn8
/5OrF4J5xT3l/b7bnwGsgD/TXz1pBLSHQzC10Z35Aq2ZTNbfGCYzhvHnV8YNasBz
LjMGpixn0+TYDTWqnZey88xDmlpNHRT8EbfFXlUmM1awrq/aAtI5L0lknf0SsAa1
KQoqfAFpKQTG5JUK3sRpNOGrfK25x4DbE81yF+j1pe+wWu4qhWQVdAcRrCM7Ws1p
vHrFXUP+jdz2CFch7OnfPnwpfmYS5YwB8WB8e3sdkAaQWrX43uv4DA4g6nbg7b8J
nORpBK6bjpcAJBp1XpPk6NhEw1q8zPbL3VkHHDfrclYj1Bgi0whI9XqOSB2ll/3t
10VtheE8VqtywQ4Tl3TVynN9/TFSQ7ool3fVNYLI0aXdqDr62VtZJtvNeK0zmtc0
+flEhPnJkPbZei9w/Kw4RIhGtyKPq6I1TQtNRBKIVa1xtQQmn1LcR7ujrivtvwa6
EogsCNT1E7+9tBjrl4PwyHgtKP8eSi6BDj6b2OV1nKszuPsllMwVDENdnIzZTuBy
/ZIl8/XifrxJVbs7orp7l8XQzN+tNX4ZC2uLSbqvuivqtcMusrg0lJVLFU21vlgD
PrweWlV/xHQiWBxrALNVjge589bfWIwfUp1EigszHmJE/1xWRAcxnhBIWgJPXU/2
7M0imsg5JE8ZL19XdULFeT/7va9NxGidSKkiZ/EzRpCAYMuq2ApXVWLwXLD6SIGy
KZVpyWo346pOwCeS+gtR0FgbQhropEbo9FQOSo7Wnjuh2Kpf3Wewz6q1rRDRVgia
P38wJ42aoXOY1vY0+UYOFc7mHt8BL+9MDc3q1ti/buf4TMzpjk88GDfViOtbZgSS
Oqu4bEzZmUv69bJKPrObcnsJT+CpZH5ydqxIUgIVJHCYHC7r/tTJH89Xgif/t4S8
UVd9nxTaWdkbfSHeIBVXZiP85hEY/ucdqyTf04LtjYQOWQth8MaOGPvuU8VFU0kZ
VfRsALOUmulaau3D+StY8CjIgUqPs6sipMooQOFsFtxkWED3XAijnDgaly025se/
jY/TZyWBLFftRQANdv2RMyCgDLffDLHUh6145RXuauwDegabwYG/p/0N8+J9rEQI
QJm3Egmx6YmrJe0qg6/kAnHaItj1ndnngppbrJXrjPBMIJkKW982mcu8f1bvixZU
7BGedn0wdDjR6BVupLfE9WQd6TkaA3XaKREA6kZKR0PuR45EkP7P7ssKX42PLW9Q
sYKuTkrWX3of6W+HoqDvjZ9cwbaXI6n64tQ1xXbJ9LRkqbKu+gwwhHhqNnCdyOR/
SZbkr9HZ/rN6pJezl/lp610udCOeOGEMFeE7nf3ZhLOdrCzMUwJ7IKIaCWO8G4aT
Vp4LpCVDZkqkkqOIlrWAw7a5RsnbDt8Kka5tfMJOh9DTabb6Ehag6HD7rknrePLH
ct7YfgUAUBn2fXItMfcwrkAAH+8FXLkDx9tUr9SqhITK/1iwKXqdwO/u3Ol9EnZW
CGaYs8+MwmhlBWoLcWxd3GYYNiglwfMUDYWyTIjhb2xmwZhNLFR4/DoEkLpfp/o2
EhqlJ0Ca6gxYOkOU1XR9OzzrcHvHeexGjpn5iqpC8JtLvds1FFgnyLO/s148/qY7
GzxE8LDGDd9G9II+zb8FeLHLGymUckOKE2+o1tdYDoAobwwrC04nwe65ZGsDWu/T
Enf68aQDWWwNVCsn8FdU+6Qse6FBmdosItNu8bvYA3mBvbj0KQBhuOJiv13MGZOq
LCwR0tDasnOqusR2oCGKnxMGy0gMPGNfzgpxBwS/4OiNg3zFYvs6GAuC5u7JZu2K
0taqtkzP88ZESSLuGlUa+E9+KIIqv5DKY2NZO1ykSmrrdQ03UdbvH+8uNPxZFKnE
b2VGccegDWymhnz3xUI8XxxIKwhc8RBUty3bxM+VXNGOS6Iqedy1khMBjdfVCDcq
qr4LwqUHA35Q/G090aAtWBRQqwc2xD4w/0zQjDYNz5olzGkuvFEkrjYVY8LpNTsS
KHaBFCJ1H/iiilILtKsa2W6tSLOLG6Y4zfRX3UcKzm8H3chFp9i7xkwvzPZNuKkw
gxm3CrgD0/879XjDLdE6SkRgWaOw9bXHv4sJRTh4XvPg2RJ97qMikTn9Uf8k126y
sYM7ufUjcUZolG0rqHXqfNVpTvPQ6BWEr0bWl7654oVxDMrw2vr9JK6cajL9ig8U
Q5qTRkjaR+8xL8JnYz5+VEcnHrNc23J1h4raEQ5r14bTSTkRqSBmtsciaEI3YHQz
9xTKCFEqK8x28lPOru+hrev5eMk5d67veFbwUvVCCT58b8l1E3JTzTlszRhTvaXt
V0hnGXD5qkLskSBjZ9urkt1VcGMtWZjuwC1sCyM3eNljzV/ab/OAxhmAXLFx5Lww
XxOBS0jKzDUdJ7LHlDuazejwPutwM+fHF/fX7+Las7SecsMHhn8mk//g007dQfkU
2rEH4NvnNwclQ1DbM5QYb806l47CVRU3QHfE00sn0rAU5IrCB3pHc106JvmYhCfR
AZXcXggOBOrTxLQbIgwIorAaA+ZsscyJUE6sY/aypk0gRZoOrBfOP0xkc9rQ8mOp
jeoP4naMUfRdvjz42RFoWk9bJe00t1vTliWtBgt6llD8sHowfA2pli/ek50zZSTZ
zlji/qpyfRbjBhuHKKp5QJFCJE5sl1ZHm5bgyv6oHDZvrmxj9a2neao4MKEymYGh
7Fn8fYNdL91AAEX6rFTukfABf3J8HKCLp8RbrHbvfKYR9u5CRxrXWIgitSoYA/7V
Z3luArbJMNMsh9WgX89j8jxdTNhQFl7Q7XfNUvs6LuR4haEzFzNmf49ki3j9MI54
2kkBiB+NPHQL8g+91dH1Cej19qZi65A2JfbJDYx+uBdsBa6es8aYHTn+h0oaPYZd
qgqVfS+6lkGobHnnm/3FRCxLt+pneez6+lX9XmHeJnOMXhgcwjDdc4vYZY5NiXtl
NLs99QnCrcARo5l1RQKyU2ZlmEVvV1CX7I+Ebj1S/F6RuMuZNjBpGqdqUApjnaVa
bpiryrCMQ0sEgl0qWmibFx1VOEG8ztqYpeg2kZKIGDwyGPWj+8l5b3hNVlTJho4J
9To9Q79zSgGshSUorms3Yvv+9juKTyyHhPqa8KUhxKHayOtVi4+J0LpDbOLdIDfY
cHo7Z2BqEEzhAPWl7RkMtMjwpL+8RhF0MJ9PLIWcgpLCbbUL4wuIICIdYPmWG/cb
/2oANM80FiPP2eo/dhaIQccIvrF3xU/+rzM/VsHMmYFmjVJqLy6yK06+9P9TzbCk
lbyD4Wt9SNRPRqfr0HyopFjBoH/AMAt2jVKlU4sTyxyUZ/YD+LaKKvy3oNChSbwQ
8azxNpyBcpbyTz5kDzdiAjAloUJfmqdRAntqLB9EB3THSzfDdUWWuboIjji55sUq
jUrOc/Wf6AaN99ATeJrR1FuznsDmPAAAxixqioQeXal0d/GBHZ3R+cXLb12ivml7
u6bMYC3zLXywaozMGlTJxowo4Ebsot/4ktbsKxjl3lL/5wkDm5kUlMTYKGXl+Tau
Yp28W0H7/taP1HzGpcZhyvkryrO7W6/QUW85NIVInl4bEvfUUs+algwlhpaXK1r5
J4PC2y8EWeEEQM6gfW5/4vYP2RKJbJtZR7Y4HP+Ls5rn/J41SJOVzCr3Kv5IAGZT
UnsxTIvCJgLfTf3GIGW+LvnNjeaNEus2ulcvIYPu6o/h28Vwix9ojy78XUFjWZJ4
7tVKS5Q2chge7vSrZpS7I4THITOzNfWcfAjLpEzK1LA5oPNj2NH+4y+hGdLjFZro
iX5vd98aOBofmNMIANz5RLcV5qzUb6fgFgIKHIsfjLFL/x/PYs1BPsshaD1eDllf
oEAAAUJnPFNjE3jAHfNJATZyFfon4ipNUBV0N59mVygC0fy87qBfwsmPb/DfYdJN
99hh1owso44mIzZtnfxTMHIX4DGAOrL7EVILJBNNXlmH7EjFhGeIrIrIYp0E+6fA
qdhvS6IZMPUfOeo70jyoITQ9hTSBG012ZrjvNglcmFia4Vcs7vSQt72GwcXVKfJb
rz92KT/+hqT+ZKKLxLrLuNYJ0z9QIgEBBW1l+gQlSTAvUjjh/ebIe9qjVtIeJuVt
mTEIwN1TjWnKfbnWx773+qqEErLx5nqMYk4ar8zUjyw4WJTnQcTL2QB21brX6OVx
5O1JLl+BT9RiBFUVemTxkRFSHQOkq2DZzIkHgJ8xWb9pSJ1AmzYxOrsLjar8aYri
LFz0PzbBMqCJgs8K3rCwmUHm/u9Y/ejRiCm4PWh5M2KBXXfewVjTRbwfEr5NgTUJ
/5vCir3IheIMk352tF/LFjR+Cbgm2pDhJ8ZAefeXTqbGOhUHtI4H6EBdl4dZUtPw
d6Bh7E5IWT+vltkYqsfu4JuR/+DYNarTL7tD5NMJCPEZ3rOanOJSQXfljOp2/h2y
XXH5nrGYnTujQyJoHXlPcu7wWiK1vCDBDy5upJfVTA+wC0jRWOQDgJGp5rpkRYF6
DgWpvCLT9GQkqBr47xG85Uw9CZAuCf1N7fV3VbEM/4PSa0RNAY4zeaXdBkSBsEex
Nk5KIYmlOV86EBnhAX3EDwcNsL2RV0b5Ww7Q2fnYaT8qyC3dfM4Fzyyu+XjU5Zvf
b43Zvpr0ayE7pPlow5fePHL5+sjtgBUlc/j4KCwUJap0L51f/eQUIJK1ux7yXf+z
fCnobEpZZzlLLYvo+YsxM/J78RW3lRqU3F01LSCwBx0VUjNZAw+hpOEz84J5Fn4g
j1/D2P6vX1OS9ACQhJ9WkjKraIHalqRKWjNtvZOKs074y5n80+QPUMWomc1tbs54
C6A6PpaIkfnFiz4psd24EKfzC/jtvYjJHyVLM950ysDG8SrIytKVUtxq9TO7o/CN
d3RXkKaRsHDYCARDvtO7NFsLWrkESylQB1FwxPRBw/Hq21mv+zDcnUoMQkyBdfcc
sF/Dz/Yg5KKpW1tAAFQV3bCdNj/+3XY0uuLknAGg1pCPbMXuCtsJBzzoHqmxSOv5
iamxhdz8gt8HyCgqmdFQhtnhlW2U1wcHJ4kikYCISYvsCtIFAHEAX4Opd6/T/RQh
6aYlRuQNGL3Dfko3880JbQenNJR0znVxF+XOJuLATwvYVZa4sjDGg+oOb+sY2hfo
CwcvJXrzD2Jy17TqMGagZ+0juS+bKDzSvKVBpw4YN+WVaJKRNV7vG37YNllqm3ks
nQpRIbm03amX81Nv6u0La+oCkZlZru1aSCXbNpNvLMN4K32IA4SZYp0+KTyCn4bq
nreRQIH/oA++74Egbqu1FpgI0FJJ1dS6ms7yrDHBpC9z7ktVi2QAyU91oxjaQPh5
xK3Cke5z1US6T0jp4goNzvWC0BceYcF9EPpz/mSEzJJ4OJnudDPkjdIYdrZvwYCw
uaOt5679ECi8apjxx0FiNP677dnpKkeMLVU5he8vvhZh6a/9t/EF/q7VDsKK+0tR
MdUQaSTvJLffLPM74Xdb/qXo0Awrt2HnILAgH44SqfuxnZI55SxYkRlVL1ZwYgoB
Q8N+g1ck0yjgH7PHkFfqPmO8y0NlocSwGKGw3MdiyvtGZiVPmfx5huGbk1U7sZMH
2ycyuairNuZcOcNNth+4tNGXgT1IWQvOCsd/1AuSrn6CAVCbWZ3hNWu2vmfoFAVC
iuHZwYK+zf9cRrq1izLH5+g8LEI7RJzfb0CAwOMHbfUjReds23VT2Q9jaGhpGy78
ULEQ9nVHzJuld0u1a6eXGNPcpWk/1mApxQeD/G/4SX6M/fMWqunEb3sDnwdRdCIs
7jAup5jhUqeYPSXtt1KxqConudCI9XW5ht9NnIFadlw4KaU0gEe0026EDwB6rgYT
/0elSfFGMK4V+oN7E3iaju11R8b0pZMc5BiQk5pO7wnR7RAzhttAPKjBLLkemu1D
w71GpSoCDFbeDJCEdbB0KjoQumY3Cp47aP0vXUOhWlaEcCzY/wqdvBidOuz7Ux9Z
faOnAYa6149LFq9RtEmzhheRc7xPmJGxfz+4O4xleMC5IscY6BFzz+DbiWGRB5e9
xRWxxY+t8sFuRLg4SIZW+4xSFvFBDAQFoDTqlvFsdxCyQcRsCDtNhX7uR5nTK6Jq
+Gy6OS+yGHCyl1EhyOQg/4QJpZ+sJe9gvpnt8fMnc2atsDp2gfw5wKXh1kxS6a65
03wWEdV96bQiWXyOrX3iySsO2HQtlmXeBa70OX3Rslaeraqi0fnE8CkfLIwE+p90
+s9r987QUC+IootrSrKzJZymR6mAoBn0LqDtDZueVSLPBGJMgZMNTReyNWE3hUCD
Any+X71iC0weWZpN4ESbmM0i+2jdGcX+GA3/ymQhj4uWLUWnKsXtzB8iKSbQMEdb
Pg4hdOt57zHgF4KIqvgO69+kg9yJ8xWm2XA202EbqbpRjNZeCi2i+/gfLHlAYVfU
N8FG14VBHUAY5KlXDD/Jm/M6D5y8mX+eWLZGi16GVE5oo74r87yRXXjX6dSm8RA6
J/rd5+7avd9QqLWFy1BrIRUup3yjDCIf7gFYy+IXMHAqeqqiT/5yXA1EAEW0PV44
CGKJJv+6ERBrfGLFwP2yvHHYZo4stLouSHHfySztxiWhzjqseEROOPEjBPXZrT9K
yq9kxJfSKz8c2Zqbpt7RZ85IFawM1QolcJqIlWxLvFG7YlYaeq1O7eE2MSaUeK9G
W/qbHC6PJUnh2q+iTBANjdWmq01wAAcBiRc8ZVJ55n4oKkOtzDwmV9pxLHWAo8UN
uJU792T186pwY9DHpseHI7WLHLs3lieajZZYVw4ndsjJ9BB8pmaFN0FfIcNne5pf
rkkm3Rmxj2TrmmhDuOdFj3bhwAa+mBIRkgT7ohCZ3P366YUZbLBWepNBrV4LyR+q
GK4eKvDxwKoLKGIQQi51hsUUj96FkyQTZrhT6s1wIKVRkPSGC4Kgi9RduUTfII1C
6NPYhHVh/S2tA0S0sRp7y4MA9IAn0NY1ODeYAqggS+O48lZZ1LQQf9vx5ElM7RV6
ibnHzV4K88AoPXU9nN2nXPTEdu6KWXGBRQy6EJ53jb/oenArpmRhkxIW2OUgz9wL
d+5kbN8Cz6ldoxH3UMZbUV2DXbPhjQoFnsJWowUWKM7Nn8SiUdNLbapv6kfq0VFJ
BSEDICaw1vNgzJsRCIMuSLL/QkioW9BlSX+ex29AKdLWu7Bb3PpZHu2PwehVbFY4
4vGe5oMNG7AT0kAUnjQ75wu22DjFijkSYcKsD78yL1Rl7X4ujq2WEapqw57SV50S
4zMhb637xoEFZhI6CuG4R3MvcBWaoA/ZNAEolLAqmwLuWiE+BjyYvgtqBO24lZCQ
NUb/pykU5L9nfkeqQZzv6cP9zTvU/4MsGtBmd5dtKTmf70BlV5Lr9Ke8HXgqlIs8
FUUCHEEJsiPoSs+aXQYrzMk+j08OqF9a7YdpUJcvn5QAyjDuKXYKgYEjyNiz/dsD
hhWWL3qXqbr1sWexUGifJdsQ3z0AjKztj/tnD4YIlebDuXOBUNwVHQGMm/1DKhhE
5X310X1SPy3py2MhaxjBz61h/slEQOV9MLI1VFtPB6bkC3KS5PtDM59BbzjlONq/
9zNX09AD+NLBBfor/bnHE4/AbwA6deXRb6jQ33IKz7x/0gnu8KTOnshT+yzH0U/h
GXGwDKFMpbIA3gZJ7nyW44jnMVEM1KNz0DWAi68uzbvg1RKxJ0IYoDo1Bw/0+44p
G5ANSaiYewJuoiLEK615RneyEXGmJ6zIwyizWXhBKcJb5Vcs/eD7wIepMFk5UAZP
yPpLFDItHyrV3dFypUXvGsp7Ip0xRiQerczDKcIXBHeW+cM44sGRpDi/zirNAjip
hgjVQ8Me3wO/YQz+aQNcBGs7oVGjPIrVLuPxMOAbb9MxuqydJpWvrL28oz/x3XVM
HvrzIZbwYQHyYWc77BbqEU2853ijJcb214cYBzCd7TJSwwmDeSw+eG4syeo8fj7m
e1pAFPF0MshkZQQ+Gz+mwykiegIGnJ+2eHg68/h1a3O5wInk+1+opo16GmGEAcmu
S+RT/vBpDNrnXWWIljCpv+/Xh/ujIxhQ38cIRd0jdo9xQKuCpSN7+j++Ix4aTb7H
FNcUlRf6G11/zYdJhewME3khb/6c33vQ3roxow7Ci3GzI5ZeKqcb/JUBGINXy+XT
vTPlreMjDsNTAW8AmFtPdDEqo0SLtaSSkuxc/8QCcy5lXu0mTTLDeVF1UxhokeWu
PUtC11AdsNEZGZD24F8ZgnGWxH+wvFh0HHqsK/OD3tqm4JygcUooe4pfIGgOKUkm
cpGqmnhtgkvESob4V0qrqfl0Nm0YIPujdJeU7DQFPzUbBx9Xx+NQQ0rOhnA5vKsI
otBhhcvphqnoc97ZrrG5LUDRmLXzvm3qIR1tgGTgguGE+V43GD8Etb+wvQrx6sb6
I0h4XcSzs23JQJX4mMkWU3vcG8DvIy01OqlC6JyCzWZ3bEueNpuXmTB6q0FlLMtH
sco6W8PwMFi/1T6yHq8IdsvPx0QzrdwxHwmk5oMqMgkzv44u19j4HD23LZVfQX31
1GXupzUGmlPPrJfSL63qwxARO4mCH4l8rXo0ZtxOZTRoEGCi5oAy2GlTPUzs325U
4jILpKWYB1sFj63HfWWxo5dySPZvAzpHWDzeZrfxJaXy8BY1JsVl+BqPg7Jla3Mv
tj43H8BSKP8K4ljMSxpaFaVQ3s/RXWCwM5K5nMNux3wVTc2o2RA3t6dehD2WaZA+
EdPE5klp85hFakAFH16xb8lzOvDm5KyeyRKzTcuWCUtfNd90eqAzdjkyRxYb0Woj
Ft58L9nHZYYHxKa94RDOQUsvIeh+dHUD2imYoFvD+Smo8JwejcSVoFkN78DsR5ps
OJLalPTlNoXJygHkPkjruylkPTYvgQrvaJqznkgBjjtJJjhDOP5WVOBtuI5iXFUy
JDz4y3rH8CNd9BYMfxEYwJMgAnZdCThb3QIN54TI/31k6l9Zs4M5wHNueDZ7H0vx
pfj0Z7nkWlBCWsW+dzAgyyel7Y4xBkNpKGciTSDd67iP2VcEl4Je3AJ8vYHf44Zx
Ucewqms3w1XOMxzRMcFA8NAn8B8pi3LnqvIh6aEmFDvpPFz+YDOOIeoPPfio+57w
J2Vjf5NhbYvRnrTlMOyCFjsXpIMEgd5z4kq4IJugLflXroKy4cPors1LYAiwMuby
fdVsH4k9LUcKzHdFoiWUDBSA4El+dARy33iNDuTttZTGFLRRwTLZqCP7z3VrSh/h
610+k97oMwoTwGlj8DS623jvCTSxhxf4Nje3xsiXFWFiHpfCr8buSi4NvKr2zo64
le09q6YYjoYkgxgwb7sRAKb2zznklTZ64Yu4EGEGxIeyBlvtDFd7NAEmTerzT7SJ
74wL+1IfqnHwE26PoTwHOX18FYSdGkaxkLxNxh5DPSZ9KX8dO2YC6dK0Bcdpdf7Y
yy8zsBz4Dvx+6+5Qb07qJc0mh/2d20Cd/HKVIEuZK0yqB5eX+aNQ/ADdY/puTEDA
OzBuhUa3xiPn/iCC6cgHPpFukfX+p3aHC/AsABiU+a4nuVDgn9HNCFk+DcT+UBHh
VBSyeDyblB3vBQ7wcsAmEh0rBxbHRX7LvNONkDGhE09bfhN5WgavX8R8CQHr4KO0
yBqCSXFIyXcOM4m8sObI+3X7NxqkmWcvomOJz3BT6YBXOyvxiIXkaKHdbzNT/cX3
3x7qc9ixgcgMErPL+CHsa7s/6guy8uYXHI1D7Z3yoLJdMSpMdg7FQkXTO002oatA
ApoVOoXQ7C7S+ozz/A3fh5vU1rOCRJtWPBTjEjc5Tb5AH2KwN369YSNncXLz9cNA
IHUPWX/MNDK0kUfigzUER6Re2YdRXrJM4a53YJjkoSSIGF8K+bT0/dHPpe4xb03I
/mDtV+5Hg/FwkBBSMumB9sQaIVf13imYUtaMv2drweZc6yECG9CxrfcYau4JyJb2
VNYENCL4MhR1HXVZvwfcw9RwJT8KbTOVPxYPXsegsJH3qjb0dX1bh/9v9zReOTGj
VqkyX+pUetJV8y8x7Iobb5gBZHNFhQAwyJHM62HEUdJ43dZf/798KCa5qzIYDLSw
AQmSvL8SIgL8BgeTi26aVqGKL4Z1+Ad5YoC0VDE2HGXTL6QP5cG0UIRJeAI32mKY
ismoHtnz2FdggaGU8rblQCfhE/PQvyZbrJ1jsJKpL2SAYAALOL+EFQFowg35vTOZ
0EGG/OC5+sbvl2IMtCjlCSCEalIZxlxpzgvM5+uwD9IRZE146EbWAEXt2BCDnHer
bj637obJp3OW/6fXa7L0dfaaRcxVHu6rI/XPdspX0zF8vF/P+90ktDveEsVTgxKi
O3PXBzxK5zc+45LlR5gQ/MzSpgrcAaWp6ybVCqal0eRHTU8gQ80tvJCKR43P8diY
CArcev2cUIN8XZv5vrCBc0FqpHvrsP81WenEawT5hIVZHTnglN0XoL/HNyzPywmY
SSjOc+jhvhbUdGvO2ZhBcgbRlNN/Lmp1RCPfD/NjrC6DaH/7na+1oremHih4zERl
DZ3AqlSCsXgLB81SEf/usW/UhHQl+HiiYff/+TIFhT6vXh29YSEQr/yp564DMJ4U
RxPsDa/7Kkzv0m0VcMJj4LLEmLU1lDjil6H8lSfA6t7+cJvu1mehiNzvOA8Mwqjo
G3p7gdcg6tiJNpRrkdm4EF9AxVlTZGAwx5bcUHPsKuMILvsZ6BTmdrYAdseqnj+F
HRGshPpwvegw9Y9+wu6SkhyY/GlSU50km3chVqmG6JJM8nGwzzBzp83u58HBW8rn
bmfY13i5arT8vUIEt7U09RGZ27ipxgLbmd4bRiG0roNVQnEmXj+18FdOT0FruSLk
FuImhin6BGZiJ33vel1mKKLdaGWRwzdY5fLbgEcmgAF9pm07PmjW4jVFw1nXFjsZ
PHw2WgrJXCipXJI6FfJXfa0CcSVoMZBCEKlWcJ4y/BcoxKDZ6dTekFu/OzfZvJ4S
AGpwcJbcdtC3gQux5ybU/US29GHN0Gl9T+P6XK8XUB55WVbYAHUentTvyjl3XDi3
UO7iBpDl6vO8PAwEh2iAjl3vsF0L/BhqqH1z9+5D58kIBt+oIgMNGDoK0uGH1466
KfgFFqTIjCVLLpcV2dmOnJb3LCETOhSV8DDc6V94JtRCt2zoGF/cBfVO58pp3cWS
aHze+fkmHtEzLelWTD8i8INfIcpIkRkJNn1xqc59ob25DpDFHFTghv5WgpLxUSG8
/EpsoOzjKNpXbBrmRdsQR8w2aOl/nvChyKGePQxQre3lac3+kWvrw+BXvG9RrFNw
gTFULgiS/YHimH0qbU6z6HkOt1xYvjbD9sEViFtJG9zDX/LuPiKR08VWADBaWeXK
vFPrxm9/NAtxiUyeSbl1Pfu1/O+b+fxOMCXgDp1IK9/qz2f+CCEsu3BZymvTDgNd
LuJ9stOokfJ0x360z+wYFTL3GJOrH39UnAm5b9WoAU6fcWix5mAPfqTU2xIiWXvC
LshvGmQK94OFMxmTl+W+mZumzG/yGnbvQBfiPbMzLYJYyXuHC4PfScEWYl2Dhq0R
HBM4GvbLgbTCNaZBNKpxJ8zTH2WVNrJVad4KAREsKLf6klFT/UXPwykBscG026aN
wFx9vIYoO6/fBf+tEpzEH2QO0R76XxTtVToZx5ibFrUnQSLRoejLYEFOf9b8GVYb
/zsmQ6veyqBtrIo3fxtttj24wv8CFYOyMaMGDnlteso7GN67nXRD6aTyJqrD/ujn
jET5++yvJG/Gj7pjPOBHsDcYm2RARON/u6bPRcWqwFqMvmcA7T8YoPtG+QYaGEdj
ORK/gMlfaEABgLIot1eZaj6pUWs9ahSci1DODSY1cMjnCPcH660uSD8DJLNQ2GLx
4dDePGhEkJxKMd4kej2fQuF1HkkY1PcWE7hCWBa2vYYa5icIgraOV00jDwFz0NYM
RigR5j6c3kRbEeqAXiUXyJNED6CmtWFCE59i0afAS2UUEojri4Xb9Tg5vVny86Zb
B2U7H2H+1osKA8z+SUmUj7rV3grW8Yo2W8CT6Vi1Cnuet8fn5a5QBnuTbpK+vz5Y
pUrTpaNS0YBMYhO0RNHGd3OS47csYnxyZ5Rkf26IQ2jZhRtHRzdqlvVyxXI1yipc
qhuKryxHgNpUThJ/ilukQyIfTriXX5eB2twAB3sXam2UJKc0CJnqdmeaO1EHAk/a
52Dp7nmDeDomKVcbz+1rZHrw5TvKoVQUwFciExzjLuxAd9DrUYucvTNw+FRVkeHR
PjhMwO81Sjvi8CRMpBDba9FnxyiyGdEyXiCJBHVEmWmVMdD7X9xVevL1q82rZOy9
PVTKVWBL8jYnBFkTEvAk3VBy5bI8dJYGBMKgX9uyOyCNnevSye463LNZ4aRMtpab
LZ5m/o9p9YO0Crs86EZON9zZGV5Ly4T0zLbsC29asiktNo/WmhNFJFtBxVzzwKoK
7zB3ORjeS6rDaoS8o+juW31nab3I07jVFvAOMwUmZtutEe98UObtmWeu0RRbi00u
CntAJ7e5JqKn+dB5q+mBSB2iUmJMHKQMh0bMWSPIWL96Kd3sGQDyTy7qEMnXG3gp
qosXty/QNIYzev5TibgbVe8FVdVaOgd15TDYl59+aK4m+u5cqWHQj2WBHT94fpgI
svdIjFKrTmg4l7SAPjlTSg2zqyPwYtsXDL+DegWFS08sG7fUJa1atxltstxCNvBK
wsvgDLP37K1sZuRGWCkQcLarPO75PL5r0ZrFsjsgQjdmlWLxmoT1mTPP4b03nfgL
iMKpvSPXdrka1Txt6RrQdHEfbwhV+83o+qFp1yQRoWoLa26RP7754/JSj0Dpm+nm
BGcSRtn9pTuudhmpTDaQ7ywypXqeULB9Q7h8v1T2+IIDkY7B2M2Lw9GYQ/s3KcbP
a9utfKy9dVHDyCg93fdxOxI1bV5JHZbLUwZtpzkh8Ez59XJ7G3BJVLF0gaa6fejK
mVuHkEefx17fuZg0N/TGSLAhJRHdtt1Dtbz4a/eMFou0jLCQKIgYnmN6/umDN4KY
46urja0VOBU/v2qIabl6jt7xz/1kVqRcBeUh7Pk3yK9CRnpOhkJIH3dmp+l4tYnJ
cBTH32qG/jLZ6g3Te6Lu3osVBlzPxDQMIj7AgoFLhgbCcBitGnr+3h6SQNktUAti
oNDCI7P6VwcG9FcufOuDDvVht0KF4LnDgAYulo6l64cw42YGI0btoSb6ZAVoyrlf
wplVSK1r8cFxhyLPBNPYb3s5bxCLBgoBsqot4T6+Z2wY65/4fAsKOK7QTZ93+OhU
IydykQZxmoNvie+BSgnuuzqmcgjGzno/iUu1sGr5+xlM/pMSp4U7+2E0gig7lYxK
h18ySYd6xb30Y8wENBjE/vIEO4+KpdQ3ACKso363/fgjek0YheVMr0AKQHXfjdmY
uOiD/zrwCVySuRZOzb4et29zuq5k0qeU00fo/ZHmvC8Ya8clI564b/R8tbJIprF7
JPp9LqUo+SxPMu5Ywq4NpERfT8bKmXknPuIL74RDzDtAEH2fYTwjF2D6N+XTBIFH
NR33H0xtocOZVoGOG6+nsjN5dbgGgJh6wdwCbj2hQgUCuUbhzcVv16iARYlSvs38
U1x64eFTTJTE/5lbHKv9tu2xREL7CwfGhqu4uvoFITJ+2ZhGwcOZAep2Zc1H11K6
zSMDRtddwcfzzAdeGVQ5R7RiHbQleGYzasH1Jiy+P85SEVQhm7QGs2DhabReJH6u
ohlCNZWzST5Wrij3quSeIZXcDmuL82Mdmuki+WzxMT0L/nifwEcpPVpF6ZuE/s0l
UeoR1yAesSISjMRGtxXJGK5KcChhNP+V9GBSRA71P82aIOr5ab9qo3LwRbKgF6f6
CTax4Hy+qnc1xPxCMPTxsnSPva0Rqzo+1ISPBt084QbQ8JTvlD4e4trqW9PlIWKD
LjXaPzend6S1FsyHhI7pp9MY5NFh0FFyd04OBcu6QdENr8jXXUOVwaGNiLdLU4ay
qvfN8371G86UqumCy+/foXk1vBu9Sgu71KXXioAJl4IKsx+QIsXUJfIMhKn2z76f
UZYvRx2PHdsgZ0S38iGzoQzPIVy7TMBBpdQtY4+4WMob7004F4+liecnAjWHMEiK
WiXD5RatjtgbDXF0zHYS/u1b36zG8qzBd0hOyens4J2Mrli+tVUCBLocnQvxIrVb
X32ux1r8Cr0QfcmeE4DE3q4PUp5fF4eJw+H5eVGMttATFGPvt8jxxscMEwAtTasy
fTp+G0NEAo5VQFUXK218ZN2QmyjrXkSEYXjrvl2L9t4qbOT+Mv/wHuzrOEQesu5D
KNAoNA9InTpQLkxOSFcWHbiQhDTbsN67bcUbV/EizGRORTJNexZ24KA4AF280KZj
6O94PrRkz93E3LQ0/arbrYxXd3zRSdwr2u0neZZP6MzuDn+YaOwUuEtc3Jz9KVqY
XgXoee77maKWPcAi3tLcRgpLpG48SFhb4zBysDL0fFxzRlS17gu5BETcE/ghYgLG
b5KcXcTohi6OXBX6D7MQhWbFvdEKezs71W40XrEZoHihykV8wyugEjF4bcG291xn
mhPIopx0aiv1Ro8szzuG/KRJkTwO5AwIrBhLH5L3nHwPebI2zPFY/CCSaLT/EVW5
MC2DyGKlArhU9NOUdegwoszgtFBCX+o7Te88Vdfze2Kks7NQpLpNrAmgGtb0WOI5
hMk2GzWBzE1J5q03a31p+5sbG7AE7D8Js/hKOn9p3giBdTMlSUTt5Cq/cxNLzvbu
6C3anMOTEWsGClcnnV6xaiz9iQcRlGQ5h1ZvJiBqv2zyDwITw1Uxvm3lBRNkz7h9
8JVvd1gTcCpN/Kd1kJLy9imDJwPj6vUk1AJSi+H12xgRX9aKe4gHtYFuz/wQPoBS
MIPBsu3td3uyIlc3Lr6ju7yehPbUHCWGqqLQReSlUAqrRb81LQOA7IN9pXPYKcT2
RZJyUCxp/S9SvkUCtLFJm31tYjpDge4VzF4HrvjHcdqOoElR0rjiBvn9bRlinrOe
6tqPD07eH7m0mHP6ijk7f0nLZcGFQ/GSd9whfSxmB/NyNTInaqFB8wqhk4o/XL87
OEAFFTDd8pnHHzpFLMXJH+QCRs39PnkEJeazuhQDZsYIDFupnlV7LpZ8VEK6xcS0
eJu4f3r0BcyuPVKTpkX8yakUyxMKSrA7sy7F/DqjCDfP/aTmLUL82VRWVegDJQdk
UHDUFuwGyaFQEI6QKnY5NC7zJ8ITms56bcskISTouxO0xz8XJ8HiVyNPvg9etmzR
gO7HlsamX5S+r4x1DYSGco7crox2lPR225vxKJEas7VxG3IxCGDqZDQpW2jhj0ro
YwgLFWyhqmxo3bRGki4FEBgKPfZALZJEyRTQqvf8Nkf8jFcgeqDQaHJFJupxAyW5
I2kh9kI76GTK0hFivhQYglCEaBW+TrOXCQFJT98taeFwQ7EZCGqGJ6wnAmCCbQqe
EenHB7KjIPm3w+mOup11yOG+JOQwYsQsH8vXPhHOJFTWuGePD9m7poQUc3m58pVh
eJ00gfS2uVIEab1bSywVCWia0KP15jjN2vQihUb7GJrx+ppM0h8mqYV2DZyCwc7a
rI2SzdJ3kT8zhl4okusHWxju7i4ICSNUW2yyp6+KyzIKLlXpKNc3526a/Pe2GJmY
NrB+iwZ3c0KRqQJGgbNMeRivNKujyjx4DQD8PaxndHgxLnuWatFIOFqkKpWgX/Oj
oPexh0oc+e5JYrkxeIM/2p4xTw/FDxhPO+eqhZEkPQ3A0BcapcDpUkU3A8GexVgT
bVUsppFQjkO9JZ2ExCDbaVIdIKgSwH69LRHgiJdDn/Lh9zoYjX5K3X7reFPbcVGG
6TAss+OEog4xVJ9V9aGTqD4xs4PnaG1v7SJQ3HbMmWyOzBs8cR4sDKiO+IAYn87H
+yK47YPMy2PH6qD9xfLQPIo63F6PxiqL6P8gYKFajkEfiF+0vUrSozjPQil6tYKV
6qxSKJnEuypcyzdGoYCR7EWARbO0afd6rXXCcUSkK4zAHQNMCeBH55kmAQv4fBt1
I4ZfHJ1iWP1YMlqL0mP84as+Xo1npY0WH2gne7E5XEE4evXoz4P/dGuOdpuUfHUY
QivIp07JW0jcNuXtfkueCGcXBFUmPgFFUioX0gg/xiQCyh29dujpj3MiBoqNA2NM
EBW7xXdQlxvZWEsObF3laOavO0yVmHyc+ujBevGv/gwIYOPgjEC8b3rvIy4v+7sw
xlqLOXTWZNSfpkS6gE9VicrmyqU7T8PDCu/mWWAVChcppkDMw+JD5iTQQuZFsdG2
wf/RnJ7/l+577RzO9q7Jz9rHTPsZPlTDVDOkEZezOfGLBcBUZhVYq9RIvRHy0H1D
B71xRfEh3iFBuv5fLAGYov+igzdZFe0RUzaNwcbYXRJr/zMVYNWbrRmLYGskTB5p
89e6LHKacpuOXe7TebGEiZP6qNS1mRmX4WoevOY1cOEQaPLCQ7xdvZjPl1ib4Aek
bgNPAnDbLPZnS5hBzjaqgEuOdSTlCp/qAi2Rqp0NPpC6yG4oHtqKCEzV2sNmQjK2
toFoH0gVmqiFE66mdSBpNbBtvCoxyofqs2myLLneCqnIC6wcyAbvoxnw8660KVn3
K2TcI3AWsURKDXvEYGY4+Zz7mAhOud5FkWBq1p9lyn6S8Y9A7PloDca3a8goxAzw
kerYG6PfOW3jjEdxDyXJ7R7rBfJWjdlnkuQKVa1pOk+me70fYkMqIIlfZi80iLIK
TE48VRXiCXcI+RvPvqqMpE6QN8wSCxw6QMqKHzO3xWWUKzQ5oA4kYZYdxYoK5IyI
93s9UkPoMZ085umFo8XP6NpJXCeJFfsZ3WqlivHkeDRwYQ/PDEKfzA7d1RY0IfOH
hS4kBjgZgVDLEghdiZa/JJmUg8Ep6NAhUPOwbfSxlE3/TuXTqygbI/pn/TD155/4
H0L2qvmWObaxZqBOQUXk9WFKthPYfHBiDvME6FWoNOV+6Z56F+YSrdjcpqpgRQrP
x3XACSWZAhJsUTShfPRRxu9zZt2JGnrq8OGnp8mvqEzkpDwA+tIVhTMxkFoRkDWP
3XVhYbt2JcjM7s+OaRGmxMoqaGd6zH9rphacXNrL6JY2zCaANoRvWKAkgGjJD54J
AA9WkAJXwCfnyzbzEhDwMS+mR8V+acJPGmtdOf/iggolUC65m/TWwyIxiAWAmFMF
nQbCrhSI2Mc2nzt/JlH7Qfc0uSMou1GBwahqbYyAc4HUXLZcowbfnSVm1Qjgr1/T
4Ve4JMlNgz0TUH1tNpWuZicDWIU/OuZbK2JqlNzspptgikZcHjDavhfx/ydPBTGv
R+W6FYI1mhFuzfLPyC6abmx3+g7DRCBPWu+gkMgvm4Ay8kLuTwNs1ogJdZVFPTdu
fwDu6k2PMREgxNTX91mzphZ5lO6VinlhzMnukBEsHIQhy6xldaYXw+SYU3GBrmgO
mG5iMsijNkpakVzZSQyCMYeVZJmEJUiYWmeNgBcCvfQIQBh0EDRXnUwZpor/ggc8
YQl64h7v+4Y82wdMdm4vZ2q2Dqf4lFiWfo+5SuTVvhU/9MDqG2vLCwjQ7d+vpxNu
wM33XS8Crgi2BCCXq9DmwEp4yYH0uethkpW7Jlxmn92adoVYLikfBtvH21pKl4EE
jyAPYpFptONqQhPD1O96HCa5dH/SiWLseuHvyjO7jMXUVe7voY7OWQxW8DRoMgYk
uQbdU2AKmoix3sHyPx9teAKjqjA0VU9cDZOBOEdqJYG3Oy7WwQ5eeSGpV6RDrGOg
zEsdADf0vZNew4A3FqAY11XWbUfW69RmtItYIIAZ7P5LQSJnA1aBKrbg2hCBk4MQ
r1AshGHEFjJDq/wgtpui9lD10hj/TVFzpvzjWqvdcklhPI2SFYQ3gi1JL6rYhyMQ
n/Xzmu9/zQExJy01xQBnUxLa4S8zgM/dyVxyXpIbNn1hfb8NS7TAuZLR0WuwSymT
Qu9aa1PGQPrf1hXt6EIvN37TNaimg8oKe1UuNg/CKfU2kCtMahxHAFxPP57znWOD
8yuC5c0rD6hyVuyOuFyxbZRj6bmb2kcLQKSZiLrHwGYEh29KzHhBYERIlkKOmPP8
7Di93/PIghC9C96h6aXSp/X/vYbvafDCd03Q6oJpWQFx93MQ1CMwMtnL7Qsci7I+
bP+6oaWvTOqUCBCt/QKTzU7s4ucvgZUx/vGT+nD3gdd1H88YnKn8miMrqzDsrGDB
by8Rw+DtMGpbQWbIraqnslYra26hwaEX1CFt2FtXMAONeGSeP7wcjtFnxKG0TZJQ
cOJzHV0tvjzUIgii/KwI1jHzDH7332pdMeokEqtR/tQ96DA0A5ZeeInny+YpMTHY
MNeA1fdqTJajFob5surRwYLnwVQWRduEiWS0v8lQHj+38IYm62TtCI+fEMIrCma8
AcjRnboYumcgSeUm2YIdYMBn3Ul9hCAA1DQzPzZQE84MKyKn6b6SNuxnY0kgodHM
6dqMqp0+MxCbi3OgpfXnzZAZmMVtNFPdJsynVBURvA6zeum2kLJDspf332yO3Zfz
yFT6a5mpwQ12CjOumExWF/dHTaNCOm2Yyz2h+9FUa7msjrOpvYOhdZ767q9G6Wr2
5eQftaUxWXzcfeuJ7q5d1svLikz6lwERgH9CxHA8AhjMtF6B3EqAIH68LrvzM8vL
ZGUNUAD/hoFLhqLUSzwgYd1gN7UIRMh6t3nTQMFlYlufIYqRJ/X1HqmoBGrKgXzR
I6Dm6uRpUQ0kEPAI8BNbqAwfWdIVmQTCKoHu/VX0h2rrzasqCHIoIB/7I0SntCzr
1HDemXTnOjRDIFbwB4uFp0AvJTZJNUIHxnzD9mExHcthfFxOQcYg+6v/4o5NyHlw
YLaZV5+7/A8q/m9+jZlhNxuZHuxjrX02zZI6Ugc8w4UErgfvglyZINrXLhWEHpw7
WjG/zwK+AkXHNeVKfNFxHxT0c4+1GiqqLDr9Q+2sYOVQ7HDm9VTYpWeJCi4se2PI
6a8/lC0ALupFdf7AnwhpWKmmNTLzTrCE4KgQvDch8WC5n7N//iAhNsvg8eAmuijM
eWigvkFNG49JsFmtJABN+oMDDmhdzks1Qzq3g6CYHaWC1J/GlYPM7AvqKidHjTAt
+5m0mdCFRylXjKDnISXezfmWBum6MRQl0iI3WIdPO/Lv8aHe3HqWGyQ7+SqDtXOW
PpbM8FltRAMiiYNofUi0UqEMeyqHlBxKItfom5NOrx7gMLRb9QImO2Kvmx3U+iwy
x7kFCvxDTCcErIb+AWs88O6AF2yJO9HX0zgIS17gufXuBa5cwvEzdFRwldHVMeyk
RAEmJno3mNyyE/hiqtFFodg4gfjIg33MpgoLYLBIsNjWUNSSeFeJWtDAS5PexL9k
6a+aC4FcZVWj535xM6dRTFAwRBRV82OVhP65XOtiZb/FKfIkDa6RncRPXQhPM89E
kEZjhXu9DLEhv8I8LORdn6WSllJFCqdZNnp1gXag9dH4wN2mtArKmEHLL8845UFU
YT6FKXlYlsAaD/j47gSIXR3X1jRLX7U1C9o0Ly/hWHk96e6x1Y2B9sid2XsqDssz
KM2dr4ZOgda13QsY3mk9dU3kL+PuCKJBIzJ32xQBxlAh7uEXUrm3w8bCMJd6EkYU
OUJ/NURb6ATPqpcUWstbEIxyFCs1CBHNtcFGZF9E/8uXgS+vBH20tUQV+UXA4v63
RF5ZfzR4/JullrbvZwgAo5Hoxbuh8RcfrcP7MqOhZs63zgL7Ca1rb+eAfguNnu8E
bb2GEsB9LgYmDkiC/LAXnzDgQITIWemrLCx8aKz4HRhM2vMDELEadULGv9c6BztH
W+EFKM+HfZNlGTNjZgj/VlE0/mr0ZNvfnEG6e7ruIfpR0/pODG61mLLCHLwtldwF
r5MEUO5LSYjJLSZaLjAvIx5pliBwKr6iPtolpw6V8wgCtGu+b3cm6GX4uRUiXKIx
3yEmgR+aWlbF72pKcdLwUXcrjQQjR5u/jIVPl9/QdnvHGHcR/N7DNG51KJu6Vnl7
kxfkFVpMPYq1M8nAOXiXAbMuZ9I2a1UAWJiuJ3j4oRbUqgSf+EbvTsBpnm0bxiGR
jgIlor9isBwcQ0KIUlqvhoSgBVd5Xz7yp9kUSRKaxd3xwNOSXkS9owRQBwFDk0wB
bcaUIGK56FwColXE7jy86R3GEG/p1bZoIQQOkbcZmBvfZQKt5pZTAuzqHue9Fp45
AL186bdyABTfwPjzB3piEU7PR+pAZjYrrkwvbkW73eblV2k9r5kGFbAa/wiEVi9I
Mj4MTP7KmTjyK2BVb7oNkC0URzAKQL7P7SBPpP3XMHp4wAqMXOH+hUEvRDluK5Nt
exShzhz9a5u1Kh5U1ahkLuJwjZ2Urqt756QNLK53KgqmqLVYi9qS6Zr4SsoyJG+T
2HtJMibSOa1DRg68eHonkTmTKxxsQ7bTGQJjcEAHFJVEVeO3q5v4uVzGL6bgQI+v
JoNGZntjnNjr/qSVHglAB6IsVqDE1NXqeexbfAMn1C567UzxAxl5bYzU1T6GwTnH
V9Ud9jS+ITPSKPFRFqmHkFYBt+GZDbWswKVDAZ2dVaLzOESLFNLF09IU9aC95Kc/
wYl9TR8mgujxbQCBH09mZ1TrjQeO/InnqOO6BZ08HQFKlGasIrp4+9DiD4xnmwBy
bRg6Yh6iE/D66WCRn4LWO3yoVEsq+ty2HAa0rkb7UKfRHRKc+cmZbfQtD7QARLNR
XYAPYJGlzSxO5KpcE+Sst4XfxA5WnIBjLYlD2GwbvwskZdz1zotPyZGvCWYOfJ4a
gavV9Cec1l9X1F33+CkdtdTpk5yvb42TZcnERXEC/toTmivEFuo42R4tB8qDT6Yl
oldvYpmhRdLh7FV0Q+4xl9empHuBsHdFE50vjvdgT13tIn/4+V7YBZM3enbCVEr4
26B7QeffYcJh1rwftey02N7zi9/oHTxaFT5kIH+pOUXbrkBSwhe+Chzfud4YDYv6
g+EXD2oP7aR9OyKbakRy7Dw2JVtvszw4MkAFhRcIa8l+xDkBS9daZvPY4hWn4vK9
kFpyILvS5upchCO/OP5A+ietIr35kR00WNXCYw/K9IMJq9ZiuRz1yN9SdUhF2QHt
1eX1UC6xfx4jAtZP1FIXX7Sg3NRunKtuaaPForiZ0XLDuAv5nrGB7Il2gU0SZ3V1
THed7o8VX0jtDeEOu0fcOJX8ikvtTcTkH17Py6HHHpORmluze5GTdWWsfMdPVv79
/nDqUG73E6/X3OBibrckUzipcNQWo0n8Wn07Shbt4jnJl0hxGjXUw/tc+DagJCzp
AdE0ntuKkLFwWV3Ic6cUcc1wpzJhgZK+P7U9h3nnTKbLEAkiDwTgJZmWvbKdZogw
wtKFRiKPUx0+PhLHFE7rwO99m1h/X7j6fwwXdUQx3OCbLD+ezIM9NVpRlVgoJiD3
qG9pwO4LiCPfbcMROTX14gs6DEad/gNzb0pMwtfdH03pgbQBW3enyJNehvTXmsu6
AFkD/7tOlbcAeRb1K4MTqDtVEP2RdikL5VmVXf//dmDoq+yqRNjqBzmSURNOGazq
mt2UQXl9ojaRHuBm91VSBpDa22nHvmvfMMdV0S9tEox6IAe7Z+eGSK3yOFEc0yj6
9s6wrmwqlmwV5N9WUHdbJcPEHjW/IrCCVcl8U4dWaio90eJKpePEY2xC5KHyYQOL
HzH6xXclIgy9DnwwridSXVv8yyT8+Ud8HPfu0vo3IcAbrak4GuJ4tLF57ZSxg5iU
+u9+5iSvm1Llx/l+Lteexeh+fxPZmgrvoOPfh8w3EDW0ErDgV7GdK75MXYx60uDQ
UwTqq6cvJqdUjCBKpnBFjOfu2hjpfQoLzgyuqMM4qHfM2Q5Dy57fQhYXsaRSpqAe
dlvpkvSMpAUCNjbkHogGy0BdfqMvzUQsclRwVhK8CT4mG7wpm+WYESxXjZw9lVcL
S38st3lkc4CqE36I8dZskWZp7ofobrBztEwwNKL7JsmkJnfJb6e4WSLBnzbh0ul6
Tm7VF1uQzdQ9ZkywpHYOklN4QfCOa0RNlr1bZSDt3GflKILInoM4rDIP0QsB7W9i
kK/7nSfGYInw5FNT3DFylWLUbMPHO87ysUZxHw/cdf2veE1DHiYbGNcHfM1JbgTA
HaPdUOqcZKhkaPQmxCC0mRHyQIQhDw/ZMht8mZ04L0vOL2S+0zSzU2TFmwJ77Mrd
l4FDYQZ79zPUl708ojPX1A8KeSm03CEA1yTuvxdmjoIOVJjbqV0b43jR0MGLQbVb
woMFW/OXwk+ZGJl8DHL3ubp0kc9HH2epzsr9ziAPngZ2PNGyOMxEywovxLCRbiyP
55ul0MYoGUYf87GlhgPAm3utsKFHe2td0jvZHbXKcdJjFwvRfWNSu6RqcVSlfL2O
QqvprIqWzmRYIHiXcO7LzBzu9vjHPu5IldYlSc34/Pi63hYyu/yf/tJoZ1zJjCZe
r+yTkyrXALCjuq4l9EajqBl2ZUg0riwgCdtO6SwoKqSHuS8vfZqJQ5L9EwZO18zC
wjN3cSlFxNEEexCfIQposK/XLy5QVCIIkesYwLk0mykIJf0xHnbSYJYhMgEmkP4V
Kx1TLN2IHlWE69AbJCnfv5tctmaV6pRUHLWosbL3QGF76hGqn/CtDhhPtVpTXNWT
o/mQ7mgxys0In5K4BwU8gM6vLT1SyfxJPhhejTvfSCHcTe+Cu6U3SYj3DfF/dsFQ
s3bf54Pzx3nKrJh32kprz1QDy4BP0ZMg9ObQQjXA+s+Yb2GCUHjMMjkE+zL5O3A4
UvbcH9JcRjy48y/C2/fBA0dU+u4ev1WtCaZy8JaY7fCDDdaQrn7MzjQKhauRZN8X
F6b54bbPS/XJgSEt0L1LVqU8Jv4iWydLtq5qM+3vqaG1GNfPFusL1ZOo7VJ4A8kn
j80QdDChQI5jQ7W2NFuwA3C63if6VhOXObpgCXsOzjXTWmM0vrzxlM43yPBpRZLH
+HYYBIdqnzV5F8Io4KqRJ6ds1UPWRmfn1FVXq8gjIf8PNziPj+o0N1xvPJkmSb2T
q5irK6HTUc97/Ru4rPIc40zPV72XaHBQQkJ1GdUAcmy3mAvVUZhqOjZqDJjZpfRI
p42NhBrQMLPyfJi6cTUrg1n5z+BZtnsWPSRVYjcaLmXsI6dAra4nB7osx5XCLrMl
P/AppiH4T5A7tZj1wGQwkb//F+kY4yzxr6M6Y87zV47LpMwuY+tPECc8VxR0g9Sh
3tIh0uYvTCYq9AUPBduHKY7WmMRM6xIfDufum38ln1gT3hDoy0LEuffIPLRwIAf2
sojGAivXO8c7uRompU8MXOa6n3OULArQ3eOAzQEEj76fLWzU1p+LrR1u3kru2W1D
qC8W0M3xCgGIAgqIYIA/saaOFbfSCrcC2Z5K94GWYK1W8gpGz2NiCMMzNdTjPG4v
TTwTb/48DmdRMqhxRwvt1vqnfwU0iTRu4YqwnVVGFUDdMRV4TExZdX1M7TejcajT
I7x46PlSMWJEPV5NkbomqFDc+UpLO+holapwVLnQmleSwu5Juj2/asR7IZ1bXZlz
Iyu6ymdDkkkU5yDrbdygdrw3lJNNLraHc/HUgPD0OWSA+CQY8xJF/ScMKVtwIdZB
XaSlRbUnHCYKInJUKyR0pAOAAOy6XJG8T72nWq6Lfq40O3zyUwNu+1BOOqZVnt4p
YwPl/b6PkAK2Zo0hk22lqW8sSOzJNnNyR+svJdjI6KW9FrHSy+6W1LNJ+71cWZ3x
Px483KyDl4vYU7DE98xasQrQwQRQIyzkcRXVeQBb8QYa8BQJ8NynxFLWst50v6md
k6jJyGByXpKc3VJsx7QMgjwTu/TL4KaDA60G+8NU5rqot98SMKusMkuJMICz1tas
cdUZbpJQ7tM7RwaRyOiLBWosEY2niGu/mtuPTnGk7WUxmzBhLGUQpXzqHEWlRhLp
miLWTP2Y1Cn58EVoUJKUaunMDxl7te60tkD7Pqzaari5dDloCEU8g7x3PoxPpCo9
bFVyAcS/ryRFLeYpg08lyZEoBNdPzBGSm2FlEjk/O4E9dxJ5vAAShTrqYBDCzY07
iHW2oln2ohOQkSzuMp8uYAYZKWPuOlL5jfeRARs3wC6KRNdJBz5KlMu2ur3R+ze1
r59e/BAg8rcC+6CRJaNi2ZMo8YdZe6uNMCR4EqqyuutVG6b1EfayPCs+JRWr7I7S
KcieoKxosCS+IUV2ytI25gjof09M6aztwin1TawS4ZquEmx+6TvwrTUbX6f+YWT9
W1/ZopEb5JWZQjsjQyytH6siiqv1HQKyu4cG2A4ENQW5ucX3qwF6KWp9w8sJwplo
7icaa/dn/FoRliIitTahOofUIzYQeaKkPsqYJNm1hLOG/JLJGwM6z3zaU3EKEgon
ZE169oKXgGlSbz3vYl1TC1TVenK+ene8l23MHNwXGWVjZxeiCVao8nc9zQmROL2i
tB9g8pKscQrxDArKzUT6oJulhmx+Z76ja8w5TwksvgWqv4L4YiHxqJbXNLehQxEI
/rYotX6MhreMAF+UeJ1qGofc55COvPa++uysLiGb4vP8pOLNwLmsw0gZUXieE4JR
xs6Own6Bk2sf2dhxSMM4W+A+UjBQZ8bra8WTeJa18FhpSnyjai9CpfhndiEcHw/a
+mUXJs4Praskz0qZtJ9Gv8yflFn37d3208EXAy3y4ykMYSijR0i4MOGziYfAnhBt
STNaHzpkXIo6OgjgRO/jm7LulfGOL2vmZ3wcnyvYpNS/+eCvEMucS2Y3+prO7g5h
Dx234uGMyXdlunqZYlmscrIa25hz5c+gETo4c2QcB3WltvwLyKR0Y0k96MupL938
wLE0dkeBU2LMKrvwt9cdquMO+rtQMGRGdNueXidOUG506SJVU8HrE6d6RBQYBnh7
nsv5JngifTFKfi17+0bbPKN8UeFeX1Fm6HBuYbFNgfqDjfg+cWfSnVMwr5Y9V8oD
Nt7I/7+SOFh4sR+SZArqIXB1GgtxSr5vXlisy3lw65NoA9MtoLgdc2fJl6OXjneD
HYoPRQi4qA4eTcbltlw4der/6Eqa7Fua44H9iTTfhudEoqjDyacU9s+ZZsAtA0sv
fQxsfhhuPrq04TWijSqMVDnFZA5+sLtJ46DDRTAtjTy1ImhFsbMOD5YefOGfbX+4
mNvOgEYxeO71SwY5B+lQVhj75AQudzH/9C/eMU99Yul2H2T49IHp9f3jtILFQuFR
cjV2CHIdh1P6MjEyjb7gqzd38NS95Tpq53sqhJnYhXckU6KFQY+jYIW9UBlp/mjN
w4mcK0NEYZVEL1s3Q/3sUFqGB5bYv+E/K20MgZ4ju3DB7rMigXYpQD797nSpHe2R
8jZYlMPmdR2OiJKab90IEsYZ2FNW/8odq1Uw2BtgUmXKku4GsFj6fO6vRLgmt4tf
grkI7u3MkzdasDpWa31bnTrAqF1RRdNaEWRkjXpsTiAgfyYKOxWhqZXKRAPuY0al
gm7N9T5qxpHm1t+COcgEu+9ocYHfQatZSLqatXV2EnV0wyk7BAv6eJ2O1kPy4Ai6
H3T4gKDVuk9GVMY4YYqLlogqYUeNaiepN+H5ue+3/WOgv2FkOzqVmv6MCYJJHWlY
eC8g7kLLt1b+mtsuAeHGGW4m+4hXXlrz1i2uf/3P1JzR66dhJ9Kve3JvkTC3hhiE
3+uiLduDlELIdX/XQS+NFgv2K8/qF0yTRZhv3Mqc4/IwJ4jDEDLU1lPx9Vw3MWyA
UP2XlUgCCEYursbvb82sC1g1zPxQHrsO+I6H+tlTGz0ZYsoo13S2ZghNgwueVz3d
5Vq/SvL9//mZf+18yAndi7mWDe942cn1W1Ul0RMfPLI2pXJFB5RBDGWba2NbvgY4
MUxyJp7skGIardC/Xb8YrkCvCC5SUcx9D5AVX6SRtqUXLMKrJPntgCXko19e8B6a
nCijzHvkUufWQ7f+UXDVfIBG0Ai4z+BV6sK/SjhRfgUJtTjB20EDO4iew8trXniP
S9RTruBIDgCM47ec0JqXhFS6KolZ7qeFhcNNWKgdcIkDSGXWZPb57KjJ0oAiJifE
mq6wzD7LWHzHIFUUTxcnH0J3k/4cdpcmYosOYxVWEPmCLagDtF1US8kw88Gd4BO9
4nX3NCtqu0e4EuApRmZ+mW2ypDCJkswfT/vlXBzEg8CTYI0vFHkD2CsgZUx+U5AE
Ht5zuUbCeiovJ3QMilvGp6oU1ynD6HMfNrotikW6/yrG0PLQDkgg4KnRs9YDKPF1
zwBP5E/l90SEFdaP7Ejjzb5tc2DOdYTGNNWl9YfVY1/QgmT3Dhq/ALBlI8DXlyuO
wrG4/gXUW3yuarem9gY9JMI5A6aVJW+kA/Qa8NExZ57uFN/eLx7Y3HZocrgzQUQU
0b5ZKB7G7JTntHvCs1AMxfnqc3K3xxk5EhI+ji7bGpfDUtZPQJQymCtLVRtsQ5zC
eSdB4J03029hpfnFWNyRzenZg2MG9b+5VjtLWf1JKraW2bHIv0B3MJlS7D6BRVbs
8+oSzKMat0WImawIfhHvUYkioRdFTmEzFrI1E0VJ4xzg1/rm7KTbE4rElMOQxqSn
guLMTz8osEzwmv9C6fJvwNmVe1rbyfyrUbNIcUBz9Xs0QD9t9XiEHoioX1THgf9r
WKNszviUo9Iep+0tOYTieU/cm2ahXIDPDryeJnJXlDBbqBsLQ3o9NvBqlntumhRj
VYGZkroFo9tBPW7Xs6/oPxBhApdW8FQnBdC3Nu+ETbVLqLE4R9msGkkWcDL/R/Jj
UYd2JhHE2Nhpn1+yiN+kS5VSSVW6nqnugQ4giAX2A3P0CBULNrnshLIpypzB/Z8j
tXXkzYl+/FN5btqY2M4/aH/QFypM5/XfAYX5pvmKVN+zs0U5w8nLQqfaBwlUclMb
NvNJLPMfWkMzar6AOzRfZEtYci4o1FoKo41pDlbUuvIlrBgalT4dklbootrYD4Ew
gQwROKNY/wKD933rNTrctD0l2+EJfqyo+K9EVp8boT4eaAq4c5sypvovOiJcbptM
5KHCe2bK5b79QidkzAl+/Lvgrpj/8h56ETHJ5vgCHwyzV5HUWlSzhw87A9G8CPL1
QLwyIGSG4HsJC/RWgNHNOzG0QNIMAgXvFUNbCupyoWjvq5UzlxBfeKZyTnFndXq5
YF4hHHIxnXoQRLzmWcsjvhfMEEaDCB7swd5dqrnRYKMxGeGdIpIIQFupuDkBsMDR
uTKYNpwVfJg+bN76Yh+78WQGCc2H/fxEyH8S2uNP9HV4tmDvyePVEltDx9bmgdwT
S4+x72CXu6exs9xGdRHsHtiMPbXVhuFcfxUeLRtBCC/x/lnftKYnMYGqIkGtp73a
7aOuirh/DmZXJ+fcLPTRbXQL1eFG5Ujt1dl/jMIouXBgMo/JC2M1DRtA0/r+v/Xg
hgtrrsuHwzL0FcsXyMqQxXsysdpKwr3AyhNqmlxZYmG7sfEcCtJdkx3sOEeaMyW5
RX2jlYzwTrsBGVAbqOX9uu536dYbvvMQvNy40DOwKuOzdUF6liTAyBCBulNvgdln
Jzdx4ky5eKBs9U79T403Q85OLH/xTvnv6y6aSi44KAOzNdrhLoXeG3uCp9SUcWrY
Ml/fjddgz+wc8tUTbJKvE+3RXYD0AnrECCgcxliPSMsL/fGMGIdJxK+yOUUX2t4K
WKOCCz/6UGU4sp5pmuje2a1FFHm8XULSYaxkVxQ8sHVA7Gl7uG+tMrvh0MgstgVe
DhGj60TwdK8fvMl9ApGWEwpGHWOJg5W6gU5NfTJPEeOzlUDzhoaX+XAF6Q4n9DGk
c7EoR0y/6YrJ568TG8b88r+6HRnUNhNR051SkAiSbnhEgB8V+r7GNK1cwhnpBvSi
RJgQcklpGySPadzeMQHjezk5eiZdfdwq9B3gjwOqS3Adfqx7EzQ5Kmkd7TPRPOsn
olsN5mmwjNjqWXkN3DdZEDEVSGvE9B0UNodPib8q6aVZJDbkoe7yGETGDeTej7sC
4qF85j7GwFp2+auhTaCaY42i5FVXh5I0RctY2EVxjSkKpCUlYtc+0FYAKk9uS/cP
i7JyiK9lcUvkvMwh8KlnojCk1Y63Z+V6dekLnzig2/QpBbXvKKjzVc3UBYyi9hh+
qfwHwnWTxUzqzQAnA1Dy4G077SdktNQ3my4gpc77DHjeDy1FG+waYArgO/XUsl0L
J/WK2YQmR2w9iQEZHPcE/WYXJ0uKcwgEEjhb2A/McZss7b9aBNC2VuR2hXjBkjBZ
VPcyYXgG2rMp4SB4j9nd5S/s71wMi1VrlAphKEqJ7PRzEGlM1uYJAZssmZWHK/5n
ctLo4QZM8yAZUtTINIySaVzMN9ctDV1T29OBgHDdIbzfH9QvUyvSpNhjEL1F9ECA
pY4SIjkZcymGA+QlIuZe0VTdxMhDFc/GTRV7v0fHyddVbQ1LKoGGbl1FIU/JAyA0
cokeQqqjMCaKan6CDh+awJFfYQ+NsY7QAWxj6AwlB2c9/coSRlsea8z0OF7BmU2n
cpbGOz2obsBD7/X0XL3hcNP1o09dlf3I9tulG/FJwm+ekSNa/DRR+zeeAGWjK/IY
PM70/MecnjlG5hKyOgACv3v96yW0PN7uxxDqKB8dW2anWytXDCbeaqnyDAxD9CyA
8eU5fMhOnFNcXC8mfsyMotCBwLyo0Jp1e5xBgRpZvSywL6CbSL8l77or8qtM/M+Z
Wd7IjfWtkFRH/eLeu6sTdYRVuLH5JGGIid3nCtWJc4xJBA6P/CBf38ivAIXUh5uu
2U/SqnYRelh3IXjlAJRZn312f+f3bSHp98JVcUUOq/zxhcK5jcwNs6TLoEgNVnkP
0kifonfPriYYaGVPTXzlhNgnrw2dCrNCxwcgH/WFD4imtpPWX6ig0ogCZgCQcAqa
Uq1AwsFL9pwzabGMHIFwp8Wc4hJf9UAr4sBaHuqvh2x1G04/oY/0HP++h1d42Etw
Nsw8x+OkLzoQ7is6fquuqWWZJhgFvTl5DnG5iVKuMgI3ZS3CJ8ekmlJh/RIjVwyT
cgUlaRBoDntfwt6BXN5FCmt+BOnHdjbVUGv1TYPgSawnKmtG22PisBd+HT9tCve8
8Wh/DUI5iV3GOUrZsGvAri/iFKk+OJKSHzky6AYdY71b65DBVhRJ9NN7Kk5NSnqg
FzZGuqRP3sx26wTW4qxrn2L797bEwNMkT84gc+BD5jIUR4czFX5GHhKfo7iA+JoW
8vwWaNeiRL2cQZ0YsCpd/kAAVjgu35mCHVHr2BYGbAVvgvB8bThJgpkh31RGMRHW
/AD+AJg9B05QlPtoGonfRJ2EjV3reBh81ZWD9C0tq5hyz6GQtfCyxxjhJjlfwr/T
x+JRsq86+jUZe9qekw6gXe7WhS4tvgZvxq35IxQNgOsuXFIfFpW5rl63GtJQeObR
38p0tle+5dm9fHOJPLVjOn1rjCl4nDevaZQW7KjmpDl01Dg/LqBOJqMXVbVjpugz
QXS29yFgAQij7kdNp56hhjS3vyPX9mJw6vQ+E+yROyfbPBkWV7CQ/ygfms+ArF9Z
WR1ZH9KZboTg0f26O1cdoDuOgxdlhEfByOJF2eRbKPghHtliYO0GoAPUGVeriRSx
H2KTxupQ65blJg9WPcfhfTlAlb8YDyAVPyVZCDILJaiQn4JW7A+mqenW0BgzA7G3
YlMgHpat6sdQD/t9DGCPj7HQmrYBuAz70ymG86GD/IZfM8/HGlIIF1wa6Fpx4yGz
3u/sgLajEpfA50L6eqPOUTxTFiXAQyMLh1EI34LwF/0FbR2Nonq/Trpns1Fmlxg8
6KURp5Oksj0Fsh16AAg6RAfQQTJsJ0HoiGQc7/0ojRXrGaLjlvS6k08l0o667cOg
jmrSScJMYen3eZ4OUpBVwyT6YSlcmWaxzJEZWYvfPmh9erfDQi7mrLDx2ZzuftEU
DXZ2xRqCz/fe0WkIwXM3CvEUwlqOulwasO0P3EIXXX97C/OYmwcTgN2699VnGBSj
Bcy7pLKl85vfgytuTptzlC1RdqYQfuYPmap5DHo5z5IM627g1i4zRY2cF1ZcSGHl
8M3klXRi4BkVd3VOLRSvmLguooLEForvblWwNd7ndhP4VzqMxpW1Gmd2FRXXq/R2
b8cOx4b0NPeQ0mALzWd3H0qd6m3CL1gwUy/goUbPvC9xnP7r082/Z4eSREP0Jrff
WUJ5/YhZHt+90p/kb4Yy0QSIgxaLng3Yu7zrM6VblcvQ4vLCapDViHo6Er4W9smU
9FQM6mfzEO2ZUrFotdZ93HEWIncmmo6Ag6UKgcC4YZNekMH6xnJK+UhICOUmqUO2
6Wr1U6G+hAOtav42Ta3pbuAMREpHsa+5T39Ul+j5voM6yrXY8Vk11bsBFHLVrOaV
AZeCvt5H3UH/z/chjTteeD39GnagtT6X1YnOFEiQTRm1n71IoTq7JElzoLUeyNKV
QtHiaR6ART1POmI1W+zgGO056oVTsuoC2kuJOHMqJk4x4qS2KN4KcSlFoy79C2TW
IXUmZ8hutUWqbOerKI6nGC1wiUzyFNXPlMYsiZdCWb7Q/IqtYlWbThQ7dqgPq4qd
hYOoc+nPOIqeIub+22QcDR7xPwCRxuuF6iaw0kmNkpDsQycTP/epKWRgV32Z8e88
iM9lcG48NXiGs864JDzsEEhwXn4bFRHyNPJ6ZsE7mbdIvojbM2oSpTJOeWE55dRr
9sTMdUrPsxYyhRpG711y7CIylEHlGHJUvplK20q7o10yumjjZnewB2Q6dTEt4vNE
05b+iG5E0aGi165zgmxWRdkrAH9e3Ot21m3NW92x4JawR5ibgGIPNfpMyRFyra6u
2J5OjXdxBJYGkCCs49vXQldHi/WldhI9hWQsCHuIwOQ4HdZKvIwfxCo406VKB4qK
lzo2XglUl24CUxnsyA76yik29gIZqnMQcye5Et6AYhFMw+9XS78rMw9U2BsHw8Oz
HUYziZW7/xMIqtbadLqoOJkdiSkFIvQ+mLafWsWU10SO+wp/jJkpdk0V5rP1N9fy
IK/n7mT19939tGayGBMDvBcl2/+pOIesX33Wx7Xhfkjft6sJrdU6TFxYlAHYFHWw
Ufdz6rmEY2j2UYvQ501V0F9bpkSFNpYHMczxER8Kw4vDNSXRni/SAZ7rlES3Bv1I
0eIvzkZAjiYkrxl4yUKCtrKa1SROHHSaGgqowLDR+ff9PDTsrZMOZ8DsSiIOVLsV
xMqzN6PsIg+WeQYtKVl+y9T9JCvKoJqAvZRYbcZvpOcQkzHdlNGnPLMzLsRNBVbN
+lQxZ2yJO4rpm2P/6YSGTgUzTsdnr3MIEyg7PRkMaRkeeWtHfW/vUMFevjoLuLFV
ff5GsWMJccyPqVBzlLPviyVwTzFL3t3o7v5n+In4dLOEoOgUd+wORHBzmeo4ZGo2
sSdCQuVDGIiV1rKNLkWXa5/+b079+sftMLhHew+ZhF+K8zHSBuR8O0pxg/gFIDFm
G1grjuIktjlzH3PkC+xl5xn8radEs2HQpSzB0uB/8SCf1th71YlTxCVa/IqJFjjW
gf4hwwhkmZAQbYga0z0GBwYUTxTcpNs8xAQnIHFdrUoHgQfOT7D5KKYYZ/KDXdhQ
r81BRr34Jo7JGDaKGKAWMLRhpjSAKkvgzkc5XD+PZPyOXV108nn1u19dy0ndksqm
utfP2SGw+u8zcj9BXWvdE9LKXV3d5JvbEmILmP1SWHDoGGnBSFzRVSTyA1G9eJIm
XKAF+e0zizP+DnqEVpGIvs/1BHCbIwR+kf6pIvmkL6eswYAtz0PfysL9jyu8GRdi
LNuOFcqYkdlnpCh10MoVX7XtDympKIQVDhKSmFxj0IdVS1SfkXzXMXb9bYu23fvz
l3HGGlzilGKzyi0sGs0tns9tz8r7kKaNXNfYqJvTJEvejdTpyJTt9wfRcgY7xsg0
+HjuQBzH9SUKYtC8qppDn3qVaFCA2a3P5b6QqIr0TrzuvGptuEC6n9IYy/vgAYpK
hCuVs63pfPXqDmNingH76FxAajjXDqh7YgyMFWQkytZoL3/5HWSOFfyy9ZNqtyh/
0fysrKSr2dB0OLLx4UHrgO+Is9t2+jug68ifi0DXWXlGJiEq4U71N5Ko6LTGrP/y
PH4ZwAmT/1YkoHbm+INqKWSwclmh+KEfDLFzDkofoeLBrHSlt3sCrCu0ITKRPgyS
lsjxIQaCVfRmyZzCQL3b+wrQK461a73MKJUUqirY97utfIZHC2I3hQYRW+XDfDcy
BK8m6OOcTz2PnNZ7Y+Lbn0hUPrcKz5qXzrcbE5rlAsDU6wsrPsrG5O9ZhbLMEvjW
mxoWK6m3v43QvJ1vjW4BjRL4B2tSb8gAMe053Id8+Ftl5Y4mVgHcWInjwWtwjVrD
vLnizp5QngyXnW1A3E4vC2dVHFxh8aDn5QdXxOJ/evWYEDi5/Jj+0kPYmFffckTK
5Im3x/CB21Cio2/rgfc8O6fgqbq44JmEHLa6JCiET71LYloAbWmO6kRQKQpJNlhQ
IBgWTzLPmZY4Q69vM7mW6USwHIA59hhGo5fR13zCYeACqM/DNLhtcBxtKsfTgIQ+
SqX8BvRu0R1W5uphOqzRymi7O9EebfyO5sluhjgVOQquobq3iurMGzvkHZcfYCZK
RyAfE4U6t/07MYtIBGv+bT9PirKCLuirndp5RZWwWteU294mHL81vYqjL64PIaO9
w2fCNLgBca0B+hyw/ogkaRrzKgkop7jTprMsxM31KBurJw7V9IZmuq6rnQLHP5aG
s9AO/2cNfYaiSu/rWqPTga2LVCBuviKnUbbkiSWAgdX8xZG7OfO8WyzgD+L/MNT7
Z8cFUCJx2kpMo9JqrGssfhps0i7npQYHAXMj9CIOGC/p3nE+kCqKcjxSLrXQQuQn
jpvC+VMe5RvVwWwEh6/jp7MQ6QPYJHjkNrtoTTQ/vd9MDUHO0VAwd9rQuz+i7NpB
fxKW1Pla5/CBMaT11Y//Gc26kS1uKDmneq8ffplAOZRU5RdyWFOviHp4b+P0fHm2
UxDKAdUj3u4nnGqfDrJ+/SEsnw7o4Rk48l5I+71dn2zyjVD40fAhwp3e6A+XAhs/
lfQl65NpTQgfDhSE/T3HCATNgHVSaSIj787RZBz0/dtPwcs7qqAg+X8pDnq2MPmf
qNKmgCHivSzIs95nVDVC0V+Gk5NULkdjUz99TPOXOmxM6phOS/qLBUzadiJyQcLK
8N8bU5R1O/ZRMy2oLWbPG7ZZxJ1VPZl2upDqrR/6zxPYQYQSEJedEo85n2qGvzLx
YiO0zlJK47RpIScoCr2cvkC1n/rIkgbc8geMimMhH5sO4g/CiKekkEgZ0uaLWXCU
DoEwXhu83gubdyF9IMNu3ljZ5K+OsmehKzyo//wI+uK734ymLwOeoQPJrq+ZweO0
SDFO3UMJTgQkHytwo2B//dZ5XojNKlTOlr1L1+FK8OAyiq325ffk6YDxHOgyErXO
Mob+b2Nlsv6ly8oxzqzqvsvL4AzvlXqS33hzv+nL//DZf9xn0gaCoQ/EIzOMppS3
0M9Dur9UZMFzSoGXSkKUk8/pwY+nV4FhCYj0h2zHApetjsWGxY+VmiO+RASj2qmF
EB7ctawMq4PVQznUfyQnWXyHuihmvWwEYsY6DwhRk+fDkUpFhZ62tZE6l1uoleSl
D6tPEqlSpXLL6accgTG0C1r8A7dDOP3687WPao4jjbP5yxwr2kjKZ0cFAG+1Rjqw
fUCoBNqul7qKiBFTf88/84kyhzeQiA1pOrY6edMbLgBCJpgeD63OmO83PMeIhlcS
R1WcDX5clvk+Tow3zgG+uxSIWwRBkwjs8bxsNJp+nkuOmb8Y6EfqCmDO4MkeFbY2
LqWCU08CsuL4U5yw7Oy1wc2I6gVGHpXhccd3F0Bkht7sD3wkYAjyoNnM9KfbPz5K
R6QwQggXqhDOjoXBt8618JVlPcYDSB2mMwd66EfKU4M6S1/tiuAU7FGdXlCXRRPM
305DMM0eTaLTFS4+5s5I16kaY0r42w4R8yrA38/tcKfuzlZzB2KiwOYy7Y3lWxfX
0j8V0XavuTaOXec71SIkvmaKCFLCyjkamRYJ/HAqkosI/SfX5L1GwP44UWeA/Wrw
gnJi3HMa1WuvNnTMnlOLcAMXILzKobHOmgY1+BUeCuAwL4MqX/zhvy5vUtWsoGzQ
1EQoPqzmrN1R2VShGOfFapyv1bRgbZIR3nPLsG0odVzS3eMymY1RB2IhRo2dhaDl
XSBPwn/S25DRCJn33E9oqlJiVfOGI17GPhH8H3NuDoCdpKLKwFyMh+/eBmaiDb4m
lixKrz+i/0QizOoovIRZPNz7e+s3U08zkmK1RAFU0pwAz8/lQtpHujWieknCGhW6
sh0XIbIs8Wy7j6YPAYnuOr9C5puUP5X0TfULbvPO6sOOpgNF25fuP8EhKBGvV1uD
Om6lzdM67vDllc5i+8ihTgTK9zTbWcXxHwJHWm0NoigilKfQfjCIyBqKV02F2pou
a/dKivUUh6UgFfXQ8XyhdEvphKqEmzN6UsptAhyqQqfpF++T3YZMsObQdaSHyQdl
9aurfQL35KCMdjkN3kEFo2CwjjUtuxJuyxDznbgpa1XShIwlbEo2b1j8k4chnRfl
Kd8Gg08dRl5rLDY5Ig56fBCZuE4CkQnX80mAATmGfGtJ8/nDwRunK02cEigwOgO9
KAL74uTT/oWSd0xqdMBg4fGC9vagA5AlGWQnxhz8Se9j6TJ88Kl8L5g0WCIh/vuL
TAJEL3psOsXherzt14/BYNqllHPAxPMRsQroHTXLicCfZpv0UvSSUR7Nbsxeimoa
RAGFpHs6LcDYm1Sf6rg2oDPjQtACDalo20pcrKgruFXO5jq2ZRbZl4EzO+eyGQLF
dn1vYKHXO1NRu74wkQYRTk/1VGwGfmJeXHFuayrG5nT2B2ox1Mg2H4eiJ2upK2NZ
snKSi73bObYM8fWs3ESlDgopEm6Hfm2vQYMaQP3dWtV6YYYUcZ8Ii1oxTHigGHE7
/4oY5c9FaEvsPlwP6TeJQ5oLfuLkSCzqFkC9uq2OgS30/dG6IZON+fyy7CefofiS
PZo2IsHLx7DFjrUZrI5z3kACgOzXkfQ7WCvyYPC7KwgUsG91cvTJV2AMu7ckT3uh
tZedp080ucVF3ImoHyYGuAt+cONOCYINKcgiDhqYPMI4JSZJeNoEgNp/6apAvGEi
CcrTMOliMw1P+9+05a2/CwGodHZ68apqi5tVuSeLWqCg4+/a89TP3CzwqhsU2xLS
8SA9I5z4cl85/7HgiI1l+QOYuNVBeFEAXWErVNsECua/loLAFvXhdjmmGDDTGt73
D2Yxdo+geNYRpgnuHrL6bgiN9z24YFAXhknTNZwpjvxMIuLQZteJuhAI7k5g71Bq
xzI4ApqwZtGy73HMYU0xHyzVvaWckefOY4xU0i5Osp/XOCaoC/BGQ1wQ/5YQNF4V
uHD09SJAFmQM7HNDKfD/SZOg4XAyUzBXqGm4EfcUF9ZFgHt4i3qcekVSNgy/s2+J
FY08a07vcYGbhKsSOK8ZQ18AAsIg3IqPc9rEEPG3y+ei1bEV1qm5yilCwqVT3jKZ
RieOSrIgE/dxVFiLxZ3+yyn3JGVcJF78Lxn0YgIEQDiemTqpdZNcBNUFwgjP2U5k
1iUED6Vr0VwIZD61oTuNitOCc507/4VeE8eaEtVpQeHnpFsxKPA1L8kDF2ewTD9X
c0VrGbxQ7oKUkvJsM/NTbfho7VdZl7NbbLA67UhMGdlI5YavVFKWfr42fPOlgsz3
AU1Ot3w5cOPwhTviaqcYcocf7uDA4vWedL0N6HJZcS5vzP7vb8oIg+KFrqN77o4g
yjMYqwcxjeCXkBpzOvQxMsaJe2AYq8OoN+/isFM1g+1wkGQ0uqGWvHTVI7QPX4wv
mQxkvnij4sGeFGIXtC12rIMxLJqQRSPksWO0dUSpaYGMOomnMNPobo6+hFqkkctj
xNEAe+JAj3gzF0Tc3Y2BKZfmZxiYyPkCa23UXQ1PaL4B0RucOzbqJmub0GsJFUgy
9HZjOeM34pHCHjaPO+/y98/O/zXfM66iOxJXP8n+Vn8dbh9tzwuQjJOetieJpy6t
Ck6+qHiAEexvuaQL16IfnXRWI3XCSZjusyGyS12+Ujmu3K4VOHGtWBrvA/tD3drP
tQxh4mfrZIMyLZx2lajY78LyElZDs2DBspsDqmjEcpOiC1cFhFBkYLvK8Lgu5+BL
S+FoEFPQVdB1c7F6JqArkbmrQnywQsKr/UQDCcyA5G9BkWYdL5ckj82rxoMIT4Yo
6gOVRdl5GtyJC9Hl2b4Sw9JcfdjlHwSec6fcuK2jDClFTKuhrnyi3nibQRbwhHv2
imi+W9hw689LPEvfyQ5X37HkqeoJZONa+cm96Zc5SmaYtZOcNM/k0JrDkelfdERH
pE30oJ3iHh2KZDMeEbx9poV2JiqqB0ufA9eqyWzjKGzAmaM9kY5pvWvHlVr/FSYA
cBnQN5Seejv6BKYkRD7drzBV7Gv+Z6KdyyrY7xAu+UnS937/cS5/SqZkuFefMdu9
SOfCKA6V9H1Q4O7oVlVvU5dRNrqEI/UaeRuryh/f5WYvn2jZWgDXqeQIKJNhxYJF
qPxxIjNfRIS6zPyUwOIS/mjGNymToyVsqw578RmY40sBQwEINt37u/fzsQSErB68
QN9k5JyFo2CeJ6Ov47LxLXjPTFASZpJDvOxQLPavc0Cuim8ORSxbp2tCDUO1qb9i
RLWUuPqtE1R0SmFd+9eoOH4P845+n83byuHzIV5+PDAQAxNWhzA67UPrsiKLjTV+
OuTlgHKCDp03ImE/+Riz6RqwvIXFwO5dg+Suzo3ALfpSy0TAyKNDKNbSm26fnfUK
3ir46dOSmJzgQYM2ZzEB74ToiTrJvv+wE7ih/CtcYfYeY/+pj79HvVwCS6Sh1UTc
sqw5RV+7nkZ2NH3ckTcmJ8Lnn1+4v9cXHHZUJqx/f+hIuC34Yj7xceivBymCHgBq
06p9RHD36ZKKBRvWN9zbaHmWVYb9iAYMCn7Hyb3u5vbC5IeASXFQ5fdFJuzM97tk
Drj5j3STmqpn9r3xL7siEjmbVxlDXqsrZcCaOLbMwglYGNzDkRgcIZ3wITA+49OD
aepIex91s45+MK9A2U5GWyijzMWw0DPKJZ2GdYw//7qTtzk4Z6KXqeFdbqw/XUD3
a+h3f7oFu1PCxvxK7cIdkeQiKEWny5rH0+DBn14BZfukrKAfExFldnhe3BRtejYS
hWt8M9SkNLVJuuhWIhg1i3cChOzeu4Z0DFQRZYHbidVpgmAOWUVOlfGt3pMGs881
vthHFpsdmAVWcIUigcdo7vogG70UapcMyRu1kUyuceF+520UW2uY+ofuwA84iIvf
ehuaOalBiErleF1lVKgjENKXcQN4OYp5ACX+Bt+55XAPqrtajfqvzU6s7mLbQu8r
4ONYx9HQCOiqMSXhkLvJLofr8A2I9sv0BScf4kDL5M1yiGEA/pVnot6Qw69MWPuI
mx0yUyOb6+xQ/VpftWnlyv88FtMgb99m7rFqTvUTHmJNbe2MVNhfDjQEVmAerLxU
mOWRqx+yyTaNAJ0bI+F2cz6e1k6JTMlOY3Ji2FO4BPfs3GARlL5rTjFMZtKG/0YD
T8FbpLLxIp0kUTBcRVzbjZYeKLDUVpj1ZDYajfDIWBgyMeR9hbeJlBgESs2SIyMK
qFyBA7xeFu0aphWSUGGc/RlCwSRKgbllEb+S/0P3e4coRQAweVTNqdsdbi+WM+D1
UfORnVrbgNQPQH7PSqcx5bJU+gI7P4yMnQPvpcoie4aKiI0Ew2WVdFGmVUpXDVMF
rFrEECueE1ODvsJz8yfY4XhIrPvcZyuixcsBX1xU/eybuThUC6n3R/7lpC89F3fU
lZM/IN2yJ5omEjrmX5CQvf2GGr2PVLOobkNR+KLIUZ3HiiaE5x6jT/rtytT6TuaE
ASO9Fh3Qp9MEGzeuAPl8F7iUqwzFaXDN/5CYoO5Mv4sWUMqPpcuYBuJN1sOTrkfb
K2gQPohvhji0cKel5kdOidnDodcoC8UCeKrXPgklRFQs8oRGO1kmtSlJPRuWuJOT
opcpMJJkDShcFUsTG+kAetC8hBgtL4SPpBaUXlMrmqqKxBOECt3eBeXGE9TyavDs
s9XJ1YGi6NY7T/du2ycON1bzwx7bgvEbGVX4rzT9XYU7PA+dLq2hJiuo+BLtdpeY
ooIeMxyhMQIpZcYyLQF7dcG6a+MT195inXVC8S0zf2yRG+eFb0u4MC2jE7bkfg/n
8RYcgPnNy4Kbv7iWDN7P4HAbzhFdzq53BT2YzdLv41tvjXHoe6ILeKzZfaKt3dDo
pIGdZ6GAKsN9fH26iLFP53oQDMI/fOnmD6QAK8FosyAjpcb0htHXHOirVBmg5v0s
T3gBKS1CrK+CnRjRMDpzAdwYRjfn3J6otWaZM7OBKVL8Io3VmgMvrY76HYyhQTU/
9y1J1HxJYCuA21EDDui/mXzZ6QkRhxzuEtLCzSqGdAR6OyJWI5XJ6ks+SsR9w5tU
3X5QSqHtlHIFF+1WSgqQHOYWGHF3c7jIw8CfelizLSivr7GlfIeF6LY/USQejA+P
c82/TVMW+kJ4jh16JzXvNUX2wBrAmcSCOz1UlpJ1sIqI/x5drPGE5b+fgJ3SEIka
/CNmlWVZRHUMX8NY4KSpFJm7GDgojN1HJb3nKrkpTEYTpcF9cQsE9ze+oHmgDSoc
j0DBcCafWG53Ep9oFj2FBChz9BqwzQaTpUl6QkR/1tzj1pnD+tzc6lpdeNlVJIDh
qyNw1RVa3jEhWB4qMOds+4FbSS5GAtc8eTmDBJRLxXhpU+Uq+r3JU7wqS8GoFSCz
lMZe6h1FTJxukPtXmXya99SpZV6OQQ8r62DeO4ge/XC3Txv+90fUzsowWQDXwkqn
fi5VhqxQ46wc89YvGxqSSZ3Xbz+qQYKfG42EkGwfeUDdhKgPVZqsQoxTOndiu5Dc
9SJYzj4jmToSJRcoUO1QtEt0dsHvoqe+/gEXJtQdO65ap647lJvwVJHrZohqVX6W
WS3cdwhICOQD9mIeZvNrVc440zQIKK9l5yCTO5wQhlR/FEXXY6513yr7jz5jJ1GR
70zkGyz994A/sOh65APkRYw0N2vGegY9uBDRTFKQjxDeAz8MLiFRlTRBRbwWIdek
cwInjWyRWgwky0N8SFCxVMxHtgJEC0/Sf1ndu/+x159MehYTlCz0C3ttUgWaf/3Z
agf4/7yeJkBT8s6JPmZZ8iGL++3r+AyNFx2JYtWxqD/ktnjiVq7KgfFCptlnAcxH
fDqBkRgs+j0oUx5btsMbZ7uwSz4tbHeB+lSDRoP3CM3CKBehrSo/T/3GHyzgpuGn
9f4ktQ4Yxl4EhLFwzacSdZlwC8RDq9dMuUtlBQ4MuEnSHk4gFnUi2h0KMr603unz
6FgQj432q5VbvqLgVgAaVxeRNcvPjLPRQTAD3OXkBWQJsIHOPnkxiQGK0T2wbG6v
YAEimhcfc8UcJM5416koHdEleFnZwDIF5rZb30wXWpFdYSJiIIQTqYb98aJA8CUP
FVuJEE600EviMRePRZfAC1NMOqTv2a4UZpIpG7YMlBLheAVAlSKwzA1IO1FD3CaT
IBtciKRj1Wca3C20C3KcmAYVdeia6ETBDsWEk5zvICz0TayA6NCoYByXONykUT13
2hOTTC5crTLToNgBNeKvC5nWgXN3UT4AFza5EbovZxHL/oOEq7nThCsVvvz1yvZu
KnSwk5ufXciQgtULyhmqP6Q6KN0Ictu+fTa0PHlFOsJZ+nukG8QMnY2PzSUEJ2GT
Cuv5anT+sRTnKr6KnWfV+KjgVNYNfiMI12tCVLE2mfCPZzjHkR10+kUGg+B6zI+S
D1qzmaWmCpRhbisz6ZcSabYwD82YMcCF7S3wVwoUxXDtOCHxfQ7bklN3j4ovVW+G
exfqttHiwLM0CUKckC5LExRBjZ557x/0d5VDUNRWUIWn0epFfjLWdgh+40RbaZ+V
V/J6n+zuIskpd90s8KVBhyf4LpMu1Yf/Ez5s8M3ibhkxmNcD/HvORuIH3K4DzA2v
D1m7Uzyzk7OkGRXNkI2/h6uEmm6hPZjnWEgBQ80ud06foewmiGeIQax3a6VYzqkW
W+rOy3PWjfGcRkr8cmAFq06d0RAmxyApx6IpFlnH+CgszA4nThsd0Kutvkg/+tEX
mGCtzJxs/98aHctnlWK4MW/OzfNza8/DlRZpeVE9MV7H7B2leCAjJ9gmys7a1Ca1
l6ObyG/KEdJLYGaW7Phz/+1iD7j1T8/8a5LAZAsVjXWr8822ZSdF90N3Z/0WRYJJ
MiyfnZlhj/kG/euIZ8VZwKT6S9SUc14eekGzW1gdhEE7Svq4roqeI9PA+lbNiDnn
gYCRnsnKi7LPKgFGHoqX39xbowVdQQBqyfaepuXCiZCl4PWhggVB9aPfWJTPCKWZ
BUu8R+477FPhCnI1etEOR151maNRCZks/jdPo9dKu2cBk/c1hXyx7u4tYRRDcMbQ
4jlxYLsNP2vo9Ah6uQj8Ycdec7bxXdRaRrAbb4d4zB8Xe2WPMn4dk5r7cKY3FeMY
FECvh09IonJl9T8XOUR3oslY6n7GcV19XjIvnkF7GOl+PxuljwwkJnjsFbLkfqty
ojVq+YdSFOweJbP1JknFLtjkWLI0KmZcWjkghYObaniqdAdf6skfYI51vjZW0/fx
snAqIKPKQlFwSZ+bHRwss463csyCbyKotJ8u7E/5W24VoFkNlLWOf65HkVhdwU0V
KmTGeviAMDVjzl4otPkTwblkDouCKPVdvZ7Jmb7Ez0sP/WUpG00Q7dL6gsu3c0Mb
I91zRM6nZKZRcE3G4qKzTtCJUNHQtHS+56fDyc3dKws6YVH9euUycvx1lD4OHGlA
v96GV8zsXpQByg2OxF363erylMCiTIj3zRkUZrBc/aGpQINdflKsTNT+/NmhuK9j
t7xQWusfjWtj/cSgQnt/M/cnpwtjr7yEgEwkTdhY4G/LVo6wlyGGp/f6c+6FxRf6
Nw/rhiTNx5MW+lkOxxZZ01cPHZQaPPxU+NL1MKKuv9EOQaFol9nwGixqaBB3rBEc
nlHjDFZ7XSlcy9gYsCECN7Web0UpYfQ0eMrwBqfX6h068tmJrX/Gn6GDNsWuuohC
msCxNeKLD49kMMWup95sbigefacHeYEIOvELj3MAApxtoerZTlocaBmvbAGv690g
SAg0G/W7LxPWx5pfZAQhxNi4LzFbVFyS3xQK8sFxY9Sfvfp86TtXq0MSN6NBOZ7X
C/xC8gDveqLD1pPclXW0xXq6YZgnEhf9gyYu6Q2pKXaBIouoM1X2JHvkRSV4m4mK
rIaTb1h4c+sTYjkTpCYAxTKc3PJsIIJq8KG5B/eMMSoIDTp/eLsIajDOXa9QZ8CG
UYtFbnr+SMe9ROKHoDL5wVipKUyOknxk/Fx1ON9KR3vZqeiJm+AwN+O+wM5wITZ/
GJCuJkS/m2hrgKcTVAh0TXNvMahMdL9otB1yUIA3osk+ZEm+QPXB5+kMMHmj2t0H
V82QQvoxOxXlLmjhQluH0OEPgtUsoKcRWHxk+bgqrQ0YQ4MkTF9QkyyFwyqiJ2bv
5rvZT5eT7Tf7m2gu9278AFch9LubVS5jtsc3P1BFzlqrO9JiGQlvQQpSuerFSDE1
EpeuZADsdMe6GXTr8YAu3GYRTBc/6yjwIy3WNjQ07nLwHsQzlaVi40SSC03wEuTq
r1RpMhp7R9DSvgsE4WspRiDmrfwN3r8okuUCKReELKGtZnTSpggECJ96VGtZL9lP
7NiWcrdOdYsRCiksrthiC/ZEAVb8GbhnSHqhhp18PztcJ9rre6EhPxZX8AvFp1Gl
7g+dv6u0KoOBQevxIbpO8cOiJTCPQHDLoJ1ma4oyyYxIuIfasVjrqFDsvwcPGZWX
VLqXc7cXaOHcjb4G3ltkAekTGItH2ZQ8SyrY0v0xW3za67qg849KpJKzrMPUE9na
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
JpbzCuslQYGpFWj9Mq4Rvo5mQHmgBAJiIDbPYSyeAgmvUNDgWMtKyaS5gYnz6AdY
7gfVtpySt1NENQJg8Nue4HouycKQx8RI8Jk8WY16x6ii6vVEGRQDookzIzrf0vKa
mbJnHf/9uaOBTzTCv31YvlTTbfiflRUbmL2PCVKQUc43Ie4oROvwLwMLzLh1LYPr
+9yXY38lRhfstVjOyWATeTqkOmBBhnfpJa3U5/NQqs9o7D2QmSvfbdOxX5ZnQ6AC
dUe5CVx2l6dXw7NC+CTAJES4z1tZCeEaIolFrU+p9W+RFYZ2Lo3YqS1BJHlXdILO
UTrh3hpZb2rYSF5tk8wcrg==
//pragma protect end_key_block
//pragma protect digest_block
P/PJQA3gnuoqlSZ46ccpPbD4Z30=
//pragma protect end_digest_block
//pragma protect data_block
9LJvuDgqhICYlcIZPTGVMsxzY7PkS1gMdMu4UcftNJZcgD8idwmrJ9GOAnzn/c2r
kwy2mV2o4FLZNlXQUgZS+mhUJwaqkwqL0OcNUjMwPbAmpbxzBcm0eu5V7bl6lSZs
zaYPOUQ7mmkpA8XpA/GsFOsDTwDGBvXdpoB8wEIIliiVnNgRTVhqfpa/z+ALAMyN
meKIThKiCnFt9Xt617C588fo3UFybM/Pp8V/Sx5CUqVB7+CDogaeHdAutp19+GhS
IXD5l6tg4TyewDPTzR3YstOPXNTgGMMZ/aVQuZlhrLoOVz0hrPZWzg2ghHTVPcg+
VimuXJyrAD0egWkaopy5zk0Lw3+EbMgCaaTkQLyssd4eV0pWCrx3MxKTxkdSWG+2
VEHnSY3fdupDsJ1gbRxgnSJ87XL5h8Cw0kec28CrxmZY2TEq/UnGU0SV43nsKSZQ
1Nz5klo8hRkh32ssZS9f3wtcDdFIfe1mvEkbBcufrjiDfzIv3oEcUBorHe9WHRbi
uIGDtONTMl/PqY0jlXRsv45HKze11tuf1lCZtvRVtV/qZP5QKaphsHmA5vwTWuak
favMeDRlEdmOLPwkepvgaGmoJRnodRW5ImFIQsWOyCuFbPyx4XyZpiFaNUr2BTCD
35dgs8pl2onKSJiqFSItb59u5uKj/sna3xq2s6+FYWOG9fs0SBMfQvSdfSKVnSOh
gaS+sC7bK6cbOEAdeKGost50VU8Loz129vZ9BnVkAL7fmErCcHf1q00lm3hm0TBm
s0t8bH9uFWAoYQt+HHrkicC4RUSlBiUq5mhnxWIxRuykGUUgdrJuSz3SM3npQcPu
njFGgRJOk17ocytJ+SPVRwwOsFtQhU+PODwzuZ2gzXVSssgwABSZ13qsCCDWOEQs
RbbcuGdydoxy8VHRpci0g+AV6SVACTIKTKsOsVVnyS0aAKpua/DBhEwW6yZOFrtF
8TPH1Z3FcpvYcPerhwpzAlT6enofpoUjyjhi0XLQcsBMYD/fvWeK2wNJeWWMA9uJ
FYhJnNWC87nJlCwWFysLnCDJCUYZe8gH9HcLAKALYkLxjIqwu6012ELb4uqyQ8SY
HUNJDufixThNLpyI1EDuxeKIAsr1L0hHYhnGxmOl8IT47iFdzeZjreI6FTsT6Rk5
2EkQzvVqR9ujO50IegNg2iQk2Z07NFisj/siOiZWVZKYUwyNNa+LuDwAoCl+nVfh
sQF3BdEIZEEhA9IywSrIUwCAF7TXNlSn2V248G2tDLHBBnV554X39vxq9GqGtJcH
e7CVfkU4qDgwzG7hMAz5gs/7UE/L7feSyOkn5JB387VkkeVqCcN43sIzzRH3YBqJ
vNzy2Y5I2XtRxYlE64HrLLuguWzP73+by9QkonUvyk1rSSqVa9dHXb+BacruJ7l3
y5xxFGr4ysxZDScyy6viK2Wc88auI9yLoAlhv7owu0QWeEIN9Bd9iiN+N7ivVOj2
03nsCp7+jrZHIycEcC1PGFxlmvHLydoFzjlD7Ww3Tvu7hKMzW64Jp8AVeZY1WNeN
RKeDhxJqpVSfONenPre0QtUeB4+JJsfTvA4qUk+t/O+K9E8ZwVqaE1Z6RT8813VU
RWOyFFPKWpkT7sBLulJO0EMVbtyyISE4kgVmJT8YBwaikT8nS4mAlpVfravMEbCi
V+q7cEMRIHkuXjbJXECJtbfNO7II5EEEQfYzY8ryQdou+YsgZhZlxSp7MO3dWVms
0oxPngPLttFkVo4AgJjKo8mEOw7BpuQxD/Ic1lX9E3pTuWd93eS3PuBYCSdGnl5U
eeVlreVAcRVbLg/hETkkf9nFa7HvkhVmJEzpdnQrzMk7BZvRKDPSLyj9Z3bHXeai
h6+RXghyUwO3aZQ6tmLB8mVKrAJZta0o3EhBSmiSIxw0UzFcyPej/1dTzF/EIRn5
xg2MoBOwwEtyKGibosRObDIHkdmrZTtC6txYEnLVFmwZM3d1+zQRlowiMTvDwmQJ
U4f61tcEtB36d4optQfBbG2G+c27fZMy98EsAn+ir+a1mzrw/P3zVEjZmQnutK94
g9l7lieuACfSeL7b9Akkai3BLZnSVQyzaxBPqnR9+uYbmJu2k+N/qzGqR1AGv+R1
5bZXnv1JrI+CaS5Zs6RPFjY+/dMtpNaR9IiZlEfIGwF5OguoUNpzGG/8S7anfSFF
XJfjfU4rcpFevAMXalt6c2CEklDl/ok2xGMNsUhuiuBVI1IEbr2vDVq/yVA/GS0d
j4hAVmct+julSSdovibPPPSqIhSpQY9/tOzzBW18g222SFdEzQCgZhnoUaJGE4f6
VG4IK/YNEV8quOPvjYKsQ1JdXX4XCrF5sH+mB5e1tG33M/M2QkCtYepWOcq9NtXF
6SGzSbRIMmF48mJDJa3h82CMnl1DsH6AU2ZcBLNMQnagx77rgGnRr2hJmm59TxCQ
9V5wbLiiRNB8Z4V8Ugb5J7YZSVXCcTvgE018N1qyEuszaiMwJ0IaBVO1UG8NUcDC
aSkgNiHQzxZVlkQYgM3ARSfoPvn0mLXbBvK0VT75mdkyvUv7NnEqyD4RCRiooPoT
Yhod6+FqyxfAYmrGggdjvJSinAOA+6ovyaDfFMlPgP1KIWF8N3G5Ok4j6BawPzFj
GWFR55z7DpJXMXdjb2GqCwnzK88d4jcNkDIctpyecV/XkholYCUNbkn8FzsOkeYD
PWG6PnveTYVpFekG9V9bUR98ok1r1RZymU2XcU8ewB9KGs0DFBN3ZAnmJqxuMRCn
zEp9n4DLZ51XdRqdOFvx60iCZorq6hmyJOQzbQLx95ii4uL0d3kdKxfufM3K9/Rk
1bsk8OCK7yFHy2dDYAZHrzPh0E/K3niSdhdx09KG6d/WNu2Zx9Y24EWU0lyA4LnN
L2ziDLT5jlY98GB562+OFTCSWcqc5zgEfrc6+E3Yk27QV1in0n92MGSZp3EVJwo2
AqvixkOCb9fa1tQIbPWPdeGaJ9g9wNXqVvqdk15/HjkfLqq01EMXxoZpE4rIP7/8
WlPk/AaUW++esxVvTD5WtaW9YfDzbK+bP0qLa900JYnnWohEn1iKIIRUK9BZ4TWH
SjfJ/pa5aVOrpKb4kANYGl6MIT5CpBmCAIkYjqujvnpRp1Mveu70t++E3VkNn+vU
pm7ACt2Kdo2N+/F+KU7SVFjruD01Di+q9hLBHG8vtSXwkyV1dnSEcnblJxhdqo7s
KPkK1AgwP0a4Du1GxgKuLz/PB8U4uqvSVBTUIQ+pDa0qnFrYbqWf0EwTNkrwPkVF
phvzcwOPKcMKD8w7gAJY/Gni085m/J2TuvkR9Pn3CYX9iq7na0U/SaD5Qt4KDM3Z
m5Uk55Qq+b9LTvuUxMok+K42+1wpNIycqgaZCTpi+JTZVLZZUbYD1eQVw1sxsTkg
drA8ytQpp0vK9I16r2t37ccZ7Xi9CzF4w7A9l3/QmTKjTFm2QE5hPJqeYVNt/YQj
xSzfUPL0fPv01JH3vpsCnYMcI+KRnWRtv8nDZzTjCf61g74Rj/4hdg/PCZkldqRM
HwdeZJBa5N+VlfDFu8bCleYGG4T5AWhAoHfG5aX6JksspQScGfYIxaPfYytcCypz
pyWoPHuUUiNisOk+APpDIRhYPMridgVkyv2J1Z3Wd3m75Y2cbC2xXz1GGRSE+H6H
SviJ2OlSbc+2o01/Uua6XZzDatSvHD7GRBPjDluy1EMiu7SsIfC0y1fqER89qZWs
vlR6sTW4Q8fkYHQyKuexb39/Vndv6wPJLROI4fDBaYkZA8wknZJqS6Q+okKFijsW
UUkbmuYWSxOUs5nTvrjjHHTKDczYodES7uJYcB3m9Uhb25PT3M12svgL97+FoQ49
9lKu4EjjkNRMBtrnZRi1REue9WjxVcpa+e0ChhvVxxVWCZSUi4iLeBacwbve+U/7
LZKixrI54z0TM23ft3VwK67FB3AUS8rcD04Swi6q4xrY3V7Xo1QwhR4IAclVCBvw
ffCVXg8neF9P6jgmCzipswGGajYGi1+6kT1yS5haaxLZ3N+lfgNbZirYMs0Zwu/R
y4mQL2cW5aSEXg1R+CiS8NGBe9iKiTgnWB2zx7eqY/iYQqx1hKVsm+LFwYjNUPUd
04zrmPGOCBSEpmmJ+8/h1kXSbDIEC45mXScrKwTEfKm/ZlXKXbQuT3R7U8FG7jsw
LQwyJ/i7ZclgakH71KdWZHZx8ZgslsP7Gqz9IIcTP5pk37h8WjkDo0I7lCOVPx19
33SPdE+std/Tgmo3yrwtW4wj7zJ2Lux0JJhhEJWFX4yd37mgpPqNu4Bp3wA2PrRA
DFh7RZiCz8eU9eKeK1Vg0nppchR5OfbBN+B45r6SCjwJDwpC+8J9Du4NwqGpe/KT
7iu7gWXzzJomlM5XkIBgZDozYFa6mC+UOx2/9L7oJ8cJkeFLRqiiHARCKqRyWwQ0
ndHN2XeFB4fsm7mpIxFFnjhStAaxDsaaArlXc7MLDX42DezV6k6+Fr8NDkj6QSlu
DEvRy695eua01ip1453Lth5dIiENeiDMAqF8Ucfw4GpmrUXrmtbF8vslCZBxST9h
bnHrfbarf210vGSnXpm90qd7xksnYQ62WL2G3qFbmgt1WL/8hML2WJZkJJVNQSIa
anSZEChPI5M8uU2gIvxtCvOnZOlzixWECMJu/uuvoe3xFMuNLZrBDKLdNfM8XWWE
dJS0AUDWrLHQT8w4r6aBRNpEydf64TNYIXwu6oTkwxhtEr+4pXZl83I7yl5vx445
oRe9UEMtMm+mAerpaQm4P3NesdtLLpNpvjRzY/y18otKLr6j8QdgkZML9+mikEzW
VVW8xZljpCPYAUCBwcm/XHnzGa1r6ewz7NUKqAe4ivYdNIVGfQZII0+IQTOfbIh1
M8K/f9143KGUaYGe2CPwF/sFhE9UyGvKMbpTEhvl9s+61Spow6FTqEeEp7IZla8c
Zb8hdXFIGIukFxjlhMI+rbFGR4/Gzz5Dnxq9p20+YA1a7eX2Ps/Rzkm+s1EINTzt
1dkJjP82G3cHiWP6nrsgcmH5qGpFQG8DJ0iQrsw4qZNM0UpKoVyvCNyNz/okW1tE
NsUqGeDngCbRJ19Bvr0XFB/tk07XBm0g1Nebw13nee6koMqlrJPk58aOlzZVKCmT
FLIiucl7RQ1S4GYylil3zI4CnahgB+6PrPcIfwz4aAVLRkxkItddbzwdoJ7HnaqU
gghvolkeN0NGlDyCR1mCejxExdvXl0JlVLqLf7B/n3LBSrbGtPYhtZOYQuRyEoxY
w5RR3XMBBLdatcS95xZbztRncXCle+kbZKK5A8fprD7SyhjKu+sgoVCvpiS1YuhS
wdnOJYSHjYmkOrv62S2Eg+RitetQnfGDAbzRTlc005t0ujjqeHHe+YoIWmSemm7m
ppOBq/SVdtqUgRn4iH0VpsQkqgrjN37ot3KlXsZfpWjyqTDoOg4Xx5r+nCR+3Cza
jPv1bS8kAxwpbt1xrkWt3LYQy4DcW2zHr1jkEAbhfB/fjEtNBIg2AxbkTCyXBGiV
8BW6HUm7Mzx4PuLYwr+4GydFJGOThqc4z0EeoeUU9z8ca8Td27U6PmJdPJzId2nc
sBigPh2Y1eHF8A9HiJVe7MxCGkJs5zWtgVUa91OAnj4NHouVaJnYv03tzWZgPCzu
9UbZUUo9I3tCCf3jnT2cthNbN89soQHolhMw3WG9PHAOAbDvFTLr491si43ssSNe
KIE41AXyorfyGVacg4HsgBHoOBM7wVxPx2/vliAiKPQVeZFgpiuSBXpO7VBLp2sw
kkF6tweAl4+YglM6/GzXMT8R2ZPFRKhJpdPOURuCDINi3kW3K+uhmcm2JOhVa4Tc
mzBR8FgotDwkLroEjJRVnuIbAQcdZEb+BpBLiBBnwzEv3Tg0bfSfefixWxljsMlZ
lD7U38wdgbKMP/cl2nyc+IBHBjqqeCFaYlZLb2TMzGccKS7K+q/qv4RHtj5Jbhnr
Azn3jTlBgEABQnsdnEU5/wDrwbqSfO/apXEyrzYmb9r0GjJcv2jReONmOxg+q7OB
6DLDpo1MuSAU8kMhCDgzbf9ngL0Wg9iTa0qDVtM6ggpvCmROjeaBdwchuWF6yoFh
zOXJYrPysYFgaelgSsjhOdEI6bARpHAc5K1fZ83CgRiJgNDzw/m2QdewUi2kr3LV
LnfReBV2Ios1t8c460wgFWYXcfa5p+uDXGDtHn/MObiX2o9t1o8arNsBBGGV8E03
G1w+QaDqQn0AFDxDvqpryZqUcmmKScY7I4/M6+p66ZSiKTGF9aM7lPKLZzsXS2hT
kg16Zyo6Jdw0Lh4Ae6t9Ly2ui06ZEt+YzCIvW2nZQ8PtCAORsC9bcdJ2LUscD/8K
q1NZILY9rnZFVjOtgAuVpvZajMr8o5NfibVAN7RZm8yysASOcXa4qfFSowWSWDXo
X0C29x4fYqEDCTq8JIxUA40AAvLZB9fwNZFK5zl8E4jM6IBN0Dvev4Qy1JgI9IMT
Vm5rt5oSiZXbiqP/xNsuBqTaT43uM6oh8Npqcop+RSzmZAu6FPmAdZ6pcKCujqL5
X9Uh+fQw0hBiY8L7AZ85JEXImMoRnSm8LRbzIsNZ4NnSvGHqqoWiEMuKhinUWgTO
yRo9HvTn+O6iIY1Zn5B8WzP3Q1alrNrf9lFbISaCzj1UG2RN7epDan5f5u1x6GRG
I9M9Z0xNLhJB40DoVqIBjGi1SBkZvq7C0TN4JqiQd0vEuizUYtkTae9p+FS3rfKb
0baK23m+IyztuzXLZKn10hLPH1o+xVyrFKPF9FmEQTpE6jMhdoePS/r75TvCyJRC
T4OT07iJJUSlLvuFEmsWxQI5SiFTMLCwEpiVX0brwrINF7PMTl06Z9g/S3u+oXty
HdgrabF5u8ArcmSW4FZf/hLCPYc8gPRmvnRsueVdrxAczNmRKXz65cQMbUcKHel+
Yv/IVVeLK/LVfYKF6+TgQPKcwtwjlzuKZlTIoOdZf5SmEmZSvpZfu0uO0cI4Tp6L
pClffetwxoDMhAsUenwTDu0ZfNcKcgDzibyXnoMpAn/zAUTI3pm/z0Lv5TbIb135
HXSwpg8KOm5fR7V+DlyXhE1DVaNsWag7RaPXDf6Exsv8eUw+tW1RcwqNNS/vfKYu
um1+T7rzs3xCunnzjPmZxKB0PhCzp4tvrEyvtLaRHYS6cNtgCCNE9jMstukYn+uu
C2xSFX0DfP8RsrQtGNKMgleVDMfNtHTVY6biTTLe6n6ZEMrh3eh3wJvfVHXoorVd
/SRd2knF1XfuHECehyhd3dOcUvJlBR6m3DROqCa4RV3/F7NkMtU0WPJzsk8Ytq5q
5VR0dlPpao0M4aH/zj6HB4C7ionZZOKM3ReXBGM3Nzrjgni8H/vfTt4xZO7u8zXD
KYz7FlWcSNcNpwFsiEVKceSDo6UCcovT4nJhl0zzgHU3ifW65lcXbyQWIOkNYti9
tuz3npaP+gi/6vJCadd/mucuHXqWc3jaaIDyMM1zmfP1eViL35U79lRLX3CjmeP8
V4DX/PIo2j0kjtuMEfPzdwhHi+AbAzU+z8n1UUamDr5ejgegjRJjZcVfWaxTlp54
b7lIazKrcVq1RKbAKdZIsypR0c94q3D9Tte8UlXBs3q1Ape7Uu4DTSNwNE6ka6RB
7L5xBxl8MpxUyqgqqBGn5HNzM3MFp/uePddYkPJnP9cq2mh534gT8UwaEDIRRUH0
zOZw4To2cK+VZ+zz/NqO1NEJT2fz062IQwJBDBCO/eVWvZoKsqXpuKOy+/YRZAU6
xtE1NV4bQYUEBgWJkmyebqckN5WC3jVc33RCXnwuqwKyhGUgSlN5veJAsmdRzCTl
XyhmXFWDmkvzh3Lh1UJ4e/y0114bEwdsycTxTPYv+q7XuW2acqKA4sLc6/ME7V02
8Zyk6h7cBTZIk6ceU32yxBouxe4FdC65+TN2jzCm/Cj5HNoIVT1eEqzqSKNJnvn3
0WSftWoAZB53O4k6f0B1MZ/sSSVbo/n7bjmpjb7s18/CrjuH7ydDqDjQFL4o+9+1
Wa0E2+n8qZNT/lzhuLdMqM65tBKis/6eILgSld5iAmCN3a90wMg1DY+pOCaoD8VJ
vzRcJFf5ngrulxpS47ayfMO8iJv3AqYvF8GlXUcS7RaD3ve9c1yhFptGVrfZBCOS
kuMkahIJgHzHhVJpYnRVMgYuSLsdO3SQY4bvOdAGietnlw82qTy3jvGqTgVFrr0b
mFlnWBt+KJx0HF0OM3eJm1XBBY3b2/c0pow0UX/SW+JGnKiLoDSbQ6m84P9yhViX
M6uMYnHJUCf7F5C3Anl6JYHnztTA8J6swfPTkmSd4VB4GbSzm5k4ukOT0P6uh5sd
49ghxm5HD5sZjI98eugDXp+220S8cd1A++LF2H4pBzBovXV3Ea1HVWj2PfTSPioC
LaryIhrj6EpptDuQlvq8W1E+zd9cVbReqOw0IcqQXzpAvt+qNSPzW56pzlQHNcD6
5lM93ReCcrpun0noGs4KUndwHLQYcXPRDSvvVVj2aU9fRPjiDSrxXWV626DSfn/A
PtoQxtwklVVdLGTMSzjEBs4h4BAOAa5kVtkWwCGnPi7bTcGjGKNqACE6fb1lWqKZ
qKoJe/T1+NbTzEnL7g0LS9jh9Xdxj62jWCEns9jkK9VKnC/wzPcXNRx8avPhycmQ
coCVuFsc83bdF4N9qebcicjslb1h8UDgHRtaTiCzAvMexLK3n8pHY1QKc+PGoERD
GEyQo+fDbWtzVY8uwQHFdQD/oyfThU00USQ2d//Hog8SGnBdI0979Tpnp4l0+K7H
9W0lZmld8E5T7Viw6TA3vHaf9bAsOASZ9EwtNZffQG78mZs6Fuxmz+4qBGMUMFo8
xag9tx4lyPkEfni32ozacBLt4SrXlGRC+r/ZDIoIlyC9gPqispF4iPadfOBFW1/K
kohEzsNZCbf+Ssaee/3gr9pwwyHoH0zBMotXsk606QU8Sn+VyU2z7O0I6ISLGDOY
XJMI82rzZnoljuvynEH87kyhlveobCQA0gT6Ygwob71HiWtrNrxeaw/QCJ0sva//
XXUSk1yXOhNVbCE0UKMwtFGHI0iVX6PI/2iAw2D8Y9MtpUTONivxz8glHr/sDeox
7LWeFuF8xkNdsTh+mBiBIJxMi6HDWlIkI+hsKQA2FipJZdYy6KdR2cmCgJyD0uXL
+ljHPukVbtZYpDHM/6YZdUhWAky/nP1WHvIyAp3yWBEkQAn5Mc9uLGLPyko+gTXq
pQxX8SZPtJkvYFBC8utmfjEMHcJKZZCs0MEFigg5NF8aycj7AjShV1M+xNsuOoyF
noTR6o9dFRXQI0ivNWyKB00BvcX//jKsWxycwV2p5PkuuEAbMFhEO1Bvu7/uJDqH
DuHeVnJZxOGipN3n7KlC5+rVCkmDAPcsh4I5BzqL0EO3sQohTSKy5OjJN7OL9qDv
EWjpu60qFLns8ooc8L8io4HYkPMf4V0iPFhxM8MJeEWeG7LuX7e6gO9ctHhbhfl/
15OipkM4ET5bIM9ntWKW/0+7mZQBMqz+4qnY6tcE0y2oI8/duNInvWrFVV9S4AU2
i7cmOgdGklvTguhbUFSa6T36gQqWSkgsdGNttMUTuRSVBiWejFWjM5hXRyljEEps
OUkoITAIEaPYH13Hs7xjjSIeCicy80e5MWG52xq+FHY96k5uwSHl2XwcmJMjh5zS
xM4QmpHnc+Pq373SYxnGFcF4zV9Za/DCXS3Q30SrRogcsikbunk3Lc7nqIAM7aE2
j1vsdQkrKLRof9Ui4PF7mPYY6D9dSMrUGOQBcfc+A8MgnzJg4t2vSD/898WF2zCF
h0c1lX3lz3F52T13XHKem7t8i5ZhfIwCRNOirMEX2mGUljBxTF2WvXEG0mwsXKON
AyozISpE/0g6OrXvQLhbG2cbdne2pVMyRs6bwwXdX0ziBC/P0+TOsuiF/T1imQh6
goAefLLC/QwiJjvTh/M6sJKC51b0y/w4j7L1uItiFT2QBs1OOIyieI6Eeht05O/v
0jRwZhokVMoxCfTVoc/jOmJ81S1Pghi8agyBEXQ4HodGlTDUH1+yOog8eHDee5XB
k/9a/cczZCY/6jhtQueaqetn57Y6etxv/vDctQt6SlJNqQs7ae+ZY1kmMEoOm2GV
nXhDA1zjKALvEqCDvNkfFS8kfuvyYMb/4hcGU+mBPvFt194y8XWY1xwkE7/aSj5a
vugxGRjzGHzvyEi+ocHGXX5X9YHgz6Wm0BQV/layln+MQld6sgvXl0BbxN0b5z4o
gnmTVsRTry61t9CmvPXExzMJcHj6dzlu+MLXuXBwKv/rwem3MQMZ6ukOAu9y8YsX
Bab4saU4upq58aot+Xo7XvKPqDeFrcUlGmUgiAuA18365B7zqaq7TDmJaACM7hyo
/IOGlSoU0g1LAJNtMmCiglWcGIza7VhMNqC9iQ/mfKY7auurYHBm1fji2/Tp3QJ4
uz1fOByYlapNuHPGnNWnVxy6pq8kQlJQ/YjkomalsVlMGJo7UiJ/xFvemHbBGrMX
DcM8SVaq9WtuLamxJ3Ko9fVScn3tWf+aCEiMrEsfkbRATJbEj6GOXmETF5qa8Wx/
D+25K5J/MaIzjarEmrr+Oj5tq0rApLp8kKefIS7zGxkT2/+IvSI8BaKdB52aw0Nb
sHmXupMBnUQcWpyTsOMT9F6Vvxal+ufu0o3rD3XQo7XMWKKEkz76cGcmPqQjsGlM
qkNYz+4ioxV/O5SMWMQjoqZMayl4opbr+DG85OfvKCbbVmnRbpThIh6VxGTdpwX0
Dd1LTeXlWa9EByAkc1pKtuBPEM9wkQsFRzd8o5Z1caia56i03uDAaI31CvADh6mJ
MZL8vYo6dVdeWFbDeqHtbK5oqZn5K52rQpCxyweWZ0XLlYEmYs3kWtOg4ybXH+lU
9axZ1gUpO1xXUtRX6PUpC+F32VPymO/h907aC6O9Yrx2MP8zgBv1u6PZS46kXK6J
KHKFsVL9yF6L6VFCckxqOTh1U+0wfLOTrQ2sJu5vS6/yQgfOd53J5AOngllBb7TJ
yqC3weXq88kuBAyA8QyxDNhBrGwIj3RXQXPOB6Smv6joa5QENKXKbuVZZFccqlkD
mn95oTAO3E8WUYNsMMUvDcnENDx9K3qp6JPQ79WiEndxZDDNnvi3LMPyaMfHlNIv
0URpVDXSOKBj1zDr1YoPIMmVZCDk7P4wMpPIFBaO4gFJrIN6Ah1jJO2JG5L8L71s
A5AjMpKHPuqGe4XCtQjv/FNATwApGG2TAGrPCE7uMTduM7lk6zWDIeJ+qpTbG0KB
vUZIhWxHoBqbEh9XWZUp1Nbg28cQreB7F04tblvY4xZW9R4yJYEql5LQDUNr0zWL
VYbPOTCOTCgeBrEMrIXAWoKtANemhMebs0RCLUu7vUC6YKMAC6RG2g3/tqtC6/Hk
NFqhePkR/DGjR5ZJSZZjeU9E7zWDNtbh0/j/G5DRLutgbaiPV4tXgi6AQa5OHoBA
dB094xCa/X+Ug+e1je9xlgrxMlLPsaKK3Tq2QiiC4cH81D4z/f0Ojqn3vC6ldpAS
I8uNTnqVqxuS7srst0UWbHukisSYYo9czkBNEc42vZbtfM3q0EbjKj6+rgWC9kb7
MTA1+JqyjQmBlKNtgLJIU0YdsU+0oM1jRNOHwbyaimKIBwc8Q5sHFW/gc0jEQtnN
GdSyS/mldDqmwRI7Xo4FkZqWD4ZwSlWclhOdWHjbBsRfUtJCeH0anlx68e+jxEXG
Hj2PeXO3RQIuf4Zlyia462ZAL1CTXt31+QS6l0I5V5U=
//pragma protect end_data_block
//pragma protect digest_block
+X51VWUOhPtxJMiT2B4S5dUwOM4=
//pragma protect end_digest_block
//pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
omQlqemSVLtADv7Xm1KBJafe+WVmaj0qlzFwTd07vVvfQeCiDr2CZ1DqxzTrJAZ/
hh+nRcn8YaFsiLhoQi0B4qeOlrbRYPqGlPY4/9nthIpRI/wGAWtE7yealAFWA/RX
E28pOc9gYpff39olQbaz9Gas/MYfLidIirWvP8/GIxs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3712)
EMeLrya8tRP0hwFeG+bgJLhGoBqyP2EzqbPQQTE49rUZoqBQVHDB4MawHNSGPuG/
dVkzqEXKdI9IN7D7wC9T+kFlhjVJw1r6zpO+yMhlSWlHNtavGIWO2dLEnTGXwVt6
lcpYR/k4xpZXERjEfxNGSKe4G25D41Mf9wf1a5dAoWMs23g2pchyaCSbsy3LHZKz
vax0BxNQclI0qQZycymfEMdHQMVqrb/PZVnfSrr4GmsGMeATIBsQR1WwMjYDBkPu
9pNBOy+FT3xanytrUfEqbqUubHol0TIEFUpgUEef++XDSPus5BBUP3FMm3U/TykT
Ou1UOTkX8YDjH/taFjzvhhn9GfRTZGb7dxOkRcdKHJ+Y/OmB2w0ul0vbyUgv/GKn
RjiM/ukwc4mtuzy8bA24Ug5cPeFY4tb3UV/TWANX0hETDmNwqyP5rdd3YXEtCi8B
Hl967wSHokwfcj8xLb6rq6lDSNrJ/QpMGbAJ872WacHcNX8Cyh/wnzFHFH0Uux6c
ZIpvHW7UOuXOQiv+S5KVOsDIfb2XvBIT7uQhhijcXqJaQ82r63X7vgM+SY8fshTM
BBclTL9KZRwWiHvmVs3o7HzqBEauka3oFkP/KwQSRqcLyOqYe4jXiTYPqFzga9Nm
5UdUdCLfiXBuZvvBC0BUdZO3TvitaLxv/xbbxGKSiCVQWyI59jAfmMChdWGQwB52
9CDU2RaBz1gtrew5JjSi/KH1tSGDh5+wMUjKWITFnxfG/gbPIn8GFt6JfQ4CJz6w
WlXdw7aZ+SrcZd7EN0q6ubzcJ4HKRvXvYVI/IRLjSqZqC3fNAUY2B+SwrfpUTB0D
DWEppyVbWrpl0qr+AG3twEuTHtmestVjiT5GBvG6NAB50RZm4NT0lKs/eCaIqB6t
dHn0kUSN3SHtKnw6Mc6KXuPxhZjgLdwEy0cpTRYFMTKnDw175nSrBOTvcBewxcC3
AezWWKmBQ3KJqAcXwdVOmVK459ZaamheD4208mmSow1eobH13EXoZuRsZxf9Qp5u
KWnhRmoJc4OF6zZyacK824/uHXGAUb5EY7r3TAoiZKtFVAGECGO9P0duAjBpfCNd
fWUDY0V24DnKl1w4BTswnVM+n2jKCPfiPlLot8rBRkoa++WdtsKRzJmi78Q2Ubi6
i/CFx0y+FcHtoPBcohBb8aa0MXj7ueqnafNRv8Cr8l5BCrmpuP8Xea77A+TqEGgW
Mn6Q8eMgoAbdGSKINQPV7OqbKm8pZjsFGmirLX9dhP0D8RUQI6rTVrU2l6gqV/lT
DmqFskvqINDptHEnzvgW6azH9vkZFYc7snfGPP9vuZ+PK1t11KrzqaOdqZadtcPr
2RFb2o/RsNQ6Is5X3XpyYAvRjCvAFeojr0xeDuLTp4qYGuR1xK3leH+MQQ5rH5Mk
ccd1xrj64dbw6KDGf6R2xWAmoaJg9xEmg/JoTpl9wvm5qIXB1YYuZ0klyGW1zIns
Cj10TkDssLAblu402Yf6qF9H7oXslm46SS5wK4KYcrJyXAik/S7tmzXomrsmrna7
HFWDK9idkIoW9WEWXpMnHJ1knjU8p2j+MO5BUJaCqS5xbSv3o6WxrnMweA0dxvSq
zMhkvFh1kmybUegIWrsoYYp8se23Ip5KAQPUXBUS1GkZ2KBzzYz+G8JBRdkNG9rK
ZRho0g2lP8A6r8heC3w1rs9rusazv0DM7BniHp3ZaHR2OPnU+6uUQoKWrUUk4ewg
w5VLRRsAqoadRZBSkdJlIA3H/4kLIJPeomumqYY2gLQmNBeASpPVbxzhoZ2C2kLP
OInVSyvFrjDJbO9wiTv7WSidfdEy7pqkyBSrQKyuqh2F2EWBVCzZ2Ki3w4SqgDME
2wjW0nLr0YWBYAdyyBExFkrOwTXSRL+/yUqKpoMP0GpN+JIzuHcpX8JoKqZ2usCR
ptF8rDDJZ3jU14fse7ZLdh1f3oa9rInKcPVVNHUA3GboDmOo59Eeys4GPo0kmzcm
gELtOCA5d0i43eCp2c7ENXwcPyk9hKznka6oN3k0MShpkQjyrq0WEliw8EOp2xYJ
v7Q0cr74sBiW4XI9pfryPii0X4x7zi01r2MDsoENFbLYSEDUbOrCLaPpxWF8nsKY
VjyHV5j0+TgNye89YrsYjGLRG3YykQnjeJH5pxNKP7Q3H4FyLSTpbWMDprU23uv4
9rYjPoRFTwh4WDPtmTjRs32yxxThuvOCxnncLur2nndD1rk+Ty4x8DgQu1/q5ASc
OCmAAWMSTniBAN70A5wtyaMi+QeEk/KjYD/oP+aVuHYzItC7ipBNPuxob6DsBkcM
PQIjtoewzmjDzeg/t28xJdGQ/hZHhuq/xL+uxLIMohuWV1q1lLZUSiS/Sq8/tXHO
kO7pOHpKf/MPkZyukRlO2rz/KyYf7RH6AJO4Nvdn3hPaDU4QdrBShRV8xuz1y3mN
tc9XYpOmJJWO7/34N96CqEAsFAVhpxURgc/5y/HvZPSJzruHNoFcIcJmjE1qtaHS
IKsxrtoLgOQHN7eDNVaj+JcReCkvLshi2l0EoXo5tTcotA6JM0U5aXDOfrqBMVqq
Zd3PL4cuDfw/Y2MrCIZTUvkpqgPwDYgmN1mMlNr4auEI29ezVMHSWgBCn5e89leN
IRSFkRKw50Mr0G8oXmO6rYzeK7HsKGJ818R8kM/r/CjuOJzJmm8z1B4Lbf4IVw6V
RIpClFc2FO9bY7/iq83wLgfi2i21jV2rPKzq/lJ94tgMeaFckKa4+GfZwYwCiLGQ
uCEDxHl+kQytWM8l7VOzvtwJm0bnJmtj4Vw05o7zCNVZqvJfGzEAcj8dMTZfNGyW
1wRMmLvDBgTyEPkrEKdXT8mUwOx1g8jPjZ6jAgBqD2Nn1+9dxhBHrGmXvTb8qSzs
1J4cJfpwZDcHi/pTF81F0tn2LM70c/TGN8tfULiEKafS7QyYkW3nrqtJeYL3aY+8
vIJpYygPojWZfmi/MIkJrhxYNe1CcaNpzXvGBISMLeaM4MeKhzVSNm6TnaDLvN7p
faCExlPVBXjvXjnXS8my50vJS9mqW9tNBKezYjm7LEzUeNErLIYjiqoU5gsIn5hj
w+Gy0EK0CuXmCXBg/iRFSbu2vCDXKvtkwTxdN6c+pu0p6+Xwb+wrZ+w1WbLtCXll
/+RxL+QozpILyY+bMn9J54YTCH8+SiOFdgRxTQAKdghiPCyp9N8t/sQD3fseF3qh
M0Sd3XxgQA7Q0YKwAUnQ1EVT5RyH71W3jhI2KUIU53RBRU2KlTnxDzSe4Ek86R9l
ilEh3etmBFRKv+otXjDYmZIffrTsSsYlU89e2wJ15kAWQY/+Kb/SvUFDNJevLJ1s
kb7G+FWwXf29mfHV+mq4aBubgZjzRTAA76/O05zTOV0j0wmJWaIKjkHWvfDPPxCx
NOCpRHmSEt46f3lWSA2VHw1B4L8vsAoPorDFeIRgLyBrcv/UNXMEM3pMEa2kabUt
P8bVMfM89F30uqNlwC0TVgBmXdGobGDVVzLDzrXoiOWB2obQC6lzKAn/h2Xrq4QA
mt5NxSdmLrKuG42611sGEwSRgtHK9AqpUX9pjI0GIT0xP2TT7t/HGkGhuzWwAa9S
1JzG1bbcNXQgPM6e/fmWWcsKRny5Fl5/D6mz825Ctmo57jUAarD+AmryeQjpqwnr
XhGfqH+DszNMnFGLYusB6qfXZFUZyqKOhPRTqvAZenqqMg3F0jbIp5RKuVuUnc2l
z+Z7Tb5hMxD+ac3oW0oxpBJdwuxgYxz+vHX3n+maSB/+YAnABsw3grKOYi6b0SzJ
4wbJJF33kFJd9pNusurrK3hXndpLtu2fSXzv1RSCmxEhWt2DPT88YhmI9rOECNCr
4OOdr8/3+Q/Nfbqmqv/G399d3yH2zSuXv7i85ClQD5c/FPc+2TrdZ7vrry6ifkFP
fNxOdmpaz0H20TbP1gzTa4DtWjNSjQr60mwn5oJDcyIHnVWCE1tcIvfEWfo/Ity/
FxZkuJEsd1R4yuUFfPvDov1VIcNuJntTV9Pva0JhkTB7L80q2q1s2bcUwgWLLbQE
uYPp78o2a3jl5T8ZDaXciEzf/5DH/jmF80GnPO84GFafzpHvjuu36uA4aJ+Farsb
v2kR82W5TXAj8I4H0hj5hzUjWjwfVmHdBiX96Jg1+1FIJjDMoiBvaoiU7GaaMVeK
jTs8SpxMkRUkPA/xtnU/3c69w+mF2c+KUXt4Ax5OfH6EWd7v/vmuv2YZOFmooJAl
lELgHDeVezwAVzXM7rmoxDBitGIl8ClfkVyn0ll+96T80C3gjGGkCUetp1CIU+7v
6V3PN7hrX4M0Ruvxo1IjFgSDzW4Q1si4WTGiHNx6f6PIWMu9pwK5QPdp/u4OU3Me
tNu/E4SK+u5wHW78tB2fYCN/749HYddbtHyDFvt8TlOBttD4ss33B7cMW0pgFBpw
Vx6/Db4cDrw8EfjOb9osYE58zSkqQoocFJlHsQhnGTT/hG5h9JC1Wsg/lrdtV5Sd
3g/gA3EVfcwYrWfCtKKvnV2Ql796tDv+L8VV6z3Eh+i870Z6vuEvvPEEwgBA/HQp
JcdVbKJj1ly+W9NfEQIRdjEiV2WUaQeKuwLJ8n1okWXeZPWWo3EMJUyYgTPIKwoh
EaG2+OdxrvRcLYqewAI1NtCqdTNHLS0zkGDG4Q+3RNY0B6AQnmUElboJtd4vzczC
+w4TK2sjRgT8h15wfRaU8mNYDKMF5PhqEo6ELEVAOScfqj3+hLtIpOdOmK1Zsbzs
uKjUb1B0KbZmYGqmFgRtXZJzTbAVgmFZ9fHAsSqQlF2eVdKDpkkyyQCCrrORj/6Z
NeiqMsIrKthWfcfeJL3aFuY3xo1onlFJq6NpUYk75Vpo1NKX5QVAnnAECAfdgmNO
UMLQWZCuokkul1/cPhMQWd8nVRV1jg9hPxrqTN0duCyqkYd3TZQD5LwFojy+d6W+
lAPU1y6T3/XrMON+e9g8vg==
`pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
XmfUqbEwcecDksOXmZnbtFXXxOJIyIspcZWB6cXuQ1d/9Ewli5A4uCIu0ihfskSe
q1nNHI/muGBUW1nN6kxU81VYSaZmyEJm2PMxKYfjiMahNdecMG0cp7/rItDKfjtk
AH2fZCLTN+DMAbYRBupIe/tV08zIMampdsJIPxLA38k=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4608)
h+nAq7l2YCRhwnd70WUYu1CS9jGxnoeF1DTNPDaK2YR7P53ViUgQlpq1dRXxKlLx
Vt9cVt+f6VCvKOxoHXm3LM06Oemv6WCNs5Keb1h2UivYeA3sVNNerGV91X4ucsuK
0TY1qcjt0E9NlV+ALi3Amd16dCaIJnVpQqLT2XehfX8nxiqYyXKiFbZTt9t/BuKz
D/ZGDhuzu2bPHlrtYdjYdKoFuDH9ybkLlVo5jGCz+0etU2E7yw9D+bV1QDffwndJ
+EcfxIXpCCQUZLSdcrFeWShC3TrqA0BTGqreYO9xxDuCdrmh+iijIKSnz+6oISef
68Mz3etwjyOSDFOZ5JgAH/LvNqXUpT8IBngLb1hbEFIJLOshMY1NOHUpj6vxxghr
NEc9gCsdfyRmxjwYurnSKabALN/GRAHmdbYpT8GOPFNpB3Tl1mUXglHkjIlFMONe
vNgdXuPRZ+/pRamiZjL9/u1O6kysExzGiSnAfo2IelWyYi9UF9xaEe5VkMuYu2Vi
RMSsbF6/avqVQbR72PnD0Nf51hVAlXplU+LOz3EUo9DuN/5c78VQ7yhxDR4t85s2
JWPyUE2+nTUBoTzOWvcl8in5C508OXg7a/eESmTh7XPq4/lY3ZZxgUQXyQToPXdG
8iwG7SaroCfuV+sTPPMp2Ydge4kYwGRPXuUfqkNiPu/kV2Hx1iMBO426AIxBztdD
OBEayZwY+7mMOXlpYVnUK7IwhfWBjGz1N43myz4jLuG8A8ELyS8NxdVIXXtRdWdU
cwQNtcj23nIwOIDj3waXrZMoYugb+RzEzPJjEXkWXrK3jTjtRDq3PCKfbL/s6er8
3bfZzQOv9J2hfQhITQIZ7squDkoASqZ8+axRrZjgZwPfjpbuITs11I1/zLxAQkIa
3Mbl4ubqNARzp/sL9Ms/99MpXJl7MCN/+g47KURDtuZKmKnPPktBx55nUqDts2wL
bxVnVSbYpXXLnNRaxsLdkeqzzHi4xr66plIttMgp5xHFk/yrmsIjnS1lyf977dZM
JXVoe7GKOiJEcZbSw2iUiJ5ZycS8M7cZz+2+BfmHtwho5VmZ3xFdBgHRAQz/iu7Y
M5/xmQY4UOV9dJOUSSUo6quZqYPdlPCR/cioTLo+LtgCSHf2Bv2Wgf0Z04rV/cP8
WkFpojYBJcIbL8SnpC56+UneU76g8hvRHJbY7cEYr4HAzeVeZgQ3KfRFiGZOhOKJ
tPR4h5DrLWJl3dRRn9SBdfrflr7U9TJZGchqizQIA2uy6gxj7DbIBXbCFSzlTH/L
3l4MCIBGEq2GJti5xR9xGP5sgSBC4Sn31txURn93cM3Cf+glC/tu3jaxziEyqUiL
nLllOAbLcYD6KhWa2IiFaDtvFHcPvnbre3MclZBVechznbKAtNfjO8z8/uBYDXNh
qysaJdi+PrKwbsd079OUrgCsnh8b3crmpK1oMjKvbj69nLwCwh8oaFDjmOZpniAO
hhNFGK9R+N0cxz9x7BsFintiLI6g4pkZCRW6x8EvXWy6VTBQxPjGxr4wkt9VNwuL
sZLH/gRQYzisVOaNyXo27LoTv7JO1YH2Goeh6IgedAvFMmNAUof+mHLH6MM4sks3
LsVC2ZA/8WGUIugE9Qa/6w3E6si8J3GyUyRqeDwu89NzQLdZDjEhAsPiNyRGI6EQ
Q/36iSeg0wiDs/w8BEHLMXSDAgKASVO0LCFxlN/VwCsZV9vJ4fs8MSOHaW/28VWo
imO74hsv/fTtPPyZkO3sSaBm4Is5AdRVUmwRdsSTJooQfC+PL/3Ny0aAdG2SC4qT
gVxHWEH4UcYMDJkfS8w/pJAJVKZL788AGZE3JktnNQgG3LGZ1Qg4jaqAsd6PCOUy
poAB1B7vFev0I5IpFcQP9w/YfPGfWe4muX621vQImFF+nyX2pugdbZCrO+AeifhZ
iJOI+f6Eoya1sMQaiKr31UR60DZpghb/3CvowHgBcWfvNM1OsxjpH/IpxQJffgsl
5+ApLbyvqqeCGpBi1ZIyozDJE5MtQ3GxEFZI/tYMSg36r1anbapnOJJsu3Q+i7bD
tknLBmlpQcLfHDosW8ZV0g26CILE009JyGA6co7Flr3hYHfmLStzKeG+2TBEhIkn
NcqK3xeo+S3PsNlwnyfJdbwz1K21YWxrlovbadXSicb4kE1y/frUQs7SOh44J85z
IYx9nEVjPMaCf/pCwwNmSuchn+EnwrFrOXQdmtZ/3W/3wh2qf0gxxnONe4pDmgNP
mNSCWUEbSW7ciONDAjdy6ryrwnzJ1V78hOK3+yHkafwocIBP/i3PNrqrv8rQVsGE
Mj1b1B+AIrrY39q001dqEO9lvlX/3cSEG5+KWjMINBMHgm0M1LGmBpc30HZ60ITz
T2n26fHcwp1eW3qISGlYig5beVWP44ciRKmEGz49YVkyoYjheHTYj7ZkYwhQa60X
cO+fhoi+PJgBUcwHFek+qHMiz2sQEvLbn7i1wq+zbLyGZToagulCaL7D/FgZ5HJV
MLoShiHOvkHFF4UZGlru9RU579naCmPFWKUh36YWF2p2T+xnCxaNocDDeIdGj+s8
8NbWFEL+2ATvaM2qGl/x+xt3x5a5D2G8nfoPH7RRWpWjmu+aAyiPabKZ4cCyO6nU
L5D9vy6ia8oal93ymrl3XlfPsKV5ZMYiokh7KS1yct7D0dxmJToHlF46VNOIaccM
4odl3E5Y5qls/St1WLzgsI3VmTfU/E51cc5J7Np1T+9LMHrd+lTPhYgYJ74qLKoa
1qr4EHszzGsMkoRXzgE85k8gH3jos0p9IXX/ylzzuzrhbN/KvwKv+9YGfDAOOp58
bOKAEcBVeUoB0PL0ljbDuQt4NJLy/q7rmjK/nvxhqWz9tMqYgit2AdtypWkVk/T+
sZmFIIvUfCayfLX/Rru8RRVc51p+iiiJEkXesFQxnOv0MlRmRRJLRmiKDcDhZ09R
Q30WErjMWAbAmt/PKVnWAKR91k4i6c2rMCVI/tX7JfChrNMFXeYeZ9JUOqWRLVm6
UlD3s/GzPyFzVjij02mAfQhFERzgI7vDvaxIdXXVi7mXAUmf97GUD/FdAJlvuF90
9n1G7TqszQVsaT/z4C/3bvrwAIpuv/GpoxN+58253Kkf7r5QYscDNJdqZYnb87xQ
3J35Am664PkVqphz8pkkRn6VCdLiTf8YhKR69AQgZJSxPfZj63YTjjIv5gyWTAab
8aB5L/PRse6b2p/BSPU2/9ZCfHUZFpN8SkdD5CQS2Vt1nrIMsJCCDFOfZuyoPbqG
+5jhXW7qygXHaO5QdM853X0aY2ZNloxrZ50CEXgS33qIP+spCiAH5n1H/uhFNner
SUHGFLabmPl6N/OPVhjHQWoFQVahnX0lpOfSNGJiLHOu6YY35Jc43cLtsoGe1LUS
EnDNDowaj0yMb0SWpPBNt4nsZfzlTqZyfb4glJdBrlXVwMdg2CG6ivd4y1uyYUSP
8rB2mKmTCQGVAd0AV6BNpYYlip6C2uLcRCNI8SU+UTHDwCE8ydiADvFaRipGfwmf
60hJABjZtx7ac/OdKHZyr8Nh6waXeovpkpVjzvaldi7n8j/tPYUN4LQll9EXMGy/
D1+NbSReETcgT3YvSyQe+Dij4tBcMVJC2XE+9OsJQwIKPVNZANVJ34UXSC32ZUzY
7PJ10LeuUYXZZjampWgMpxhI1r2aibFE/yk56CUxJ5PFwkd0UaLa1X5gm89CH60Y
kBfTdVTdENTd2GVD8v9zLLnPirC1vOAU/z/91QHnqweWZCKBUIhQ/b5nMOZBDPLa
2Eych4g1gcDaKkZRlzbx1tCTedeHxM6qb46y63Ptmm2HpDjKNUvuPa2iPTL5vh/P
ljrxasri9AWCLj/DohXUllTeoSgUHPi1o2wWHvK5RyvnDcHPga5sIh0gxhxUyd47
aMR4befZk604TcnZuqS9SPh+gyKMahuJ6qxP99Gipxdvqihe6yFNH+l6s8LOC8LS
BATIP5hDqnKPNNDvwWMSzAcgmlBSMcoLXgDLBY1KRVNafl0xYi3KjIs/7N1WlPcw
3YbG/P/lygtTj0hvWh9Q6kmJ7l6n+NKMSp2qt3gVhD6IURF7zN57DsvXhX5D6kNp
2tqsxUaE2k4gEbmEyYrIN0VB+bwS8HTblSNdIcplLJ9wwq0lLB51q4cFbEurJt2p
YTZ5wSIFDwKxbxRUiBThJV7LiB7ghBj/0K6WRPBY23bUF9nMeekKJHF9H9C9TvtG
PQbJ619d/wHSxT0TQShzLC3MTV5LrB+l2mHyuFe3hJwD3sU+IB1HIznm3JBsEyP5
rImMUc23ih69wiJTXTH/VqAMZxXR2vl/S2ZBxNYBh4y78u1SnZowQI79M2SAbW06
qaJ/BHCpuxcWt8ivtcM0USmw45d6LWmJlqp8OiArGY/AqVkdHBS+q4AgiDtuiPf8
EQZUQ7hhaSVZ04UO+ixYLPYYkNjuOIBBXEYnA5mMABbZo+F8/Y0gjrXx24OJLAXg
r3enqCVP2tfXW4x0NoJ4cgz/fm+R9CCLP78W1HyKTKGjUXFBLLgX3CsDpZLQ/kCC
uZVLN0ISY+KsOlHLTJpb0uwHSC6e26F3LKWeVVaYwXfMibPSMIxNfNZ7avq5iuL/
tGui/kY5mySvG6AXrR/woVWVdMu7DvHtPxpQwPF3JZOLFk7A0CxGqQfYd0Ywie4Y
CoHyBeE6kkdp8tme9eSYs3lUbjkAygl6/Q34KrIG/oMqzsSIllw3V2uy0qe4EbkC
8l+DNyAoPWeQl2ZFrgCfV4IgrQITqa+Nvv1Bj4cPKrgqekJCXwzmmaaQk0rG/51i
GTxQAnvl21GnW01v9VH94i4xAQych3nV0NOe9Nr0vm4ZheXUFkY2rYUBeJDLzsmt
aH7pitE+kqVhmiRJJW63MMOmsOihuizkm0yvCpqLJNBr8tm5bIf0iauADNYXEvzS
VdN2aQXOW+1K89GaivmhCGdUH1rIOmGlscFALB87EVVMRUeqCPK3UKeMjB0N6qwD
6Pl70cWAhU0a8xRPtkIeRFnS1RtyJZEghUZ93QXFFcbSC6f8hA1LyYwWupOLqMCt
FtmgdgQFt0cvcZCjPkdEgqYDvLKYWDMvmZU2Q5ardyqgiPj3YV8TvYfBmskZRte0
S0mkrz3pbLYtfLTXXQLc8f5rCg3yGtJ3rMBczQV/JPpewJDQnyO/PmR6poF33Vb3
GDL/zoIbVyWbJK9UVQ+R+Vd7Y43LpmGyU7qaHNGL9/nmbG0ZXN4eTo0ShV92tdac
RfEAPW5rhqWPiheil7DhcPjytf1QyjOuUJtYTs77OT4Gfek7dArtFJ1COQEftbvu
dFEHa0GOB1ln+nvKnCSv2hNmecbj+f3vZk6wC9TEevDk8YJOxTo0Qe5vwOJN2f5i
D0MfXNSwqQQww0UlPia8zRklegHTmEGVf2g8VqsuV4boM1/l/ObHO8dYrFUlgCyb
Ta8me6o7aQE1lV2vWspXl+qYwkjuCrtM9bAZEqC2HnkG0LzTR1+ohfTKc+EyxqOE
RrkVKYQ3fN/l8523gCB2D9HqM7EeEoyhY9KcpXrkmRQZElJEMwqTz4m5ENdF+M6W
yW2vxqtLqHGTFkPQZH7AvpYGAEQkkPx3ESxbD+/jUx8cYY1oZqOwfC1EXLOZ11db
9TcCuoqhRsYz+fgHi8bmZx6dbD0cT1x3VQp+DgT3XxAMUe6/lmkicZAEYxX7Z8hM
qyHI0lIk3b9D4lm7dRSpwjFsa//XqnqhvqGicXBG9XGwbZXiidJXt+fEFj1ki8n8
gPm62Srn7oxKN7ixLceERq00fKUD6jG79UmrhfxY0FJQTGjbesLpVL+56D5p0S1T
4IokjmuYP+A6dryvtENm40/lqTTkvLMRfSjRQgnffMWA/yciz5bUqyARJs4HMYSc
8uccxrXZnb1+OeDUcfX5psjKypSrxQhT9LtjZeZHtK6V4x2OKXdGdiotE0il1kFO
URJT8jINpalz3erW5NiPSdZwjr3hrKtY+7kJRoM6rFGXgaZskrdYB+f/YqG5qxHW
cmwGfan4Y2XtaswAmhOdeZQeyAAxMTz/OrmlLXXeuSJU3iaLbxQK/B9qdhvpAGYd
PFQWOzBSo6cnfSO0m7MH4e6Sv3MA6NxO8Rvvyd2vTG0DhPoiZfLXwWOHQqRdjf3X
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
s/TNZO/cDcfyrWWpSHUvFdHQK3xqs52pCihUOGRcN7++Pi00G2oDEaBlC0OQewLFzU2+mDB5dbbw
A/SkDQNU/7PmE7SL8WUJSUjRcDrGnmsiUjh4IKfsTB3KHJ5fPcv922Szu+xd4jatX6qFISavtzB0
mekgsheGN4mg/p25kKhy1BP/Oxs8awBL6rSuek+l18VJ3CLrBmIYEJcs3DsWKxzr5jAFLvF71gse
iBUkUEO4jaDsCoaZZQVYHKF7bFV2O3lYM1xUwyTKhm6EcFronhe7W2AHcdRbX+tgzEZxz6ujCwta
rgBjmbX6UXDBtJsPjVb7bAaRG/zaaSTUvX7ucA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 6736)
0T/ZG6ATeZMXLlro6fJdgXHj1zLpbXuf0WOVryJF63MXoM5q1+Zyu3eMvTdUeMGlE7TKNkvG7Ifw
0XoucQKRPHiByA35yUMyrTg+UHV0TeQCpSIVQYlyRa9bhC06CSSd97iAB8AeZdydK/58YZDv31lX
FpKQr3LGFWKy4cbPPks6ySKxzQnjmS6U6mWN20mjMJIzOCp7aU6BMK7ipG8nyNXYfR6McgZtMrS0
btQBqwtJsG6nxUoWiR5fAPp+g//kHgrpeqU9RoHb8827KHBV5ewZyttSO7W+Z2Xw6jimdx3S6qKR
4LkjCNgW1iQOHrHqyY19mZ7qSbN6gR8rsfqVkkbDcXNZ8kOPR3KHL7ovAhRn5hZmczjFiEYcY8sF
ltan87WT1S5lBFS6qu6Br+gemw2W0ppqXYQg2vzhnXMyuShVIwqKVR2UrnfnAzQAvZgOS61GERS8
bhoKO3iMS1yE3W/yiLNLgL11dfUsdBXCpiauOwGod+1lnni7VKlk6337uzXhvCXwswP3iMrLOlFN
dYccsO/owU8+KwzNf8+KSskfhUL6n+o9fdR12Gvjwu+BsCSvyJNy9A9LewfYyrkgy/njN+UtaoZk
HmdCBxlkC97Clecj7uSLrYBicgogyGujKLcWALWYH3neoGs5P780P90HBp6UPYtvixIE6srb95Cf
zwZmkM2uS4nb95roZo686e1MuKRzNLi03SzlzIMUdQpltXeKSlWEQXafxXCuybsPQ4/tHtGxgJRq
tz0T+o2XQxs0X4GTqroVHtTdSaGccsMUxIEMW80qFWDDMMzbGISUyDV0+EQ8hSZHS4PoOGS0yH/t
rb/KSYYTRY5v5ZFBIi6ihtvz+2trOGH9wQzqDxQyX3Kb8htIU+Sp5mIE2PXIQA/ORUWec0LDgY7C
KNkg15Ng1TAbLaT/FuTvULAn3GJkGOoizOPpR/FIwyGybugosS22KkekHBN/KdvIVKcBz6o5AhE5
DJnOLrrU/ZmTqVSdVt5dYbA08wxBeFiOFBt8GLqS8jFHvrxJ608eAyDtZQYOO44uapxeg6dL477g
NUODOVTiG621TrpE3QRI9oxwCCQ1xhDURTBOw6T5Iu+SU0X9Gtfj9Pxtt0fi/g4YskqO3+qgDYgX
fKW+m6KBrLj9+xtBPOvd9+PTc0GvkyNFBX3RleSZtLGhx0d1X96llJcekSFRB0jxrtWIO17DBEPj
wPmGRQT+v+o8gZmHvHLiMvE9fYcQ0qbP71QFXD7iiIiaKKoFd3fFyxwFp2FJj2yw8bW2tOGa164y
XzX6sG0KbMcnLzQRkq9avAsBMJNk847fcRR3GItyuQl6Dx6+82j9ouTseVXlJykJxY3UlxjpHxz7
qwvWKT5m+V2cdrmGyiprsrFK7rLW0/vCaVc095KotTWqooZXqW43I46uHX7hlUSbr4kuVX7M4yyw
hlmpa/QSlPpEH+oAVK2+XPf073ly3PdWor7xnqh/gL5JKdvIYvHV9C3A0dEfkOK/SndrtgZwUmqR
Pz2KPZcUOW4oioQxEIe7uvNFuMHKBgcZsyCP327uokdE6+RWimaJ0bQfg1o1ZJrAYbjgnYTaYtYD
F1SSP5xemjSc/etGvjxnygZNoB8MJKKqGPmwuHCWaoy8z4AbhyUPcUhQHbMK9Ti0JXh+n51HPQir
Begvrj3XkUGvNsX4ynG1WCtWfGl6AAD9QHDojZbcENE6SXv6ujPM8xfCw7ZqkWDVK5YM6wyhketQ
IH4YxOkclJPNsyfT/pWskM2TtZ84vPJev25iFOmBBTKoGB7d45gaaFp1Tfs58jEiBJ+uPvkyMdlD
p8enYI0UvRVOCnGLUwscFyYjVPF2jlHnLBl7kcyCtJI6jlgg616OXJUvUaW0tvxzoRTqNKIwYJ9F
ON4pkD5vx4dyeiqC8PC0UCSPVk1erExvIO5rwttIhDi5FvEsnqyQKVFP4ONbK/MNAUMTd2p/iMN7
wP91FhuDMvRu9+c3Q5kwq5TWvuZUwZEkm0TZbuVr8k5bibidCI5mmWOS1b+xR+PqgpDcYymzKNQZ
76mJyH0S8teix+/eZ9QMc2wSHnovE0sUW8Fmxxu9Um0+PgDPYU2rxZuWZ6rJAQehI7tGVrF7XiOW
4+UVY5KGDgOHNhnfajZfrJZsqscDxJyF2TiYZcTsQi93I7qkUTUmvXJzsHr+Do7MXq0P+M8oK1Hq
zHLqyNl750LLuM8VE+Ro3cZxUH/NzFy9uzC9aMmL1aODft1N3dRAjCI6cRyl5long7wvkc8s0pIF
lg6QmQrOLYJ0dN57spqjnQ5QYW24xMMyCZjEheSU3cPTnzPSrJEll7bMTVBpJ0WdfXK5Jzi4Wybl
gT1curCoRSZHiGPlhGOaymkVCYvWbHqhu+0wSwAA7LJgOUcSEIyD/VtExgGXjr9OM9tB0L0d1/7M
2D4RfdXUJh7cArzMSBkH7N1eLXxVJBhs2Cc9XajIhOtBC8hvMqplysRvtXB5sRl2kJ3VeAPpKZSF
bj9IY3gBM4gfvkcYTdKoj2CH6Ajn4/Atl+rDfhzSc1GQnxshlWwglqO6bTKoqw9CIlw7UGUbFlm1
2RzBr8wyytXH7oYX1MAPvdjEqUTAHmhWd9K6znBG55BAxvs8M4WexqZIZB4mn3RK6Sv5x1L+J7fl
fUdLo9rl/nM4vZgPLyjqTNeUEkPfCk7pURoFC/F0mPHUjtJaXd+rM15lD9YTUFQUPr3+2t973Ysm
aiRKnK/2H9ZUtF9uucfgxel+bxdtlCxHTWD+QtOsB2vmJ3UV/1e+8meeUfLwURVmmm5oRAF1hE76
99YBsPwgGJAN9oKm+1SaaZ8PMfGCFJspE7z6HJlB3q23vb/OnDB49xgmwTMjprsBAr2SvkdoWzS4
V666v6UXuW0jisVRLVpJST9HvdAIpiqgi//++cJc3zICYkggwOE50gf3GjF8dTFxHTLq/SrC4F/z
nhpmR45ZQ7axKBtNYnH/HP5y3LZgf2k1Th4r62YFOBUwjDcCU7XscoJud3DWbn2qhWXEvTzl73MR
zV6HFxb5PqZxBe6367k0/zLnStuDsBpuNPXMbRPrwI43coxBBmym1XbdYxyxd9fK+UMb51Jb2Si5
kj6qRCAqDZ6Mo0D7f0OY0yb5KtQLkXj4fmOCx/7pryZNwG/cA84iae6fqAJfQr2C6CK4JAngTZOJ
EkSjoievoGFh54xruAUswhJW2r8TZM4Eac2MAQr23XZ0Rh+X5RyVUxpcTrJGTm8O8Pef/ELGTey3
TdmKBZ9q0KN8dsyi+lTCv7gldugLYq+6nX2W0gEX7HkzzfBaRi++40To/cNAjf/A6nh2Aq94eIv7
YebmZyARG216MLehv0jYtNZarAn60TQjmuZhgn10lEyyi4xxsva8mYbu08O0enzesdZu6OPfHuUd
blxdWCIg8c/4xHZPzgjXYi3V0j9vhsar0FIMk4ziZxu1pNyCgcgoUPGWxtMuRyUHy5SJxFDTtPq2
TnJgQvX3HjezyqziCrIutK49VfWg5ruEmhhMuEU/9mHdmW9cYSMgUElsK5ynekVPAeXeU26wdn2P
XhjDJPwj5Mm2WeVOn1FVeLvGTSRW7TRMy2fCdudrWEO98ce7Wlc59U2hGL+Q6cqWx1BWg+e34S3b
htBYSkcswS7TeE+e9M9sL+yETfFd0FTud0gJkJn64AusJ3rfFlq2uzno1O3li5R3JNvXL5xqkoWx
6KyHFFjzWX0PEutHI3G7/sCSh4eK6XOnrBX5/Dw32SscyKYkhkuNA7RYM8j6yMpSA9c+Fw+mDu8H
UKxSoukgNs3Lu5uKfARxY+olavrByAKCTm0zIRWfX7zwakuRSXjQWUqRJed1u1gSc1Hppa/+D+lU
l6jrugakqdJYI5bDMynuRMVFhm6cDLUa0HTVRGZbTp8IzISMHba7R47A488tD1y1Wp9F24qBLY4d
NVdMB3qbx2lRmIqDkLsJofG5DkYSuD6TMD8/pfnmmgZwDtNEOsbsdyCz88PVHLLkFCoE6LlhEU6W
AeSfiDg4aFGWAIP6JX7ug/1SWhl63GvTZxKDHUPewkz8BnnYR/45h0bPzQfo1+CT5wdPR0z6zo7C
i5X6yAs+KRg9rRDqWCQWLiIrN7WP2f4eCPWTo31GTGeNE9e5pQKVzQSIBoE2zCkn+PCCloKRy9v+
z1ts2RBBJyNG406U1TNXvTGUEoSH7V2YT32Q7vyItQXHQD8GIsmZrd8/xzuoIOwUTKfokjCfwUK3
9dZ4LwEe5Clpb9vWylyotbcH3FzjL9ZuHOlG+26e0M95HVdFRQKZDRrUi5AzbxkVCOJkg/apgtLu
hmY499dryYNtNm2aY2DzUSL/jh+R7lw+jAt+vcgHRCHCtrCI34zd50IZJPsIFpIDFrKU17jC9MLX
QZidrJmxwbKVHSiq/SJydjsy5GxfBD6S3JzU1OUI/xjj18GCtxe8gV+b+xvtK9pCf4hbcQQm8NI/
wUzk2JGJ5d2bhXd99APPY9GWKSva5UhC8hk70X4iM3gp7es1Gu9dw6Km2S53GJX6WyaxsFALML/4
FW9J3bW3mqjZfsHjghP2farix8s5KD9FcXUOohZtl+FT/UOwcj/Gi0wSWQX2FMwtYE6ZpPGC78Jw
lECDrixLDIR7wmJrAAeuJ5Lhi4QFsR3IB6lx2fUY51K/Wu6qawHg/GfF0jZFkkbblpgX22Qfd8ai
IUoLKAUOubnO7HV3Qujy52bJxyt0DeSeI6PnmQkOnjDMa453mn3mTmTMZmQ5kfACtx69VLGj0FZ9
m4iFpkPwodClUJ37HFq6/QNRKxtAwFtd0GGS2mAPFM/x5v0xaVlK/Nc/osi5ezgAB4BS7iyvhPaE
blB6AH2WNjtVlwcw5gFxZIK1OwzQeTlB/8Cn0wdarvV0APT0tPk02dEli8jLHIs19p+X69OeatPX
mahFmhyHeAWq8MnSqlaUR1RTyS69WV3zmSFV5pPMUs4OpbeI8rXuaUzCl1vfaaxWUsEREOHVA+V0
yw6+11ZNmlqclszcNzipUc6lXsECgK0Rfs9qDaGSo9R3cJQFyzPvGgqkUaVjwFpKPEBBHojZAowR
UCpFI/0yvO79v2F0yYlNN8HfJ+pRDbe4Bi2ZDXwQf6r3o0NIJCPBOfjIT3rbQY5IBlXZW/4HxRKo
FfyrD6qCyZ4iPIh6ZdADuqSWYwig6qDjB6yMpqrzi58TPkwOpftTXMpMmZkoDH/Zd2KkDsilTfP4
QXd3zxK+nPT8cq6d6gKkb4U+ntKcRK4uUwePoBVKGEnHWjFmGVWgt+Oma23OPJcrs30+ngggrcw8
UK6d/9VxnczRm15YAetCs6vU14euI1ug9j/WcZbWyD02Wh5vdkMbwUwLVMe5tEsWnWbnvtEZSkbo
8TKc4aq+XzGfbAisQmfLCGQGU2R8TS7RA4Q3WjKb1osagHqo/1YE2P+YS8/9W0AcSYt21D+flwXS
CXZXj+eMs116b+Vy4jO5dMwDZGlK3EUR2ZUSa7FKLugaoWVG8HjBhpeQGozslcuk/YNVPo3glitB
nu6F5tdu21WPqZf3OPxiL+wLLT1XMo8OgLySrQazqQLMrs6DPzjY/0JO2b0bLbskF2m7/qT+hbMt
yoqZxNI1WVxJAlS8zcACAe6n9QTPpN/ZJ49VegBUipnALRr/Luf9taeCa+BaqInlAQGDr59Gvagz
ktRQ1fMnhBRgIhISOokF8BOA0DsTGh9EM+XObhsMby0cfR2E8Tg7t0MDYtHVNGSNfF5hoSAomSry
17HcQQjFXCg+MjfnGhGasoW7gQcfKm0uDzlKQDdPapFx9KE2jD/ypJCwqRwVf3ITcRbh+3TLf+I1
ZyyN7Fx/7zzsp0tDTcC7BPk/LYHxW3c9mCNp2qgU2AQS92jtFGhfjcCC9qBob3zdsDhwxayC6PCB
cFw3CZBYD2PQaCD4LvmnJKhrWTMfeY57nci7oMNEPCRUgeYhaxanz1uxscqrnxrn8Y5oR3hGMrpC
OXaERqLPpBhMzk6VrgITi6idGNIxe1ZutWW8SfCm4rAv8Vbh9HLSXZN8KrqxfrC8JOm/Q93xPvPt
p4YJlUouUxZe64wiPpg5Ejs9Erv7viCXur7W5HrpxFs6oMebQ/lwUUXBqt3fiOnH+nKKN+md7jOb
dbGIBbPP0EiCdmBLXIDi86js9SvXKIiDfpUtTu3azbB4L4j7UDlnxPVxHs4rcnSiM3f/oZ2sIv9K
Q+/ZE5nyJNdL8aS9omhB1P5XdEfcwpzAbk37VyNG0v7W8tdY6XEt6q/JlSagaSI3/kNRIKVkgJ+2
LT6JWtYT7o3877YwNl5Msyk19HIq+nv1HSU6w6tXfm1SNSqf1TC0AZ5ZOIf9YqO7R4wcvBjBtx2r
sAUtGQc699Ms1kdTpvhJSe3PjlJcFDzBRDo8YMwOJ27WBd5VK+V1HogSgotTkvaz8dCXh/rFv34O
9ITPwgBXseT2/GrReagX01TwFHz14HbEbTX0mOV3AA6CQrmB6mtqmP3Al+1o8eBumUS2c7XcBufT
UICdINlQy1a+9BUAoED3gALbfrhYHsmI+lntweAUNYPYyeTra16zSNdX6ROhBN8p1jVb4AQu9qTo
hfX74wFBRO02HPAXYG7r7dZaBVIQEW1KkzlIR4glrhO67IXkmm62E5+Tn7b1Y9GPsIsdPhqjpJpB
yKC2hNF4DtvtKD4I0g8D0VrBFwxw4LyqGUXH0+iEDTAHu0VFbwZ5lCtdylpV+HdfQUXQqmGyy/Q9
2szUymQwafvezgZPLN/LunrTr6mVbZIW8sPl1OkBfz/OALaex0shJwTf3JBP6loBN2dxId1SZEuG
eLMzD9cAVtaiZvYgHPArw+YP2k8/0cIXY29Yy1zmg2IicLQMZ1qKgwpN7ZNp+7ZR8oHoXihiQUZT
jbWkm8XfiqwRpFef9cmfJpGNH6n6SC9NNDmCEYvFgR55TKvnJG9A3jS9u4GTTKtZEddQ9se/yvZN
ZN9G9kVcIKMjQuzEb+EW4PNrFf/A3sCzMYQYU7l5TkIl/gHutq4sz/ZxsaD2xIPEdqeKqmTQ1kFb
kUTecKeBd/NXKUFeaEiC0XXNVgdXZOrzcRXl7c5gw8kEn52/hTuhS3aOwNa8zgdiUWtqmY0YLpMs
8FUNcVV/XM1M04FUqGosFF4pxZP4Mfb8aQo9yA2SJduFwDvKDW68kzo2gv26SUmNTSDApfBkXVGq
tmB3+pVwC50Yn01pWuh9F4v9DpxKXWPrsHQGuAizy1n86K7IT19Y9JumR0tD1auOM2lw5D2lrX62
QJPZWEx67vL/UgALMJNV4NLXPnmY9yRuSJx3c1tQIC5g/fbxWTYYKN5AeQVPaF2dWxrwE3+LkM7Q
xYwqQ+uXlB7mnyhciI6lg8dytPdvtqi0hoTj32f0QYjxVHYimghUgOJBmRJzSkGVtd6sLuBXGrDO
tWQ/0m30JOo38Bp+I4fH3AzusKVqXEdc+G/wJIxHMsm+uV5FNFqUZJ7VlzZMYUqXvl0brINCNG2a
marzrdOBhdn/jIPRKFDuUpyjS2iJ3EvJIxVIquWuvidDEVoFdGCdob5CKF7g0FHyjO21yapPXynm
dstY33eAmO3zTV5qg/zlL1gJbwZ6aBOR6gGvIWRXVBPg2nEGL2w31q9UYUVYyf7zQ01bUYFoSTgo
ca8RvyIxSjl/mYelMqYQMx5ol+RFogpDlH+bVTHYtXsMK7nFn9+sfrcoN1zTo14wwib68lmFuW8y
+wN1aCKfntrAuxyL52wQy3rD2TUi3HfA4N6n3kzGSLNxDSCbYsRowOmX8psmru9sKe/VkWr9XCRn
gUyco1aSdxxlLEwIRj4bhvx2+rTyFxs8eYb8mztIVaVs3ZfXfTXwVZOomwhEMk6EJIIcHzg/WEVD
wIOd876gsqIKj1DNKT/5bQZyZFV325aqB3Fa+PvhuHSAFwZZnJ+IZxnGRA62myVMwPdyhanmTjzn
FUkIf1D9A6Y0l3YhcAMwH/ZUwZJ1izym9C4eCm4DEm5KDqy/0gsxWR/32unFSITb464sp2HuBLDi
XKazuy27RPpZNs4Dxf/qg7uERimAPyjwV/iZsrXy3x44NHF+fV4qQscSuiCLAdJiX8wUuz2TVSMK
+Jt7uStGgZPFNxo2llrWHh8IYUSirRuMRxi3WypF4VNd8a7M9h5Oey6KZUk+sCsY5MLxjCmcxMpK
mmcvmkBZgjfoqe102Vv9iZ4CeuZcmTvRJxlJvwnA4HeaWt4fed8HcfaU/c9dlkDV36aUmor0kbGD
UGx7+3wcHXtTTLwUg+E9uxmg/sCsjr+M+749HaoJZSObxxo2V3LhcZtfGOa3bemSrkOoJOjZCNjv
KTfy7Gz8rLmKDuuUH69nvPgEn5MUnw/HmSXm0LMfm8xMt99x7l3v+VTvinwpKvz4o5Rr0+TzJW8y
FwjuL/qPcNe/yNC1/04afPKRdy7UpxNU/nwAxKBd172OTQjeLFClc1Yv6XnwYdYJf6bNQDg/XWwY
QlF0IoNUm8QyxzlfwfPLI4dZGgHK7Z/NrIhx1P8nLFPDAz+IJsq9Fuje1oQ6rNKu/sUM4RIdMP4f
y8rWJOsVVwZYuRUg5ITbtFSmu1ue9wpXH5nJ9QbsiCW0YvmNeBltjYphmnH1jI0xp1v9a4Oo9TWx
LGZCP/Mg57nm8eC2prV7116TZIIHOPPI93rvhYTVnRuMp6GHozbd29eR9Ykdl2UhsijY6k9D241+
CDOvoOlWXz8hDUP/397fUkymcELxnM3Q2y5RdKTxUzCAbKRUrY1DDAhPvtU4RZH2JrHrvLKvAIEI
a73Blcrej/626N2K/L8TwyGWhhnvv1bPyWMv0PO6Ocmp4hT1TN0FZ8OWAkhX4NVOSmzDV9Daf4oI
7PlkhxxotpgEKLTw++RgCHJuKRq8degBuuYvrHCi5/B/jJt4erASDipon4rw1zQXBl8+QTxNETkD
d0x0Wps5iBsHZQ==
`pragma protect end_protected

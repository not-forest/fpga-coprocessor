`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MLQV5vYfsIK2icDnLa5cBO92Vg93XXLwPqRs1F7ZrUeFyz3VL40ntRiUhRE9lNwM
h88KUBkzwqkFJj7ECWtH379cmVBIrHtBAsiEtBJzn/OYfye6Ps86US/PQbbmAiKf
91IozeFHHaLEd/FAQetEd1i4vZ5KScSiYjHQYZYabZs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6272)
yYkKmdF6mooHqhFybSh4r8I44fdXFn8cSTLnJXUOO8xDARdLjY09upUhaCofrvd5
pjBgIq5yZ4Y68RjhAm9mhq4NSRmfKH80grEAv7OrIyp2s4k+mr6RT1fL/uqmoRhe
I2ZzgVZ5Li2rNz2TKMZqDoJPTfQLRXwBr9Knn6mVbhfLvRNBb02ZaWFuEpCUXvl+
zsiqGDez7nur/uzw0HbRqTB+SENjvb5Dn9YCTNXzE30QqTL2iGbGZ11q+MtdPWvr
YqWbQ19Gy0Xtv1DVYejooZ5dzpmeRMnpXbqgiIP15wLpVmzb1EiHr7zUYryg7+2K
VgoAsmTzj7WySKtj+W/qRs57fUGdSlcpiQKabl4QbsNmt9scW/hZaQ8bRe08XZl/
C9DO0aCGhbInlUkhcJt+cWQxMeOfu3Gtg8jbq40+QzB9W3Gxf07ePQO5ASGCNvob
qnhTCMCKzt08vEWFKvIN3CTVP0qEBRGi9DUTgsKFFpUVjgtX/JMIWJ+LT+CYfqke
2Vm32nnw5Sh+S+N6zbtOjaawDUlXRfrzqrzwufstnDSBZOzfeEUy2D5pBzgsvUbw
DV9IWgE6RgrM4OsGwgzOVTbpEwp8MWfJXMQEk87K7TUi/BVR4P7K4+YdoQLf7cb9
nealZ3BvL5DFMbu1FeVZ794tZ33VpOSNk+BExPKhItnOU1npTXlziGwcnndET5FG
nwYsCcBx8M/hFIQZa9VviSzAij6HXuMqDEXjAPhPnNmeRuKriBRWkZZeEmD3bjHr
Xasuz/vjh2gQ6Zho3Rao7Tyqr3dgFrYBWlJlP/Ty5oID2fWPnQM534x14B5HurNe
45wUDq/QF0IJYu276WIab8ZhKYb2GJL1qzdFBU7KTsbzO9GOZDxiKjfOMXk+0+75
wZZnYuybKF1qHO0z20VHL2MrmDX+J0BRaw34MUZk4E+i70L8jtWJG9HdaFrhUC+I
yiybTkEortZwbi2vvDfzsYIcZQf7CZeAR0G1mMshtjx1thBvlWXBpuUOyyQ1PLpe
Hb1AUpcL77g5pDfGI8mpS/+0FrGBJ+h+Hc5HG0NMVqOV9MvaxHehQiyHRCZwPi41
FjkjkdivDdBw6vaUjXQqCrr10hKGXl9u/oJheDDAG+qY+7alk+rm6MvpcJbcrUYx
VmNmIlyI9k2PBj6EzsTFDwYrN1/iueW2IBzXTBNloEcxTn6QKgfDljPMal0KDXHK
sX2j0EvmmeihAeVn5RGKyMxJZ4PWSBG2P8gREUosqmWsOrOi5l63+a7G00qZ682o
0IilsthDahHutUGHX6jv15QqJsm0Ml1MwkUVP02C5Vyr456LDDwLHLgoHFLmEVu2
CVj5OmiJT8FQxfuwPjLBWbuxWuXHX4CQlDEFH+MYlrzJZffGz8801eWg7pNLjsEq
ZlldbirJuBdlDUDQLk3Ffa82or/M2lluIQ/Iny+QMRdR+Jd8Hp/LLycQzjL83SmA
bQdoe/n2DaateIpU4Dg9IffowY+5hVxMBfQdbh7l5YcT/KGTZgO5wM3vI2PKtXba
MGDGO85KIx31JyqFXxZuqDa/fDi5z0SYx04ktYX5dVepCu4bmh7DGp7v/dnaCLgh
GfJG3zdWlZ0DZz328Vjl9ZqUrg4Ug+XyQ1gfVEnizmuc4F0lwKxen1SfLcnisDeZ
U6fkl/wg9NfO6x7XcYk1YHTlLq47YRhShicgYam3s0Ldpc4bD+fF5kYJb5JpkANz
QwY7LpFNcU/SHBiwKkrU1II1TsJmvKB40B7Q0tvCKXAQYggnnrSVl/VECz+HoDU3
cEMCTzQ5S9GovyHLwj4xi400ySCZaADJN7obG5sEXSNFt/A2h6ddmigBf5dGdf0E
6mgFvUNfiqIf2vGC2cRjMt0yv16fVhJ3Xu0bjHrqDCAsUlOSxOq3oEDe94cerL7+
n94wPNDa6Qr3yrdY2H25BjDmydb5EHVfScJy1at6iVHfjS+U/UOHFH1pfGHkUufi
xIsasKdaAO4Gp84ZOi5BtLeBexO6w+RZdy3XYEQYFbPTigkVkAcC0kFJfgxqlgWR
Ptfc6J9MmkwQmCH9StxjV2FNXH+9Y6OB4IyhHxVl62bBtFUcKPLiN8i2cW8JvK06
bO3xlY+eDgeEIg48JZZr5qeAzS/GEQgQf1jhUWv4PWf/lknUcMvrkSp7Hgvft8f7
/at5Gw5T2RSbux5O9U76xlp7cp+XMwfYkIIlLDiPhaUDkCNrlKYIEPBG2TWf0zyd
OIE3RE+LTJj6ybh8owGlc4V0NiG6ELT4Cj8yAi+DjmGOxrnQyvG3BmE/g5p9jJuR
NXX2tSGWB02uIa5bbrljlwrngwRiLGbDCvObPy22/nRaS5IIPnwVfGEjkayJVPV1
fRj8P0QQORCYH0cytyDcPcE6/pG+zAriny5Gc4zIXmXw33h3vK/4hapOqvaTc2HL
OkCah9m9jQ0Acxn+0oIN6LyVgJ3aE0/2ChG9lbWyKqDG9BtaKm4GoQzuoxQmC+DX
5bJc6Ta6Rsjad6G/qp7gqDIMlSZfVLgviHMowEdkXWUR+BAtWbkEJqF3L7kTgtHr
Tz5G+w06mntyFOZo5Nlozjel77ud1YaqKN7np9EjjIYyZaihgRsFIPfbnlpfGnLv
qv83XTWsCeGkQ0u9bwrGAIgX4pU5lO22rIjpoJ642/X7bWeHvUzuOPm65Topqfxc
t+/W/dcoopjmCQhtPxSlyzV6X5r5kFOYRpX/ynzatvHYRVF48yHvABSc4Tes+ivg
xbr4peTBh1NXsxPzAdS0354cxKIuUX5zyTlBKqTyKuNWymQ9Vlb0Z7Xl4e5GcEvI
6LgjEwUrnvnQSfyvJjPMRR01bn4Qq5A389EP7zVM/5HNKq9QEzUTJyJS6misEug3
gq/k0FH213icN6m91AIMYJ5Lr1NVEjGUMhZp2BilUeoo6LnJaW1M5NAwhC+QEynY
mnyF8MmgK+VYmImf4qmPVT6o0HzFOQrYslzTdAxCk8m2YGfoeFWtj7f8x1J2unlC
486+R3bJukNsK1TbGmm03BWmCiKNG8ZgyMI0Z058UFB4SUvNr8E8Og42VUpEsdRi
V6gNwSmuRlFh30UQRgpAWGOgPYlQe9nmX2ThCbx1ewsdR0L/NXE2duPhIpF2Y7Ec
pYofhQlNNEkVzTNxqklGFafhA7uPlSHGlI2MTGCqUrNNa1L+8ACDwEth1vo/B24Y
sgYDz1Sfwtz4FTy/jUtgrut0B/xWl5fseHiGt97VGENQeBmHrAsNsBcgsuHiUelh
v+y9H2wCMYclVKP3jal+ULXoF1T6JPJIBpZvM4+6TZ1DTMUKvYKwNL3srbCKfe6r
wbApHkQUllEl8cFPHtrul2EPo/xQVY3Wvld+FISdXrtpLaMxQtBNzoEl4SR+PJ8p
xzYNFOLmWIK25uJfo5drjKhGAg0ZaYJ5S6ObNzJuvH+od+RS8LBympdq6/1IXBXP
U1oiLjdI0ingiglL0gm5HsFiSY+vcwUb8AEDSMx905xo1f0w/6V9ZacHHdkj46gy
3LA7rgsuNX/gGA0XMLFdUVD51IAD9pnW4uyIfRoyBaV1hCvFI9RyEMYLIIUB0s7M
u1S2+l9GJ+8uBKsJd1z079jw7xCROtUfdixQvCWQyBUx98QY40hWKj2Z7bSiZDtz
USQiM8oLFEN+jAPo5HfiVWW8ee/lmLKUZfSjHsBD3gHZzf1jg0RXsALvNcBPW6sU
c1Q+nW9AUaREeku3QCu/RiGJ1BL6MfG87BDtqQAL69pE9xOzpw6mbp3ZNBiTMocF
hUx1FVsMbF9F0m5uNKCsqlGUWfhu3lLPyCF2uTn6Fw1b5ukeCCIY+tr4L3lBos2O
oa/ZRHP3RJlp+CpNbkOjF0+W38NOaHmSSPeM07FHcrZM6KdCvPVXnx6XfrqE/wLe
RKs7YzGzbtOOUPo4tRBYrylvHFOkieiTwii467sfV21oTsjTN1EHX5MT8NeCQpBk
DbWuECs+a5NDlmyc0XqBJP+lu2BFNCCfAuCHvjnOVLQXahIw12OtDORE8W7O6Qgt
qH1RLKIJfMEdcBPJCdT5xUMVuhOr06I9ozt8eXLqgljHanc+LiWZTj9OW21pWOKC
jjhKC+8vBUAyXnT0MDMhoCnOcKUVwjngzQDZVIBJ59N19Pr4H9NMy2EFOQ4EoDkm
s8LvVBiCFVsdXLFA+8W9nFXEc9UK/cXq57NtginsHYI2vZBevzI0Os2JzsSPLI1t
rpevn0T2XAlHNYhpETWEVgsshCVYLVuZgLUjX49P1lz2gZXq3bf6W4TEFKtDM/WB
ROpbYJMM+w45+B3Zgiw0bShLib/qCswBcxSklhEiGBFyOEvxsBXHO0WO2VcGwUaG
s5JJ8B3C9+MHtCP/Rvgp3wmQxiltD/Z3PqkycLvUih+Vnpe09bRIekzSZ2CPOy2U
hDFYp30ONqZnzUHNqt0bWOqUM6CuF+A2KiFt2Ff1k/JUZEBClTk2CqdN/itSMpVm
ekUSZgvGVUOmMSC2pI+Hccmia/UC+lVRR4/WYULcRMOX21tJdGRRpp8szmyIiNwR
J1rsK3fQ/s5AzdcqaEYx7JJlAQlY9O4mVaoyOQW/v6vDE+B9/sh1qrf2/wdR5pjW
/twCwCIHZpJzyrNrQzMxg36h4ZHMkQ1nnDARk5q7AK5H/OKiD3c4Y1noLYwMp81w
vRZ0FykaGDYACI394fHBQrjgJkd9jyTCz62xE61wyclGKWDTon6QBgI6W4w3Gw0B
4lL/3a9pJMZj2WkhFn9CHCtvL1B4CLpMzBqkWDryTSnM5cT5eyLi1EPnHrc5Ba9J
4cVNzco6QE3Q3FoY82bq6Iy2mKDYY8T7l5EwMJ3F9qy9woWZtzFxCPx3tY/qWhb6
1w2y8VScJg54GrNJ57X6lEy0BnbgmuF1kN7dRssExwhfpzc8pBhzk6dFE4VDYUpR
ApBwoFhT5PcqLfoJooa2+ECrt1gpCao2eyiD676ve6TE+Oo7+ZCxpiSMbz5hSeHf
cJRFTx1UZ7edyCGepfB4kB51vpmbLSqpVFazVDyx8CDV5mYDGccdq+t1rE5k0YIn
XwvXjjb8xyPu4fxub0T92HMAvo6TnZbe4o6tARFgew7NlcremEi61Siw0Ou5i1Nf
QDAaWIXYTqjktgubKY+368sWYV/ksSmIVctNjJWIdw74/KLE7ivbQN+YMuuRsrZO
MBTLoAJopWCmYo8oIuqlrSPxYx5p7Cpor22H9RHOoKw7GAwK3v2FaNH18ucSofFT
RZHzmpi8qgWmk03PUhZmJD6Q+B5dvR4H36VdFch/q4YbDl/W0k2vdnxXZ1NMp/B2
MNaCOwYNH+eV9a/RqEQZNmLu5mh87ozwHd5OUVit6aCs/XAsh5ze1VXrqGf7LLMP
oZhgeeG+OngGcULdgVwlm4S5BnRgeJkZErxFlkcdHyHxniBlfjTA7TmxSKG5NlJg
pin0tu75b6EZ2eMrZIMIq9TexSXInTKE/krLYDXitq0zGJZ3a8ZDkn/Sz+dZZ6k/
mXFhtu3xDUi/GN59brEjChuyric/0cpd95mhLCoMzqqajwN7nA1Mn9LCYz3jdWrD
x+593X1J+t5h7ziVDlaDx2hQ6Esh9ZHWD026oiwNPOy7GqpDpCXaXaEej1nr843q
YzI5yxenHCS8sFnnVuq7dRJwe/518QWHecLYWCIv2KB4U9njy52F6B5xEuctkQQj
3/1V5/rK2ocQ7epDWj6Xcgk5QqZ0Cfl9sBwN144OEDxnjG2Q4mg54z60MAto19xs
7tGnKwHK+Xg0nReKB07ln9welNS4H+p6AtTZqSuJCuNFBLyFgbhtGEbN0aRczTtC
/NCLijypDfBpEj0HILs0Mo3bIG0iLnYdyQem9PAmbPb7vk8t0znY4IrnhaWL3oMu
AVRfOePg/PHyWgdta6BuoLK0dqUC0hp2nOoBtszCOWlt0vlTyhL0v0mnK1fKfYy7
TYl937iH6GmRAyvarzkll40j01D9KvUOWCkseP761yGqNDHO50ZXuJcJnnUPDqL+
v4Bsc66jKoHLxa6H0h56aZoKko3N4kwgsGyJQHXoj0uLY8QJJrFpsOIVHUSHxFSO
bLW5SDMX9GZLJo/CdHqNwFdnBwzo9uMSgDK0JMwq/OD7XwwWC56q90kQptbeoy8i
qXcRtq0w8PMA+HcdJQwq2o2HDoFCjcl/PwqCEHvADJz65L+sDKwAkYjOKVHmmOpz
D568txQTw2GNZYtQEXiENuV3L5xMV5ps8adIK/MgNWbBX0huneVuvgLRexZxR/Bl
csk3Uk+PGoHwhaCi7VsgW1ngbj/uZY/aE/tkfNANcNdmeGwT1+0NFlMXzQW6c00i
xUSEOnPuC4JQbNH04YKlGwcWg+ZLSM1q3YCQRTf676lac/veHmI2jLc/vUf7fiME
CRotUfiq2AG0HfUiG5Tu/MTQfWqLq9J8GtRTgbv+EfFGu9pgufSHKvJbF80pu0Ga
gqtJCmzIVFjKJWg0WgYUEiLMCr1dfOs/Ifmx3Nr2ASbHvbQNraE6m0NWUccodZYI
mt44J1EmwYkua2q7n2EP4pFeQSpHLf7sRq3Cva6WaNhdJlOvBG/9t6hhlbeWbabT
Nyyl4X4cSCxLFI/Bym//WUsXbYDb8HzbHvxmyr0fthby11BENXXW8LIl/dCHret9
OXC/lVtCUSoANoFiNhwxrwb97jBJOqRWG5HtPVvxQIkymKCqPTijdaak6qnv4Mi1
u+LsMsYZ4MHeIEA4deiJwGdqAjE1tpOWtHH/QOflHIr1pctfM/2fNKXA+fnMP++/
H0XyzOq9i+k5tQh81sYTPoUvMi+VpKfH04GPYXhKoP8HpbsOkwShv7i4D0vsuol/
Iyh9aFRER5AFCypLk3GpVGlZ8+wwKSnF+ed1gdhyVD4yE4DcPegW0LKK185oUtvd
+eW59lN02AnMVCvsCBfZC7l7RPUgkMoOIhnOM9OcTaEAONBFQjzJlhApx5igwy53
e/PnddDzrjg6i19FpH6wgAU9u4VZ9PNA/tjgHihd6LkHxoudwB8YnEpwuTDImgx1
cPjpiLmSW2Ua7ESDOZXS/WjSAusyJM29Da98SiX4+eM0/e7rOYPt4uCUOuyR9rPE
pSlNRQ3KVUhXlWGqGfgUvHydHOeXdl8L0k+5IFcm4IFicQ3Ulk19YjR5xV03SziH
J8LPqBGuVUxzy9ysiNACBLDiXE1zQi09Z3zVh2rJNRbECqSzYa/R2Nax/vPhQvnE
ocvQGpWic6yr9WmQLqwiaC3Kfao2js/9S3bMUYgd1LceN/QBRVrseAyFK+GHySM2
b8e4lqfBk4XkInn9Mho4zwgmKEPmdgQHremGk0B122h+A+PqNcA+aveIHPjXjbja
IPAwswiK0gLqICt7Mk31tKVXPwEJ0Lo5ktl2WoeyJlxrdmxbayXGsMpoFimyP8Jo
KdGgeDLIAef8uuTv1EmnGlxwdWf2ATLSzDLjlOKXUTNpoX7zVIQJUBM8qKFvCIzf
ss1PIRBztRHRNbwc8By5GGqk77t+L9H0LX175NctbEmERoihq0kmMjqrTNQ2Z8Gm
DS13r868uHR+q7xrk5OiTQ+wU/ihIqYaKm6PmPi3HVrXr+7BBC3RFg1oz4eXL6sX
E/5Bph+PvEiorq1W+IxAPjeoYplcLWbmXemWHyzV9mQPqGrTFaXle77IzN2N1F8U
cjibu5WGMPGgv3bJ8pWYr6wkGD0cxsngJBHoMHT7OZchXuRpP//3KT43W/IMQZ5o
4pel9WzUwyE4RlkSO9Nsp+7WQMj0TjJXKgyaoNLaW5hkFWofdx2GfkKzFZ6muauI
wFzPFTnjPGqOdDI/ce2wqrauxENhWTf+/qZXGwSM68t7+yyWXWs6FWImFIacACka
5kKItS/xQwyrQBhUixEtjaIoii7n5OLFBADRCQ1A6e+2rEzoA4VwXunAr/hCzjmc
Y+AaCOD5fRyX2MYVkF8D7s6AC1lotv1+QuHt58t1JpiP0gcpoI0VPWM0M1Yz8MW4
JhwAowPts3c/gtcT2crgFMgQmVnPReoMBqEO3kNXvEk0jaeNWoVZDSUPjuOR4yyj
3pdiLhiK3cvS1daDZ6keTtikHX7j3iiqJ5Y36+9p8Hzjun+tEn0g0IWiRjXnLhwq
VEwxlp/jkrYynRWFG6psig/n011vP5q2ZplKLdpHkKo77r7WkfwHmw9XJwwqyViU
5D2As2gCKil6mc9jkUOK56UkSEidXErEOpVehWMifYMSo7GjsFdvD5jUrKKDeHP4
HTkB+SE34oZ2OpckvDTd9TR3clnskUsABX8skZ5UX83gBYhHhLemsfcboD+plU/T
fP1WmKtzDbnhap79hr96O+rIV5fME2kGmwB/daojd8U=
`pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Nhoy/YNMxvp1EdJkZV1IRqZDSVZbcT5rTJ3VUe97zKfXPKsxhisPr1VmlTPDCmrT
EM5rvTY1SDcAD6UeHF/Fvn7U9N4iHj4cVFnouMq/+1PN18/sF7iNqqfD9TS0g/ib
HNTTNIWBWYFFANXkKFTKdVsGpPuwi71t19FvfChm+UE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 36816)
JWuWJ6l/t/KI/47G1xIem4KzPZhtVgsrtOkZQ0bCVchXJuTE9zmw+saAnDd0JIej
Q/Xwi8RkHiydQV1Qj7/Gvas6viKuQtCfDJs3BdHzYksi43CLiu4NvVHHSpRrMiVJ
9XdBiYibEJodhs1iCuOfCK1SKLZTAxaWl9h0IylQOSY9CJqduEORkAdrRgrJH0FT
lfQ3Dyx5sizf+7oJJxyG6YOpXz2R4Ja2gDPT5iGH++BF2+O1gijSwDrbWj9fiLvg
dZK76dGaVqd39SbnptEo41Tt0IwXyJ57QJ3NBQ91rCSM4FUinHKbkFb25ZSs+WGv
kVN/do1KfNr4e9ZHUM1FL2fp/5/v/haS6OiWEKOru3GygcIZUgbSU/7jqEJl72Yc
opTol91ZbH0vAikz8MzU08AbVSCUzVw0TbPLQO6rq48QDfoIEPiLMzdb3N4a40nU
Rd7+Tu6TOSmIRaUh9Zb/dhmh0e0hVJtA8YJye5MJ/uV9U/HYOJUy4FEZqHf7G9Jl
k/DXZ4n7kZ7vuztIJxXct3EfZPa7bd14jge7O9XYi1+c0AUTNxG8DgjHX2u6+rhO
MFDbHKyrVYZ4z0litE9iHS4ggR5EiO0cOONENHln0D82/IDJy09Ctztf7qrWphcP
bJLLmpO2h2ayCNl6IVGNnqrYJItEwMAQNNCMqB3xZYOS+tgpHXfdw23ln+5lJP7+
7rOCTBmn9nMg68sscjcrhIkjEHn4wcDOhNEJQS0NqB46dZn7OqoA4M/+EMQoi0Xy
kmuWEVJExM5uQYABTqPp8QrzkB2t0cZe3RyC6rw4rJ74hK+NdRUkASvFuNSe084H
/2gOMnWeyEC0GG+yEnNMu642W5IFu9UrWRP8hDekHdgJGh8byKWs5skTyol75/5j
62dnKrmRHN+TsPUqJjHKVLsRjq1yurYpf63SaL2ZyCriVOEOLYj9EnXMIe0GzQKW
Dwx6yDUxDpHZG8CORtlvjDmqELHG1KM4ouQ14+maCLDuOk75NNtJa8bnIm4zaKVz
YthMeavHDmm14t4z9rO5D4h0UWZSWyE9wMYvexo56Z7NJdm3fJ7ST/QGElkJicnY
pc2xK9os29yzN/W175bHz/m/HJB03yyhXN5aMOX/iU6EWaxUtcHp1AdqZ90MPg98
bnP8tbL+oVBSXoIKBEZwcWCZlxX/XcuaBKKxyZWoB0N0PwxpSxaFFCFuNYP/1jSQ
ot7haT7TpaiW7qeXONl2DDEyAQw/xUV+yOjwnjpbNLpso8+Alu5BGwge4F4KaZ2u
7eLxdCiWf5h8nO5+55S18Hyhw7si9IylS0Gk081zBPRL8yM+UpcnwPbek0xNbqMp
+vv9glth7A5jd3k2blLVOV2B8vb9i8jZ3GWPpC0uKedrGfRy1Qb3la38uiMWX1Wf
G+vrDzLwciv1/hoMrxHwC/4nY1shGEj5kJ2SeYwYh/Y3M4AKGN2pU/uPoAXyYOFx
OL/1WgtMZzY2RrP1VGozeuQ+/ZXoyw1tF7XulU4v4buwd+SzWcwS1D38e8Jj/cKl
bFsu2MGSYrNtM761P7PQBfialPNxoSRjJpBza/R/Gk6aTZ4JqZumdLahTCmQoUR+
cfZdij8Akn2qlK7hIHCbwBnPVy+Hm5X3o9LDcA8+b3H2hvQpGKkhAFlcplY6Nvam
3aJm81/rApSzXlpZd4Uk3FGgyibAsHkSmYLg6EhrA47qwtLQoY/YvHK4+TpkAnn/
e5zxzb8FlkAVVwvjQRpK6Rkm5L1IbnVmCW/L1IvQSXegvZCF82LuQuzeG72MNq9B
vGi5yg1TC7ocWk/5fPVa+8YH+UQ8uYuOaCPviSDig9FVn8q56f826wcG/SN0hY/d
Vcu2zbeDuzDWkddMv6imq+6YjuT5bW1G3Npmnd2IdvwEMErIlaNl5A3aVFneOgBP
ex85U1bDN2DpXUlV+fzox7enEmiJ3xKYKpdWb/H1dxFBGNGHFzJEpoB8K4YFhsOG
sn1EiAbKs4n+6iaTaDxOKJF4sFSjBTPdPezzTzknQBpz9XniwGSKrmjhtkR9qlm6
d2NqiPbBimZj1gRKe/jE85KSF9xfjhp35KW+j3Jg/1oz7JghEVdZfQbnuIFmn0Pz
2Mk+w80ZY7V4S1YWQpkBLUv15HImSls3aJMJhdH0H8QIqtc17csjb2khtU2oYAQ9
FjdT/QUsQ7nhNESeH9TVBxikSTESCq/M4VNoidqBeQqFlKa8L4ygOpM5uf7D+GXj
oHdwaP+npPQHxkldSkZQOiUP7HiC+ChmFqeUv7sNdjGabOoEXKlu/2Wva0q3sLHx
Ervb8EwGi2lng/WXnU08U8hN+wSSpClS8M8ciPjZFKngTyGwAPavNpy2Slzgx73v
fGaKJJ69uggfCQmzPCvURseOcjB38wf9dvTdbcc06kRjC1HCTASpem+DGNU5El+Q
p8P88t1IpDoU2pPNJBBAikbsGcNqKai4sSNT0xmNOiSIWJVRP66ZaGpJGTfyySFZ
/OwQbL/OJWjozXhfvx2S3GshBOFvmfOD9N9nQDYomFXQfvbBDNSDkmmyzcfjSnRl
DuJVyEUth98snNRYP3VSqYMe17HkWIo3mMgT449UP8vEs9ha+fDynMboJgrZGLwV
qRMFPayZGMnM/4wByhdoW5Q5Y2UXO+gHXFV6Sj0Zu4FUqZDvXNYWBYo3rkcjjaUK
3H24ujDGoiLeiUz5hSzBFl02nqmR/vr4gzyfizkaNSmre1j36Q5FzKbTlECxgW/u
Vmvi6Fm4x5ARk/iFM5ClCvLEUnDG3x5CK1ZEdFcD74byMs3YYoESDie+TIECsZYU
letLVpYMN1lbNxFKMAf05TOVuPgpn8skhumnPmW0LjIG5oNNQcPocZ3Pl+vus/l8
SxwxrxbCMdI1TrbAbdUO3w4RCGpxjJvxpVqOOMMMs+qY8WENTMhZMsYX4slBpF/j
O8len9aPdinAMHOPfT1cr+wBALszfyR7dDsXtGvcSPMvXlLp4zU6P7wMtMP4Iddu
sFNjBzMSsJuKIvcYdkkfYEZD4jiZNIVAotgqZjO9FdwhFbah6fF+YEJodBkS62dA
nOohFGeO+KiczMYP1KSIO7RhOMXmAzpHz71XPKDgr0FhmmTTpOn2GF+bHVGXjOOS
/hI37lfXupyJL2PCRX49QZvy7OvmJ/HcjCOj0/AIOa/u3ltGMfLRYvc+HnjMaO1H
605pQnaxe5jEAGx/B2qQg0MNOp14HThaRrbgF3GBm+hcQna4HmFVFqWUay2H7bus
eKfSkC0xP5MWmScJT8dv+HEiLoj7j+I75t1hYvP8Mno1ai1MstK0W7ThPafCJv7k
P+03ncpJDhmYeYR5hnVm1l5h9fEFrWkoFCD8epOaavikBbVxwA71o4m+97gqfVYj
rwbZqgHgYivpL+jhvAx1IbwH6qcoDFYKhrXJMsh85mcdtFacPe7FcwLAX9McbGNy
RxV7Rd0Plr2MrXar0X52zqPfN1/Qvcc0NgnJaL0Eb+Sbw+4jIbnPMuJyB4H9mfZk
9tl6bY2Ecs97zmB0e8Rxnqiag9eO9scN/nAR1N8RcaJUVMy11LVLthPijmnOZGxi
zmFy66IFueS27q9p2WEv/TLYURvhgZ70yMV3xCv8+EA8HjYOsJ2vacheHhTdxy63
beCSUvU419BNEq1uMhL4HQlQCPVDwgJT1NhpOaTCJNOw4qK1KgltQGq04SzEDtBB
VSf/ZRZFOswqum5331r3sL8bSa810Czn3wjOTP4nUuaAuKnT+g4EHrCp+PFxSaFx
w5rx675aSFHZA6qpfe/OulCY5WLRBn9Jd86OSy4qoCv510entBkEhYxqCbZaxtYM
Lnws7CvJPvZGEMV9LntMHtyctlaBvFjmn/Ite7LZVjgyG/mlKHQ2g0Bs2UWbQA/F
7euJMqQRhZ4GJIbcKRPKl2FxK0KZXorhlwo4gq2pBqDslRE+AEu5l2UVW44RYz21
qKITEns39Iiz9JtdgyCSExgxvdoj2ZzUmaLUfJMUEnKQNcX6LbEVgavlqYDoBp+e
D7MUKEhIvIZMUwu61ozk27y1Kd0Cz8fWo32i81D2CCqqGfjrz84lYLyrza7eoTYN
6zknxSWaXe8dfCjUbv7NJvQMfkGJC7ZonreFvlTYEkRUqVAVrZz6dq3iiUEuehNU
bzf4eG6i+IAXq8VI+Ft7fQBEg0sZTSZHJGw1Tv8Q/363otTBqM4RT/a76k6PwFQg
qPis/R5HpThWaFHsx1OsbZdIEst1oSVEXH5DAEDXsCNlsRIyHo/VXVG6RbriZlhI
UetZHvDeWIwC8IkbH03vp8wVLBCiF6bNcuwjvDIzDk/EVAAj0xUUqRL+7qigL9mu
W/1a5sylPBg67osdSB8ZvHshkF+a+2SBDzY9YUIopCKGAtu02ctEFqZLsaMZxvVe
4AHEQw2IWUjL9ATsMhlosbpGi17PwP4SEvJPEk8kxszQ4KJiySOcB7ggT3u2APxj
d1DwcdBPS8lCnSE+HYxYM6JOzgrnQYjFzYMhw/+mz894jc2/dHjEjChpDB9rN8rW
OnQVoRxWoI2OSVXv2rfQrn6sroQefq2B8NqjzBStBgR5cf06x1Bqq54zyigPSjOJ
P8zT2CQHDZfUbnQWU2ymyijnwyvl6siVyMfFWkGcc5RpDPc1xdRdluv/a1jK0OfS
yN7qb7B2+j4tljEZ2Eqg5v7aBXb1VhyaZvYK+Nw7spoHypaQT9puWVoS6T4TltkW
zXqk5qA1U/CZTm2snmi8AXy7htwhcVdz670efM90ZW9fcA4CqJmLuLZIZ62QoWEn
AKPip/Uhn//trICWkx0YNQk2xz6gyvqVHSQ+scZGkg+OvTUFRe2vv4YgB43Vzg7a
OXbBXVy+A5/hOLMxXpByboLyGV2oJv2Jtlflr1Gbr2eJaFm6Hu1Yl+y0Jyv+WcYC
dpFqTGDBwZsKB1qI2CgAG2wPNZInhppZEPp2/PT4H5cS76dS088K3wlZ4cAq04nz
l7dTyi1L9tFikspCKBk/z9mb9FcAGjVHppJf5i+ts3DI7KTa7jWeNdreB+Ejmbi2
5TfoAXLHZxigPw01JHxk494IOjU3QaeZHAf7u0IumcpYk80qtDDZu9f2jGEuBk46
qmoXtGIJfmOlScwoqHOSYp+2vKpBiYuMd7ZfbGplrDmPSBOJoMY8vbLfoptJAuHA
Cha8mMaDIxo4AyOhmskiizWA5xwCtbJj8ruabnTHpddxhf4doMkcnblPXJzXT8v9
cxQ+Pk8pijkp2wkBzTTIU7F716Zqbu+gHIYeCs2V9oGCnx6Xd8Jzzwx1uBaWeI+z
WLsNIyUT4WRO90zdlC2zPSbT8M87fl3jLW6EmWDg6oHiU51qa5i/ov4aQm2L9k7l
PT+Z4mPec2d5An7DAcwUpIu+iv4pKo8s/pR0nRtydLou9bPhkenK++PZtNktSByx
eGK6RKXn+rdTAQLfIVogGPzS57kHQXgBmsy+bwwu31tIg6eOFM/Tkj2mo4IMGM0D
ZzlvLBktrG6XdTe5axRRR7mPkKu9Drsy7GIiq2rbI8hCnUru7HaxQNu6g0DVSwbk
kYT8eUChxbd6fZUadz2w3thq+978RqKnCzujDTE9RCScp7It5Mr9UWbbKiNim8t8
j7kV1teJ7nSQgxXPeqA9vjX2x42Bw6Itj2pe3hOtyjK6yzJEUxq03FbQ09yOfhPn
FUg1Ux7q0oHvYRfAht39iiszhSYbcIf2cu01S5wspNPkBpmjts4OiXzVWc/33wwI
2QuIHrZOH0ywZERajVLWfF3W7mtLcPuq7Ian1WJgQJ7Eb+uMjxFeUdoXOePV7K2F
Cm0acpKx8C7c9Q5Y0zMAFWcbKfSYLcUqNnpIQcvBg2mO1PkfPm7t19FY7Q8HP8K6
aSiuMdvBVqyKv3+9BH8HeQwEcQS+KfXzq1nXIm/FTy1S2J2Imf3zP4+rkU9+Vj6W
LLo4nHYItiTiAcqt64uBjOkhYQZAHKhOLzX030F9xIyl/WftcCP0/kyIcZTcQzQq
lMlcAC57+5PEs3y9D8xOUKF0BWAXXFAAci9IoqyJzNWNNzi1artTgHnXTQuZy3/s
Z753ImdsGCf17lL04Kky30ux1+pt+xHZAvNKK2ndvMLFXtCEZ848wnKcs89GmyDh
61LGDWlEuSEryAYm7dre1c0n+5Vubjl5HcY1JJPzHr4FaBzmnWWtSyzb4m0HWWnP
CMsg9lF4HrEJDW66rt4xHWPSIX0b90oA1DwbQKlP0g5nGsnXZtyPItMUeAh47sEs
cVmUx/3qZ1TgtdNzstwqVJkmjGmBieCPjPEvnFCAsGFNOtACM5UswyPB12Rdsd6Y
DN01RcmsFaeguWXZ5qkEM2xmsNwYUy2EHvx4PHi9NCQFKsvBcFkP+/uht+SWpohu
6Dmf1LU1OkBtd83EsPK+WvC8Xi0CaZZw5O5jrUf2solK1imntckzZTxHfZSatc/i
dNs2KKKmvK8ANAApbLjD7ZtbRC79/+FRjyUIO1IAg6+dBeNhdeBs7VrfV16NaHi3
VeGqJN6nW+wcbfOTaGwwCTV1rHNgWeCtQ8kg1gOSJt/fjemp4Y4sOpRqWTRwfc7C
FmKhX6kvHH89HZp7Ic2ZSWIH2pQByC22Ekf8X75nZGJH3K8u4WdsIQsWDeabzDkU
ZKGmzBMFvPpok+oky8lAgWbLDeUnXW4+/6vfH3rKwjQNwkYW8wtpRRSb6iHuW565
MCqTEXIGdFPIIpJ3kG3YYffTjYrtXCh3tIi6/D/Pad1e8DH5AOodTWSElgf+a435
943t4JTrQ6HtkW1KE8FwoQpxNyjWLMuZQKPlIQTaGzo3YeDTrcu1y595k6ddOjLO
YX4m7l8m/c491ZJgSev/xr7mqSbjy8m+fe1uU55ZDAYOkr+m474rbaEWF8a4zkMm
EsAVHIDQYwj6h3Ytbz63ICN+PwhaBiCXg/4660JJt0dobaJ7gOMwYJI5FYQyTRoa
UaIKt+hPsRKmV8uYOU4Ui7RpA8dtamjHrWCAI6QvRz43u20t1oaESRBFuf9N7Dih
10w1MaMMr9sBVo0/I1aManIJqLxUQYPJnKWgQUbrC4aee+StgRFljHVmykcHs8GM
YOD6WRg+BQfDYFX7HXqDxD6hjfHD65kcrbpbwV9dDWo5va7qA+4SfuRAKGTaXqZv
2z2mbzJslOmCo5taEltU6oOFbquPka8gG5EO3e/18fXjq96eHiuzKFlRgYqwoPXV
CruG7zWR8BvhjDpFqPS9LDUyXXqkaWDtYPEbXRRgONopfq/ySd7RtZp7Ex3eeMdd
TcNCtp5FX9nwjniaiX6R6MHG61PsfeQNj0335mVGJkdC9fkFEnjjO5eA2+PtjiWl
jIkYPtYaSPiWBtmYsVqOPivEqvSB6YkrCSJQsfssH/TtIV1+o0wNS5QpaHv/fvC1
u1cNEpc7eCdWMrEU3Cef7RPgV3B0tQmYxj1mnrnIPAZYVBUMcTVN/eeaU2IzyVfr
Sd2COznT1N0ynhEbi+elk+c7RlEVVQJ4RpkDmXP6JLvDb1Hkqn0yIjgHfZkD6ETD
DiRJeMxyYMwYdMTeWg7LW3WZ+4YA95nBhQ7WwQKaZss8vzXclzKJHlYu9sQYD5UF
6Z0i0v77dwZuOG+KdoKMpt07DWrMJ5DvbnFEgBx3epykXF7tSeV7Wc+tDYvqSSA/
c1wcWyR999B/mS+hLuwI81UGLi0dMGFnNts8TY4yP8daLtHw+Q2vb6ETFLEyHZtf
M/IAfUdbryI1cCAVbezY2cQfrOOT2pvXOyt3gAwm1OALoSPgmqgk6TPqRoENZCJS
dTGVxuCXSXe5v4jqOUGgJWT83jcSDOcaehBTO9ScmQ1vOFouMjwojbkH7wLEajeA
yoAiKlirv8/trzbGuzHDQOxpTZax7e91mHYYEgKg1u6xD7CohRfkeEy8EKfZRmbB
abYHLAW0hI9/KobnDVwUuDzzGgxZ08UazEyMu5YuBFHwvdDdDNtKKOZsd2OTzfeA
Cf2VB+9gKM8XdtV72aR+gZnP602/9HcUFHADA/A/NqcIO70GTrnGC7ySMEc4speE
+2k4Y1OtBJpinPhKT8q56eO+nd6bOP507EbUdw8BNBOvWyWuTNCJbVDVOInuNC4G
74Cwry7DlZgCGyAhGDXb3KOWRWPXc/e6JydLB8SgrjJyK8XLGe5fR4NQXfUdKZAk
4Juf8wUklkkKAijy83RjUbpiiQGA7GM6Tn466AWQPsUlnRZCbhk3t2bHGVs33TU3
Rkkxc+GAxgfA3OP4q+ZrR+ZPfuhfWJP+E1dVd4M/U96/TZ7y+KSpKphQ0ECb0aIm
848M6OOVIPboG2tGzDJLcsWc8A8EJ21qkks7CQiY31sfKmKrN496cRdiDo6kJBHJ
r4PB0cml1NX+HjYmEFoJ9/hh0ZQmHMzc02eq6ByGSF9lRtIXjPHQqtQwzwKL2fvR
iZoh24GyjGehUq7QkWlXimfQ9uVPcgPTJeXryzrPTXyVpY3qQD07JG2TrHet0Vku
11dFEmC+xSor9ZMNEUb3bmHd/dqW4WcVNhc0el7Fnc76/doN4qMD0QAYFRYJyy+0
/uZUNqGPOkg+52WCRMjpXf6Q1d1DmVVOIo/KyqNTvIOP7ttyxvwSCmroBqIzuoPC
DrVAemweVa6Ytwmp5IcBEWRs8SQG+8FHOA2QFwYQI1iwdJTPB/AcKkDfKUSTAyon
P7VGCDtMp+SrAujqXdDUzLjVQYzYMmS7laqsueG+gXaDvTaHQpk++qzpYMbbD6YL
7N4rdCudc15sZTmFRAIb8eedgRR0WRudWhfnVFTO+FxD6ALKhrnPHIIEfm+ax9rB
BYdZUE1pqbIRJ/qDqx2Gl00SM4Y2lZpm3a8ae9zGK6o4gZDHfH7yrYZJXtDk9OJr
6gSokqmA/pBIfxxm2eAvC/SNNI8OJR2HLy+Lem/JcQdgbCaNxZCwz+3htPpDnc9N
ciC78PUUrmoCWguL4D/NSlcJKlccQglxSiyJ53fGsNW2ElERlGNG4UdzOXiBlOSt
eo5Hlt+mZbYSMA+RMuNnPPwuJ6BdcIQbbGwi/yiAVQDA2AYhJOqjd0TWaemj0Kyj
PHzGjRP8KXtM8GaB8g6j/zui/IKn7BtBM3QhfOanbP2Pb+2spf+u3vXGTZAckQEW
65dg8NtTY6kHPvEYOjXPxtMxthkVpeYhKyGwiXkJKMH8xoeJRhpqGfK/nFltg42Y
ZTm4E2nvweKgVSpEmKXwcSg6pR/dOdQxWNrZ/xFwGBhggVMYRSrRij79JI6WSd0o
7nPodnTRqJiEd5mk9sv6okDRZ9o3uEzavZuwFTGv1RQDvPsOVJBwJWp7gi7AGnZd
LrB7pJS3CMNKOfNz42xVqmSo7xl6uU1koEM52FpdqAPxCGOynqlN7BFyyp5xYkvr
Y1/+Jkrgkw4xhu8eyVd02lnqY20FOjM1r2DqMBQwJlwWY0sAvoIEiNUmyqGYsMGE
ftUvbM+iKspIJAv6g89SI4OFLp2ShaHeKrh1KjsDhZrojDMGrzkvx6kcjD12Sere
6uaeSnvsFIcq+vrMJJPJ3xVjkB7OT6bUTfMmU+kFk6dn9u0vDaEA2GhgW1uSB1Ag
84owOcbaulCBwkN619kLuIhhIhzAWeJ9pDqwxCaT0eTCH6SEVtD0bN5X0OIu+itW
tJeiqfVdKqZd/w58OovJXKRqbrx2U/N3MOIqvji59W9HAGkBTMXxyEKECwPFZkCO
J0xhbVAzvV4LXypdZ5t28JRro6v5MCBMtndO/WRhKVVx84HFAYs1QbEpKP8qwPvR
BG1HhuJlnzStUsZ9M/VU84h4660TNyaL454otXs0ZAsuk19Rdlo8py30Q04AM79f
sPsNs0re1bl6r3QYUq7frMT66Erg+lbTPqzmYi5IQYkMU2Y3IurCFDBUS1dePXyx
zOK94EU8rpuLXRmkCMLuCYM2eOualfIvnJA9LpCi1jVEbnjUOzvCQfKdx7mNMkhB
ccLvnTZT0GqNGPSllfFJ1esK1fm0hRfW5wjFhutKcvAOoEJ92kXKSkOlMaopJZZn
YNVGgXuWRqO95Bo7qLA8HxSuHuVyjAEJG1uDKtJFCyR7hvIAgoUu5wgrS2Qs1qx/
bI/oDM3adpnWuFxKvtMOEzQGtEou/ZT4j/zrU5uXkDj22yrPPx2v9/vwD8OQCXbL
7zuHWuSQo5OWVIevfn5MNFqi0gS9N7JBu89twH33zCk4R6qyNnpQE5C7BhtvLJif
NYM9Fxl+6TUHMe3M9hBtR/Q4v5uQuxinHHt5K4ykn8ntA8vgPf2Ecmlvaa2W46Ks
R0Q+qHiz8AljCB2wPD1+8+Um8yenQkJDeE01RruZlf8iaPLaoTpjtthJz2aPYJOO
b47wA8HSHu8euEa5WxA8wNCXpdSNpP4YvpAAsTHp6UP6t7GdUiJywWYRIfJqeihm
0tR2gLaZ2OGsXLxNKW+NAbb5dP5kHXPqjrvrsX1Cvn4U6Q2jPPstzBl4ABDODSIp
izHpGDyV9tXyStZVModGAfDAsFAE0ANYKo8qvaKO67WXJXvZn2uvD0c1qB+eaYXQ
nMoJEbPJLwNIQ+yEP60ozLRdgFRbSgWghNJ5d7gNDmqVAMWjitUSWsb3dch5SW2o
dX1ttgvJ7scSYHj8scJHR+JW04vZBRgqaD+A3MhFMVQCLGyPlpaW0Ulb269V8Hv5
56L8NZj+hS3hLwxTC30hgpGwREQiezp+uTOlW0vuz4C5GCX8CbmM1zrVb+jSxGMQ
NxTJFU+SJKe4r+LTg4nzgtsje0qJbjEG/JaQYHr+gQ/c+TfN0i3J7PF2YjB3g+dk
awSwluRsyh9HaygOaMdz9hpocz39NAt5XkIjUzFeWoCPGOwdhbr/ZN8uxPFFGpCH
B5yc96MqDZUeJDCUi7pE+wtTng/PWnVf/nnbQsPTDzI8MoZNeGcVLh9CbaUIceAx
KG0UZDcjFEnSS+hspkvLxBKXe9moeQixuU8IM13gnIo/Asfya/cj0HX27XmUQXJY
06JsMVQX8eeWSL+vSyEun3w+gpLbPoDS31nR8pneTBzv0059lPuYEGGym5uDkbkQ
WL1VdEkL4KoLeRjNFcGvwTT5PZYLrQCJelGMUoW410tlheYtm8hxwjZnoVKADDub
7NuKxyP7VmSx+U7cgXCNtDQp5YcU6pBg85Ki1D7Z33G/gqfs34jHpe17YhWeuYxa
gay6DLMDHJ3Sd7Jgd52LXqdxg5Uhw1Th/gdO1UiPRB/taWz0vqZVH8sME31Yk4hb
D5X0iGzO0GjcfmqNF61kL/hlYuxi1RbhdrYzRsL4YvpRxvrOSzzx76+4EgXl87oo
aVU1e+CBUEkOxRVLlqGrN/A/7tM8Ymc+a1zHXbOjA/ddvoU6Xid2sthgXTppDK/f
VN4RV+o7r0+GmR7HBPnvxViNRn1V40289mL4zw6/YYybRDcHHMx9laLs72QGwlSw
PV4DNfkxGzCZkVMCwQKREIYT3u/bd7eZl4V61pTRycWHkIXDjktJpSEBU1Krgchy
tDyaKxO3baTVmWuQge7il5E4xT0+XxgsSDYNEg4yfiDgsbPaKndA50ANpunOrGfw
sKNoBTF5vpKIwvs3yO2KPxmajjOY2VYjfAPJ0bpCDkiX6WMH6N+1T/3MHAiufXr/
6g6URZKSL+9LazYvuH7pLsa+zk2ZygQ3fN/RUTs6Sxr4C9bxxjHjLy0amygxGuNH
f4K5qB0eK7IMehDair6nqdPGzbWFdf5ovyhHsJTC/9ZSzJDpAInEnlGughls7uS+
nSpfc8KD2fQZPhHrXGwa/otMVRHrL8R7memGOBb425ibd+1JUfFLtBne2HKazmBz
TJT59heIyw1RR2upauvlK+rH4XA6dzebMZY2YGpIuSn5vy1UeqRHEde00lekEG22
8xCAmVSXCeedNIei+c54lfNiIKK8DGLzeU/kzRpuDwZquHEl6nsf7V6nao+X7Zlo
M7YZjx5Z60wjGaMxyef41SKQ80ieH8JMxM/8b4XKvTmpgmRgL0YWV0tQeHduD9cM
edbX6fiUybIyVvtx5tuDDsv5LaP7rKvFWnvMsm0GNoXQgtsflKoxvC57eB9k//yC
WEcNpdy4U/Z/CJEvTV1b8EYu1DuALQ3hx7CU6cda3wcZD0QmOVmp+stdQcPCnul8
T/pt55DXd+WIfPUNuXr+TBlnIKVtXLXSuAAP7iBit7HY+rU9ILn+Hgusn0QSGDIS
PQXFem2FYNRL+fuAXX136iA11H1+62T4INmnDFhbDWkSuLRJFV9lJrNKtIwInJGh
F2mH3ygK+UrI1230NzeHWw3jNezb7u6t/+NIiD5qJmRR1MVb2ELySfCltbsqoUKF
G7btq2eTiMysPk6hoR/kLNHJrSpQAZqz89P41DHbeXdeBjyb5G4bfWfW3dR0awoY
MXBev2GzVIDc7VbLW6t03KCcUHgu7dCZ5tK9GOJOYOHlU7AkWid7SFdoptKxv3B8
THpci4GsNzH268gVK67CpYS4WbmhFno+i9ElTt225WNVJbNdy4Efj4r5s1WTGLoW
NJRBsFz1wfNL8dLiA6kCZTcyS2E4Wn2MPRoUz/G9NiHbTnsM0eA5jUdJDuyDXlyl
tQvPJLSrqFOA5Y1Q6o49ZL/v9nZgC8suH4JxTks85RhnVNz8dQI8JNjN6ndtiVoh
8Uv4tBDQsxNnUv6qQDr4NoVqOrOtzJXs7eSOIFJ6HHUvP96t1hswxzKPugcAjHyI
XM8G2RBmVBwN6tPflB6CSlR4iXA3lq37MSEj02cOyBwidyOvTrbSDLyIHGaEFkDY
i4tooCN/t6KdiV1Daif8b89IHi465sv/PVJiVuceBkc16M8NpLJr4d5p+MHgr3tu
56jybSm/29Lqza7O/KUbMwMF/YY8MnJkFB59y+sXv8IGGP30arAbPHnQnbXs1v8f
MT93+TNAUhQBVSRzL/S+T8e7z2b/meafvKznH3mjdI0s+kpmiuztAtVNKNVK3CSG
2vpHTrYC/yRgsPqfhAyrWlRfbpE9OOb4fBfuGNlLHf81Hc3fs/rOI/DMj+2Dpxai
SVBG1k/I04Y4Sa8rans45ap1y/3NHzhOOD3BT5PvyLxE9TScB63fxW6EZCPudlEV
9THTpR2Jzuhm310McgBWVyfmPUuro9j5t1O+56Ln7WpMUTdY7SXeSVqzW1WqScF3
bNsIzbhSW87cUlx+TRa4H178kvGGbvP/T2Gtj0bRQSjHnuDB8931MdE2optAY/MZ
xA5jNoMYvAyLKl7Mb2+uPzYrHAhML/FsfsP+XydvYPr3VHla8NI6xSqq8+2m7dZa
tPMlgYE3chmi9JZl7/zPSjrL22X6bPYtWOHtTDdV9aOh9D1y8lT6RtX4jwY6TQqC
IjuFN6UKXKIS1rmPIHiIzothTggFhT+ZGXLbMsOkzltQ+Wft+TdZQjVVX1XrcP0Z
ZAkHR52S5Wp0kJZ2J9td4a51W8dwmLL/MxpBbLa0HkfcFwbtmjOrBWCvVyyhta9U
rVZeK8ADt/IT93CbKneqeLJ/fG6XudUqAHHWsUVB8ilVfvi0s6Lk6lqEL0I4ppTd
9YbSVKr840mPIrIFWWzPkjlXrReJc7M7EG9OrM6L/KJtWFt3faG/E8SGYtX6dlCw
/xeq6lGtwrLT/Px0JovnGa8d7dx+OZk7h7HyAxFa1YDvMoWJjXFRgCfwDeFj9yYe
GQ4Nr+Ry14mBQGDXTREu8JhmxWZaEMR/zyuXkzsAA4FZ2/WszvbtCLOVijlQUTon
yLeStlrYq2uHzQCXly4g6vtAACcTB7QrT54YLoi+5wEsW5qCgDwZgz7S5OlwXTwZ
AavyXtlaWRnDZUzz7vzsOEnS/0cN60fGXheWQNU9FwnnY8G09SARt3WwehR4cBcg
qcCiCaY+7UUzE+oakI8uwFHVfC3Wooc6/LvOQET9Fnic4zOFNT5xjyW3AfaL1ez1
Z3HLvWbkV9Zc1qTY7g/rYwB/SSiyMcZVauXUWfObtU+CQBeeodZjyUsdo4uKrJAY
q/EfoDEsMh7+N0dJrk2s/6MH+odOkd/iDHodXsvmpKSECeNloM+hD1cK4XC6VQh4
Gj6lG2TvIiKCpMfW530Cu0BAqsbdl9vEXjGL4iol5LeelAOaOfd5BCYdOokmsdAD
gZ2bx/dl2T++8j+ajx+TbB4xocGYnhAmHFslqwXEplyW27OBzzdujKoRcM7SXH9u
AabXtD9AO3+891TUP3srY6IvlA37learUfFbSd96NIJvmIN0dhOCLmJ8UqaWUcNz
utKlHgFejwDJc/sMY6pzP7Shf1OnToRrtvpnvnjKirTCU1bY6F4nb6yjLHjUhteF
0e9VhqR35HkVHI3qs1Xixg3q3d357P4LCa4dJ+4WQFQh2bP3G8zs6anGfX8OeQN7
K6BvaGmSYoeHrl3Mt8rZfsMKFbu0l5rsoHUUNkv2wz4DNvDlZgtxiC5MlvqHjhnF
9UTeVFI58hChfqS8ToE6HPDYAfjY2ntDE+pNczWDpuaTkloJ0eZxbx4Jpjr4aj82
mlUV21nG/LXiGMIvd2f8Axp0vnpr7p2MBu9WoEIJWufe7JRiqg4Pd9FDqJd+39+e
PSct+dVFic/vWqnKpoyRWZrzu1pjw4KL1Y87zCAffqbTcPq/LqxkPR7+NC1qIOV+
DyiRi9ErfQ9PD0lgvwSSqOVkOmWhO0dvr0XgTrCHLtcIFBDyuJCWULrSqUZQQ40n
97Yf5o+y9K+SSndatCGcMq6KXWnLLd064CDQY7fxXpadhdnP/Rp2lKnpaz++xL5j
MB0o8KtDqjIofcUMhC0u5pUsZ5GspvOE32DYi/LxpIy3amp+fOmtYWMt1r6OlgIj
vpbuyVPtmR78IOCjm+3tRW3a/b09vYk7bnurU6HbWXJ9K78IS5idDzRO9KnDUX6R
mQL360lh8YUqw432rvjBNtpermgBa5cSSbrEGQMGYauQePQBn1+qhPDEtV1hkUx/
cJXiwCbwhHum4i/BsvF0VLsbuLgGLXFsuChhC4oyGPZ4SXK2px2poU49yvu18Vam
a0/rpPYSlntf2OvciVfT3sWXgdSdjde7iv7ydZ5mbao9jLEWpnl+7JAemQjefZzU
ri563dQ4fXk1DEkv1Nkyl+dmMJgflk/kH13PT5nktxcqkrmSnr2wxl0SS0KXLpli
h96f280jZ/BbfbJT5TX4Dk+nwTj7kWaEDE7aeBGMPYaJFj4FWG9SxutdKgSKVFuQ
hPXcM3h55jhvvFPMyWNUnePOOne83dfWCxPsYZyOqw5ZMtggfF5eYagqAJgMtmRm
JcSUXDW1EvaxhKiSt0nHwp9RgIb0aOXOyaOm5AqcjHD9BLwpvCSUNhtmts9LnhSE
ScoiXNXuNvjyI3NuwcdA63jkXwcAX4We1Nq9J5zgpNiv9OIXXpCrHvKUhYITyR0I
LBZRhjqWboMJPr9LiHNSOyVyfkuFYGHHxSWxyMWfnOp/gwQ1WNnJbDECtROY+K4w
OiPb0KnsBOEv9FA/nAYXvkaQI62EL2iBm4N6VYwjgfeekCR6j6cZQTEGFZP0fbzp
nfda4jBjLbLxCjxrzYW7IL6Z0e6UeSvQaihIgi5+AQIdBVOX9/CJzs0uJ44QIGz0
12j7nhdhwdSvfJTNZ4HYIJKWDpSOw9Gsk4ol+sqvZyh+Ejb5Ot00//QmcU8vu7VL
BrOjWzhM3CKJRqpU9X2s2i5tkeD2OeowOf+dpb8caohmeqOfTKZ/w3pNCHJjSXmz
/5oQHCFzAznFjLzg0uFyb+QZ3QrOVKrwfRLrw6TPjhCRzdZAVEgNEcesnFvb7iSW
IojUNDWkN74CLr7JXT9qQcYMw6tmJLAybqcfnB21a37tKF8Z26u3UpEm+yuWdffO
pffiMbY9aU5Of7L4FYXxkgC5ZoMryC7EduDpG6K0y/FZAETw/utDzszr8QBpcGOy
GkgSd98zLFsV8ek4NwShS8OzdsuXpr66rI9yge6pIykID1RTKJYqKRt2f7wRkqi5
WleM2vfegfU9+L82UV/Ci160Z2ddLYhoxK5UTIQjgjqEowLT8Gdw52caGZTQ0Pfz
l1To0RLouf9oajdqQ9adstWwrUBxnCqyO39SjJthw5ae+2ZP0v4MpiCOTnmrNnL7
VWBJddKtWJ6boiaILujB4pfuMO2Ku0W0tSM0gW1UbZpn8mv/XTB1r9cR3mWcdifZ
5nV5N/Hk2i7aqbkR4ow18jMOwuZufEy6gLm0fv3cZVnEwykFT3Ub9UR/lhFpc7Oo
DQwLHlB4UZqvfccVq1+zH0FWkc8qFZw9iY9IYGdYK8UJO9AN3isBTJ1EAVNBS0QR
djqV4hhoo1dh1YnxZkz/0UJp8I5dTx7x5q50HXdhWvImiZ4ee5X2HiR1XcN+KDEj
SA1Twj9RWcVUU5qb/9DywuzGbUwM/yjOzrCb10VKzOXt54j2XkvZqoZ2OXeNrxlg
VhOtaOHYRu0T0RObQS7qgfMkbh2IOF5Wq5QDFchfEk+1okrp8+NOXWKfLzQHh1Gt
5rh8awBGwYnl6HidDIUx26GzpFnQiTyfEb1RMY0h4dSiLLMmrPkAcf+7Pcg0PWl7
XuM8wbjsTahlVRhslWIRaxNx6kzPZ2YGI76eDQC/9uCOVFJuSsHqrI6/7ZwELOiV
t0YcP4hJ2auM21b9w8nNz2uzUH0DWDQp5zwb40J4adF7sJ/MRpaX9c+c5EiFwDDw
VxujMiE5uyPuEAbZX2JesSHVYa0oZ5bfmbEGvAj6I+LncyQo8yEKXHV55mL9AoFc
c4UIoOKDSc6sUIfX5vD27RqWx5vw+qPsdfkwVWXbxX+k+qSmXMA03no4XlKZArSp
tIBlGz14VNIwPATuKqy5iwZSfg6vWfTaDri/HWAfcNlp88sRQ6V+KJ1na71vox9b
YsNE2LPX+MgLjbgeiYsabiiIzFjuE/gUUZwa2gh1jCzpcioiu9uRNcV9B0n6Sbc9
tAxrA6shD4wwnfb3JqaKNqBvpUR97ClvFPViqxjA4JxbHSRm+4Pi56Pj2tuUTTZJ
TnbTaxr3ZSnv+O09Atoz90fifmYkhz0GLzeGmqNn1NkV2omS5DI1NBInXyTSoC0Y
X3leHVZ4h9ed0QZd5i9RCrTUugoxk8DOR1Tv3a7FP+mLnJsgH6EKk+QLw6ouTsip
dQo8v00Tw67dYbIjVoLxo9MzpCDoxCjKoxbgHAWuK/T2AS1pfBkNYNv3/SpFjtcK
pA785yJtWlrvsFKNIaPEvu0D9wDEA8aw/OTF2wj3x8N3kzD3o9ESv81j8YVQF3ZE
zE6IZXTEQa4H40KzxXdHBlsG7FxVjYnwh00wrOzuERcd91TMUn9Otbkf1fJT6uhA
LEW/OeN6ZYp9unZ0QRsrnbyyZFZPWaoYrrwu3/IOLjctwiG6eaeT0ez0NHIG2uK4
bExB8opqc6T2HaaA2urn+R2WlvC0e9vd8YuHr2ARDnF+A4S8FpsZduxN8KL5rbQE
9XNf3qndJhRtfZJP1MvH6rOJmDbvlTprHBezLwnHWTljVUcANoUo0XgLbYdWxnCm
+E5RoyZkn4Z3IXsqpz32YF1Sz+MwoUyzFHp+BIrBuZyw4ITCM9wSlgQ3hxXh8Uqo
oQnxaU/5LPxtjQE+auC1BQ9hS/LcYDRoLJtP/A1ZD/inJoO8JuoEY8/tKlRQ5s4I
UoQyc2X+u/n54R/Trl7kQdcoDYCehSuJpqc76ZuXXOrs1hclz31aSM2fHfSq1+BO
5iwvQMjxT6juiH4AabMHKJXhKM7GlKdJhAycEeEL0UlWXZgLwq92djZXk3B1qJ3a
WHwlWpnYu4VXdMD2lJEtDLVaF5jYmcTPfEnQA3N8o+d09u37UEIlVlPeKtF0rf95
P+nUW439auz8zvRlZG0TM9HJrRiJoWvMtxCViNxrFFrvOPLb6/XOFf8XSrISwoRe
211tVK9frfaSCASH80V/QzJ7QINcwBeX4zdXdRi+0paIkC4WKDeaJEd1XbvrLhhY
P4fKZBVB/A9EPGYpii74UEf09eUM1TFV89uVjaT6OCLuPBXYeRhNRcUetLCi6Xrn
Z9B4rM7r4qkBzYPU8gVDc0uv5RdUZszrGuWm5YDZTfYGYI4Xd/aMF5BK5oMow/zi
Nx+dO5VLrNdaCX/NLR7Rc3uqqEtRQVKWleof5Mr/3Qp+V++5NuPmMfjERQwqimQX
ybKcLe9efe0/myPtOaqkMr3NcSbjmMdv+CKGyhJEZ1V1YzCwUEi9fw5Yq+Kd+F/D
Zkit5NR6Ozv8rjld2cAkuXZDkdvgmt6r8XZBP8r0iRcvDPQ5/yZ37T8/6v0Yunzc
vSIou/j0bDV51FTSvdSa0oK4bZrxsYepDlp8skRU2xPQeRX/2Aa8bVllij7KriIk
yW9WAdBMMj54Srt8KFu0kkyKgJd7g3ko2AGejsb2Ps1fCJwAMNIRZaLs0NDHrN2q
zAnvqtAjur5J0eUzUa7lF3zboAvW3mrMM+RGz3t5Plt27Ua3d2q0kVfd0zBxVIK/
BifMJJMYlCLYwHmnwpAyr/Rk1LD+RXuyp8BmAjf7wqI2BnRVuuieVFwslRvv9P81
Mrh8EaOC/g8bp6wVnZivtng8YHhv6fIs5pG1wRcVHgByo/LDOqtkW9q66NSsILHW
Agrg3JOSrrnID44XlwQ00JB1V+ox+CBwWGZuhlPYrFIn5HiZ6LIXwlNFjlGpdFkM
Umrwx6JMhvlgkG4+68Sk/KEihlTnrGrGU6rCBIMnhMFau/ieCjLpWeG5osLgco3T
mIYZoGkkhJysjoCuoMCtjwvXVWuS25HwVlH1lqsoswYZuxGHv5E3pMTW15qyANKn
b9dzRYYg0N6LOI+pSj7AzOib92Z3AXffwCm25ugXOQnIQ723lN9cwO0YHEngozA6
MT9vo7Ncn4utkbbb577YKcznLG66TpQweu0+lN09ZSze+gy5o5Bksp62/b5yLdsU
sEFqhleACjZIYNM8I94ujl/1S3ATqgG34bgEimQnZV7B/W8RoHBPb9wbwQtYCSD5
QB6JSqdDctDm+M6dl4kqJid3m8E32UUOOuu7CxTxXAyJr3hGF0I2LPGD0fgESAYN
rmQ9ohJHITCeCHGi+MmPIMu+aUp2oIh7ktGPDaVREdB4tzOiiULV6dhIUx8h/8+U
c6K+S9bcUGHiBaF4BGvm6gd/hqBlEYXTOk2HxyzIJn56fAA1YfH+EoMm79UEEGn0
5Ln6hdP/Hx1VuijRA0Pw9Jh+19RHlxQocoGh7ocmQa1ZWNkh8GIlXR08RkgkqfaQ
no13Lzv8krkb1/FEtLd9Skr1FNZQx0NbPB38fghhatPE4B3gLv1iPS6HCqL8IS9P
PCpOAvK9hi9TdMTSlkH7Q09rhlXIUsQuVQY/m+OZXgs+KXfY7fEtWOFMm20Dy3sJ
ZcrlHAwPnEKtJ/MlcDtlPbMymdsmtYuatd3J097zT9q8+VFI8uH9XOpSrn8lrEn4
XNTvtH3Ez3LrigkVsVW9+1L0p0+wSwXdKBAfc+bBGPISFj68YycBeOdNqV2dqSIc
2uu0j0TKJs47Bt24U9HiM6wxc8CIVz0IMBSbJ6NZWYHAhow3vR9b8i8Tc8FapoZb
Ip2ICLvSZcZXNCa9wRogTmy35YNrt9G1IQFYOMf2BQpySwSUHw6ajnTE0SHu2rU5
KippvEB4kRRlxNPanFemO8+MwcWpxYUUBltq7lHF2mdpIa9Kt6xT9Boh4xvBRplb
guH9FjSXlX9bP1R9uVrnwGmt1FMwZDCdSCOOQvBWbFyPzXrXQPzOjSgYa1+xXu+L
fodaBqwcvBcHdhz6rI57JKeA2ggRaHh2ZbdGLe45bqdMmQVBiAknlQjixitzX7Zk
CgOMcsOCJ5hWPstlHLX40MyBeluVDK77gmpas1oyPMOm4KwjbD4NP+Lofi1yaWmM
tjOgspGzn8HzmQiPXRRL5TOjZlMw4Nch1ROPeh1c64BRuKl1nm22AFD4ioTwjg02
3QVLNVyjXF0wVGUhcUJOt5HRr5kuIXeHhsZCq1Ui9z7bPdMSNSeVpai9llyDgIHY
AlihIEXM03S8TvC8yKH2cJP0XvIQasJdk/emeY7mcYZfajHyD/naEwWPgEqfG2h8
npsCX9VMJaIbuRp65cMlBwnymJwOlA+DnT/8suV8oB74F4uxYzL9egbWIwo7LZiN
TZDWHcqLw4agzbgI9cn/C1h2HJtO4vTSxdMSHfgYquRB295kK+qqt1dyBq/9QNUs
lMaBh59HJ7z03dQ7HgHDFGJYF8wv6m32abMza4kBBoFQU3xUOLVSPI0w/cg7Q7d1
gVtFLPvXY+EwCkEdaXKSZ356a6l59yLUmAM+5uhcuZXF3MSzZQikMYazV3is+ZrQ
wruulR2ljYka9YPI0shOX+hskb/NxR5GjPMHoOPX9uW7QpNpML1Ot9LT0aYOlt8g
KKLjsGS8/5CuY28gJdaoi/f2hyOF3brCuLI9HSxyWK7UmnCccRTtbBMcqh3LY/KC
Cm5CdTE1QEdeglEmjCp2P6okdaZ3Nv1blDOUZhsHpfj6cRUamwOm6xq7tPWd0QOW
0eQVqh5KU4uSzZK+ljco65xGrwyqP4EiaonWNTvpQrGTV4Mevu39Rg1pGDfNdH6y
ru82LkClHCHqrijkQahQa/zsY5h4pBAUb2mEoSBpdMAtMfDmG5r+9eO3R5Pz/ymZ
1EloAVB/Q6PaD8BWRBLXujL0lVE36igfXDjbWg6717bEk3ouBAOFlIEmqA4p+9Yl
t4RIJ9z7HrgKjrrtjQbXOPnjtYqQ0qie7shNZgnovGvli0rgEcdW77K+Z2AM+0r/
cpGbo3sFJ987ZQACKWtE1l6blbNQGouS0ZjF8NmnZ+seB5HImPw/PXkO0m/+7tnL
K/mhmqmWYtxd93UQQBynIkatHVH+3Ats9dv1ZdNn/qtNVflFoylNkn76aWdFqlwK
APD1BB9+sxwfbrLf+Psj/5sglR7dZZbw7bqG+aHq9ZbCNeLyp5NK8JkPcBopDSIc
f7L5G/HHn9IzbYv0/S64G5V4PpjlE3uSonYRzz4mRwd9Hy47NlP8p2MWibw0inRi
5A8+0sXn0+ZErKocAHQ8FQsLIU7kObER5i0lAc9b6YavRi/i3pAilCf/PoNS1Q2d
IpSjqK2+wMr/Bcoo5UD0WU2dtzaXWgKZXtOeWrEmIgFoS3phsGAv34g2/Xl49bog
PVOJztfE/6w9+V1IoXNNc9+TUav8qk9/LboFOu4M6Q1lhO0mLEpBnLRU686Cwhd2
24/nPVdEMi0MKu/ejoBCSwUBZqZbUg6L8bBNWuciaJ0Qp+lBxd1HFM74BXDE11g+
sFTTc8D/aFBQmSlxJR1CkHXQxfp33zrfCj6pFlpMOEl06ex7aWYAknh8GrTbajMT
h/ggnIelSzuNXKcOTz6w4hKCHKm7LrpAzn72B4/5kRXgchIvjmf/nNGjvtVXcutY
cCwPv76YCJlPaFb5lKv6W5gMfihtYg5fBEY8vLCxuVN5AqdvtdKOyCfOHFKbmax3
3fEYtn+UUSuFy5UCMjIVngc6pfwar+ZgyrZ9HQw0NXRaikW1L4W4o/OxaUj/95M6
b7/4wjvvSLiKVFO5UOZTBjioXrjoRuOJ/KSjIUv924Gvx3wiv4yHANfb8D4+nYgr
VTh+IyClhtTpRG9Iet9Xgfy/dPRiMXgE6GBtO1TV0HMLvE5O+Muw3qBX9Gtz5NCS
eAa25LVBoEsDw2/FMJyiDJtnRD/HmFIEUsdkXE7wdk0MUv70i2eAsJp0S/WjP0CR
Bsc8X1ktVc7c4Xl4xuY0JJRqrTVlzfsxs9lGrUBvIKFrFIYrtsbis91+Xq3i7IYP
D67K4DAh8xrGQ0TJ4cdR12glE9M/8wGpk98cgRBGE7kLzdCI5lfS+m/nf9Dki87v
Njlk8QONK4/LdbLd+OJ4lRaXWAtP1MdPeQRTpfc0kvkOgx8KJTq0sGGl0pOogRS2
SHNM9Qa1TyBvMyG8bYf88FDi/oQnehuIiaFHW5TSmR2s0VTRKf9lAaX57KDaXJw9
ca/lBEpq3LjYBOWhsVvTyf4feU0cf/2d985M/OeXzFAGOuI7TtFKW+O5S/kMb57S
Qk0+YBs2lTwkxwx7tiSz8ziOXgoD1ZN8zIYqXsSTVQrG9bGGNPH9mGs7cpVMnetW
W6D/ztQWc6i6UyofNAIfDYm1GURdUWvcFfAR6zD6A81UKdPVVJisbLfaGUAsF2ol
eANIkWi+99Y8y/Dwa/bUl8BoASOMGhqVyg0PoxLInlIzkiJ0qYlZJos6NH40dGje
LCanGktjONBNXo77L+ZYz9ZlsY1Rr9g3H4PXttm46x6K8rZRj5Y2BxiyOWFchsKt
3z17CbGzkajWPGIZ0hEz04nnwgldIWDPzkOT+dd5EPIdq0BsATuR4i5JaIhkahRz
nSjnCU8+H7wlmJZkQrnztNV6M27yF9iDVRbl595znsqkiPWBiwSMnQ0vKrqNLEtJ
MMxNNjvTTt1gPwhPXbdRSuJ/T0RtPLrh3y8YYBvLnp5/eGss5Jh9c+Xq7UsLUbZ2
p5uRSOvVtKEnlZP7NI0rW/q30axpHfDgkO3SNOFMBoKd7Q7fNMJ2eL52MPnXBaYn
TsGseXH+95jOt23zGdfYDe5aIOTvAKHABh4cw+1VlC6WHHSWaEN9/jj+uKeSpeiM
7mPZRGGtKbDTcflAMVnNlMe/hZ1eeQcGMNIXtmi7mRDBgVam/BvYBAuo1ZX7zzJk
CRF/ICevZhwcaXbG64XozSQ1xTZQgYMx5C0HtaBz24KKnd1Uolrker3jVkHpNGZ3
7jbDCGu0lOY8bin9vXJg2DlJQ7VkGwruMZ24VmvfPIul09CoKAkCjasXvwm/LNbT
aPCdYgt48IfcDlDUm8lItutwuJg06QPRPxCiPE0SXHEnJRZTF3rAJHhRjJTy2hVj
Iv4wrQlSUxj5AUHhLUK7Dgz9mEB2xi3QTUnw4sOewfCYCMrcotK5JYRoX+vesSpn
UYGdtSV3zZyLaD4R95B2mJzOLn2SiA7ww94ENLFtFfmlqiKK/OlAU6R5EmzZJmNd
40iUd1NBKfABUcy4fiYWxTtnORksCDxVj/AgxWW/QyGUq3f/k3k0sa68CI/C3PEt
jNHUMA50je13zL0/hTph4mnvTYDkDQ5Se0BzSmZLDhLtUYTIurq/FuYg55NeGH7y
1MFzDaOSYoZLZVLb1D+p94qzQSOgvgtCDB9v+9si3/3Mx4qwSOSB2X3qTZc+UH++
toN61uztJqlthfhmTuxQMpbOeAdxBJG/AimrsqdlUgQKeoWcpN358JCDZMaZ4NXm
ig9SyotLCBARC43JpCr7+m7CNWGYofeIgfJ+UYPd0tGiTWSSxNAEqtv+WtCI7KVm
hAq+4NgPGylC2p8qNtL90UjecTAHmXPkgDhjlR0kXYPppFP7/+SyfEW9Lm2wzW2u
tqkbI4izn+joYpEObvSWC5Hh70damD77T/CMzq90PYrfUhZheEJtvpNzzFKKiTbs
JZkbl4T1/jdxgQ/Mk9j2qBVEV2LsIXq6daQUp/HaXaC9ckeIYJCZlMMGGbgysQW6
YOxzk0GNQpehCPMRdu+flEYxhwAH9gTmJqdqRjbsoQBUP1YzPWpz3iOR4NII4+a/
QV3QkSffY29BJBNyPF/qEhCUiMjaF+cCyHUnayzHocuFgqIyKQSQvFWYAFiu/DjE
FkVZMx6LsCWgLfBDgbN5FnKFuJ2qAYiKxS4Lxecsef2sQgJY1mQ3/0r19A9HuO/A
NrD48HufbLG5o5HWACwNR2VroSIXP8hZhtKSd9QOt2i/VH6EpwfYevOp/c2uODCH
DGi6tjJ5ptkvChkSFKKH+gRcXMVMdpNWSBgP7jU6mbHHDrJHb35BBorlJp0jZwVR
SrRCt1tB7PdSDuVNab+Zw4qSRM2DCcKg5gKOT9G3qazES+uKfI2E7xLcxdw0ab6V
xrjcPN74XXp8z4iO0q6R4GIkjWbWZQw8VbH9x+WRf45lmzj5Zi4kpOeIQG/DuV2o
J/Z11qmRHJ8IqyNClkkcdbwCcDpcJCIt8YlbuSw5Pnt9TlI3Zz9NTuS91QnpNYEi
DVla23gzbGQDNz++ImB0PoVSN9zyZlr84QGT8rjyparlLIP7MRWoq17PrySxqM6k
a+OzoINP9jqw7HV0DngYAdH7UWTraJBcqOI9/jw3ktaR+gI94tQYE9Dm6XL0qQQI
k21ui83vaPDFZAH2EffqiD+J3VmUEB/BrLkBw+msjroI3jvWets5YiH6R0gERMWw
Ut6fqDxmCIWnUP11cB84jEjTPdC5/A18bEvHKfMoiNeG+5tgTyzvY3AnNkD+7hqp
ZbTv3i+OoJiUNmuoG9iW91yWyMXFwyKL3u5Nbov5F1eZY8gI29ue7JOZRabwL5Oe
K593b5I8pidfRLcWbetFQktQltWstVP14VhqKmwzUq914VgAB98BdWiuKZUMZPoC
b6BklT4mMEopy+U2lQFpnAUasAP+Ll4k0fnray1jxS52ie99TLsdCI7Vy9vYRBuW
mo03GYSyUOlkjJYh8iF9s9AfZOEkwb0NpJb8rhszfO1CviwLCl1+3cV6B0YXyQyG
LWni9n1OAvoGbqBAzp14Ma2esICU//F63cVTkSwsToMNAgJI088dodDuiA0nGIug
UPOYtucBQbonD71ZG/o3pSmXJ2pwyqYiNt2FqNMkZLPNOmZ8qyQsNCiTipLxahN5
KwdcqB3W72qA2Tz/Tg9Tiur+4s5UHU5dehKPM96BWN1+yYo4ED0pZ6qQyzdZtpj9
0/mLho3gOi1F8C0GtCFx3eixMaTAaFHIX+ZeVjz2j7nO4Y2FKSnNHa3hECkYeW8f
myAbtINUd0B5KbxCUm3UdDgGaC1axeOjye1CRlMF7HA0b+6tCUdLOuhUg+5ZKTCI
xd/INXcvw4dlk4/+YMFnAwJ1IesEDBLZTyGAf3qoG0LiwJ8VWPWzi4ia3FQTPFcc
I4lLJtti/QVZUkgvPccy7XGSjsQRvYkWM735Y714jJrDWdIcTKMlXP61svKuQWAx
y2R10l7e/k+LL1UoxXQidbonuFANl+gz11zI3UyfIg2VJj0zAvmTwOaOs73D5VA8
QgMDG+X7EGE1+V+YFwGKMuvU7RsPRjlsh3XBYr043t5zUvt/IdC2bRHyZmrGvvWa
POBkiKh21P15LytH086RkiLMMeeaUeZrf0xT8FLLok5NwvCQlA368U4SQ4kUtGiX
euy8dgN/qE8ZoEnRuaquCtLZgR5NBSdQaCbk7HLse78xXHEwvFPTMU9Yo/APiWir
KEhUIB8/7c9pmXk/r7ik4ZJCgMr7bA3Bj6G9O4r2Mr6y0ljtY/LImSBJM2Nug3hb
+f5ba5iTUn408/8X3ieCDMzQ8XFlfg0XzCXahJn3ojAjY4t221ePHtDJoYBk+Wgk
xOjWb1cc8eQek1SHW0ozFzSHXc7Osnw4g6avtCayTJoY7DBNm05U7jvgFhcIOw7p
XbcRcHe+H/h7Le8WwCXPed8k25w5vQXCNN9YngINuqJOEIutSUJZN8SI751VV1Bf
yrI5BjuvwLqJ7ymyCRYt5fhawwdfkm6Q/7eZ57vBx43AFdrY9XPp1i/QWaTFlXXs
fdY9bZqaBkfDmDFBViiVNliFCeygzlo8FVmEuBwuekOLqV+ZEERBqecdYIHLJWQy
0aj+gf061vPtYHvWJpGWONLWfJN42eVs/bjCXTWlJ83UMohnrTaq0Vd24CQjgc+y
7hd7fkmaEXPB3ylkFujhNumvq+xFm3Fmpmgeb5w2yDBeOJBRWBWBamw5uy8RyUsz
Ckp9IDo+IKh6mb+RpnNMi1ykfNqxRHSlaEWJ01zetXL83j5nK1dNdujIdlPrI8dD
cfoStH63XW03NRJn81reG2VX9vD1l/dItsl0dHhHEa3qUmMLmVTjPQe+bYCIs0de
jiSbFGDVGehJFKkrPDdfH84e8VvguwDPkNPbu56edAtk5kGsengGH2TJnLIzK8Wf
apBRuSejJ7tyMOGz8zHv/+dZ3vPchstVUbdfl0QNVzaoDwgxX2RL0u9Fl9NQEQCq
hrp0PdpERKfZtBh9Q4VljwMIh08l6+RTPyJUGzBrv/lUTLO/PnokRav20PkCveRX
t/KSjlSLBU6ap0T5k1bDlON2nsQab5SQOZOrnDGdhpSW83hyVGhIjtYuaoOg208U
/bcfnj1ebm9zkIHW6nsYpgky4RiA7XLuVS2JQvoL9J45Oyn9EealPatqNoWCxlge
ifaGb9BkB44Z/17mF0+tOJ0Sdeg45InzA2VmO8uhhthediTIdk56ua26ncFxQjcP
nQZJKiQFj5y8jmk9UZ5+Ne7mJ+LTJSVfxK8Idav7CVh0I5oi0Jm/Dam9fgorHOF0
LG7NM1n+HA9v9ofcvSPwvq/kVxW/jl1o+OKQsWU3h/Gb5a2ryaetzWBzseS36BWI
NljktGhjSgIlZndS6JeWRPi159CvcWlqNpeewd5/hvIvGrhHrPXs0z7Hakz2gKBr
yK3ziuP0hsuSIBi0rj6deiHqTzF/52LMnmBfjJ5MhI9RwNpImzhNtvKUzl3fam0x
gNVycJtTQ4lXwEEoLkTI7caLHtL9PUkFN5ocufQ+HUaOPEr+WRPIBgBbJud+e8qd
TYmu71ojZCfMOWIL0P1WLwJBsybzCd6MxWkCu1vgaHtQSneU/ebhdzQ2H8htSy37
WtcAZ3Mi7o07opspuAsKK9wYR7Xo0BTfKDflUTSn27spAoQLmG5F0IuegE1h/n1u
DV4jgbJZhQhKP0mRBUO1aeRNmLcMvRYPYOAzx7M3KM63CCwcnmjF3/zu6JyyNO3g
5MEM/2io9FnptymwMB+nRtRhe/kbeXHrGFCffP4vgpuGxFtpwNEU8p4X5Du3I46H
4AqnuGnt2O/4e9tD7j/bN1fS6kRhggCtoyfwztjOmekUOF4B2fgSZ7IdSaWftITJ
YKkJLfYvGMvMreWHzuM62ymruoREmAGqN7/xn8/OUSiUMMH5x+qFJXT2sazk6HPS
FyNu+NopQvbY7f8YJRhLVIf2ZSEQSrhg8WftTJoAN+h4hP9AFtCsONay/sKo29py
nbXAy5iLbU2K/lHV6hFWVWgO8jU28490kgKGVz25oEvDOWS5UG0RZ8KYUc/NkXMf
m3GB+Vl0iJka0YCr7IiCEhoiLhpTkLycqF9v30T4nwwqXWgTF+Ky4tdWWogvb2y7
tqj05e2b8mpz9h/kK5e/yH+Rln85sRqv0KCE+jn37rl5usjLGsvtk9bxjs/lYfQA
KbzCJc9489t+Ppx1PWbtBYuV8/fxZnmpOVn3/bD6LROZG9a6uOAPwpUnxAtGzh69
C8v1fCqbiGJ2Vwx5cAVFPwiEJa9JhXb7HgLxohCWeTbbDplr9uWjvXHniCXH8v2N
tNjnxbrEG2QLuNz42ag+hbvZO3hnOGg1XuF/Mqcw2ORP5I1BquNsBNo7DBtVXr+u
Reu2j+Vxevr3MtJjRRqWu9FS3TkWLM5nzDKtptYYF7axe/0aSVMbDJkQALeRIVGZ
NY4cIJlvq8w732NLX+zmQcyfsZrvmB/hzdDfwzHDj77Q2igE2CBXEhzaDwl9v/Ri
dq3pZA+/M3u0sl4HrJcKNmEkpXOuE2TmQOsCGOd78E0EvehGtnu38MHPlfQQzoTd
fKCPCTWufIc+ge0dMDkL9NZHw5rIYh3lAk0xFwAnqzZ1Suucq77QWrKRVwpUbGKE
/Tr33ELUrUfNhnm9lgTfgdcyrEOFBGCmh25hXR6yw0qbYPfZYd35YmyenlxpeuvM
yoFS3pcQdoYOZ3Kkn3aZM3+gnB8pdWObnox7XpHB7UY2FKdjqC+0Ao0L1+7lFcdT
IkrLrsjvT58tdPQ5LdwPdkV7EKykldCx2w+O0qi8wiSnvhjah7DJNvAYFxS2jUKM
Xjgdm5MO2eWGPML22DOMQBx1bh9K5dms6Mh2yWUYrpM3PgkzaShYcmKv5dskYOrZ
ze7CLReRBnK/pmrjomv/Z2Sut+/WKStXE354BNi9NtHK5r6uDBx1XsGmsPEC3aHX
vnpavVgSszdPDfC3DTXK7G3ux1F1c0r1h12iUoDnH9kvdm19lkmy1gEHfkSQbmid
yK8+hO5073GTRKAWo11itwGkRfCf20OW3nvNs/t/N3sLJA/YjSki/86SM5PMMfOs
MWwQxyjsHOc6DbEqvxYLx6bbbOOQHX9HOVjBJN3WRT9dC5dvdhcspJCspzi84I4j
S+1xUdnNUqfHoRwx5cH7XO3LhwCeHdgpd1D/ETG/c3OknOw0jGLpcDH/SASLa7f2
08k3v2Vmtqvws45zWMSxSGNhgmzemmAbtNJEmPn/vS0vCsvrhyZYzYopA4WC83Be
AQca+RfdLZOdY24vHEIMf7s/PLwo8mOTfoIzxM84RCHGtxvG+qxsWc3CpstsD6SF
8N6ZvYmJXkIU3mXcNwYHCaWUP0WHqL7TKy1mKfSrKm2R65zyjdAx8DqL3XQU916Y
PHlvXU83sQPooOlJK5h8lVKfhePpo7zeBsYawh4cCEQQXFTDyPFUNMlCsqjNXsVP
E+rm97XZfThQl/pqzka5Rtv4f8n29XWHz7oMwMU1VXNvd8iXtXMF0YlBUEO/QSzQ
/HXVsvTTkEJeVcVTA4m5Q7bAgtbold7/lPv7AtLsc2y8VmC7WFSMD+H/CsYtIRUQ
5aNzN4sRczywJC9i0orJu0gXBvPJGAmWdTvuEo1A3deoKq9nO5L5vX82Q8hBfQLt
K5efwMg4TyCxLSuet3x05qE44wlm5VVqlS5lFLtdoo71Ms/aW3i07av+3y0jrUjs
t9IOw5Ba5YX5ZJeFGePOW5DLwP0vUoBplGiDjWGmAvgRzdIZoj320sNHlIONBEcN
NofriB70OMnFrPFIXBY+Nz1CCtNFspIHu/pa1NFJ1muE8RP4KZcMiRZS6qsPR3SH
be6A0gbV1EGX/oxjgtJqHgCgRmBwbSTQOJLQWs63qhLuRGXbj+Z8PjFhmstkwm/l
gTFwgeLVpcoBDS3dZyCoPKA6kuPqnrVkm1MSLDHiez9fEtjloOOhCc9MbwnS/Jyx
qYoajhAd5bd/IUsQAcwagzEIDfAprwQBsPuB+TgZSwYVcGH/CttCbWCizqjkfJLG
IyfAvun2yfQkOBeve5C6AzRARubgQoAadm0gsOD+GHL8oGZmsVzHoioQvCNjeLDs
LgtoEFkljHFklCVNRlrLHVzxaXiD3CQr6OJW6midG/rtwUSGx7Hpc9xDndV6mKD8
XwFb1xDHltAxwT3xhiw3WQ4l8uLkb0FpHu1CGxjd3Hiqr8L9JzIqaLRO+d1fXJvd
7VeA9n+jm89GMpKXQlqDT5WXGQcdB2hMR2aAowY9a1Tx6TZ3Omq/HC24DQnTtXxZ
2DQNIazx+AHmBFnWtkacav42OSLDnZA39orhXBwYa4B4Z9LHT3BbFe5WxIxnuuiU
c3dExV0lw9B2v4x5ev/LOBMqn1nmwdHpI8TMHxgOsmIByRuZP15AEtbH/BJbZArF
sb6RJR1yHLvMPtFebJwj/8bd/HFJSpTkrRWgkOA+tO9clmYg54rSTRbIM9OS+QGX
sFTLqBFXA1vGXaVB/GLwNINWykFpEpHPHvPcNKYYwggLPvpsBt98AzEStX02Dhqp
HX73xkniXDYD2uBaJ94i0kIcXST7WhCoQ2M81K1GqiNk9VWqmHFXQlTp3WpFTAAi
uH3V+IjHKYfTPPSkEdq0Sgp9VgCMTsV5eeOmylUa6/dhrEJJ8Ir+XTcpRuVAB86U
xxoxSncOonWVsRm6xBjyat8vkh9dvEnWOmfNgKLEaZfSYUDu+1ewNk3zhfXmwytN
tGRBSj//d14FLaGqkb5ZdujwNMV8+qvQ+aLWMg7LX/yAm8ZaaarvuX6XpEA4kdgN
XWQhec0kssPuR6Zz2Cr3dMc5E7/cHUwHoJzBLngS9mGfnpu2GDRL1FFSjCgleBwy
vYTSDICoHs7xDhQARlUw/SRoty9N9uutIwxMd77HCunUrlCcnYU8uNsVOFSmF7IL
UFLKihlZjaMOospkJdMQO2hqXpE74WO/xoVHoa+U73fi7ktRxKpRhKogn2Hs7HlG
1fNNxjgjcMMmFUhI+N2VaTlvkTE5aYLhLY2w7M64zLy56OoiJO9xNRCkkWBfu13V
YGQBegUZHLH7/9wirld0Dyix3o1TEquoBt2AHieI9apOSido8BY30qoKwDRQ7TQ1
U6vPYoe99oDovGY7gm8u35ykDIWTR1XPpjKOb/Cg22mP7+NuuVFI/UWRvS5j0tjl
TNUO5PrvtHtJyNGF4emEUZ2H7algl53VnpQ1YeU0pxJGv/cPciJFQ3dcEuj+qgo+
ox5mFcMXCu1iPfCuJpDNHP8zGj/HspbCIVG/DDwq2GY8LloesZA7GPt9tIRt78pQ
ueAkQezkDrfYUkTvHYUvxjr5fP4rKnPW9c0pVF/Whl+fWXQB1MOMnEapQ22a+HVU
ZX6w2YDAV2f5n4jX+wDkaoUlRhzQvZiPRt3bcH4kJMV5W1RFF6TYZIT70S76Zxmm
/PTbimA/IaV3dcQG9Gn5rTuLtzfYsjK/cpNsw3B3pMyieR1vbna24ZOUwqE32jwE
ryG8MZqYe/K520DKsiRfMPGFMbsIvTC2uZIhaiFNxcs9sNkDLhCQVFJqCUgVXeBL
qFplZMg/b24amdiWdBwCMulyxxWVX1KgTYw965FbUjfBpFf+bdA+YzfrNID7s+uM
eumWBzqsbYP2p0bJ7Mbl4ooJlNx3sezFmWuV3u7Q6/ekSrxSgEIafPwK2nKT2RGn
oOJvQ/rHuJ8u2M+cwQDrP2nsTw+A8/tjuoWqS8xRVU7As2JvoEuJN5NTQ99Lu+q8
xJ2hic6QSoQoTgueMBG6FUUm0MlaO/Ki9hCQdt3YeMPkYuNYSY2k+Ygyxddjj2P0
1KAXG6vCPP45KMDW8i7S4M89+OHE0FUMXgpZ58UdIwZ+jvQ8FJqGmAfwlwXpAEKR
9yto7Vv5X5yOlNAP6HRrQMEj8FlsUaRYELQd31fzusGg5agTwFbzticn0q6/Evp8
xwYjSR+jUgsXa5se/aykFYzylnc9VeEMMtjOx1p5ax4uJk7JFAZrAEcoW+fdlnP5
BUKWv9GKIveNArcw5Um5FF7dbk+IWzfVu+Ilri2ZQ+ne8KautcFUoVH490ce4//0
s58HUE6En2MsHfg7h0X0h9KZuBdRtHzpEweipMsiWXfxSXV4b5Vw99DMlG0h2dSE
i45GgcbSblLYnh4aEDwzjrMin1Z9v+68Fb+ZPnuUkVT/Bj6EQH/hAaVsJp2eoWid
qYQfP3RXc1nJ8QMuvV08DrtyMNXy/jgZ0ZRQJk8NPwz1D5A2wjfcTkOpSJtBVg79
Firm/BAZjO7l4hXvO/TPQg6O37W22o0D4yZU2I30BjwYlfHMUU7XKprWSJJbruzr
PE+40E2+4kbtbued6fPwSdgS0i949euQ7LJX4/muQrnBpC6M/JiP4eNAj3TYtkbq
WJ83qO9jBY6kgei60ltcxBfUIA12AZox3Fhqlw+dBA7/83+LEbwj7uyk66hnnU1U
RTbKUS5Ebzt/KaKQILutZ8Q5Dh6ZtrdayvGjIChis8b/jkzCWB3w4fxeYPlrdW9r
yzAgwlUAACN0jfPohx00i2ab9Q3B1q//R9GuZP/MTwz7wcEZcOaNLuAv/E0Fp6xM
X3aa7s+qLb7dzGfvulEmzl538FWWqkIT1yxW23SKW10SRBhRI2xsq2KzeZF1V4Z3
yK44dGSJLAWexfYl8x9jS6Qh2CKGDyz3hyD8V7Ok+Qoo2wXHcfoyGxDQ3SxsVq3G
fXw6i4cxFKGc6I5W1UAREnSQYINg+2w/GOTSguEZpvz81OEMhJTsO228KSzmrc+t
MF7QHSljWIIgqU/54kIFeShb8ro7qgbDMFgsX0PmWERefu8/k9TudW1wfarTozrj
oLcbAa0v5N6L8ntR8uKDKLPQPKxnhI4Cr0WBOYOFYhSzIwrwU+SiCMcMyHz4NZIz
Z/9f+UMzCVX2XrgZrNfF/O7C79AuuTFF9ZSzzAB7y6PBhfXkD92hHttwdRNx87Sv
1FlrQrpbIW/Tm1+PXqeO3JnQnZjgdYdBZ9JWa1ctxJ+7pDQOyn2SUXppkkiwN62d
xIrwRU6yRZFyrOmKOoSxZ4uRETSBs9dlt/eiwfqhd9NsVAZext0tjJr9iUiRW0uj
Rqt3KdR19HUBldKEWPKTfbpqIPTJs+AGU/5UXMaiBBac4pWs0/xVqQ4XeCpeCRJ/
LgYe4AqPQ0+aDncchx4Q053r8qRbs4hEQmL0GVUn1nJqGICoa6c7JbhcUl6EzA2S
L6NsBF1lJOLmVxiWMov+d4zN6Rd58ZxyNjSPlXSoGRfq8jUmsHzg/SA1XEgBZLe1
WD30uJr/VU5eCUFRJpmjr/ykVHCkGN9z+Fupi6szgcwqtl/mGvR1xzJppmVqrreh
iNYoam87rDit1TdeK6OYXgMEem2inbZC50OHv7BxD0l7QrS26IvXYfTu1SwTDaSy
mwNp/s5pvZ5auRsG0wYfA2bsCFEVOASQgBY1f5TytCY0eHr/s7bfEHrGXrHs69u7
vvHCuJpHy45zqWelufQi08nyeL2fs6DoPmKJ5bEPLiPi1+/wN/mrn52BHtp971y+
USnVQGezAOWJlch8jB77J/Q4V5FdKe9nczuZ7m48dJw4MU5u4XZds6uat8KFMLfq
m0u7lNJ+cZSIUql2X79DVeFPMdi0e/GONXwKf7wKyofU3IkqlRbSvKMu6KLGHmXk
812JMctvR6RvV7UMcNPPTuBU5mlwbvvfypZ9k3Iy22ppRhtOBAGyqaZgFY8Vzxbx
Vatv3RYIPu92QY1sJTo73+khU55+LmbooojHQKzLYCG3681kLyk5rDmCYU2TQ1Dw
X9rjAD+2eY3vi67euS9nzTZNRBlX25fFqhgLXVNxLtpBjmd0LpjZBA3Ei657MvV0
N6kOL7c9MXeTQrMIFaz603JB4sWt48WgDdwNs52FjsH4hrhNj5CH980a44JFy/7n
F7mqdMQYA2WhnQ/DhPV9HTsdqqrQ4mBeU4aRaNnq47B5hyidBtCthOkLOOxb4gaB
CiLl91l4MtqZDWbQUgxF4bnDJDzLtxfqvWfxPXq1emtLkakI3zmx6Y7qCcDvGaFp
xdWn7KVz2v/z1szVltBk/5NOiK3xS0QDw/fa0E2Yaz90BELecgODvnPrWRQUGslo
rrouy1FNlMTQtgUbitF8YqAl00i/re+j+7UmU4Umzlb93r/wRNgHJwc43WE8i/XK
GMtSa0JXCs63k3wesjehuIpmlxOHLMbXbX1X95jDVqv1WqowtTpvoO4MwP3olUrF
//ys0YIqX1FsJ/A9VX4xnw3aryWEeOc4QPTAfrnc0t4n6kAZoMFl4hBi3+BbQf8Z
fEPsZVgBgCcPlYoA9AD5osl+jOVC4xQ7JtwaNdTHFjHWERiyndcMwrQvAfQS9ioM
g94zR5trBUdc6aIcPAY+2AY63hw9UaTQ7fhdvtujWU8Ul0DC/Uz3GINjCH9BzAZS
3F7Aa7oDHy9ITTzhgcyiUZtUhOBn8a2nvBMpL45JzGdJ63t9aDx6Z7uvtnVPP6+e
i5JCHM7QM10nB/RbR6QOsgkY+/2YoqI0XZ/3dtKrKAAXHDI6YzEbS5UP0QotFtPF
DM6Hjl7cJ2zvHGBJgRRSXTS9/WNEUHR9O9E5l6ulWeb09JKTLZ//Yz/Hb44B85mG
J+v9+gDmQdKrJR5g7YUkLN6gCsfvPBhnydikBew1junwN3OD7aG1wMOlpbAJWi6L
+/upz+yUT39gztPWcTzTWhn1YX4vCQgcPF6nyFVZxJfCOiHGiLBx+8LNriZX/Ub6
VGz95LKTWSZn7YZNoaydxKszlN0QEEOpdi32PBvQ1UFq93u51j0JpsRhJje8bvQW
AFWHsJ9IzOCufSgkBZsEeP3DgXRE3V9UzqB30z152VhJY6/HfFBqdFsTqe2+YSb9
GJxpItGlwJ+i+BgPtGAVqoVTtelnSwx51SfSkJSLoXqeHrMfmKKGR4T5z+j0SViv
wZuOmFIbU4TgYgqIcZxFwY/USVZUp9UVXfISMpjYOr7jAIlkzgh8hMXLewEh/hlg
HfT/0Bg4RQe28bo2+yJ9F/fRfyfWDtz1Zv/aBK4dHkG9RL6ipALMxft6L+z7Sh7r
cwGnM6bJsI4XeBAT4Pnqw/EzoXbDnQJxOVbsuXzqH/NoNRXuPut74P2OLukQ2jJG
kxY/6Oah78Ti9CjD0eRC092afP14/ysatLmyQahjMo/JoTZf5cjNGIjCyLP3tYyk
b9HOUoNPbuGquSpdd+TeYXLZEI2Fuz2teCKBvkDYDRmjocMHE3W2Q4F1SD/TdiKO
5eyH/SUysH5Jl0tQYc1pEVo1m8DiPA15Osfts7znfgd/HMYUhzWMYC+4+nM0hVhg
apl9qVP88jBB6PGYnxdd1vpHXebbhtWMU7beYrIoOoZiKXzYqXWOljXHMen1Z6ZL
SupsvxciOjO7exg4kmecBUakpb6K/9jRRRVbFPwDxiaP8VEbDI4tAPnXYU7FaJW7
K1S6UINLz9sj47qokFvPrY2Rc+V6SqlhaK0SJLt73UwIb2yqNLxuUfGuDblPXArg
lqcUHl+FAgQkiVSkVVMjgWcCvOIBdWqXm271y5YqJLPmNmZXf9ZUS1zVq7jwjvrv
5rVK66j72d2PnKG8jdmSBaAoFJs9iBf8nNgbA6Ej7t9QCnEfRMFVeiTu1+Dvm/lj
vmbZlL/IGfItlvouv0vbLvJcGQnMB4QrEyi+pX/GvfMnPpIE7HgouxyZpXhROiGZ
UhkybjPXxmLy6mZZPw7+K/T7cc1wCHLjFL9dO197NgBQMl+r/dzVqwd4s6+yOZpE
yk4hyvrpf6TfQaxoX7nQbqwCen0lehTijVHZp4d3advCF1uPaBJLcvc0G87Hrfxj
kcLzP7ELd2WYO2brp1xXEClWLoCQ3Giev0/zznXS6oNKNJwVqJJKL2gaZfCe5pTG
sTZXvki98DxKdLYiEgGEFEDLcWPdOp1xkMJqp/7MJd7LmXIpH7X3wzQ/UEIm2FPn
FMTwaVSraQ5wUFarlAGJEJFSF8C+HKtCtvctTDsgX6Pe4LZ9H33gqgItVoRcuOpQ
w1yVf5n6lcvY9bE4CpjARJI7oiP779KPEd+oDZH0nFfG9gZTlO/RS1KKK+DMMTYj
I1jvm4XWOyORsOu7eFW/NFv52eyuKdYIn27JMpcrYwbqSAr1RoRYIFDWB9EKfHji
PV6HEZkBoghqPbh0AqSqFz/74I2tx7gddQOdkLQTVwCSYcBhFGUpuyHyiF+TswHA
aTI3roMM+EqagrkalovigNCtXGke7TaL3wmXf4i2wVbSDMszpE1Wjz5LRe84AtJb
uPWnFpoFyJzUOf++tYWZHcI4GltKEKro+GahAT24Bj6IxWC0koOn+E/Z69Ufp8wf
1RZPV7lUUiOJgJAUVsLNAamOOio7049zUSw446r8B/Psz9a5HaAXaJxyu7WiMNiu
PGRipkE1F/DJoFmpS5+VbtK1Ojhe/fdmAGIemoFtbUGQvGL3CqOKsmKKxJZ7Wv1N
kdG+XIhY3vt2qAEwAjqTrhRFG/G+ulNGEqAcrvYttstUwy0/vUq1cvZ+bmUsjFnt
jshfC/EZy07+IqqUG36pM9m2IdJdh6M5zvhtSAP7qO6eF4rvsC3T9cp8GbHK9pXu
IFdem/BQv+GAawPcaOsJFPSqcqGzq3ysN/cPsqyqxUWyjQm8Xjz6Tkq0NYq7dVtm
PbSemxG2608Djgs0q6408oUPaphgrSISsnVPHg8TsdGFlLmlIVtyMcdZsRDmboa/
vyrHJOEd6IjmS4h6EICQaFVf4okZjgpGxvQItJc4Ph0GlizE/S4y1eZSNfArdBao
MxHn3gKpqvysa2v4pB9+Vnrs9GOrhb1GcGT+ZJP3bnpNqh+kGrtz4sagGYGSVjVA
lxu61CPeyCpbmIsMUn4oEEOVImprXxvGZd1awvx+lUq6wvCfsf7eRRnuatu78dHf
0YITkUmYZ3DhD6fy1N84m4uomv+VIIi7gYcL3JgepvVVWU4J88wV8skJB8Klijn5
Jyt+82oHrMFqRv0wXDxwnXFmzOsckVMQFNyPZEcvlPEvyjZ0McIp0Cs00GJta7Za
NLsQK5m+RxYpJOMzruPFLV5bweVQOyTqBsyQcM5/23nknyiLOSMSWv1EK/yqpkdU
2ieAR73UiuzsqTK8azdqxKz3X2TSy2GV/Io3A+8VjLf7t4upIcSBufXk2g4cCrbU
90tsmWxDAbPiTV+2uDxsylHSnK6O2kvV1WGWPexgEcejB94j+gjnEd1sdPsOIrU1
LpW95l3Um1D0HSb8UbL8NvWCP/HYP7F4hgij/ARVN6KViC4JlMGTlEDZC2OTc+rU
eFYRtciM/9zTtT8pPeqpT+YEPKpwMTIp1dKQFaOueifuiG4PoGs6aSQmA0JqCe9b
tL+onIxwlWApDvOLiZ7G/WU2f53epKXVpEBNgk6lHhLbAQpgbtUmSPBE7a9YGbD3
lb2BtsnNLqZSibn6RH3BuoH3aAf4M3x84l2j8wYd0RQgzAm3vjT5VpDdd0cKo+i9
KSzJIkf7gkOVg3cesjFX5ZTcU2k6I0rkPkO+PwYe5kkIcODsUJHeYbg7hs3lMb5E
VN+YKS5KZ4EjNRyek1/SLbw5ZYnebwNpEdsPqowhKAPH8kJUzyEL0NEGLGATOUIq
RTOUWK9xItcGvvPw4J0ovX1dxQ6Jzy4J0Q23ZIbuOVs/iJPtf2excPMcEK9KZn5d
S+KaO8GzoUOkrPUJ2KmQjsHINicWl8I4iHRohHFOmjVBtee8R79Ximct8vEluzja
1/SUyOk3XZwgbP4X6z5hJXBt42XO58sHgCLTnIw22texet9iJ6Ijh3NiHB3sSyxm
2O73FIeorDJ3evJVSUjdd55l1dVRxu7ebuit2evBnAagC0t9a5282sXwuKNHf6vW
X6Grq50TxOUHKGBTIOPXl1rND6UbPsEffA9xcDxhEg7ittsLg/9wYK8nYgCpO0AA
YYJ171Mu0ZrV+3R/WXENFsAxaQcElmGnrtvKf2yYy6cZW2nwBspY/JopVJfYIU7I
TRqN6vUpyM2TAPaOYcFVCg0PNuEXoxuOiVDsmJOCwEkHGOQ+CItc8I4/esY7TbIb
8sJZ1dlWpvwCB4NnLehuaH9kcCSsTlLekAu0qn/QJ1JTCL/eiKPgRKucdhh8pnOh
yHLFmV3vV/wylO1fmqiQJDGFqTlIvReFkgYOOMobGwp29pwc3vqNT1X+P9prHJSu
ViEnPRh+C69LKJqx2OXzTHXcIJoDzHEVCNNSyOKClOjF4jY0nX+nlgIvrkN9Bk6S
9rV21BRrr8TRAalr6NRChDnu3htDq3fbeCEbfuO0RR14t2R76LwkNrUN6OZA7HKE
XGJR0m7U4IRMtj5g1Sqa2QMhQOMUdCamTxcDdDa/oaTiRdItPQZvM4hhrqt3Pez1
x39Bq45eXxssxadhpBrAHj339U2lgxzrD83ucRCYelNntsO+tzlt/eIBMZMmqAy5
0y1ACoRlec2JkmUbHx3BCKzG6//lGTR6CFT03iTXSzjf69/q2iraPH9suuK8q3QD
uY+EFetU+iXnKZ39KNMp2dnyb5LQ3gdMfTzVzgdkGWr4bDjwV9fPNCKC+dTurfqa
u5JjGKYgTzEm3dGLbWLM3zmlyfOSKcVoxy3Bd3Yr1shx/OU4jq+Ju7VO+9aeRHZe
eVCA3YtHVTTshG1kAL9kM6dtCuXYjnsjPnyQmg4RfkoAdA4kkwYcGVLwrR178qrl
VUCYITcIrY2tcSkP65qOM3IZzGc6qZF44dfnU8yCoXsDKNbBTog9WCFRYXNQhxq8
BRpXQZRbJosLpfB1aDzKRbO0ZSNQGFWxMsWaTGsxh77wSiq1jwjNDmdT6v8B5Ug6
G+BsNXuL/1u+LfYCx8jeDFliQmwALLFMdiiumy1qrfUkN6ojPALUavGeyJIET/Ym
uNAMxR/zGm2q+HTxIPfL70u3VQVF+Bz7ZqaDhcJ4Iqp59dXugTKlgS+64kRrN6SK
jTNnbAQMZqmqq9BGga5tHj7StufoZttt1cmjpJjId/cPFatza38ignXIZQ6vgJiN
ZuB4v+sR8abuogmmZZJDCfoPZUKZYcs+XDCwu9xMC+xDKJjaoNBjVz3C61B3h8j7
jATlqASZULvSGssmUBWqMDVdJzxqyutiRUWrXdwxlFBv8VanAkxqXwe3tpkm0PtV
r4maYUkPwQNmGjleCyEtQWKt8WObTGE0uoHyafz1Gyw4i0J8CV7dGG7fqlqNcb64
HQ7v+iDX4YHqYywNmh1leKe0i+NMrGrcvsVLPTs6yFE1N7UryCVc2/FBHF1m8adI
ucbXJMJ5gnE42ZMMmGgN/oQ1MYXCaxGi2ST4GwfoaMvIEaD0S322p6PvTr4hfruK
+HIJ6B6wQD04xwoy9GOKxO0MQx2flChRodMEx1pldiY5LzJ5sSUWo458gko8K9iy
GgJO9/NehU/W4NKPJngB81z1ncAv7VaR1AmUI2e22+uB5LfCo1jZx6vJzazw/ukI
tgd3oum/BlIiCiPCVGOtawa5PhnMC9zc5cQOMsFtRdxEwCcKo1FsOIXDVrAPeY11
GvR614Sp+lHwK3b6KGCYAztJJCV+sVR/RMAczPeoFAoSDRrnGtZUwDI01tM5TdeV
krlgcJbi6xF1JOz04lOruK3qzi8/WKOWg88L52tPlZXWNCs18CYZGk5C5/mY5E4n
r3QaOdfHhQiSid1N52/DHvmaqODK+R0LwWwJh+JhZChr8n6g2r55JXeMDaINrvv6
g4yej69d5CuTEAhVsEJvn/sz3/73ivrdBg+Qe4DMZXeL7YEMSpCXnYbsqJECere3
TN7vX21yO+W46ge34bGDHzHwWJ4YzdEvzPq9WsUfRlq6OLPtVNjXacdSAjN0UqaX
4TnuBVp/Mlios0r1evLIS7N9ZFdldxWI9+m1jd1v3wA9rmP5PxyXJwxgIPWgfT2E
OzYNyMSGUFIVAaiRPX1A/NBxcbv+THREA3DR5F2f565K7Qby7N/ABOLxGXc251Jr
P37GCPONL6xwJopJkJRmNXm0c9ZpH0N4e7yYq+b5y1oLcyv+r4CNuO8Bn4RxvBSV
CvUmc3QxC7aE2sCfxbwK+hcJWNmXGDx/nSrFDOSMr2VC0FndmVtw0/Hvod1lHBQZ
Jhx1T67XxdgiK4kmXypOHxFK58lZYcaOK9VtJWjQYv1WiK3+j7yGvjv3BY6IOrUn
f+S4lb+HzDdolPZSF9TJFUSnRC6k5STT0CBh6FmhpyqscNZV8O5y8/WOYqmrXRBc
rUY6NFcmHH0xWNfMvLD0vEO+a7M/v1FNoavH4iomEu+669XcPZvHH0MnYHRfGBX9
hs/kuKDJ8TTGr/3q+CsQwPUeFVFfsoq6gPZZM2lammBaUS3+wLQE640MLoSPSH2b
MJnb8twajbPQQAsAYE7/sstwllD6W+RSMqZ0wcpSK+dPQfvIKcLJ4cyzk98f2YmE
0ZdKhnooycjU1MKhDtYGcKVWlZKTQYx83vpFXV4GdM5QziLq7k8PCTrbghq6MK5f
+iSB99a71IR4FGB2J6TOLYjSega8RQfEq7iJjjQvhliRUCtaZWbIodH/5YR2mAkU
VGcFXpgCUJODiGsL999K588Sft8Wh01woWeCmTXdE2fq80uLeO0K47Qdm+XWMH9d
wLyjaRA6OH7UFIpyHfaFkWawwjhac+LV4onlxzxEFNwrbeSY++OVK8pYV8MhIyFv
hsvKNHVwFOaeDXND30vcsRentWklmmGPhSCUAhld70lI3wAp44AtEorV+iWjA+IV
46CkDCN0c89dn3S1BOAMEHufdVzZq1YNH+v4WtNsGiXZX6ONctfrywCnRP4QX+E1
6p9z+EjvCVP4+WjqPZ74uzU/qchYLRU7N40Hkhm6u9zjuyHbrbwEscdCGUCPGOkN
/D08iiER3j88XRrOQi0b82ABZvYAt1qtPrFspcglqpCyOSMlPAZCAGeuj+nKdJIo
2OmbHA/G3N0mb9BHcL/o6WJsxT6S3GGWJxm3BVJMWwi21uFg2uGE8vPysH2NNoNp
5UpCoLXt9XR78f2sjHbMGUizRoQmNCvnuuOpRuK63TKMaU9gELvQ8YTpnzdXeqVz
NvmswfxwbUEwSInlt4PiQDus85sq2EYYNBbhrr9NrIHZsGWuYO15GpDpoPZVE0zG
LWdzPhbbhw35PYgHJUKDJczSP8c0YYqidlF+SOhmLKbfr610KC3rL5OvSmCSuTDj
jn+p4nrgtCAkiF7aCmSCfv1pLOFhWMMlTlV+UwCy7pABYG1zmrepA5mgbQ0HoGqT
fufO9ydBdUrkXHbutbBcIC0uifMlEWQADOK0YJ7CJh+yFQ6f7T1N33vxU5WI0LZA
LBjefmtoQ5SlZhjgKpopUa+cdjmlPGve1UVVosEwAxYnF/RpZ7Imbl7txz6UcSnj
Ja5sngRHBXYoUXwMLteLGvlUVjtnzxhcCAnWawlxVlOEM54ikEHf4Ex3oCXL99I2
ZuYDK1r0dWQvk3h4zsilk/6KXHP9kNNEt6GQSZmXqLpvZHD4HyES41QTlVkKocua
+XLo4ZfECaZwVtWjkMvLOUAvK0yu4l+E9ntzz9jaGVHSigRfp8pa1Gihje0gB6aW
UzfRGkDF9rJ02U3cojub2Xr9zJzvriAVY5n1+xQTTz9C/nACezwFce7knYfpZ4fR
m0DyX5FWblPFScHCEU1ZzCF8C9s6TOHZRxk+g8Q7G8C+/TNTxb/zLXOwLCFecmG3
c0HKHKGQFiMfvTStck3+EhoBT0ofrJzLk5KlsK2TQ1p7x7iYNUWf2vV9c8YYWJsq
Jf+c0gG79quLhKBJ5FmarcF0AeeYCVdAbd7YdMgC+ldrFVjfBopS5kBXHhKejAOk
XDM/W9PY48DlfXyllk+WCRiy6BDwiWt2wgS74EtjLJ7aWU/sjWlK2SPXRAFIt+L7
MHW9gkDZKWp4O7Hdka1/FTaql4dQ01v8mhnSsusMElP8/+fmXSyL2IEF07iDhfYE
XwnFrnEhlvwJea2iwdT2MW7Hiv7GK0zEyrHn36AUfAJxYlh7tHSIFiHR+Q4n9lq/
A5sXrulFJOB3v1gvu5q7UrcrfbI9+V2TxJNw3BOjvAP+5jzKwLn+AJ+sT2mkrXBF
aSTxPJkaPs4sAPuG/l9dE9WRqM2JLtfCUlx4UjqVsTJDiXG/n0vyn0gnt/iwv4MN
U8wbtEwO7ynyfFJG3HCtxXCO8Ah8yrBuq04YDzV0VUwf9CDQbZlktVl4MwIuqDQD
0e/RiHuEwVNSJOFXb95a64zXXsrhRrYqjgHY6YsVuw2SgXnfupVA238Y/ZdV3L/l
oSrHAhfc7eS/U9ID0+SqJaqj7cIQlK8yoAsFnLOzLf1Vo60rQSECK146dvr3l7yx
/rNQUoFsIDNPiKoS2hxzFncO6DvzyQ8iEZGll6zd7Eg9nKzT3K6Jra/IKh8C5mAj
we0Yzfo0+QOkzTrFRQYko1qoDt9dkr3us/zs71nWD0dWOy3j/5bk9gGOOCwO35r1
KcjQ3WZ3HnE5qx9nVDwf8p4JggaahTcRnqWp20rul6eV39WwQtk2PFP5VQf4YRyk
W1DOi7UJpD4i6fh0exk2nsR7QmayyBPZNNaANweJ/WH5BQhxCWQVgJ/PFgAUM0XH
5vO26/sY0KAzby9D1cyz6Xs+j90QlCGP4LR6ICFuDeygnJgvRnYqCHJv3j6wkgba
cksJ92Zsgv+jS0bZrh/IPKeHMUPMU4tGzyMdCEYzIeigPk1cOCs3tCQRxsWLnPFm
fsYwnZHQywto9JPBJd4PHVaJJ6LzfhbeejxSZQoBOA+G4XH8yPbjLVPA25b5acyN
v8DHivLxEeQT/dmH8+NDqXtuwMiHK/JBWylME4mkIfhqxUQDLPp/0ixeFYi7KKWY
pU3L6eRI07vKkGyectYEaZeqVtqE72/m4SJWR6l15VE2cQ9EDJEM2ekyE1TXFwYF
R2sLsAX74ihUgOz6mQkq2YTlygnKvYEj6NLUbFswkkNhuRY2bZTUmcFDcyeOcJiV
PbJ/pp+QpucIG6y3twHvXz8OlwzMLHEE5txL23BJi4laBoZnWjokuMaDqob4HL33
01dDZjNMIMLYktM9FIigkXNIotLBada6TBpL8qykkkG7wdqFQqdDNSjglCJv+CMh
SgpKRIfZcOk/xxNL39KzfyP/FNDMhEGecTR3pacEx7Xe6d0hkGufVjTtPheG3pJQ
gwJKfPMr0hSIArjr3sxnk5UrJ5rOMuqEO5NN6TIX9DkVe8RMbJqkpwTtrCJgXkeo
D/bHzKccwr1yBXyK16EOBolaDVP2e5EgkJ6EH9fib0BzJQSf0mWlIkrUhmgiDSmY
DOOyuX1HCJWafap9GEoUG6SDm4PrJNhtXEmoKKsCON9qopp5govfWGRdoqtP7a6J
TkBO6sjJAWgR2oCGXPOreN0LJ3xL3N9zJIIrVJnil2XFN/1DOSk0bHcm+sqGj4yV
kGtWAEJNj/uu+2O0ex5ebtJP+fjd92zOyKv2ZPsR5vFXWH7yDgiCi0q4N+gkL20G
EvtqiZFehGdA/woCNT8CbuFyZKlCZCnt+LfSqtlaiYdZ3MiwFLrQncj9LRC88Jpi
XPPURffwOQlFTWoGxQni7rqX4qzrsqjq23+4wq2vYuehTJDFH+re/K2JaXZrXFRw
XYTg962LtKQqjBlLHGXbDCv5FHvtAakGE+bU4ymmez7tHlspnZyf6bcndETWb5s3
7tCEI4xcPLyA64qVSm79Ta7s07Ef3Nragjox7G5Ikm0BDxmGXzhGTKL3ArCj2eih
WV2w5Ys6pTmvCPHSZkc4V/J7IWcmWlnWk9raoOPTSogxcnuiGjqCN18xzT6eNwq3
8ns5cGQAaXNhl+7wWPLm7gkizhfmsyqLDYYGV9OxGRBfzym7Eac0LYLfptl1+BRf
wxs0J+z+i5a84DCm5Z9LhEa5BI+X3FJb3ObkP4OBvs2+LXasjLC65obRAr9gy31e
xG4OQqqpCRDL9ZWV/46UtzhYY3FEVyYE6bnD7oSOVrzM/xoQp95Zo9aKx4HtIJfZ
ApoKN7KxP/AvsmKBWTw/rQB5JefiJlwh7i+QYU1TqdiQpyNHVF7m2QC+hCkWB7jP
OO20quYmUJq5HKZhQ0/aRxCO/90XVkZhAXLcsBeuYBMvFe/DGRPHiv7PWQt6s8YN
2BrYcXBnWpFmlXwDOgDUpk7SckroA3NhbQ7IzrqYEJMBo4YZiIoILSZ0Madcaxfu
3Hyj2AcdOano+fY8BDWtgGPIe4f2hx/6g6VHDVn5mkroI1fOtUlG1K+nCx4BEuod
swbM2yHfZ9FEShtGmMxUh4vkZ3mDsz7jepQIC/dL6ljp3kwWcsAl/0FRv0OYQsN8
xVbMS9ZglmCl6eGi4oWsqiDqMR0SdNu7J92kmhREn7NwlN9aDyI1gBhz4RNX3rlo
KLypVT5ApYpdr7ui7gug0ob4nem2VH6HHKHl4ov/O2kki+HBGmnoQfCzZQHAf5LH
d+n9GhQoaCiyLb2OOsK94k+ou8w3SUAOBVCLH1L8iWxZ36Ng49E+88R85ehduHoa
/Ht0O2LPJsY3AOhtR+JtkI2z97TdX5lEe929qnogwLed94U2czlhdke0DK6Oejhq
XG2W8hVExon9WLwzk1v3r+9A5zBijxi7ywfWwxjyXFHL3AzepvzTozFLL5As04Sz
M/DCMWVWCVXqHWAvOJwsNtxqobQJyzknjCy3SJHjCo0j/fHwwRaETcCCk7m41M9B
5OqpcIxDp1Kj89dwh1ayMj5JbbNewOBGMYl3J4af2eI73ZPFsXjmSQvvd80Nlb/h
Pk5z9XL3BRNeHuloWNmW39uSBRo7br2dDnugUSrping/GMZZPLkF1VmYlm4weui7
eKc/r4mwr99iLgE/CMWVAsr2+/YY1gLkbW23KvY7rzEwi52H60C6c138cPY0sFF1
p4Av+lei+KjG9P68PpZZHUBGOk/a+Palrat8Lmg69+3SDowFa8TFNehI0ITLfxG7
r3ec85fAcDrZMo0EzqNUDKwB81v8UdNE6XS0py3NbnIHQQd5DLH4Xb+xf3+HpcJp
pk2hDVUfUNSzcchYNnstinaIHV4BNFWnwsevLBA2EkPkqoRiLBnVi6m+icF08ypX
VIAF1KpFUoP1QPt1dF/+qwR5DLlgoDA9wOMiEjWllx7aKdQs9PsvHNPpLvfu57fc
ZyQ8j79aAu0Ak3yTfzOjdxYGGdlXLcKGf4wcWrhQdIOwu9GbYJj5+X6SyefyMlzP
JMkTxzppvOwww2FrfO2dSLOt+UZL2ZclajSVTOt9u5R9V7zk9KbhdjBQkUu/WwGi
MFJY/jY89j4KhsPpJJajxYglJMjuanJYn8F5BMRWEAqupcGAloX5XGpVYPDq254v
lf1uwg4ax3fE6b+U3sFLVdKJk/OiMDsKPD+hq7vybQy8HHTFJ2mx3VAfzP3zGytd
MdgU5QoUvPPT3NhoBbAGqJ9Xz7GynktpFrrosYq7EPjsQvyxbK440L8sjtfPhEwh
VUmmnYaiJKoEWFkCpII5YaeaSkZjrN81mtoZSfXcY2biCEIRgZljade1iXXWrFjc
q038L1OxVskGxAwV7lWtg+ThNXvl2eb4LJ0JrqLsCxhXJ7shQm/6590FJuJi7oZx
snNq52j1CnAbQDHMTasFnF8jdZHR5uNJkIfzMTyEOIu98gp65aBB4jSwdzZl/Vgo
QQkIDMBy60kNf4sK9Hp7HGxsXxApCQPAV49X92QVmSUfeHFT6c2dYS37AxY0FAde
FKNAqDyujN66vbjisGqBv2ShYDYQfM30IgzXacAslsy3y6XlVw8eeLqAarQaxbru
fQRf+zad0edZozWNW6pJum+ZvKwExdZnxW8jpA8CedW3a+ramDXqxJRnAj5TYsZk
QQTyAeBmGcUibPgyq96lxzDl8xK4wO4Bl9m2Z16TK/LRP2NwChA+UOtyHVkzcYDh
1n/enrCoQIe11FgJFzXciSwWd/x/7JHAkUYf6o6760h9iuAa4YU438OrmF2MvXn8
FzyBijMZenQF5MjdXlBudJWyT2l4WC1DfPt8skK2eD8q+Q1hWvcJvqXd/kaHZDZw
2IGFUnIlv7af7bUs9yHweXFHaAo8GlMsVC88XGYF+7WyZXZJydfG9JZTyzjhOyjy
Okn+aXO0KBs0RLYH0P/6xxCMuvTHqTN4zT5efVvEmTAqtesLX5+SgmT1Q7Q2EdBC
1Afg4Ngc3HNhufw+M2Jro2d2cl/6cxPYYPexkex7EpcV1JtejmEr0sDY5oy7FeQf
9/oIU5c1NYilwoG5kz5GtrLTKLmTTCokEVaSsA1DwvFShurZAPu9JiBRx5nrhf7E
UoXg4PFZ/K1ZFlo+FqLm9laFVkdFDsH7wnQH3vxaNjke5Udht3LWcJxpDAGRX82/
+MWxV+U0cQ87CT8KTB/qpUCJ+gDNN0aV3uMxfjdAqR6ZTa3QyDbO2TKaJqBt1w6L
bOyyJdCi4jB0vqZ3M0zafLXt/oqspZkAF6Tv4/YHOjgCf+7gu1NUttNEOuP0werg
2ls1+1Dc6S2Yp1W/A3AcRwuY9AMiKj9dIZ04tYOvp0QkHzs+ey6jtJ9KKB31+t23
Wh/QXKOInwpUt+1+Rp7g0uHWJ9C1ND8lTSze9LHP0OoNnbKWm8Pky9sHmj7TkSIR
zxiuWSryiaOeU++UoXWBT64PrmhcVuyV2EQ7ISDf0xAtmQ5I7/mPGben9nzb+AFL
TBEc+uRsbA3k2AOCMqdTxQjSbxgf82vsNd8SQ+i+ILLcVYQzjdaIrjbJ+uFscbWX
wxIoHD0yunmcKOft4DW2SxG80It34uk6xpdwC+iXzZ0AKmo8FKsmWHhc2RnqRMDa
SiJradz1MFUdPfgqWUiufqpgXscNxFrHuiuJfjU3oaH3+OAHEpajZUDtvkZvcOP2
E93pdxTrtoYGo+vVSHnP32mGoTprzx7QAp0mZpOGikVq2JDffDtaK7R/+0jKHVpu
MLZYjubQVxKvXCdc9HZW6GzcnJ/WMKmSCkV4USmelxASZw5ESuu8uYeA+GI0f8Da
0cxcDA3aBWrU7tqLCJtQjM+ayDSsyZnf76/l+044CLdlgd+oh5wBIwNck8OSimme
0Mbhw67PJpkkKpK3FwtNsmeGf9GWQzAfxHB2kNgjimPzjmoTyOQYRKqMxbthhwgz
kNJmhSAm0Dj3JtQVJjPTXN+LSkEmxN/CGiOXxAkoT0gN0pCacZch+3PVaCW7aWY4
YhbfKeyUFIWj+t6Ye02o2k7GLm0w4VVygsLkxMjO+DlIHE35E86K46VIXErYqQ+O
WyUt7yUWYtjw+kd1ZeSmWWK2LP8rz7mA6DTyjiglK/6Kvh83cUhjCj3LXJmBmb7H
KqdJsOVMs9wAqI4m8ABwXjVeKhX+sqyxQj4nuyDgJJaUJwMdEkric5GBEcW43jPj
mdLp2z9pPswCYbub8YAg83IOMfqFQXTe2kk5tHFhYsueb2SGySatP/PKbDUkBUrA
v15TfvOKfo6uFJXx0R8qGLIxxq4/FiaBv6CKfMLoXNFcE8chIiqg4LckvBqstjsT
Ju7XdVsUCpyzmcLw8G5GRYRvVJKTkV5b3zA7jVGwACgVG2jfmQN7eHV/Tqe8Koxu
EqUBSRgyyncJfYNEAtt2jtu+NvM1SNW1RurbFzJF6f2QgE2NdlfWTrFCl2BeGG84
c6c4NJm7TmVfMEAf6vHOXwlAWCM65Cj0n9LOc33KeE8rdahSbAC6zvKoOXyZW6/o
6K1BFJ6Ap8CJWsugb7ltGt9Px+eBbCCbpw7GCKcWc7W7wJgYUvd4gCVhxG7UYaNC
nw+ae8Vip594KlNYgMQwL5c031os6ayEpD/or4Tb2yXo+ZWolboyHe/pML1XYONx
g1OWiir45PEeLxrI67mf9q4aWQFTTTqjBUX2doCGl6jlWYShfZ2WQUL7SMwy9k2u
I/J6Nuv6LHZn4TlypXLddRusSM4NZlcHb8xHTTA+ABeKel1ztCDHn2qGgGzNCKGH
lABwi5K20Fhwkb93NtFz76mGvgsaCR5Mx02j+TLiosnKZRoekI5Kc9sfRhpjcZa8
JuIs3ty9t16l5IFWgo06LN9f9k/gVkv+5rlbn3FlvAxZBnqZSIZe3HRIMH5AFSGW
cQr1Rv9dJdvQy6YgZFn45Z8h9NIELC/+NkLF59isRicJ3sbBVY/zx/irZzfSOqJM
kBEjzqzbejpF3+osyYoAzD87JOyoV2SFztd/h2cN1Z53yOV4/fXnnHQWB00Ohqt6
y2tg8TuRtT+66XqC+ek0+qCzhpDDhzgWJeDbpcA+AJi8nQbSZOn5HcdJJJhJ9EaF
3sXV1q+2z60ese1r5tbojnI3IlgwgcvP7SCzQLfjcMfSEF2wIxA2KsXNAIe3/9JY
pIuSUYDIApp8R7D3GkP8qIVkUNBzCN+mfVVNDdeVecSL/zNSGVad6g+JMPcJuhll
wNTCSZZdDkfMzUgx7GbPYnRNph7QulWbEiPMm+NsoZYLzuvFycNDKAW4ss/jio61
FUUaMvIIDRnAusUgB3z1jKwmpyx1klr8buW7FXBr/uVpo4dcdH1q8YDTl4SRgPcn
Hyys+Jj63ZLhOIIBRW2ULHrRgXL9r7+rkf1StwxfnCRjgqWdhXMHxYeSVixOEBzK
NW7+/0Kzm45e3m08ROoL7QXZJpc8p1+oQVGMhNVDOLFquTd59Rln/SRwWvBhByUG
XmRnG2oqCHIIEmJv3pj0uQMVcW6iM7XcT+jF0LBS4bjqiUaXQmXzMlfo4vF1ItRc
A4BXPbjPCTk24XZ7QL5/X+Horb6Kb8oEh9FJThtivw7cejCP5Y8jlm/tPS+dgGgk
MESzNGGgiAs9hoFg0euhtzy8VSNsL5ouUl0BaV53TJmAuGpcuNoS5AkD5hXspvX1
ukuIUkuRCI1+56F9WJxeAAHSGF1oUDdrz/3/wusW5IlwV9E2661yfrTKRDWMMyh4
dGZRS31vYx2cy+sjUSyJPfi6rH5PfLsyQvE2z35OJObcFVxcxhu/ddQ8q0xwpTdC
/ZInN0OGHG4YnZnRWJaz9/WDD269Oazq5ibBXaK49x/SoSe2xMd9M5bBA/uhcXGc
9poWaoDbc0QUX/dX2nk2wvJy+fNmahwDaA8SzcoEJZgEcyP8NiHCh/JM6yW7Gc+f
iSp2uUc3EXOPAa0+H1yL2WV8hqIrikAm247cBb5lKd/cueFXNLVH0TXh/D/JhDgJ
Tqex8hx1KYnGQpc+QMAh4/SlamXaldZdBEghrz8PvaSAG/1Jr5a+ZlN3nAh/KSJF
EJ84RQhA1qtpcVfHQxn9aX96S98KI+Kt44ZRsZTii0Wu4ctWKPjmaZ4BAePHsuNX
XehbiJw/qrIFft+fM/FOsDjqC48CiUP63fFWCoKWA6ksu/sewoEfsYHqELsiMQrP
LWqUnsvk49W0BBldC9qaW5Ez2k/6H14JqAXUrrxbw8RSAwcF6LvYdZ0CUVGPce+j
I+z7iGRdamqCn/EGRjBUBvt58DOxayfYxuCftugoqYuVgumdADeCLJwZ1+nBRYt2
eFBGYDDyG6hy6vFoZ1x+avgyIFj7oyQDZi4jnvSKzHLZzv+o4RkbJxRdecjnmoU+
ORZUVnzoUiza7UQ0S7Gjk2iVpkcQCN3wsw10z7uLxzQKtQL45o2WvAePgo/jRBZD
qcyWTfXr2q19USSZCF+IrE0QtSDt8KEG/1wpaVhI3diOCFrIspK9o1+8WoZiNyIv
QgjQH44EVgPPS9HT4fsPre0nol6X19ixJibyjVhoeiiNT/XXfyq/naUWsWnV9u2M
qGbZieEwtQOcb2ej7tuTO/QujvWeaKn277E6uKCpH9+20sBifvyFMw5asf/t9LqA
TvWFZti6IXXpOK8onTleAxZKFajYyoAGWXW+RW9V8LAgX8ZD5UczTTiYsB/AB2cb
sK9YXe2sT2cisuoVqdZOgXcIdgWwCOkzzn24Qm1e9B+tUJnZSlX6CZdEL446oBnV
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
lDP7/JwlYqU3T7FW/nQ/rqbX9XHjMeyswJILuEAlCyuv9ecSgnQKUgNvPocm3kLbXO5Zl3W9yNz4
n6pdB3ElompyDXrkzSzfDia7b+MXospwEHzJNHO2Z2yFRwiwKr1AtFD7YwL7nomuN968WznsQp0Z
fsmhNnpRz0EG3L+7qA2mRrBaHPe7H8HHgji+dcl0TOiv8tjTQEjUddGVhHoLQPSRbuni/Op6wLI0
qOYNSoK+0XLATwS5oYSmGHxkJDDCp+yQkM0J5REEa5l5NCHUFxvUEVkAJFoWvKgojuMdpr8W8oOs
k/IiRnJ0a1Vu0G+TMQWMyORWYob2axPvfhSdeA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 6128)
BxIX1O+Oyo+MbrURXbSKsFpR1wS8Lkkf6nP025SYyPalFwNlrBi6/oa+xMzs9kapkfDISwAzAWND
eRxagk6YObbTfay07V2Z4bgpmC7jGW6aUw2WHGYDCvYQS2fxA15p9OAgKNB6a7A3xx2Rni5RY+aE
NcJ6FRC1XVe3RktFWfr+3xXD0Ah9B2LijiwoyHowcQFby0F/tWnn5pAcuxMgT5mdAuL4AzbG7CR2
99zbsLE24NBwXpFj3rq5zgKApKYbGBTw/rY+RlfOUauXrDBc0c5iamoYguf/nIMAxlOalIrCWtA3
t7JYp44R5f4NfUwp5NJHQ1OW148Qs36p1ugYiojO4xFQcwvmmq9YJUGsk9vKrkNpsIGp+jB3krsr
kOZlyXyuXfpULKmGMQljPln0YHIXmSdLkBWEfVj+JWVbdZR6GDjln4TfQV5K8g5EGaIMJu1h6xkr
qBkP0gParuX8rNBFLJrdT9VSgZvi3GfHYBngCpstGznTJhi4iyQDAIIz0EqRZZ6Jpmb8j5AjJErC
mDoxcFG42Wi4SWgAm1Q3JwPKfWecFPwdSGQ7cN84YCmwPvjpPEyG2XnyF5bmG/pWGUReT09N5Jl7
DscjuZtj0FfPl60VcVJzycURqoWqj7UnubEZ0N0jUzlSxAO9dR+tSCs9y+bCnQkWErTBqSN5Ov4H
R/yzR9f9KlmVJaR2wG0o/mj7Gk/F/+wpZrvuwL6IKikQIiKnAQqvcoM9irZjB7rqTWeqegIuEobl
CTqlR8nllbgyuGk8JnWJCJP++jog6WiyXHNbAS5ZDKW+jC+YRI2gGqFKG1KArEjkrBMFGVZ4NqMW
+QneDm4rWwWeYnwVZJjtSEA3wYjjILZLrD/1AnwIwp1lOA3n3AKMar9B2dnfIN0I4Fc8+zSghgKJ
cwzBjgBCzb5NdY6g21oo1ZK4riNO9R6QHrTdq27j1b/m1EHHsfbPaex0hCFvVvZlkZIN6NmIB3IB
ZPkQmV+sHxja5X6Pv26gJbn0CleI7RN2hNfEIqCWAOleQKevUiDNveehTcUe47LNBQcxtGaVQrSI
YKIWbgmZ0oXBWSCLYEWYCy2tFoKfFfejiWrBhwyGJued8NoG7AUFlHM3SYTM3e4Fvj1Ad32XwlID
R5+wsYEUBcFUFMUqHaBbc6cWyc7nSJPulTTbr9Clxk/ZBss2xJ+7NctJtjyrisVcdBlj6DIjnMww
dlq8vuyV7znd6q7RDxUGxUs8KyVt4xNd5/XJDPas8FzfaVo8StWwHZF5LGw1j1ma6uLlTQieg5hm
yDe6RSwf5WifqqAPZeuOay9R8NJavPKJAzZ3t4SV71bjk59r72X6p7TBo63Yd4oldpyGrugUhdhD
/mHHG3xc5zfYJpd1qZBU2oeIPsaqvOkuCtxSx1iS5DOFre1pcO8WITghSaUhxHDTnWeCu2YG68yq
F/qa0wSSWQzXiYaH41jaYEu7iSyWU2rsm/MmxgXJbEhFKCTwcUQSsLTo8YQJ9WpCIlX3PYVHYqUZ
OWUmEQlX82Pg0DgTgKkX0t1smA9syrHX+FULlQy0CDKsyogP3fQbo5Kghnbm57/OjTZv2o0r4lxN
Vq8PSKfEJ7T/pgh6ZuLO1x1zydw/u5R4AjKeVccUWtwN18knRR/6Aj+RXuv2Xx9qTugnJrtClLWb
M9gdZC1El0oWPeONkbfZR5d0VBUDwnpK12bxXcF90ANJ1OkNchG1AOBalEIN9nWtIsX/j/IGOKbu
hWpvsZJ168FoTbzBKYiMPHGLkQ0pYEQjT6F58dO96+Hse6su8moBpYRhzrHd88XtXauOGjNAXbzl
E6FKSqlL4uyYtd2LmiayGPAuXK/Hz38hPSi/DNpG6RokOJqNE/Sbaz4s+DyZ8u1PXNJk/lmZWMp6
cgvHimiozKu27dWWH11GzfWZlpb0ugwDN9HuBNKDZfXmEcO3KFeFZv4zAekCcvWjQmabAByP6DNg
nAzTSzkOmH9+PHJrvd3QdaOXn/k+00BdrudlN/fmBSuK5BXECu0UKlhluPkob4vrC69ckClmDxUx
ZdJa+Ifdd1uQ+FJu4V+pIGn3zaRvie6k4XaSs5iAHubL7WhpzO+vmVbiF1Nrn+OW3K1+GZB1ohMv
C9BOq183V3OD7G1FPzBMvGEj/HrUSIxQ3tHMOjGQVF3DrjnX0/FkPgu966FzXqo/UGZ34aAu2lhp
DxLuqeBKSbxnmrYw9ZKeLxM+mhfG/fWhETApebmD6H9blWPnNWd9rWHt3700+7MQhuYHMIY/HdoR
ls5earbCWoPRdHksqAtLkRJtJty/lmgyDQkaYMpSI3TMOQo920U3l8/gUsoOgquQBZ0259FRq6ud
S0LuCQ5KZS3K/OdWK3NGlWpyKelbRk+goAPQQIGdWJiG8nZonLc8NqN6NM/CCju4C31MajfojzvF
N+qXDmRGgSkTEURvK2zhIC9zZtSTeCkfb1zm+4V583MmFySlaDAdzZbpuSsVaZeR9nw7zFoSmHE4
JmyO3SMLUzxKy/i7dhXFDPJKXFWxFHDME82sWKuUFCY6s4QmH+dIN+yfUfN9xnoBaCIErD6wgBYr
QiY7NH7ZKBTlz0dq9FoJRZv+5tZaUMS0Mu42bWJbzR7Dcs5M6a5b9Cjz1AuoPUyGMc8Est4VA9wL
Kl1LU74EQPQSu89n3gKWQmdrhxNsN+QRcpvZMMpzW2vjZRIdn4+E9anaTPL++udAGX4So+11VM7t
tvhgO/CggtkVYq77hgCW68Ak3ub1Szs7VAgrSyd7/ZSK3Ho5tXavv1K7PP2zb7GVqXUgUI1bcXYH
/WKPovTOQ6ccM8hTNbxzE4zOOunIhOyTqGoQDhgiL/vpH+AIgx/WPbzJ/uaUjI+DM8pZYlrh0Pc4
2K28WV7JbEq2cQyae6QUiGW93JLDZJ7VyiOK4zr2if/wA+JrtA0cNTI5WPNPC1WC97zXp4Z0+j6O
0n2gLzW593N555O/An66nRabP9O61Qk/XigM6krl1IhsTV7qiopJkd3xYHLggF4H7TbPwSSy4Eqg
KjRbxv7PkD5xE/ntuEoUUY68TmM5T7lia7EIaZq+kjN/3AIqhfrmgA01c0yziksGwwGzPP94xgrX
nj2Rn74aH210FaYNiUsgKt6LalAOdB+sEScheosKLpUjXzdrwVBQEXQNfCu3V/Mp4mwNhQgAtQ75
XM/yr3q31/4gItU00U8NUsmqCYpMFfOGPZ3y+PNoJIEEqRD9o44vtmTD/QGcbO5CbOu/m5nxFcu+
tvLJ1EgJPKRM6JqRGwshM7uNzHWbD/3dEZX9hdle27ykL0X2/TgkXqkuI79unTlHirQ+LkXlX8yA
VvlILikAwKObuFnpD7aX4c1yR1CXXHr62+Gw9Lr6gaX72kEWXKtZGP577wru7aCyOW5Uoj/eSTt4
Sye5PjfUsRn4hxrc7upZ/hHojcubbnHmgfQp2tnxl+qwcvHbMAGH+vdk+/fa3uJZxlREocENGgW5
AsZAWtrfYY5Y8jvmShZzRYXa24JWc8IhbJHT1zpYx9tkEzOWp935i0igB9kJXLt5rV2p0kSml0VE
/U4hSyP3IH/DV4CYPiTLgqQejdKKWJ25kFw8c+YThX2gFIV1X2HPob+QT1cprq13eY7bvrI8cnby
rBHqlq6e6aq9Is/kmhCccSxJB5gOZveumoYUo6e8izbEBjulFftYRyRjKMCBGYcVfh7vk3PqwiOD
lkzjyNZveMEPZleevPdAHnQYiOtk+HQKPDp8SCAx5FMG7z0yv39ocl9fLN3GckcI2pbzUoBbo64g
aZ4KCJuTVmMk+2wwXu289wJCoWy++cD2uiECNvEf7Zszb3kJ1ol6PsxTpBEIcrlKgUz3jxjoGYjj
BIemMH+tCqsdmCV/1++8npovkcFFvF+VdJ5Ew1qdhdS1sgOcmrTZjzUATmA51c8mXgPpDn1ieU8z
mtZKi+tm04SnUK3oa2v0Derr27bAjYuxhYnY5Zn6XGOdQkwz+mnf/RVwwprImvweuwCx0fcPqKj1
rrU7xb4LmRH8hFf9o09PaAX8k5OHNIbTYDmYzNt/+rfI4dWX/6SnHHZ52KyKRDeUnAW9FxKaG9Yo
epFSQ62MuQV3lSrFgRMBgLip+qjPdjpEKobvEpN/7TrSSnp1ebys9lH/0yqM141y9+zT4iy0ge00
qYBlaqkhqtimlqIqFvYqhI5DLnqvuZnIO1Xn//+66Ygg9sBScntj7hLCrULn7vjUCTYdbrAUpqxO
Ua+zFVocPGWBO+UTXhzgI3QWA6yjSkMzYYSNJimyWKTzn0IU82oTam+YlNmAVGxexEfQ8JM+FUxB
j0L9b22IL3bqPaUgXocH31x0MSj/7ARc9lO/UV4tljfdjF2NzfU2Ta4PEkztkEcYZQwNU5eUlmS1
MngRhFWouIKwkAKZrRJXClfCfn7GA8cR/4NjtxRAYkZZr11lh7COAmHtzx2L7e/+KGAbqJRufj5M
ja9ig5P/KDFyP5fzKrgc5XHpi3QscCNP7mZx1F5tlPPkzaFd2+FTFJc/v79A1KowvmN5ySAzZla5
GAmY9NnOTKrEktlf9E02sb5/QkN+nPdF7StGjt4LOeN6R/L9FckbbyMqZlTmbO3/lw4o+yG+FTRH
14M6u33k2lmqHkjMopIienrKxXdMrOXsN63SmCKyS4CNHZ/zYZAD237s1L8+ltCMuf6KgIu4n5FG
zfOJqcedqeQd/X9lXCxzhTBbYb5Cqvne5c5TgNt7AjH7Lxiip+0wdqfJi5kLeFfKsAHtxTb+Tpxr
PF4G3ko2IAzwX8slHJO+ebsDJzxr8j+T3W6E0TS6S5KWNhs3tmBKCDbhSrFGKWSkTNNTespxpv5c
mmgJ020iFLmbkzuanSbwZ+pDwhBZgbjmqJCJ1xWVmB/AiB3k2wu1eDO+U4Ab2kFI5+dKZ3f8BzA1
hDc5KaiQwuP+fhuY8RP8yCv00vgMDRF+ygVTmKpFZA1XIFR+fqsuyAG4iLEKcIJqZTrQAyz5BxCc
NHFBzngbxZB91vv1roAfrN9PYC8Qf8PuEZwx9breWc9JkOa6AE0pDBjGgrm45gz2VKKSHWMl+2Jb
JB0I0QrS+/HT4glQ8uCCzKXRp5szdtmc9768sPTkAva7bIEfnWHooZQot0Ro+9kZFxRLcxGk6huj
E449vdLBbl9a5t5cW0BDFdZqGYdHB9it/TWpH0ryKjOxKwXzHiCWYGVzTCz1oOj8GJimUblsNGRO
kcFxIEwzTeaFyDnN4yIj4phzOTNi8LIHrMxgiK7SiWi709OT/wCF/OVBiy1kdnkKXPOniQA4dtMI
oKj/0Ocq2DHe1LG+c4bRHpLPfyYyAUSRcXQa1sfCSJVm+qC4q7XkDl6f/vPvNh/rKCidJFRLHL8B
enOSs4jgE1G2Zw+pdn5Eiu1+ue7gWPZyq1FMb152khKcyuaejqxIjLxzCV2T1EJkrfMPWhpe6C7H
FyxE1Tl1E2PqUq5UHp5xk5GzUqaXhyeZvp+6U8RurEvI9NFkxisQbJtOxEewRvq/poybNP5W6Axs
4dw6xeT/jpb382zVSGY7dFXLHdPKIn+UgydEyMrpW93Kh1vdMfe83NZyIbDb2x+HrZODsXH9ueS4
Noz06IFI52XCH0IgPnU+YfLvKI9YR0pRQ4/kE4f9a07bMM16Fd7zSO5q1KUp7TcnR/7e3LukRCQM
fU4CO42lOIx693RU4OaZGU2ydKMoaCkg3yBHv/XW2hFNKvPq1iVdIp8g7mmPOkvRYNDCPr4aMYVc
DKDjaDC6XIdbUDgmtC8rbzKHV3DhiuzR3QI+HBAkwewVXsEVRvjidgOiOzxvUxKs4wJUy9c45jkT
WWRsRv/tox8o/ivl+zNIWxdltrQmvRtY8sQzigEKe1oxHuXJWFoueenmNIs2Mqf+7BSuKsjKbcfV
9J/zCbZajewFX8tCTnAM827sQ8CeAMG8zTj5oY3GtZ5YR8hhjFZ/YLu80DxreQKBhr6O9urG0Vqu
cS1XQIIV/IulwQO0gVYJpbjXj0cg76M4c6IWTdXSjzLJF5Ckq/kNkpg+Ai7nHfxNSnvjRDn16qrD
LFq2Axauk/+Y9OjE7/nsmtUWIc1SDQmXVW0IhhoJDGOKdne0gwGbXiN1yxzFtsCYT1bXsIlZ0OLI
TT0pcPhvXh1cc941mVaA1cTm7ulb0490p0AyS2Qw8ip6uSWclYuBduH5pGOxcSPvbB2+FiW3pIAS
+zth3MTC16FyczY/nePxrTuI44Dwi1T2yip/qJJgb3OFb8v1iMeHixC2X5g4S5ZhGRKufo1VqSBT
Q2lAsDjloTVw9LDnM7kA2tjuXc/fk0kg7vkbrrsA3RbXpwud+L/YvEDu1msYMUDvMkYb6d3lRC23
br643mlFy9qX4Fhz1hPzGndhJrREQ9uoujkWeXHayP7Na50HOh+YC+/gB7tnt5pN6H/UMkl88bSZ
zGQtHpGO6Gru5CCwjAIR0qGL5g3cEwzjZ4034zIwHrIfJvuMCS/ez9ihRB5tZeyYc1OVQke8EqMy
hdYC0OkKy4fX/enWw/CGeWkRiB/Jzg22AkPMuw6+sdE7TvGnbDcrRrLtD8Nn1z1AyYsc3Smb753r
Y6SWgk8IUj73Eas5GsBva/hZfsbPvWIDXmBkvxSKVc4zYs+DA3WSA9NQU+FwnJMyt8VO7elY+9wb
sZG0M3Xbfp3eNcW/FCC2h1hVHxwW6rrzKajy1jEM4otNsiRALr7qKPAx0GxtabaebP30th55rXkS
x0f3B3zAc3o2FgJgHcU6s+DvGSJ6ckkUlBeIfWet9fVy3GWMaq9AM7A2hz0KtG4A8LBApOWT35fK
JwaDt2zlvJ8/y+nx5RElAuLZptijGak4iNNelnAynLnmxVfOoRvROe1VdBePYOmC2Ovlk0/2b0jz
dr2L8DOXQxkWs3om60NFCtfLATEDbJ+HdFA5pz+key4T8si8PlHe+LlQsGkgg5mJD/ZCbzHTAibP
488P0r/vCTMXTR1+03HNNzPMOiLuaOXgSACSxeVAk8HA/w2UFi7Ox7irgb9qa/lES7F6DT7E08e+
yZX+N1yrk58CyViuGTYdcZrQtYlGM1IFdvFUs6wHaTnZzPut7OKJS2+NyLvTNZSNGyB2FPYlx0hB
esiN4k0M+Viz40i/T8qNu4GIk9F6Gtmrq4QSVICDYw5yEthwdva/4WD7pYIpvqwHJm1uECWw/nNJ
/d7lkCjgvGhSMYiSNyVfBqoYM0KTrhVzJAHcNqZ5enT9w++1XBp7+cXppANd7byLuTPyeKZIQBKc
Gng4J+hX1Wpn6Ce2b92XuCLuGLK1THFLhY2LDy0IcI+5RB+AtEAYVly2NR8xxCCB65OwASiDMwLC
DsCr1crA+y/8ISrgwF1LsXWtdTR1ekoBq6uwju+zzKIXnoH+kBpxHctQi7VIx8c7LT6UgPyZPkMb
fKT+/ZsCe9D2cB5GqGZsmW+UY+VgInzISiS1vtmu4VnLw9NnILNrIc8hP12QJPpFmswyadCJyEoH
VWW/EmANAHAEKHdC9QZ8NSjMUn5fqeOtcXD1679467uQ/ldjjkD+4D+u+DRndp7msODWvgStV6RT
Nej1oomubt+aDRmcOToDdKxmZe4UMPJnw3btVqDWPNYlABQSMsUzdLJEcLBmmVteDCYPxhGaDpf4
zxeq5Xds9x11bJlEQiExCtcVnNbOZhl0ogBXmqyZIRxMK6q66aTYWrrI8QqZ+ji+hLYpt1Qno5Dj
ZnofWokxae6PGRROgNIpMChZ8OKDtou7xbBTSUfP8wagx9hrIzZ7WuJiOanLW2xW0kEQrsbFRhq/
KCXOdGeaskWPyo4p/h30MH+Bw/4NXfGFSvj+DZG6PmUxFLWR7QPgYxWHbmPfbqxZsep3B+IOYBqC
9wf4fYctxgY/26XrxX1+pWBAPbnpHfcuzmAapBGaGgU4Wmb98g1xw67u55PGEtlZUrAda0sokvo2
dtiNIc+ZqshWHrsMr03eKbXtD2jg05Mo0dwwNxzXUivZC4rXtosp19DV6/3hwXHIGYoqXGBE33wx
F/cGIGdkz8RU1dhT/Uy6bh4zjkytJ/CFAVQdsnFK9ZvFSVTed49GYJ4XU4oLBESLfs3ArCJS+rK+
oQ4zGhYBmZkZzRm88AVqJGmcCZU6xElo5sXvrJs=
`pragma protect end_protected

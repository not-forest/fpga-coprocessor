`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bbdpf0Eh1X3B8nJfwnVSr4ybevsyJ9zUAhe4fLBrWGRuyYD0rVKCYA9ISnLZkvEy
hoCEaXM3KEi+1yScjPrDFTQUOs5OBFMNfS5Jd+muK4fR9XmqyYZkJSZF+00c0qOM
BTNOe1izTwTt/5zkgoAnd/leyCUBHWeCY/s673bLyUM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13712)
cOZTUgjS+1n5TJPW7F/wRYqpyhUwJBqOj0fmUe42vf5FA86R/NkeKef5zCy2E+86
4fYoISnw0gtPLw5E1FQ6g7k0QqTlpdFQb8OfRAzUSEJ+CdaX5LByAFl7YNDMBvtL
Rnp5o244d+GgIrj2GmX6I4edZOjVwCDg71Ojn1wLg4hpqUKvWaG0uy99w3WZXz0J
g/jthH6F7A4EALvvcH4Fl4e5NB9cPancZnfE7KZOEO5LZZCGlHF17mwq0qPSeG80
ZMOVqhwbEmPw21sGHe/iUjxu9BXTh1ashHyz9p/Qtd6xHm9w3DyQCoJLhebr11b8
/81oM0dMhfTdmMxxPPPO0roFOQ4kYPYz4AQnF2bzw0aeFB5be1CET548fZAuyL8h
GSWNdvwaNoeif6z3WydmgWLpinbhkBQT8IErQjzZd7X/4xczMBHX9DwxqNHkKjoD
rQHHByzwHSpGlQQhCt7/E696YRcepc3WqlWRBmjuHodSxwRc6B29MXww7R4+piWQ
kSacy2UzhY92LJ+s2BbobcMiUGG/T3oO7iS4NjTYIAcl6QW/dT07FrNALUiiNevl
T4z/irWB7gGrYfJiJgcN0RxD8c/apCUO4IvI5YIWRwaWS9/e3OGRYNMBZXgpQspY
7JEsySayu6q7DFbQwm0cP7WuiG3s33Ofa4+Od4GQYS2ac4NB5+ljkU46LMFyKRFk
ZSm0MWOtEI1ej8cm0FVB2zocJ0l1qLeV3hInoA7KM/LApsTJVUDTlCXdNOOSQh1x
guuNg2Czx9PeZPXv8DG2Gekple5UyJW4wK19yHq4M46QRr25I/qUDRe59xyx6qDm
755JQbYfGemRqDRyY09sGLQFWYw3tTgRbgUGR97VdZNB3svwNj4oRb2KO8KlpftH
eWoq7e9jKNkjxTvp5BPuHUlF++2KT9iTr7LKUS/j2TRY9G/CN4MCjMMmVQu9fioE
fSRex1Xe5fvqb9D8joTnVFA9VtUu30bcachCvRRbhgYTYh+bIvkh3w3VVkKU4TfP
Xh5iB21HHbADOUJV+TZjSkY/e5B28l2kWlYA/eEOUQJ+yG9iJOkF5FrEqlV9YPfp
nzjNJlIicfnD6S76deoYRR1drAJQ8La6H3YyTBMKRIxtBBCXCV5cu4siamsX91fE
upL25JL1Xa+fgImIDAymt+ezF2J5rPaWlA5yt94FbJQ3yCc5tsL5cEF7+FxMSG4H
u8QqAqZ6lm9OBfLUsH1Z6mtHB72j2JYrL6mBgI3xL62ed8gea3PtMmXCJuUEeUjb
533ynRBuDnxJgVUU8BDoT1BIO92RRxahE05p/LxRRE09ikz9aFEAsbzkxwNQKcV7
h0CiLF07ZVnoFBYP4U8KtzXF1QXlPImdXfMfIHRegh6wDB02Uztsxy0p9KNprYsj
DZSJjnDU98InSmN8Zk35rp3PnuUG3Z6Pkekje+i4huyqUeaLiN83vB5EM4cZrNsv
g4xlyB4FxzCMRKVF/XVsErUCWPIxWfenGgAY7YYJL1DkwPWJAVDS5IpEF1JYGkRJ
aJqLD/nPqe5CVB/D+R5d4XJH1h5c9QNPr88p+WNfPmAL5U2+yzWBIZj4lB9sLcIk
Y7tOuxB/sJGAmWRzoHniMx6yR0Rsu2DUSKKrK6U7BdWqwwMUoWq2zYxkgGWnWo4g
cLBeSxwGeQ/qtipOfG0ZR/3hZDfzRBCCScslH0otfqIgT02s6x70OGpTA+mD9t0k
BnZgEhOT7EKvG+0ZroriqrfVYpI/+wU/fVCZSj/PWvTwy/zbnIbz+JgayE/tk0UU
CK4Xq7GzBTN6CYfdD5+KjXqAjl6NprGdzrRcIUOOY7Ai1ENhVUX+d/lG8VkTdH77
Segov7UE1qa+PtBZ6xrpqhEtPm834mvUjipLEniknvocCEJQFUJ8Sz2IloDXK6D0
/6Nbm/OTcgQBBpTf10K4EkTeuldXu2e4TEJxiSU8TYb4DD4swl5tBD/xJ+pXOnOe
pLR5m6H+c3UO1M7MZp5NQ6t8tDAZ++eVqHHMxWfUuBPkcALD1t8AM/qaxTbfPLsY
irjsmoYiYAgQT1IzkD8xDZquVCEXbKk22iXvfcWA0m8tozLwag2mkr02UYVhgGK9
1x3dSBX6I5iDKotnrwFmXDebUCexNZIAsmnAl2c+cT6/kMqeqy247cO0bw566Ug0
oxYo114QuRvC69YX84/28n1bahop2gOfKFzIAMn6J7FIC0JILD4gaJgfMHX/I7Ql
gQA2Yhb3z5TWWjb5PN19CLYeQoN+5priHhkV3J3E5wHk6QHTis+gbey1BrpxTAVk
J5mSroubjbN+fX/HW4nFtonzlx0kS1jCbDGX9yEB9uWBTH9fnOxPDt6vlSRagyIP
cucCGMf6zo0oEHgYYbeu22HmYDRgfY0xgTCKUSKU9YEeo173C6Bx8MQMYo+zMZrJ
TmPKvJ5/5B70iJkxBEt4uGiBlKFdmHXQTOvl7TBx7IDo5yGCsuuEPuuDHFk0o28m
N/Z+OUVwbh3kOK9B5/o9o/HtZ25UtdMzjl3hZQKXJMwqNxrPjdzuGEv3yREIStsq
COCT9CFWqgnrWN4o/GvfP+w/kn9cZHSnYEfuX1uTEz3JCv9j8KXesOPF5PSmROE0
50yjwCFEUwnIN+B4qsgZrVZUJQu6KSQOWWtTJl8AIwpxrgCnAKxiboIsW/AczCMJ
eM7gu2+FMNzrVZ3A1YxV8OaDd2CrhQVzs+gZ7PI/VG5wRvEBjBn2MDeSnGY8jrzI
RptCMdw6OD+fe6GTgutcFjRgjLbnoQGQENzfPoTXM5Jp8YF4ZaZfdPU/qguN+95L
fV5O+HmE4efch1PN2CBKm3XjrBXBp4o1mUso0DMRmJdc3YYNcMKrgV/95bni5fie
Zo6Q5haPakrj+2tzHr04VlIV/CBJRGMQBG/A3mD0id/5BLSX8QzcyDnDhGhhCA9/
+E7IG2pespF6qwC3RRBkDoMN4+HnhU/jvbGHqhBwGkS1HsLfu/gRAJ4/F36y1LXD
p0NAXzvMCINWCeaEz+rS2Wq0XUhLDBBI11rz30HigzmrTCnokzLY8IFaMnMLlq7j
vtrC1gn7j64gyu0ni2WlakdFDShAfujGWf3ms+MPrvm7d7WqH2OwzRF2AHLSNNTK
8FItNZOU/zqw+lRbnXGjNMb4pHjYf4j9nAANcgduVTfzvMUa3QEWQkmIgbd15LEG
cLJii56cTAo/p6omNty8ETaiSND7QcoUBWBvd7WLGz3jy0reWQwTQkYmf6ZWJK4i
flLtkfZTu4ie8uHrNZ3VuvrBXQeWACVcUHdYTtMl69UM2OpD4RWqN0+FFD/0KeAE
EsVZhICuvyAX+jqopL7fyPQ+TtD3L4RVLMNALGYnR7LJS73Qu7vFuQk7AKUmfJ7T
gRMJy9G5UizKnyRwQLrKs2Q8/HYcUmCGyaS1ncTY539swUvDHQrKHrAOfKMLRoeY
1Bd7IN56Z5BwddoG3cdGGcT1NwRzmyT86yZfyM4oWqYc/9eYUQai7yAFQ1cJmmpY
ps2RvW1+RYf9s33KnyZu9+PS+0upfIczzH5ChzNYorqfWr0C23C87ICMwFdlh3Fu
W+/INqYSB+C7B7GDHgMx9CyXNbt3X9VXzOES5RdLuWSwNRZje4L8wbz+5emFnm9m
/wznFycj2lROiA68hC3vTn/cmfhSaB5TgbpZV8LSlndEWKjB2aoP6ED2sKmPHgyF
qGz9WCW2uu8Z2A08tqdUSry4aQYZhT1dacHGauEIpQx7Yb0wNBblVgMsI8qcrB1M
/riZydJwXDE5IEWnCKuDmvCdjvmQZphRgZFlN2/N4FR6NT0ETni36lUyXu3kx12B
ZRr7Nayy4EqlSIOy715Sz4hI97m6lMlZ68y8fM17Nurxqyhg2u/LtRKlbILwVR3x
Q1muy2lmWz+slgB1TK9ECKlcnSM6Vz/GwkpmY/Cvi5fw7LGGBXaRwga2pVQ0ED51
HE8RMxwcOSh389zjenqmuU8cdQWUy+WJ8hQk4zVBwGnKPP/fv0136qecHI6R/PHr
268HliCO6/DgJYC78e7bUnDNgMC7TJFMEtHmBhcSsLoBknCOC8jKzJS04LcWKvF8
PPbmcbFzSOZtau91GFyfXvbEohNL9WhDbqoTEYQpsAUcc/E3ezVwTPbKeSHRJiTH
JbXrb7qNNmU7OpqOBnlzhKEOiu2tDRT2E2RW2Uz4B/GnHtJZei+qo9Vmh5u3mnkO
3jfJUIsg2BfI4zqS44+p8q5tATC4LodVzxrgt7/D9TvanmDV0OC8W1hdF1pVp6li
yawcpiEOJUBxUStf6dbaVATDzyoY4N/gjDcG9/NiZ9IdLsFFl08rFCfVo/Vn0tOn
FamnkJxwInydH5hmVpPlRaxr8LZhHsIf0e0AgUo/0FTeLffAiHHark3uLUD+itdN
7YxX6RMwu+z5Vv3vYsHds6kohWZgcZcDK9z0W+VlUaBWcPcSUXe5lAMQqMjzyVAy
MrBLqQWEAkDRt9tfsxpA4FV/wo3E7kCMqzYrHqwLH6jCviGdnFjchGCYgJbfXWOI
4iYjLbz+Vq1bYOHou4d3a6aG1aDbcAJyAo2qABuJHj4h7sqY33Epr7pJuV47B3+W
Ff3Li00JnvtPklpj0ZvYbHMFMhqRXr2iMoQo+lT+IkgkjJ1kZSnRjQ96rTwm8+bA
rST+2IHm8hOYJJ6DVISqGGVIH4UlJK17G6g0bt5zyEc+Dpq55HxLWI2pR1j9aJTs
xd7aizyHTXZHHjFwU2207PE4GKTwHEVUZEUfVmZ5d9BhjtnNjwp30ZKnzYO0U8hN
18Kofhea1u4U2/rUKSp/2bgX6Y4GyOOrAIE3At1kO0Cmj4n/Av87hxGvRnlwj+WX
26jHHbQBhRZmr6Qb3+vUReqSblrDTpnk5t07cCbrIKVCi4ETsN1N/9DGGcoir9+p
26TLWgz15P2tXC3ER0kSoybnOeyAF0NTpvEwFpyET0QEt11HEH/mdUFN+QiMF2pP
xjkQ0QuQ6DCh/g2sLC3uuPNeKI27M4TOw9iDRTF7iVHIImIUWRc19kRLyrTHfrEW
ps0zImFvm9sO5VjLYyi6VYTCVvEZiHmnb6Z66ychqZRJV8w1xR0yMV4WsEHj5Qa8
xc+kC6WOAN3oTgcq8PuYHbQzKTu4BDTSNsdlrDr6Uz99yHHqy1OVHTfVwHZUImSC
HYjxen+mrXHlHAWVhsMVgcX2CPv9OluniheChx03L4F7e8SwQntYlsQwkow85xnL
XXKmlBc6+zSme/l2fEF4cCk5hN2cbC+144iUptjseKNRQxoFogkbyiZW+L05QglM
QVuKhonWHAFx8+UtgNy8h/facfOf4qpEL920JU5zKnVyuQi8lRMdRzHqi5HOhyn3
IBpH7/wNOGE/XkYIuQNSJTAKBr+/mhvS5jB39fkYpEQxoV9qWgUIhqKV7jUEiX3a
Io2pzsM9sNBhQ5kJhU+3D1dm0bdqbTi7st+ISnCPzeJUWgxkNQ/wwfYLx4UtcaCM
UfiPsRPC/mIiyN6HBdY89pVnHi8hTFXNudjW1sassgV8uufNvM+P9/iZ73c8bBuk
CUF9fTA+HM/jr8kc0jn5k+hloq1gbhrwlhVX3420sNnBSgpsKjr1cmmEEYitQVtm
catYpKDANZk72AG9ylGcjwKzsqkzT08UCFqAhXSzDk935bp38JQqgMUUZ39mI3WI
7fiA0JSOPaNbHcn4sjeUU/G5BNoKwNrdx9v5jD9oNZV6nEWNX9t+J2H8Lrk4NTkm
B5PzcL8VSFw7oh2hUHmENL2CSTGjQpbyHz5B1kYKKBeCcYCLp6PmliICA2t8SXZG
Tqz6NAPa/kSs8QPBwqpqORz7Hb3Xe9FGTT+ylGjWZRlfqQBa54MMjyZnx0ZeQzN2
QEoJje4p1BmDLV1qnU1N45hJpV4TCfKfyzzPMUdmyYUrW0B6o7Ff2YgctDAkm8Tf
+YZ1o0n9r7bq7jCCTvi6r3cAk2SwiYDmLOAcetSsqQW1cf6lWpc0zQrn6QP3JB2i
UizTUYIEBC5uevvq/WKrHHLHDWMepF+aiDUh/+b2CuU/JWTXuHihN8m5xL76UkNl
yKrjea3yxAviMsTHhLdpJlM8TuPCtlkf5my+iy3c1nHEETgNsALQCXxDHeJ6PgF8
yQyNXiMdGVr+hzjyxPZgGmEIwvRfg6mwQjcxH2V/OH7qd7bRyQwJsRtF8Wm7aC0V
9n59OgrOkI0Ba2QatXXwzb5Ooa4AoLLhPKXP66Io/LZxmzOWNCjhcW0mNLYuhToL
4rw7OMcejnr4NGIGOjHWTmaFf77olGtHxvXARDlEJLpBNZuUNojo9e13uVNe5Bac
elNR4F6ATeD1YtZ/ZJXe1KUlKmYpqBeN12b2oJND6A+MMSUyWZUoL+zeKWC7gGuA
WmOKbtwogrAqDi6BFBoPog3TbliQgZ5UNJZU/UxoQYmWfNANPHiPU9/PFjO2pi4F
fgYgk9kb+TULKqELn5vCVVy+BO2TvWHcLuW9OkVBn0QQ/x9LRrPudX4lhJGe79jF
+fup5CpkEsiJByZAMqsgrvYuhtEjpE+6ZayVDkxgiKl4SWt9g0myUegaN1qrGsV9
V/+PYW+WdFdQ4NTLn9AWgiHwSa5AWvyq9S/LBBsqF8TdbQAachCsJMWHXB1Bmd1O
z/zVChOSudg3A0KSflHdU0uff82e0UaG4Xkxz6sNYxlO0E7UJjs+m8TK/qpLByR6
6uGZvcTEW1ee/NZjN+lasLWp05jJXWuh92Zj3worrBzRmq3suExBLFBa2PnPPDFZ
SlrW9rO9fCb1GyXObBcQaMl3sxFMdCkAB7p1Cej9Nm3rXbeB0UBBWG1k9anVDMzx
ynLZZU7DrIT1QuxGivsyNTBrynwKY6zyNHo6KY7WQ7oviu+HkO0T3p3YhWnn2twD
/oSNxr+1geyNTWEZOxifegLz+8YCHTKzDAbBe6lo4dU+5Rr9MLh24Dnj7e48GBOW
TuJfU/muSPV+yeD9DV9WEFSnuuTIYsch0Q2ICgr+aqHX74gpdNuBybuyQu3au8jb
1nT5YoI5TQviCf2t4Bkh0OYj+hQ1fDEn5smF397kWuEf9iWrxJUoTObZKkB/a06v
wG2vnPD/8VyKApVgMwTuliPqtQyx5fSI+la4GAJ9sNiw2h0lPEJMQ7nmbdhBpUTV
wuFtj7rvTBOEyJshCVE5i10jVHhSo8FnnHsxYaYg6tbD/jK8Ms+Ip8wS04DlTwjq
ahlvX0n/vQiHto6xqh9fjpLm07OKSHGABDYaPP0aQQwQaONU3HYUciMr6hHESV0I
RdL5VQJYyx45719Ji8ihkpvtOZfJogj+B/hLajYyWH99nwwhJE+q4RirRDEagbzJ
fkJlMjmbg8JpvtcyEwXC93Xpx2iqPrKxunTOWMmh3z1SCzI817sXXqQAa4ipmjXL
NMJB98IVLVSUtSkADptrW1OmTN6Jz/V/v3hAvr8JbwlH8HRQH5RxAXVn8/5b546S
Vxeh9zeomEOL33hc2wXe+Abj6HbUfRSbwswxstb5qin3QrRmRyTrV0U3GXohKfeQ
44nifR0JChWMPEBTsNDh+FQnm5AscCu4SyNz3GywyUJycwyn/j1pes9div6bdQ5m
dyW6QPIyjxD9VLjv/2jGvNmLmyhUSMrohJhwIEiaSkKBCcGua4qllyOAltXh3HdN
WdMrTjg+p7WwzHCCvj2cBPETMZJdZkXphoErWzANeXapnEQLHNK32MBdzDb0QoDQ
misNuc7Ly3eHbhSvQnoDDTDiFEG9bCm/vpeCUErpmsmxsFRjtXgOZMMc+WMb/4d+
0FZwq+eLRZWt2VnsnS21/tPW9igQ6S3V2Rik3rREr5HoDAC5nVDsalqgFnXND7vH
I+8MGkuYtjVKiMbwpEjLNpgfPbGhuPo7YZlzGCDKYVg3StbXx8QRUaa3pDkZSEID
F9+LZK0rbfDeWrHPTwraMgLeTone4fIXdT+4w7ATAWSXNp0TxOKaxjnUOULbJq2T
esTkYkkRfJGfzjiZ2qFhUHf9DyBPgFlGmHDMaWObEKkzwSzGSx+V6OUfOoTnwjgD
gKK6LUuM7dChUbo9A0j7Bou/lSY6FaIzkUsIlVMa/B3lmCBZ7ZsyHOY0tb3fb/JV
s3CffyJkigBBG6aC9cK9YS2mWvjsAMf/LZL01wsU5zuYiJPkvhfYc0FFjeSRmuD/
rDwQCtK3ln940I1+YgEUffX9bpMv/YTKTI+RzY95iVEy+mRLfAPAmBXianFPmKi3
jzdn3SaHXBGaWGrrVw1aGUmnESLWgxwVDrNSbjAi0Fu+V7HA3fFQTK4e3MYJP3cV
dnIWpDqVD7HO62IvAdbadFw9+wp4cOYVKSIJbQAJ1+PkjgdwXvGexHe64sKiJhGC
0yfMd5SvfCYrbY1GanrPAzIqR3LYtyIepv/5qQHx3hBG4znYZqhFcZBSaVJVHUHh
MNP+FKoJ4xmF1FNIZBAmtwlTK5aFUuCfa1dWy+ehAfoXsmTpGDqHFEwDf6Bw25v7
rHsuBhGAZm8FVwqjOTQ9hj7fAWCiSIJrXIigGo0g9Glp+2zRoLgNdCtypLRCisCl
BQ2nLs/+8eF6gy8fPIwZSfzd6Yj5KWfGuSvG3cCioVo1S18H7f3mHP7rNcGicwz5
RVvnOadZeT9x/PWVUyAwbrz60OtYVjpD/a3OL4vh8OLd4nfDUjQvilWY4QEzZXvh
GcJJjfysqtcQ64LsqruKbsVKIQ1IwHPwr7WwGyyLDY4lAaHzSukOSYYAXcyjUSdF
yu+R7XFqAeJVtn4S4kJmTir4PQ/fo7uSGz+db4lsOvx8rb9xLbuaUkZSoHUrR2Og
kiO8NELDLI7n52vLFvxr72UPi0/t6uILiVPvVTCUnB6rLvpMmQ4/E7GDKI+g5one
DAmHCUC3pLMTS0KmXgAc3rLFkF0ut2oaTjcjfHkBFF80BQDqXlOyPWu+aZBTxCtH
RfhvQ1dILJ5SCqvk/WsbA6/pAizAfCiy6gNqF/b95A5Mj+8DRGkeb/MDnMX4/lTA
KIL6QW1OLYduQEGXODccbCCOY1JHR+p5UF0hyTQbjJOYPd8usY94RP9er7f3u3Jt
Xg5RReVAL0b7KQj/iJeWj0TY4Uj7q50ea2ker1wMqScg2WQoJjna/c+AeCjUWQwV
Po0zZIvNQt9bEzZd5qUBLgqIsb/xsICZK+ofUQfSTXmFGmXe9gE7a/sI/2PSmHDw
QDPzMUrPq6vfhlaRvMPrhm1hIGIdnOAmCGdeYS4LeQ2JKzSrJqAH2Q8tmqK4tJoN
I3IxGod05jbze+b5zndb6F9X58Bsba0toGT+xMxMocU2283nbXycGjRLYTBYHYz2
cWev2ym2SVYMFYopQ2je8UGr8sdlcR3cwop9d4pw7/m/1nnMdv8VxW58NdaoJAym
ROqvhqK4YBVdUHxatzinbcwHXAK5dfCJ1NeMSg9C9/j77AxnjaGgq36nX0umVklv
R0FaYJVkiMK0TFl2Vu+F/oCOMReQXXXi/c/pnwPorHOCInBXdeY1ye8+b2KCRTmQ
1Oy6LG4xPQHzWXNPR7EwTkseHpmzYL4JfQp6hH6+cPfY9jewDsRW3vwLrN0lXKys
0b7hzzo6arV785w99rzMWRDylwqiOkbhfZl6qQBRHr4o+xoPD8ZIpJD5TYyAyx8K
41t4s7/KfNG444zfZKx/v/vaN/9yBcG1/531ZNQscS+qB8a09/ybdmjSBCXCoZVj
jaDYM3CZTKLzSafgL/5kNTJ9hYoBhwsL+uIvqtl6refZjS7s4bGu7N/PxcmEum31
arvU8wxkYq5LlFcaWVXku7cp/V05GBeNwQh4I5gdUnb8RTGdSkwpgxrSdeCGeBhM
c6wS4HtNg79IC4xkD53d3cG0uuyU90xdWw5ivMny0Elu1QTERsMSsN2eqe3FqJxw
jlhzDUpB4FheKe+g7PGz+ljQ+/SOt8fjjrKNpDpyRWX2a2Buny19w74/CmbmBhW4
5yYmVZcxJtu/ZWfR9jmqPuGHeWCZfDSHK6KQOr0SbAXJwVJ5gfq6bE5TKMP9s7EQ
gQrAMncswLtwF0iLu3AP50zeMingherKV7L+8gY2pQ5P0Yn6DSFZ83q6OBG9e/Ei
zgc0wWaGGfaOOO4oW7tiq6fYnraIv+8takQmzBTmDXq8bufdR1bZN14XErvv48jr
CL+ElwmHfk7ebGY7qKYpc4baUq3DBAvAa7eQHyEX4+GY9Z+MqQ1A9mVMAl7niXIN
OM+TU/G9KULOcLWSajon77M+ek0p3aZBc0cjCFo0Stv/QTuvLFzSDLoDBc5EMLwA
Wa66ht6T1RgGSk1Ngy8haHvL9cFE7HssNSGJ3CVBGMxF7SbsOYJxLOJTlJjalrab
hZG9gr/bRBgKOfnD71RxHTJy4IKgf2QVEIzskiobmE5VPxEmL68bTSACcdD75nR+
hjuiEoEJ36/SR61BCKAfpf5fPirVyloO66zgJvoWuxTSZAW97lDMlWcieU8ppPIC
EKQkwOrtnuCYhTYkxnVbUpaqZPmF6vyhEImCQS3VQXOvnRvLRyH5fsMMYDySm/Bb
L1zVF49pKUwzWFk89Io6+nNQRRX554uKAjrHZ30US47JdTkXmpJG+4YbiP0uBRcV
f6sujOVHDIfXhXcMv+OHJBAtGwczCmYYNIub0I3/o46mVCJEM5UFM9W6v1fdvHYe
BEBnzXgtuxNKwKHcqzytbg/EYH2632Ro7BhjOLQKtlJ56I8t3BNL3hQ07O96BjTX
z4jsIUXdYmyDEDvCSJV4jDXoD5nniEr/RV9H6VXgiOw/uEsvTadrGq4kj13F8t/9
llcRJWmFUnQRlg6+MN8LsdXAIZvFIyvF6JgSVeRhl4LQmzBEzn3T3Sa8vLoLjM3N
xSZp1iuXdmELJvgQfbiwdfMrFC8b+naWqnC7HANe5xTiN0V17Sss7m5gVh+buEGo
oPjfbjyfVrAl0iCs+dB1dnvuEVoJt8BxMTeAvwj1ls95C+QSFw+dBHbnOBJM0uqU
vU5whv7Aoll9qi9iNmOK+H4uIjFCMOdkEnT4kbzjXxzq3ItjuqIld9bpo8vvbaIu
AC5EgE7r/ZDVAmYyKEb1l+i6kJpwWr8ELKoZmh1pe3Gr9uGhL0aUORPfxiRSCH4i
DGhc+I1e7k/20jSX5kMdn63dZZmSdeCHaRMMtxB/HMy8QBG5kCdIlWtoM/xQ0K1H
yO2+BDdiMzxsKe0AjJ6nu51S3H5NyAIz8HmbTsA0+3vXHjUzR5T5rAqbG2rs3BDU
Z+GNHBe4RfNQD9YHKhV53jVhs0U/V1TcEF5rrtUS6IILUYf70RGJXADlK8MFonpN
BXwFr/iRP2VctpXyFMS06423sR8K7RPucB8u/5FzG1ioeIEMVdQQZsAK9oO1oJAN
HwfGU8AlWHvj3oPBxKRgqLRNCWb0O9Xloy+QEdXdN7c1ZfQ3WTj5dDl+XV2cqYHv
6WrlSedmtVCmvqxiqsrFRZhGkspPhwXDCYT3iInJWHtdAXtjBfOG+ssF73XGygfy
Y98nuk+TA518oOw7sXR+lDtMLqsc/WCWU1P3j5GLDee9IeB7pxhQJUWWo+PXXQdk
LVsKUHvmJCFQH8l9HPqXMLXiO7Aki6yKWjOegB1xdHTw7zFaB9Hp2JCrIvILiOgk
dO/E+zoHlEVM3JxGLLBoz0SG2YHOzj75IPHf8oOVznkP7lwHqIdREVoBZouRPe0v
HtbKBJx6TZXk/nLTB63eY4UI4he+5kyACATBN2Ou0w5SuKDSHy8F0wW1PTVQBlAx
dLB0TCmNMmgkf6lnI5nPkcoMYHeu/lLNTByl5RfaAtLrQgYsJLQCWpRi6S0bHLvX
xlp3QzSbqBJdrBw/7SxA/ymJlECV+l65H0YswqqxNup9irwuR4HOyhH/BEauQHGi
kbLCwRcYo1UiklfuWPhRlXFuS9QepbwMq7xEqDKww6QnZUWUKiy+A+w96/ZMjjVs
Qqoiu6m0sSoKv31VFZ+Skca9QGcuMnMf9Bxj68etqhzhXGCR1jGGNV+4S6wbhhV2
5PG1FD8664MS6Kf90yYai+JLTh6IEbCUJFYh/G+HNN2tqKvULebbvX7g2JdoWK21
Q6lxwbFAfonG2j3WX3AqJxOlrVlVmnIARCOVcSJhu0nuqAZmQrrNo6+FBqRX66lQ
gcV1Sw+qbDCP/dCDwqDWfGQujYCxl0Qp1OsLKrVYcwFkGFUrkRL/Lxfx9B7HpQ7L
lrPE9c0rLKeu09J2X0ihkimZjvuHDUPDjFECYvN9ZJp9icU/05ucxiq6iXGBm940
ZS0kRKOqwL7MMH610fhYcXUKWpdZ7qASlORBYTXf6MDQwUszFwxzAbq2GTkdb5wL
YldNcfEyK1CWDFkYQzpGxRmM+xKqGEtxvifL4gYB8sS8HpAmwNItWJP25RntuEam
5BwNf37m5iNrjrfqFTeD1Ztqg2WjkVRpJDv8Gceop9ZWMrNb3bjqt7g0tjS2dw1w
twqZ/9nuXlYbj2/0DlwP+zIrBRz5ALRzK63hgAQoUWGcLhH0VSmbJxMRcdmPTqB/
L0Ssy4s+acjfYG/gw+yRs4LCzaYwD9eQjXgWa/hIWVzEFLGVbJTJJ3shMM0bKAVx
vtUUlh57C2TkCPI+/Y1saP/D4ZEOv1eICbuOFlVsFYbVf+4+yOdmVm3ILkgPryOo
adOxo/J9JDlV7CFCMLwecaZVU4qx4uzUHW71w2WzDeJ9UuUeCbqvuSCDmHqzZF3i
LrrZn9CFOatZZOmSBBmM0kFptxpzp7SnFwCTubhVZe6jYnGzcOGxhA6qVLLAXc7U
8xMgw60APv9aExyIdTBh7L/aQJADz37EoknAnuqg9Ls6XmQkpTW3UNBjZp3gaw54
fLAU3QwQxXd7hcrUAlYvbhap0rN6uuEWd/JRoFfCGGZs68cO6mS9QNuJV4zmIjpr
PaFFE4SSDIhVINBror4+BT7NJVpqFoqxEsV/6d6yc/d1Yu5FSeiXwfxCDQPS3+R4
SWzRn9A4viNiB2lusPiuUXU5eZQsTuq94XPKaXKJcj01kZpa+2XxGQVoqlh4zCTz
qBx7dBsfwkNfbS83UV8sc9CjQpN72IqOXCu5PPSZ8OMi1NmSIqBsqPEgU6Z8ZRof
dGuylVv8J9zgdwyXfP9UEz3c/BoDp3RweVxRwXgNIhtg/7ftC5MEVhG3ZzDThagD
IfwTbZUWOVAjvjMcJy4JF+sCuNLUCNAudDTthYaxLWb4EABeG3eC1ZItnH3B1EY5
At2jHFsNWdMYtJtsMXTQedYL47Fw5ZrC/6KEJ/TXIOic3HYhU6MMSyWjvAOziXM0
Pyhn5Uo/DAMY4vTMvENPdLYNeS5a1R3XPNxe3NsL8qHePUIc5vmvmC305MqralA8
EIJSyoYY4qEq6ukjVeUlkd/5HOd5om/3o7pPxII/pAZ3tvArFz1IjisIguqsqcoG
ffOyVdSMVnunPGQ76NKAGBSXCa87dryuNveNHbE9u1yfZY+lDXI+DOR7TGALh+7J
nPkBSVx7uRroUM2gHfjWf+jtz0BYlJ4el+kSxz7lAH7ulkywtOhm6fmYxhbnnsh1
5OzLt1qgliStvE26OtATmOzFNvGUlP+kornGLZvWKeYQDwXpUZtFhpA00o4V3TRl
XG7yYcLiCz3q4aYyaH8CcJqkSgruPMS0PSWcWzO15BkvdWsMfV5JtGavTQU8l2Ew
qzTC8TOoAH2OQCC3H8ivbbhZFW/5pJ2AmV8XoM7EMg3ks+Y+rnEE53yUiVMK9Pl+
qBBVL6W/4sv9oj8Qsw5o9zMehnRuxNK2LrgVAhmOFkJ5deQjo/L2eFGDfnPWiGZo
zTN1gjuidQfSfSHrLRmx7rgg4ifieSVPf6Qhqz/Sbson3FOgXEowyDCfjFTsXQIe
CSzLrzrWVhqcf6Q+6BEnk73sha8UTkVeL8kC3gfHi6lwUsk/0/L0PwcAbmzi/JNX
LUoNJccqVLuYQ5S29PIbHG6TTSssXWQTdjw0rXJVGWk2fPRMostheCs/Z0VK5vOe
TDBCN3aH1dab6f5UR3jEjbHoOQp/20mKzP2D/lBmiUx3GejxN0YWj/SVgqkP4+go
J353hW4o6Tare2H+5h13gF0jojRwK10pmN182fbt3Os9YuAIdRdaTAo6sjAlLwPM
skoU0FMJyPM3ZOoNs+In2tSEO9Ro5trtJdrs3Pt7SmJtWVqWo4g0et++I0qJqlh4
25IJL3EkPZ4N/hpZjgr1hfcqylnZjzUUHsTjGhjA6xYVBYNyLGyWzydPgmrqFgLE
xIH5Eef/9BIyYMAnrQWUHvv8fs9S4lWXPh8m3VLUarO9n5msvhC4oCEYZRnm6bMJ
gt+th9Ikf9DwB7Ccu53EoG5BciyeMwnNiRxbpTu2/Rxl5X9h2oNev3alzaKEL89t
4j/XXgiH2eSnk9F44TpQ/70OVkUjIqBwtEEEeD5zuJZrVw7gGKxeGSCwfrMTmVwj
CNOBGjBtdTtB9xJ/2PqYPw1ss7aZS47UfrGedacAQAajP3U6R7ATSQhjtH/oE5F3
mn5HDCmMBfkNlAkZ2YH0jkJMOqv8Ys/QcL5eEaBZT8ufyy42cpCCeW4HWNYgwgNV
Vj9Ezx4fPqRqZxSsvNog2GseBUju1bngDGGFsZBAZTaKAC1GxY6OG8U9K6h4gQm5
IHa9BXlr46hBfZwJxWdLFXVg4ClX0ijgfZeXZeNB8SEeZ4J6EjTavnS3bC5Pf7Z1
ODyh26Qm5fwwNsfrL45PrSFlIkPv7FDXMin2W0QLr0zczQEjPZn3QpZH+e5BCpJy
HEq9vSXzVAowj2o9U2IXcZWXOLoD3LJw+59b9oJaVChJAw9OkILgh5D42hNY/Flc
sm7r411AqJ8tEentW7B8ZnbrExJUvJ7fC4EVqlRt752koVqJMaiUXKDo7rMsDiWJ
ankVIZ0VOt5jicwl0P6gdWJUZ5pJfhxUpZlHbX3mmphbFF+u+GHCHHeA/38jHopq
bjbTmf4MiCaGRMs7XZO+a5RvJ1fdO02sdKuyHJ+qakFRjkDY29wa1U6DSQXIDOLm
fQaGqFutFl8bfUq5awglSSZqup0KLjsBxu/nUzuXPVkafiZw9AkS2a6P/U6a9xGt
8cmwktj2xiMvk6SY4NMFp6O7xJMdiL4M+SUUf1sJbDZhoTNct4BnjWNeVv7B/Dm0
qjTmH2Annb/j2ONaHWYeZ81MnSZc3QWXZtCBKft2YbmV+HJHmM5UaK/CMsOt8rT1
lFNUANKUg+WKby6YA46M7Swoz50J8zKZRsCrFQDGLz4I2mmoTTHV0XkB37J2+f8n
xJs1eAEpWiK1nFOdbVjiaVe70rals9VQ7i7aLqqHxUBuC+Vde8Bv/sfsDITrRFId
jfkOXuIa8YYHrmJwo1ggdsY2JQmtGo/9EAjPh5N1VsXh/SrAa1W0cvGUPbMIAccJ
KwG2f9vvYkYuXAdihi7+/LMPJ1161yHJbJK5pVJCfrg481A7oXFEZ+sc5iVfvjMs
SxVzUck4/LxQHXB7nuIsOB1W5cBaUUxOUDO6lXCTePaqLCq1z4lPoboXyRng/KWA
Q6PtOrZwX32ttG8ehQNMpj+cYYkvpZsJMKB3uLAMAfNe+ZppubO4UOHEoJqgrOHd
yYbK+Cfl8Z5yW8tG2Bhd47bbCiU0sYxRHRyI471vaJo+UVwxYtdFD0TiWBRq4Yh8
yme4pamQdGSXCc9Wm3AOonKp/Gyb0AhP/FSI+PJMfV2tnB9q3iMpjK6qHGjmHWW4
fjHVcmNUUJRD6uhd9u4q1ySpZ2ZMuqQnhTTgaXJqmn+0uHaJjQ+DvYG/jYMMz7BW
8bGEufHNB6Tw5tOP/1k/oEHTl6OhqPpriJrrvhb9AeLvfXEIUXcMqFs0to5A9ALJ
KE+7boNPr4PpNgoQSshdAmI3nlxFe1sJXhaix3b7280SevK7/WLfojdH+oQzobj2
4yptwxkucqkFAxunu8x5aLHG7+s3blEcFdGlk3+lPAbHUj/Mxp6bliRsOjlW09xj
XKTO2nsF/6dKjQ7st6KEELzNNnjfFABYRcZ038XL0p+igNPFhWNl1srMXluDPJbo
05axGdt6vN9LBt8cOMNFMNZjSoiA6+euqNx2H0HJxa6uli90+H+WhZdLN2eaE7m4
mmtRKxZAG4+nzEriuS1oBI2g2ur14k3Pgv9Np7iEyRizy1w7HjyDa06f/cZUZUPX
KlFe/zEm9yvbbGHQ/OCnTS1XgCE4o3u2VFtWz4cG1xxuMO/+VpNJyK4mUJ13n98y
aLGLyWiR2CaF0C7xM9LO0W8NuiyJYl/P9XupHuG9gFuqbt0HbiwfCGQb6k4f8FOG
t3c9bj/DcSI5M2p7wx5OoEj7bOVxVI0AFrOWudV11S1ptOapCHquLbvxw58bTBb9
CUnh6xSaE7gu56roAxBMfvDCmzbaCDydsckhzi9Z4tHI2XLh1ASeLjbPLpg3jTcE
uyN1qeRmWKVE70E58l3c4eEe+xzmGMRNP8mvpgKeLBSiojRk0nckjbcyK525zjnL
Hsi406x6L6Ilik6U2LOdH9AE9KS73apb9RmPi/jZrE7Y47u30hbO7x3nC6EYcqwD
sU+LcT5ve1O6hnwOnAE/KFzjM9d+7TwMFUeG23eeYlnduO89mXmXs+EHiMoDdk78
lKCGJ0SLI63UWtBshd0MKBvNoQ/WOpYh32n3/8BsP1cD5hCOsejj9WR7FLxxwFqf
LZEmx5yXK1WgJGaHXJt9hcURZDqNcVBAuDXSaHiWXkPwIAzvzo8QQXC8YWxYe4o8
zZvpCbp1w/7fv/dVlK2jahcK4ujM35/43u/JLMmkBFclLUB1uWjc/VVewvQFYTlF
dZFMWj0qOquqAvjKUPTlCAu6tHspPM1TfMmkDQKKDXjjvZG/TRQ0xSh7Lc3QU27s
virZTzxQSeU12KI5WaIiFmJEuQJftJ12AKM3mj7zJFdPBD91Kmgva6hHWLWuzTUS
Dn1A9QJIm50//hMnFjzj/L/HM0dWCTBbCoU0j70hhjlQoWxuuJVDuBUCntmeyZOj
sH+n1JVdbiZWRAtO33OdXp/wYorBEKQKHcuHQbxKz+D7/3k4s/t7f/QNTCSBNhMt
1W+bTO/xAVC7ER9sIQSnLBRLnyk+jZBERgOhvWCiXgIEZFIq8pv5pDuApRfV7CcA
fPGjIMFxRxEqFUtUSKfDKblkIjf0AXrSSejeH+Ukn9K0HgfH7tELw5Xft4ibO4cm
hPiQ+5clf7vMiaUUYA7vhMA4+3rnHOcBnD766NfkyneBUXKv2wYL6Xsl9TE69HFc
TAa6bqBbqM6g4HzU7wq2C/FJ8Ec0gF0wBLYqmE5fpw+P035Rr32o4QGywf2sP169
cr+FJfYFwCvg76aVJQjvr3+TVXJbws/zgdr8oHkrDktTOn3gGk/W4FWW6PvbPiaS
DFZVRwuUUAexOPnclgBQL6NOyLW7YYRj4AqMdLOUisG3J9w/LsuM6nVy9Lp4QSGj
TbAtxdA0Ywp651CvZ1YQZ37To52Y8kHtaRpORD++oQvsG+e0hbzkT8MJuETjbaoU
59SHiATbGnbOHU9MyEU/vAzVLyz6z00KPHsH1thbaWn2Li1slj+pEjOhJvP/S+Fr
eFreOdfA+85Nm7Dz/MPUBnxBzTXd5d1585i0Jjka4GzUK1pgYxNq086MEmMFbYsX
AKZAl/9u8fD412OW7SNoKvBHXnKrL1wCfol7t/L+x1EDo8eU0C+PeWBfFQnnuHws
rDdlhQsvp/CK+U4LKRmzKuJhiIOsHrWw9F2RskRh+dJxsVWPPe9Pq/qk8uOirTHr
/7bx7pPe1z/6zKdBvLGO2mCU71PNAbz7BYOiBCQGXI6qCajuvGvhIH0eDu7O0FVH
AiwPpTx0SgBBB6eDXFK4Rcmn6OmemziPcbOHJu7+ELOQv06mkp6nTDE6MbJfQxup
an7R05WDY90DjBB9y4qan1Dv+E1srpFcSNT/vn4922lqBZv4T1bHGJG9fzSNXko0
EAfdUGObd5isDCy+FGTAIXKCd63NAxFnHS2Gzs/BO1LkHPI1KpKtS622TPrpOcRt
ruGajvjugthSZXjZRSP5gB1h8XM1iw3LkdNaA+/51DvHgCVR/1BWx/bp2/iRXYP/
S+ERdyBKJEYXpx6gqojHyhe3giSuQTk5f5ZtHHj0BJ1iJhvzjR/dRnnQ0sQo+aVn
kmkKbG7CWWGrIn6Zm7xzA6rfOo4sF7b4KNOKcJkMJ4ag87AFuRJC3LvGMLB7lg95
dtrvTRqhxpW3oVTh3FKIhmu0JI1Yek5Sm4WaYTVQtsE=
`pragma protect end_protected

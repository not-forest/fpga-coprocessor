// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
cXr0KgsZccPU0opaf4rRvq7R9YU6JRaB2l/GtjD4waAz7CqsfRuEGv9qtuCYuVZ0
bAEkrQC6+QsucHbxQUCqva9aEx/6XPEQ/62Ih84+CII6zAZ+R9Ef6B5kWpAep2a3
EHBgC3V1uG7vk9+pvGsTQn/rb9uvP7/QzYLtZi9OBibXDnktdZPYMcxj91DqzKLW
pyhxLgIShpslwnkGqjL/EEiFtrOpVvzp4NwbVksJ9ILVqj5mtU2onK6RsNfrG/IM
gU13frWTzFCXnXcsItodnsMAJg9HYeC6DSPKlbIzVcd6ahQU4uKK7njtxkSHsbq7
qqf1TX7Rxl5x0aFxMdxY6w==
//pragma protect end_key_block
//pragma protect digest_block
6G8I5rkxUfbCseTF99ZXALIVsGo=
//pragma protect end_digest_block
//pragma protect data_block
jXj4IGAwJZdDlbcr6BEwXoQMy5Ctpo3q3Mut/gNp2Dvv7eIqGOV4Kq3v5vXzIuhn
BnMwYgtQbHHK92dYP5Sh12kxpffX9GrQpZ65/Fav4TfjbTOtvaCoCbxvfqRPpkcm
vngyC5XuazJK39mSmTigBnJxzphHYq4Kufwlrnuta5S+q63KjWECFA9IlGqSTYFN
lUdGiehQloMqYfp9+6yGHq8QfKt/Rgxa/EqLJtUPoGUMlyQlmG6Slhx2uKZL3RBM
bngc3IO6cBqgn32p6zbpRF2oGSdr1lJDMB8yDEF8OfQduGPpnjKDR2pUnp4KRIo5
hvZTyk0AECldRTT3K1opl/0mbMOadflKgfxdJ2vuslOTlZp4fvC4Mpba1QOtgizf
DbptC5gxVj6qfphCWjSfedUTaYwAALACYp7uuqZITEXv+cVyxeZXv0tJL7+5pzum
RYJkf9TPca7GNMmLQv+B/PQEBy1Mycf/e0vYRmSQzPbufpGgxBJJYummkeTfXVWL
CN/BS3+jahEV98ZhACu+oQ6KcXuthQX0Jd1R6E/oGA+VB2N/cbLHcTIyP6HaX4YX
//wXCyayaSaDbajdNngNE0Ph5JecWFk48assUZseY6RITZ0JYsmFbSTmNOH6Uadl
auF5ypO5TqL0ml85QhdkhhnPz1JDS5tIdwQ8Oh2cmUsJxsFq9rbePKzlo895cDOo
t7dPi535/lUyNrXdetzLd1s9yUAZoOfYI5ya5q+HnORUxgPFPoVeAJF4m4cjw5XN
WP3BomzVV5Y01s7D51luMh5/ulX4Sm4VGjGQqtLwX2Cv8Qk4e0kcRzN67LlH9FnV
x+J3vcXNBbDz6ganL1JV2BVkpx3dN1/IqGeWm8grnLPyIn/Kee5I0aDRyLKP+/IE
vWQy0M9Uhi94XMMieGiHMMzQgQrS4jfa5qhYm8j+PfmTQUxOZQSztoi9YPFV4Dw2
yV+U9CaGD/KD/if5QwKMaU6PzapGne3dYw9MMZFlmGVjIA05ZFpoIcKwGcKWIIJh
9R3i/5Y60TUc3beDHIokougkA731vFJVDhQAy2ooeFuOt22XTM2p8zvrqAXH1kg5
ZAaP3hLKFQ7l5HPGt2cVWz+oIQHuSA6hrvuyxrgjDISyIR1AETrT4UFkHbAjBAn6
JHKhKVc6mvY4hsG8mpU/wx7oHFvJzBU8MEgjFvsIeVzqsmqrynRtzmZdfzRqIfH3
908ha5C/UO/xH1sanMxEV+uwNgMiicuI0fWOBBlx9oV4+VWhOmkH/I3cyTlXbSjD
NXNX68VIecpBAUSoQgg0rym+wyHrnYb6NX7Zh6/1danfenZ32I3kjC5EMG0H3puV
0Ef+pL+8b2d77abWf+ry+G8wygiZGAjJmATWOfpOxIStMrSmVq8/tsj8RbgRsuWI
hEUCwEZtmu54vg+X5uOZVY8gJ8eIOtRj2u9w0VNJ+m5I8Gcl7N/05CYb0cvNGO4p
j2Ca7CGYq1vZUYdUMmpRWD26OCk/Y4z/XLE/F7jS6ojG2Qh5ki/eSZ+9s0cq7zyc
L/VLqLqJbq3GQZQ2ZCvqX7oKJfCSjnIbAC8AZUOKv6NBng2msW4WppisVcrp8f1d
HkZAfH/xOgOYPsHEYByxtSWjrlJjL+4nS6WJdAJKDz+lQe7xrnaCfEBKZB1J3h+s
dbhLcDpX3mn15kmzpPwGPNgxdcCxt3+ZvDfCUF8TkB1sS/hkd/6N+EWvslIDaTg3
2Wpq3q6EEFhh3E/IPDWOHcyMkuQPe0msjZkI3AxTkCq2fIbQTHBjFqexoe1PF9SC
gEwRuJlSf8jWIEpEPwmhovWqS203afdxJVua9iwD0JsKCMOnbqzhwR6IiYnLy7dM
zjr8pELCUnfIGFl8vvFoGo1TjsCZq40XhIULOuCvKf92NOpvQAYcq2OY+djTl4/X
9Dl3Uh0i8Lc5ZQdaSZmsstHj/7msFKWMOtmt0EfIjptEI84kV5/l785cw0UYiN3/
2K/15fOIPPwuoXYFHneQuEsPuFRh7Zb+5pu4xqRp3NrIEmaYeNw1JuCg9dTKLrLv
bAHuLEFpyHfQNhqu8ABUW+VDDaTbHFm06I7bwuOYci1w3WpH5+d7/kgH3L6OQhNL
DRHh4clK7WFLnxT7g/FkhoKsixwu1a+ufdo559mIwDzp/bsgMw/+JYmOH5gvNZYi
3kilPV599JrUNlKNKSGXgvhhB19QpRY7tb8hiJ6lOrlZVSRnJlGSBO80UcUsMGEj
0jrWKHQCE/afNTnFVr1TsWItNS1Bh6vUZUufWbcyRqyCXDOysYLPVIdmWl2cpjcW
5H8rBrJtWs7pP8tilCzMt4zD+EI5fQEShmvZFgssQ2wC/vkFto52f5GlnyqKIi7A
NJNr5HkB28Vd+bJHvVbwBzF10JYQV080EY66SUqupMO5tc71uBIW4nGt31n0Ecs7
/dCHzyl22FR2bqkmcjsZA5gaZXGbs/9Q15h003bzpNeKiOh9l0qIMqnhAz7xH/pX
7//N8UxyoUZ9VFUTAhQOm13FHbRzVw1O3Ietjk4D0eXGB9zkvSdk4/V80gzkT468
99waulgSFH6613f+OntjPnQCpgtjsUGFURdSD60JV+Ix3cCMx+rqyzvVcnUkvzxj
dna4/h/zgEp5RXhw77B3WGqQknkKtHC994jahrardyr3hAs5gEHySlxdrpH5ji+i
nJOgfRHLqCm3vmfMXTMvoYsqotV0YcshfUxbnqfkaHkR4kEHj9qFKVqIbQ+ibymn
ms6IKyRTk23Kfnye8JXOrNv0nifV5r2K/Y0w2fzu3llTVf9pcM7XSnWoZXHNpVDu
WjdlWihGBciZTkfFptyfWr3mmryIitJ3iWOl0wMxNss9JjV9TxP1ZwNKuzzrI0VS
P9lsv/xE/LSYmA33oIUex3NEgqXP/senKybTp0V+Ww6wxhYhjfgkilj8+r7tQC4X
1BD94B8UQ2RGCqP/FrxoU+4dnyDWnV5VUaodYgX3IPo2bkaIw8EW/YkwFkLGa6tR
751cwf3Dtel7yoYqRMs+OnH8Cd+WLG8MT6cpiYFUdN/L8licVA0TdoQTv9r8jFHG
L0at6RpdFvEci3UMDJ2SRa8fw04NvvquWmVAbpI0gSEn+VAZgXZYWAjmoJUtDiha
6IzO65e1tfKQeFRsN1YboBD1GyOM9TBTiHuuzGIHHcd1NEbYqQkmWCMjMf8zY6VB
qgxMK/rJgmDSuheoOQHKZB4k6e2mVUprusITjH4mLwR0qqNJwd6d0xE65w2w61jl
WOX8XPBN7TNXss0jf0x8gNw2S/u8c2xPr9X/O7M7YMxXYXi62borc0G8+/FnwN0t
ik3ftZcYBqaoTxdwAvklftRiXJqYhwM1f01YkHtwoZcGKYvn0YWlV+JcYL816EfO
o3U1gRDJoBtCZMlYCpSq6HqQDjTQsX8WGtqh2bkZmb7ek4Q6t4QtOQN19Z0tu9gy
XQGa9mGtffF3hZVqG+UootssByYUbKAdJJdXG54E97VPQFGGLJjQEzAi3aKxU3se
8Xc7R8rgJv63ys1b5a66Y6oCibEdb2GFbIoq+N4Qy7aJ3NEw8cRrbFXeND+spyNv
x+J9/59w1kohVWFvbW0New8WvCpZT7o3VVCQp1XMK4Fw033MvcNY+xGCtbDBnOZw
0ckJsOYGpeG9fd5rBuVE9cvHlSfIzkViJg/xlY78VfmUfROQdkaaFgAoROVdwhnc
Nfn1VqS3EKD/3wuUNLnyF2gZJfbbx/i6ZwapJURUH0D1LRlEdkYfod1b0MTDvGut
KcDUrvySkbZVHzKg2g4qY2fThKS0j1AJXReLbOU9rWF25ZBehfg0nwerTDBxr8e4
hXG+zbwQuT5gZZhqL6BJ3zPAwsp+zeB9OA1+0l6U85eqgQEQM+fyaO/N0JUnUgeJ
nAlP7Sn4Wvow3wiKTkUEys827Gn+ZtfNqoqI0Sdc8VJO0xhRHJQ2A/usCfaYa+it
QyySyDxg9JdSiH4+2wL+BZm72gTS9AlflP9Gw6iRxvw/+/ZSnCCba+ZipYZNz3oO
GUt+C+jGxsbjlO/je0WBLnYO4VFeGlgMR9T/qbklNOnOSmktSAHcjokguxTs+LjA
r8EHoTyAgAWJ1u+l+nlLKSf5c12cYHZKWHc7l+pYp99z96wKiiznR7r8sBeAgURM
s3yNTbWF6dqFeHY5JsFSmrqZj13ycwj1PnQa+8DxFYNOLa6jPeLIrxnWJfYzC78Y
NSyo1IF2x0DB/43k27B0xkkEBxe2uRvqq6ROzRv7P0vQLr2EdmArtHVtonf9JdxA
Q/LHVJ3DaG6hsYovbvMizEvdIA1iMjhV/mxkA2I274Slk5SsBHRBTbHAZ3WTPM/G
BGshjiJOjpowgv38d2ADzfcrsRGCTCFLhTfWz6tuiy2YKxaVOl9LYbtmm9ixxVTh
/GybJ7QZkM3ttHJp2yiTEOsbZ5chq1Z/3f9NN9FmzfOCbqNnZcADqomK3wGGG08l
vWFuUwAN8frKqu0knNSOAN1gawoDEbSGakY7Fx1P2zAEofOJpIAUF+UO8ScDUp/H
8QpHjLIlK+RXBAK3vuHq1tWrbBC+87lRw2wn7apCH/f/MQoALwJNEqCh9K9qLmv5
ShZHwmM2K2OC3sz+VOcjVBqKg+lrstRaDom7nxbHq6TcaoEzL0jepTQ1O3k+ffO8
ENmVbF8V534T1GvQpg8a+8TQB5x8xmC+lObQl8OZjeYp1qL0wQcRxwtSBURJp7Fq
tbbP+UXDycZcp8YVeQV/n9g6Yg75xgz+sLkZ/B23N9Ydr3BHD6UREqs9nuIdDQvS
aAHLA7kAdzBN/IlMa6y7cLbHWqjvBW+iif30sDb+P2aM6DRPtIbimRsW45EDACNw
ubTwG1ie8tyjtez6ZUwH2xcqf6Vwdgm+JJxvM7+sfnpeJFalJsuEkM6iNByNUZgR
RIawyFSREbpRjNJRj+yeVXy4feFbcsF2I9vD0SE0QgKzB7qswfwKdyydZmY6A4Ao
6O7m2Lt6tqbJhG0qV7LFE1gFvYVT2P6TnkaAebcDNT3duNqqVN6G4QtqnpsrjG+q
lrPHZUIxcmILAE9kzqUbSaw2VI9LcGvkP/zzninJSxf8nu+3Lmszsza0bPWphUHX
Chk4xb33D6ltU3DNRwXOGfmAFwXN4GG/6JrYAaaQPMAjfAH9sLzKWKLvIyiYTkVA
WeMkGthmoAVBWl1cADdlmnlqYxr7311O1eYSA1eLUq7JAXHRZLqj3HIVM0E/xtGD
RFd57rtPAKa8tPu+nBnCIym9OFZ8My5vi/m/NO1c8E1mcwDXjzac/HF7xFzmdyaR
5C/qg0zuwhcJ0lQszHAqN7Wz+daP50xHmvQ/wsuFOwxkCnIGHhFaThPNJvt5QGPF
J8ryD4gNxCyQ14kEQz7cMG5vjtlVkckzm0/5UP9TdPw7uD/quOeWrVf4Fa3QSII7
K6yHa2VxMF3v3mrbNNCM7gzJ2V87948vAdRT+lS14BUgNKi/y9dV0uUwDOapcExd
iKOXxwes55EpnIYV78BjEisbT6qN5CB2KGFVb/bzsiwB1Qq+XgE0EaadB+Q/G9px
XK3liAPxQuYuXV4y8M1HxSTYoWUrbFYrJzwZ0c54lfWX3T5VjfBVtJtn8sO/rjJf
Z/zReJtto6i+8elkHTRrov8vqINatWFv22cGvG/7eXz9vxMZYZeqvyuYJB556dnc
Uvc7X6kgxTiSU0ry/UC/EqJBtfI/rVahsE+Qgmf6b5i6bn81wQsHws6uhn2ciiC1
xEsMBuQq7rGAcVMHTOWzpt8GSKDSQuUFnSjk4coWfL/tGWCDOKxsC7NjPFwAOma2
akeUvZ8YuD0njT1UxGMqGrxekwZSd7PAarU+kOzUS0g/r40EPWuG9c1ikA6wZ9sX
bkaWt7B8p2Fc2Z81YJqh2+X2u2wqNGDvO8Prs2h3VzbAgYRAkrEvaQ1HzYOB8y2I
Zue2ZhET0pLN0xX1AS2Z0VG6RMkMfH7CG8nBVt4E79gpH4odQ6s5ShwbvLX+9vGd
ZT926g+DFOnHiT3Tak3NK2kdbQ0jyRgz5VR8GjV4kr0qD958aO1JqaHiNWT1QakA
cYI7LImR1F++UMGupl66NwCvLgApA/mjhimDStQ4KiHHFwH7a8ggP3hD3GsDMFgT
g6S0VJnBf+VgM5rGPaSm61Zt9PiK8A3I6JRbAQVG3+ZjXE7fop09VoYrkGGVSxt/
7oQW6u3NH11ZSi53fWLxKK7rTTGy6dPAgqCQnhPu3+WDVAbUTYFgquSWz6NK3naz
wiAPXj+J7507wKZCu2UHbIuMIIG6S3RNVF7WOOHv8uiyAc0RiD4NHlqhzhYa9C7L
mBXSDPALDXK+5CrNwSl3Spd66iqcrvwgn3uUvnr13ue7uGX1sBuM8HBjhSQCt0NF
luVRYttbiSSo3bQl/oGLOG1qSGizfqe1x/1m+hMlXcBgKmuVAA721HMroI/wBfxA
TMzz1OZjznecSzxSQ4V+xOLYGORGHKQDRACoRnpIkVv30fHGozhjw3BHahDnOZdP
ilGG7EmrTsqa2CZXW7mbPldBYYyGzgModpmJ6Eoq0XvLFetjc1kMmCSkX05eDqa7
OTyg52ls+VEbuuIihdPvr7TNWTgkh8/i1brO4G9wzx0DmvRc4O4rqSyDGJbmnW+G
tkCnpyWxMyRgLYjGWX1d4rHb9DV8iPW41jh4IJeu7fUAOfcFViJ1xyVWz5YDnPCZ
dPnbtyA9OigVQlU0HWNfh2EAbk5pJrQfcnpvnWMXbOPsbiQjTP+gJ25chXaa2lQz
Jfqv7u38qAOG3RTVH8JOtFGSTRHrzxbg6uFZQHk8h9PXHvtLojrxtKlZjDhdiLTV
2JaHrsP63mOZuXtI2vmRptrVyTkKBQ3A+loger9dOHSiDaycWCDP6pNYZOJpsj4i
9mpxaTud7de28/Rwgjz+u1Hutrg2H5S1uxA94oIwCRbrWf8hDnFavXO0jKm5FGKN
gbaMycLg7UmsY3j/L01TAsOixve86p1bpVkLoqs3ENFG7W2B6JEMJk/+1zSa7xC8
KzlN5nEVvZ/sKq0M9SoEyB4lTlHzppRphuE7DIY5xZcBSKE1bzCnk6L7aFNBnl2/
8Uhdn+1MOGPTkp+/F/EImF8NGU5ZJO05wA8PUgeEKKDGHPx9nskvw01vBCl2BoZO
LFTqITntuxFEXXJfOPwKARR6rd+KuYoBsBvQqlx0nDA50NfqLzSJYKrCTJXTHd/s
kMRoUMCkWlmCrCJYM86j/MdLHTCoBYY++HoUS1LdryAFCSPRTo+7VPE/bUcnpjMK
U29PmNtt72CAjhEqcYoV3ZiDQNYk9hDCBJCWj9kRIbQl8XdhbPRurv+lWDTtaH33
vH/lU44sC71wus1EmvBUcWUqDbhBsJ2CucbTzHgxGaiOpP57Hw8ujkMo65v4jlAp
AuOWsUaYk2wZ9dbZ4dQTaILrpBBqHwOKfpG1uT0c2CqKjxWV5nB92Q3T8rAdrra0
jxEMtJ5ZlJdCHgJxkYHjU7lonKkTAvysWTDptWQ6p7j/QnYIJeuNITb0RCaeVo6z
HJ29Nt/l6O6e3i62ZIdwA7m5QWHiiMhc0FzBDiGFRcVzXRnDk7ZgqMB4Ivmu/rE+
WeYazUePKyWBqXohhXIbkuCpwGI+G2A7dl6KJBQJ/O67+jEXMv5AT6q+JRWwjNdH
up2PxF/XE2yXo7tkYPAjHCkIMOgC4aAwdgrqGASBG3/ipYZ/Po8GHhv8zFAcmPN+
cZux2in8sSM6G+oU5NmiHOpYT+vh5p8Csfap3OdlYATAIQTunf2kx2w+plZmXppr
jZOWFSZVR2ax44IjU/2kDH9FtsrWbMHSmPJ9PwBKlDUvA6mE1LAVsg+rzUeoJ4Gg
boAx6u5T1vaOSKxz7htkujARJQ6LOKzEwOt5+jxs3RGFOwUmJqnZJt7iJosN2Jwk
dTzx7oUGK2L6yXl8QSVRKkGFdfAnysyPMUxMsBlKFCGKgDJgPP4ImqZdP7NBRRQw
ctLeVVL3QiN+3wwG5MfaGd9FjVQZaMfbq1I6YRenmiVauvDt2m56JQLbPUkdLvHd
wki6FLKSgHildUWxCvTGSdUd3TLNBRkDk6LTl9zwjk/1ZeY0x4wicnj9O2OWsZFA
0dlYZSG0T/VC5jkPG91l/IsZ/eDEB5RceACIbTXUij5DmYztRtTtrD4iGCgGj5pU
MirrvJWBTLcXCAy28jkDuw7Zhx+1VD+8ZEwJyi1uBUzb8kyQYN5logiETt8SBwC9
BGmTr1LFL0ouwHwE14CyJbzr/p5Tm7zhOf/9/SBpBBL6yx5h+9Ib2JUduAjpj4qN
nD9Xxv1ZYkcd/Tfxg6iHDOPtOfhnkMKr5H6B/zrTM2Q1io4K2m5xjof2Wq+FgGHH
1DHLMKhiECBMeqoA9k8fVnnRIEsyriwIcg6n4iUU/HKHSc32lryeFva+w+f+CP8H
/mU1q42aJm7IM1nOB5SCNGp2WsfdT0HnQFR+gcBCf9fWqIr7iXKx8ujX/MStFe1g
P5h8Xli7V+Zo5uud1HJF8PdiwkXmz+MXWkVRbEHZhPcGyg9XxZUXsJO2W8f4Oux7
KvZgpuL+qGqZPhhiclkaQudZvmDXrlMhAaJNawrMK8lmg9RrPL7lkyrPiOjgv3QF
kWz7laubOevudLO35Im9kIKoJzKlWbSlUualQgIRsph64mvRGnM1Trt8mrgSngEE
+Js6Gf1PsokICUrEfMeNKMSPH/soJx+ACKwGQ6fbxdUHQ6ZXgtiyaQ6WAE+2E9DR
MmWYv4Wp1zwy86gYozXhuL/XvyWtdDIKfP9zfeeN+5vOsOnNaJi9YAFO//lMtB7A
sXjZf5/uA05ejDAdM6f4m6ixtTbxTeqw0NB4pRIbnZCaK1VVqs3r8bizIQyTJosL
vnCdQ/7gNIJgeVhSa6Naj9SrLuEaGdKZoeRXGWiCqJkhq2KKUMW2ZG+y+7a8/Mr3
coXxL7IHIXjr1df3/7N5pw6walCinWUY9FMAyqiWY6z4ZkDEE5rYh0H5BbgBrPP5
HhJxyjkwqRzdpwqzPCYZf4aO88meZgRO1NqJssios3g6klxqdyLVy1mIm9EP6181
MQCv9yIcp3/YZ5nSAHBafqEtdG4mBlFzbBkJETA33W9ijBXs4xf04h3bJfWwhdFN
9SjaEl2hZxv04PjqyEIDQ8ph5jTGROkqE6auVHjNyJJPY5qhF6KQtWagimcXs9yD
s+b8sy8avbZkWv5TVjbVd+sxwCEQg9wTt+BII8y7Ys6HR/xlI94xfGMozzgsTESg
jsqJdgtuvOgYhbl4VWUw+mDUMbuq7k6Rw724wVl1twa57414KeEqEqvph0ErbqHb
ZTML3NJTjpPjz5G1SiH47R4AmitycddWOcug9hR2DcQbwDTUKPjax5veVFjj8UPw
JDhsfDe0aO5s9l5+6OQ4hdTAJfUbaH9RCh7VseYNQDs33rqmYSehbEFn4cXYT2q1
24GEzZvOP1fcghPazLjtFO8vBH6O8CQb1W2NAIuRHrAticqIV+RS3ZRLZGcCGodz
xgbagM6e6rXk7zmbhALHcwsdXaFgKHItVBSR6UyXRH7H+JD2VSfWoxM5Q8wVweLm
cCLmX3qVUww9/rq1aQq0SEugXxihbeVsj4FKDyP/Rky/chl1ilbUUUebu+Idnpy1
U/lfN2xbiS6Jg2GMT1pYR+bPWHWBXOZry4Ml2Db6lwG2xBqIemW41FFmWs7HiizA
dByjYLf6Oa0TRxN/b8xIznGPIPAopq66G1WrvZ++ldoIItiU7mKQ+7Z+9+2jMIJD
BRSmwHso0pMtVgx/Aza/5fJb9RgJMMJHkwTdRWdcKQOIUF/laLRp7M83y42hkU7f
hCU9GqNEUK6SJLl+C5SqbJgHe723I+G8HNRzJGnW2QSq2PniYLZKEumHaUW9VB/W
s6T2LxFF2568835VsvBDqWadoZzhvodPtsO8A3tfCpthnIipPbqoWAZbK02bfR4I
+kP7GHyqZUZlyCphHPIjtEDFYz2ANcXWsmZdmHqlbiW/s+F0RmTH1c0NkFWpeYE5
iPyr5LA6WaovuFqf2hIatz75aQVHiR3nE+BGUEdIu2+9tW2AFes2rDZf9zqTyVGb
3UoVd3Gct42PtmBYam++5KnYVTU67eFs5bpU5KAgXlLPrfNaX8O+yMHm6HqaMYZu
o3jhcYcQ9laFyJccX4lI9F1KliRzY6f/6kcZdlFpW+hHrqoEs7PFtsaW2H7AhOP0
+vAGs0bfyuY0aga8coBUmHP6gSyLGBFyYQwSQRaUxuY=
//pragma protect end_data_block
//pragma protect digest_block
/H0223HWb89pd8z380ZWFIGLIZU=
//pragma protect end_digest_block
//pragma protect end_protected

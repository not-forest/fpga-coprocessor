// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
oX965AAhw2X5pjSoZLJb6vv0X4tHq5Nx3+f6q17I9UznEmxiEn3wjp3i2jbmaUrV
LS5IB1z31oKJLboPC+UJP8OFwkjLmU1g0BoQ2eSBObU/tss7sepoYUX1MiA/87kK
1Kug78YQ23Dezb9f/h/rkLfMX3iIa05f9hSajWHNvY2CCJ8gL918JcsRjGMw7jdU
pyLonavL3/bReI3gdBItB8warfPFKo5riI1Ifh1wdOT5QqMU0K3lV70JENLuORu+
l4AAMgl3IWgkXZuLFTm6VuUbxZgOTmMUG0uYbHES+at9VNeeb/1BJbAai8lIFBoZ
fmlJ31w6GW5ondpQNUGbQQ==
//pragma protect end_key_block
//pragma protect digest_block
GcDRVHsXu4CUc+YVH1PJxRHi6hQ=
//pragma protect end_digest_block
//pragma protect data_block
eW6ZGoRwXWfu2fvQeu7pMVgSkJhRMmBdIdGiA3q0maWJjCx0Jwx/PcLKv7XbUXJ0
ZTJSMlN70wPgty7gEybn8LOZSROiM72zDZ14QP8jsWxj7R5/nr9itvJb1Xg9ine2
hqLB2cIqqdC6pg2iTUlom23gDrArkLiHZkKCft+fMntOpPTd0UwnyUwjgu+LTeS/
i0DP72v+aPOhndJvZ9hAsXm40FZExkotJ53c2zJgw5kRX9PW8d5QsN3MIsUBOWq9
w6v34YtG0Gx0QvoEqZ4/AAWazLz0bdGRhd++8T25LsmhigtVfQCZ8iYaVwNgjD/R
FhrwrfHz64/+/vMkpDVvydJBeXRMjVyxh6on/+AYFB8uP6JWhQ5SSRJnTG3fZk3l
vOg/23Pm7EBmiR0FE32nLgF487T+YVPbJIkpt3QMBRCenNunpgWhVLme6UEEFl+Q
mGWxqOzR5Ts07KsQ69x7uGgipd/4k9tDu6opdUZFuXBmCOH1qHpbHoVIEjSJtNG9
NT9+nAauUEqdIeTWsBH+iblBEJXLJUX/9cXgAZz76OZBPs+JOQI2oB0kyuKUbLA2
E8jfAZEFQHSB1i/d978toblBa4EBvzbylvgx3f2AZZqOXpXVFrkBMzMBws2oEa2B
ZX4Zft3lDXqlmV+KDx3yjG07YjoiL90fFtez85VFtam1S9vJg/veOWAl6Vu6NUte
2KU9g/6ajm1Sckt51EN7tE41Oc2f29XZE4bnSTFcDHzo3eL6A9ygMfmwTI+YQplU
x4XFNEsKQITd2AlNESowMG15pK0ZkEe7WHbVagT/JlypdnEtDGhPEJqV8uWWvyUL
XcpeHPlraikebJrzCFpzJbgYWgysYAisRbUqjINXWxzfNvHqi8GUJTjZW81dwAnu
124v+oZqQoRlgYnxdNymKefp6tDg1f1PFpwWRZH1JeZp1GcIkN+6CbxTCXhnwMkc
CaCfokRk0eSwS4cNZvyzyTcCpPJTmXRIem7bwdwVZzDv/Hb0gyNzMrWfpXQPb2S7
gIggoVzMgpv2jkpWMrjfeO/5FnddDIOZsJppHnRmPApXg2E7a4B6rDX4kSg2wEwC
k0HssVAaVgCnRxsnuVWpUnahPa1Mqng54HsDXZqUieKDvzqUdWrkgc8Ekw7qLkIF
q1hZZ+FtB3fTANH9tl169vLQWSRsyA5QCbG6dcZcbZjSeqMF9wQgNrghQVNi7ePJ
AQ6Dr67aafzl4rOw34QgNnZ1o4yOk3QDipsR6tSjJW/04OvBOOKUdj90kxOS+9ZF
y++G9/8hLQVXTCrSCacn+y4pvfAurE/EfbF4wHY0M1A529KMMcl0dRvfYWpMitn6
JtfNomhSU6cwUb32BeGgK9fmvcrDLUzm/2vufbAC4eswUhPctnr2uAbFNgffFtim
I1ZmS4NANtZ9ez3VEU//EmqnXojtNi3OzS6PMtlviKUxHKgMWgGN00fcwb0JweXC
xtor/DeQ91JLBejiwaakFZHLmC+po01YyJRETl2JAepe4G7Z+c+RwtxmI9dqTyXH
XMWfTu3773S5lF8i1JWWNyXtEfeSEGW6VgIZbVm14oRmvITFw4dxMGDjGvDob/g7
gMo/l9jqUIJMFdYlYR/6Nnrm/yjjLebdggCxfSbQHHV3vSlWC2K+ot2+25/qsSpc
3NKdZUM7gIwDIS33fPvxQibxskxq3f7Rd8f/y2Uz9iVwS+Lnbaox4YyMQDW0UFox
OaG5M0/V+z5HUHo+pGgKFhxs0hT/7qF5Gu8R7QcOy5Y/x0iO5QeDZBDjnTgR3a3h
fa/oBp2GREXnXSrGgAiQupk6U3kszaE3PsjqQeAOw91dVl1DDvi4xdlJj22TaZG6
9BNm8Lh0XA1DnRaZuAJTVUKxLLF2C8T1bv4+LyZfVPwgrIWP2eFD3CvrsmHEgYIB
z8clXyjqwTQtNga+YEjwfg3+U8WM71OdQ4cjPW7uwIgRjbQWyeFvQu94GIaPiMbu
Wm/acubZ2mXCvmdsgYuJLprmgWCErNIE8dwBuX6+ZtlkKvkRQFQk+RzxbBE6yErX
gVRtJZhJ0+1qu/zL4QqncJzD6I7i5Akde7nKrhKSfs3F1oxlyDv5R3vUZvl9IUZQ
76PzSoU3fAG0XVKSovWMNs558c2WpPoIL/cKumoBa8mtK30V+P90iKgBuWAG78vl
/Fywt2mDv1jCUI1oOerHpOcmsxfOCvwSq4konvsidp3q20eHmKhtGqU8cqKzEZtO
QI/XhqPksx7xSFkgdHo9Yd7HoHkN7tHzwqG2cni87Aly//BClohCCW9tToLfEutC
n5AaRY87qSfUw90kDwyp9J4u9A161inxjt6xvzx2eHCoS3DvxPY8KNJmZX/7/KvH
G2sTkwqQOYD2CjPgRwTgDwV5hinic2/QRADUlTZLef7L/4QHBYjQjs8ADpG9ER/b
zhvIbvvDFfh7rxenmyKMbIMsf6lKNVM7J157fNQ5+OoIXxncs3GqRGOiaEWnyaYu
8/AFIo9TxtJmLpakZV9x9BKrJ1sq9t9Q7WbPN13trRcOp3bSEYzvgfngfoaC+JVl
pPrBJTXgS17u0SzefEdcWjeSXdgsX6LNG7yMQp2cZM+uhmDlxgLs0rcY2sjBwFGQ
PsVEWbCUJSuHHo3yDQciO5cTI4yUiFJjOlVFf9AEHT4zNsTVdRZfIeYEFmMTxCD7
RhH9RoZF7Or9G/OWdCEjL5ZN4e/lNipk0OzXfDXMNKRRtqPjsCKl+QARPzh8DsVR
/WslILvHUn0dihW3HwyXgxip6qbjeCiWBtIYhPCP8QgAOsFmmsOTSuFiDHyZJ4yq
z6GXyCMGby3JZ2h/P25J2HMEi9z7cO8wQZn9EiwsPbfix+vGcCJ8Gi9xz2+r66nb
QNjFE7qQRgkdkqvRAst7IykFw0Ajis2TGNKK//zRXw7kYiLb24B+uQsY639VwIHv
fSL0Wjh91N1BeDjgcl9TH75LJxHXftb+2oYnLEzmTAwLOnD2yOf4ErChBg82OmaA
GPbAU2dJQaXGAYnR3qHo19/3RBGjn/BIKMlxvTQnrf8qGHA48L0c1IwOnPcleprp
di1EwgySh46axnm8tks4MSKreM12qraNaqa066oIZWn7bz02RQRZnVPHcNO240VH
FYW5pABsZmyNhpYZTDsTNdMgr7zx1/cCg6UXjdU/HHEswO0J++im/ux76zz/zI82
IHe+yEplUwwKOPMnBzaYMEJYgqMxHqQtHwJ7qoaH9aF7bPXpkDStNlVAs2hTbrpB
tH8NepnpR+EVhSd8CoJNK6zBYtcJlx1nPHAXf3npTzxe9T+wpS/cHqPw8s/Zpqr4
mBRo9u/feJ9SyZ0x2FQ9F+2LZGHyXYYOWl0vpPopF0Bsrw0B4sfy0sSrEp68+iIz
INBy8SlI+C77MUz+aeBHSecwRNNMAfHxyKQ38GQEy2kfYXkNkorg5YhNFggIWFxB
Kw53+hyIH4b83S5NHv2kD4tOW0r3Tiz2gpYvuxVYhRcFb9q+yB8tKfmsUR0LOp+X
SBWntSxhzgG658moAJOe3ygPwNqcB0FgJp6u/narqF9e/ubvLi8G6k2U7AoFFS9g
SkYialCRETScJRIKDixy1e6C4n4njJfWTBjYtadKRiuyRmkjYuvYOLCv+d9qvwjg
E+5jIU2zjODLB/zhzkRIucLXyrQlAn9jynGEpOHpCDwdKrugD8iN74kI5aaZnm36
v+8JdmSnHVj/svui5CQ7vG34TOsCsBqwV1FZNdF3TPiwC9urKinPT09fMxynlgjB
LK4FOSRE1rfbGVpUNKcwdSnv+nYDhbLLhm/gmJzEtZf4cvm1IpR6fKdchuYXLQny
jq282e2Vo8icorL1AuuqtoCf6y5pY1km9XDvye15mQ2eU2HajHE1Y4GBdF05wdci
8w4yVd55TmL+24WuEWHv7B65e6Z2ERPJgGgc2EoB0bfuzOEyUrONI0qeDrYPvRqW
YSkghuof3WVuzNuZIf5qWUPRcgCklgoTwdnkg4IrdxC+SgUWxmG77+ti8hw8R7Op
RQyfMORpBu51xLvlQAb6EkytOtoa+ryA4jeGHbNgZFwKzkClUNLKaMv+Dvnegr4y
2mfaUnsDeJvKhknQYauCH58xYR8kUmJ8KKwXtfd+3Sgk9h3EY7al+25ioyc5CeXj
9VQNomYRzxMuxoXDfsNY6n9seQR7KOvA0KYPV4as+94UqRKTAKzxr+rSjHiY//K8
DXtlBFTam7ej9JBl3GBFY/fRrPXfjbNEEQYYxSlkB4749ArcXupR1LSCw+iAmFUA
q31z3JBlxte0kihnGunetWEVQFDNrPrguFltGUU4/FOTybScXn/aKAUMNm9MCTyn
cf1z+aHfQ4eWqNRwteULq9KCcJBOJGMK8UesEM2PCaFuFUFHs1fx6h7Zk5Jl6qop
IGNXjJHliWLQSK/LWypkwZlF32dShSMWs2XZJr8qNb91XFeK3TcOxJm3dcSJ/TgS
jzwVtf5cJV2rpjemAJpOsDrYpUXGV5tomY+9fd+6HZWJTFNusG3Is5ATl/FFJBol
HDD8hKT8sN1sP4oGouJC5MOrJue6g0cv9ukFz5xpVo/Bb+3JOxgmtzh3k9AWHtgR
XHk6MSfvc19SnXkT0JXFS4mgv+IIF8RRtK3VWVEKp/kI5ggH6ojCW+u7Q66sx1dj
X5uqY5d3W75K14dNoQgviefauYjxawluJAckFsDvji+2nVlm+zNe0fAQlsT0YT1z
ksM92Tb+lZnkexPtC7oqlt9sG5jxV9BorF1EOUydIKgkJ+MOZwGrvklmM/2Ug2CX
vXJkk4A6mlVLiRFcagPZgiwlPfNXGF2k0+3UaD0n+8VFPp6MZ5g36egW2WmHpOU5
yOE8qaXJ0i2gBPvqRd8kkhIS38dMpIkuDNjjv+gaAN+sf6AmzBEm8tdrHFtFdKKK
ZWBNszwbpzJhENaCxdhRJp95BBt1fdr9UErQm+g+WSs/UPlY3ImT6qm6Z0ekc8w0
mSLLu53oJirTToVM/wzGkIuRmZd8Rbrx34OTENWWzSsHnlmCX6PE30MBZKU0UVi9
mk+pFozP1HNPq280iE9+Zj52c5VHm0PT4JOmskFG0WbJaR/zgTbHAneYo3FCCtGf
syERUjH83Ryq8m6mkQw1PMA228exUq/AhhSXPdAWFRCNyBVaFoTvORHyCPP1kT8A
r4iMNmjllqpzHa0qwJ3xx9ffJq+nqJ1grIXNST6Eb9GkmwxFARVPh5md/XOwIfeb
RUDA+AsUwxxr763InUNbCPKAvViYP50Lrnst7lD9fd/Ikwu/Y+Ukna7NLKDigrOy
cU6MYXU+yCgzcrm+/XC5INS9NCstIV/i+9VYAMXqAfXV7kIFuCKgP8Nizm9uXkyP
r9IUUp1s0+BzbsKwjnN+8ZhzlLlpJfVs7sVQfgo8YswVtggVKVYl2iwHldjHN/Hr
nWhqa/sqW0YMA8+i4dSYTu2qZYO09bOjq+WP2+2uf+0vbwluotgbYD6w1Afelcig
Cl2b3WxaTVkRaIOJXU+77DmnAKt385oFNuFShzS0o+u0+2xb5yvVhuO1DV0BgOUW
a6RHjm373gNfC+jhyjLG5KXh73s4Uq1ztKbR8Ia4ymC4EgXAZNt64V6+RNZ9cFPP
8D4TpwgMqjFQ1oPzrmHc6quvBzJ3pR34W8GJF5Heceu5xW1AHfGdLyQ4ouA2oGU3
7NLXvvv+n3Co9lro7b/534//qSpy9J1jfzjP9WFfYMWC60cQMgPNBhBGgzcSqASo
ZxNJ783EUU3yphZQjuXlSLsj/4ZDVOl9Ww8nkvxsEUKV+sLIgh4L9XYwLMrjeBZ2
kmR3w5lKkzjpLvaFzBdPvNuwWRbU10ttwP94fsEDRDE7NrfPc94XoVCAoJp2wrAt
j9aQDYxr3XDmnNb3b140KXotANnNaEDqTWuB3WGXqpf8uO00nQQw9CLqLjvnKW8F
jrrm3QNpbzmLZYrGrM5Fa8qTdaaCtfzWiwAjR+5XQvRUqn623Wfky4USdnLVc29z
DY677lIwUXUpKb6/pGXssflrVWe1Xm4q6uPYn3knaFqNHJuVBdRBAtMehQcwmm3i
h5mLWbnOJLYIID16tt9vbV3bqlHT9uy/iiK3sYkbWnqd+K+yM2SVzYmC9Ybir3vG
vj43owrPenEeLOU9XVjnssEp+BTXA1vP2vxo8R5v1tQtxzFzj/19zgCCBF33cfBg
EB7WXy2ecGUnHMBlynf43YcrHVWm7XuNtp6u6u066IzzPjH4FODANEMJXpHn6XGZ
DXpi+8zxz0G8sJXTtr52X3eK9gBhIdb6Uy+lnn0MvPbazE/pemtxOUGyhzE+K+Nu
Sg9CSll6cYuaY4qGTOprQ/OXtyzYHHz+CvHx78UJKV+8mLNYIVzDO8HDzJG/zNnf
DEBI+r5GOKkRTOV1ux7yEcIr5TtPhll5LM6EWaY6EnuQivJRNJg4AJ8aDaK6fD7z
3aKGVTpo+4IrScAsk/tQJ9iW/SP9yHjSebTNqf3ktrdbvk0/sY1hWVtWr01EI5yW
xVqVEGS1NWd5UzTMhZ6hG0muBDGZ99rqWVV9FHTIL10Ku8gtgjr4IcAps/FV8X/v
AenNfUQZKiSPc1gnKvDDr9fZVlPUeIYnqSY3HfPW6OJtdJwqiH0sKNgiSErMihjf
puwSD12jn8vw9IRwREtY1vGq+mH/zpewg2cIpUWpJlshwLxrdbS7CVifJ/3hLQGV
BBokyRVQAfBAWldTPZ1jU2biVrr0PXUe8BF3tP/d6iagN7HdnxnftgFO0lS2mCEA
IW7V+B1t/aF2TABhjgX35Z/zT+ssGZYYS0tSdDg0qy4yvvmaply7XIcXiR6iLkyS
VHKrXxh6KxKCkFTBRK8eeCYvBlKUfVuUqdkGWfM/cRgy92cWh9WiWsrO0OCNjoHx
lu+YO90Yp6pTQy4iG4kgPn3XPQp0UC1uEKn0pultaomyv+F8yuzn1mBJg/yRrss6
TRzFHlt+2HxSVU6oqWC92b30f8rgSwkRgUw5wYFY7rp4MVBeYXYfzKljq48cfTOC
NPpU4EEijMk4NqezzV2HRpRWOmLKN+uwaqXi1O1iPVwEx6+90QxoL1ZqDMjc6nd9
M/fqnlOSMGvlK5f4nhDUBvpCYMg+sPttsuJryoNWJLQRsBqg2+s+9YWvUhvqPFkh
uDCC7LO/rNRMdXZU2Bpkas1umDO+618XlAxDu/M8CgCOgYWVImkXxmZaweW0JG8V
svEextCPqHnvVedAu2Zmbnx1KZLeqW6BWtslsv2DWbzqdzJPFaSgcwq++tqTaXus
t1TOXAfQfOi/ycpDH2ERPk7JqQhecVZ6wHZKeIzQ2ewDSc18cNSM44lhFv/IGb/7
Uhep7FQxliEp6UK1O8GplJB7D71ArEVzwD8y+oXNZDa6Fu0baVRy159cAoIA5Iqz
Kzx4nWvydYxiAR4M8hz7DxxooeUBYt0EBYOlrSsethjLdkKS0HJyuTHXtbNpNYMz
hROYaVLTW0OkDs1bhqwzyJC/b5GtdSPViLhmfDE2NscH1ZLj4YObgQ2sjdgsAcQd
t4aJUii7vgSpDd9ql2MvDs5MgjO+xrhS6mfp6kdhVd/50BvgbyHQCBueIVi/Nhpd
NEiyYsRRtpEl6nmCVW7E1qUyQVAiKug2t/9N073LSDkD1kGTNEuKGVNS3KDOjboB
S3OqAJV2oJwH/2OLzyngLAhZF7c1UNxEtMDz2+GwTMGUPvJnNl+lnTp3qf0dn22d
EiuF+LAHzAOITDM7Yjxi3U9i+lNwTjOpU1+/7AGHD1GfHetoI4txUdDztVBa4Fmu
3rt9t8rKfv+LSR2GuWjmFpECFSjfCr3/L/HQZIW5Q4ZUTSwuuqKeHWD7f9qktarG
v3UfHRS2aB4IU/HpHBuzejmv9RMwKVWN9Pw6EE/dqb5SKP2NhmlER96rOEn63mRX
S59A/HEc3q0bsZvT5AQCWUdyyhQUTsrrwJUUl6yu5aGEwQae9eZYRJoUL2yzwcbu
0pX3H1wZW05WDcBZnQ92/6XgSLyueNJ/HtD8oNrojxOL5AUXhmehoy+toPcGvQSj
X3/ALFRGBnjtE0zrwQ44xnFpiSLqaVGWTI1up0dsjej2yow9Vdg3UC5FBSlBX9LW
c8PtdTNNGEKmBaphr9xiOHeUAZGd9puhTXHm0b4ZhStTUeDBhcRPivICWTlo5HG/
5Lvi0/vGImq3oMne/Fv2hcan1UlMmJhXx9LasEc3FbRo67IZvIiZ7b9ZCQXkfIhd
6hVJI461WTEwhqHERQlBPRroXmvf89czEGY313xFP62O7oG5JsWs0QBXgcJWQWws
f918zXUD8wC6UulPDE+havzIRRN7wMHLIFscc0B0c0wMH01OxqA0hQI+/U7w85dM
FMBOI3YApiqNM0EPq/lhjyAJnakdOzVyS/aL1Ghr0ovgN6b4Bn+NdnpUCb1j0hO+
HrpCkI8pJmh2Ft4x1T/AbEgc5c1BDUH3R8W7um+J/yhJplgfkeBQeEeXw0Oy+M3k
y2EIy/ufFqfDbDlBQvoIhzShYPgLYHLckjD94XqAIuOE7zDPNOhAAtcbqmUqWfJP
PuIRafKr1Z9wAER85sMHAD5kIZBM1Fl8hBL7Cu5kXEKxDRZzr04ERFygJtK45k5f
cXXHrime6x7+K3germ5ZDw8CwP0JFIqoNLMoMIC22LQNF8iWe3wTZBrHydUTFl0Y
WQPwuI1MEIus95coecqn79+ZmqtgNesdTF/ky7i/6jaH9PYZtpRXzUZBXGO4PTOq
ITKLmG0BQ3+toXQAr8CGv9mDkW4uhqUt1a4v+7fcZ3ngOaow6I/AC3vLZZEvuf66
R0hcWkDykcN7xy2J/59+kU2Y7mzflxGatGykHg+xBFIMzv8WCaq4grYFwaskhaSV
MePsMzD7SPSbYAtOthbghkQMMdwWl7gI57+A5EOUFeH1GVpvbWHcL1jHWgWRq5yy
cahdFV2jFvbnNM9nJZ+OOgq3qE8yjs9HcyZiPsUoU9HEzGUvwvXROy1ZwfEzjkti
GacrK2aMlerflQEbXt0xydYeFyWyZby2ReN9QA9vY3erwkNfXqYL5TO7OdVXORLJ
BAd9+3TapVawW6nzJvtRjxNlQ+JGcn9LkWo+TetcK83F38LFOkgZfKfH9F0QE88m
qc8YDMsRW8HS0zyVjWqIX8+SrpGck4NvW6cZe5q59dRhjEBARpCOr6WkY4x0k8Zu
swOXjJxTqnl4OATIgRDXvxMQ7UDQ4J4S+PbqxSEv9kPJy8lH6dvQu5u+OTra7Ldp
GpDMlLuuhLRWynWBpBLRgQ4p/cAmCwzi/3VylcQdDpdVVGXCnzIzqJL60k+8o+mc
yy4zJYJUWdrzFoMpuoXGGcYsOb9e5Av6I7Eha2qy+3F3AnMfMyi1gsNhzwVJj4Oq
OEx6QwSLcGzRguEnc6Zt7V2xhr0qfsZ4/AVX91zN8H/1PBlAX271WT7ofvOFrtis
7VxMGCkdGuQvFOVbslHule3GlHRLCsxXGHg3YvrE21uq+1m1GmMYMQ8urMiKtHUD
BVb5FJbpCAhouhADoKARppRk/auaRDSRWpnUigbcAjr/ExvZnsUI2zLPc1sMbx4P
Wd8JvxIpLbdR5yejywO5Cw/KGZtIx+Hw9rFeFwD0WOWLPS20oFbjHia8vvK2kbGv
LRVM2IcJqu7P5LeW30zMCjtrotDlCGxGKXbtH33rxzsF2w4HrlcUiB0AN0pK8wzg
ZQd82EN3L1AUu74vTJskuUHBitGve3yCmv/LksoYUfeR+tzJQ4ykWjsshmBuQtVb
7rdpT5hjCtoQIL+S3Bg4+qnzG1JfUlJuaSVRR7QsUM54bG97qGy9W+vi1/MTU/kQ
9yj2X1oUovknftmwzneTXoAsTFZHdjQG80pHxT/XeaCfNg22KzH4RkCK2LBZjLkp
z0j7NLDSyt+GIoMuIDimELuTz2a3xRqVer43AqubS6isizd6E3UJCrxCkePDe/IY
x+R0zA3OGm9BpxPUfV6Gp6eJHXEtJIxYpQsFReMCoGimB7vtIk+uYcLWUnOLyjsd
fiZPq0NLvjvKsF0sQya2tQDut/SZidYnSVCkbYL4EmCoQA3iQxSvweIF8yv8hpAd
XRYWvr1LlNbWtAt5hrNR4wV/BbJbuCaiMomXI7LwKiyn5V07awcBRsQowKwLKtdV
e+YoTmuLsc7Ga98TAtZF8i1rm/TOsvV4/23JmDsy8ZsbaJezVbbfxwQPWeS79txW
DvbzN5Bc/GDEMj7wLBNyyKweXsTYvwWDCxyuVE6R1rxot8//LrTaCggrMkt9agDu
DO/c1DnyGcFchuxKRIr/uJ5Unx/ntGv4SzZDJ7h+SfurfpbYgk28KSD9ebSaTjz3
MnBMFfk/KuCPPvHFVjnubsYg3FskdSkCxl+C9XWGZOc=
//pragma protect end_data_block
//pragma protect digest_block
KZ1mUW2jrWIF4JhiDEwddzBqTnc=
//pragma protect end_digest_block
//pragma protect end_protected

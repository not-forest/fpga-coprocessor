// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
YZLTWfl8i+oeLkEaXxOkvXhwE6QhGTCyn8UvrGAMTfyVl/nh0WoqYqiOtjZa6DkV
ysZBNxj8i/pxsx6r8pHObp5eZu1GUZfSui5h5S02NBJ740Lc6QgB+1FEl7t5wQDx
bpAKTM29hm8lV9aNF7XA66tgjtLTo7wvKcM03hn9Xow=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 13840 )
`pragma protect data_block
PY3iomlN/AcYrl1l72Ad+NVFKNQUOT4EUDSheX0+LTSf/jixyZacUSnFnOzoxDWH
Er7A1pv12xcWDHfZ07V0y4EG5klTy+IPZ+LCT4uQEDm5c6OKzU80qD8WUlA2L14y
kCYss+oORGzS4VLrLv+EbWE3r7tgDE4RcnEEXCbMfsjOERLaEPRknIZaW/j8MJcl
3FQsiAiuHge2D+4GVeNYi+ZWfvPvJP8rBiYR3ORQUHlp1/jCxe47w9bEJlksaIzS
+EUtMefbn5MJ4YcX4kMqpLhzLUVWhogcY9tOkQRL5z4vllMTaLd4YOaxU0KnOO9u
WixIhvRmaT/Kb+2IEnTp6iNVqFqP3v0IpwYzyflbHst32JJFfhizzM8SeVaPo6kO
HU7no1fS847xcFjWwp6ihGb//o7MuoAQdCkYseSOLHzr4GNaHsCDB8YUda0rfsYX
pgPal0DcKawdwal8z5EdQEqSm5qzOyggR3KZY4WbpuJazMd2dRtHsVjyW9tR7BWn
W5iaFJqQYQuK3kdKvOhOwcZiWvXLZ/k7cLT7g+/+4VkdDvagOAx+T4nTJShEDFur
2VQye5OrelW1/OD8Jy2htXZf8b3MreIxTeX/ld5ppFQlNaeRqYApmJFmBrdpDbXZ
lW8aGz9vuDHGBtf74xUBFEp6zgH11z6UJQcwG5ebhG9dacOVVzsefSmxy/iIB9Ig
iJgF7MoG03ySf28JTCJWwuK87lI+jb8iqWqf2k8dJ/VCLzgl5YAMhExKCzOjbGmu
pdCk3V32NHi1j2UabF83xzyrLMCwi1UV2ZH7Tr6BAKnLjP1Fi7kFghN48R9fJ95p
JV9YQ+CfXjb3QRyhDCf1hg+ZdtzOi7UAWs5NcY5iOnqiQSGN9pPWof2dZiHCT+2d
6/GyDNaT9GK6FIn80kd0RQF8EciouHOtT6EO1jXZIcEXwTSvxfzROkVA39CheaPx
bpIlKIHuGexDmvLD6/NiOQAXP/MoVzZjfMn13k6G0IDqD9Ja0l7TKmVmO9jNT7QX
hLy90/SHg8tWlXytf3LoJU6mDHzSNkcAGnNoN0T/RPlyY+pVfPzc/nCyrdSyiu5w
gJtTDGxfFO1m7NvKFpdjYai+fOJI+5HPM6DdZmEkFZ/7Bd9AMGIkUES9vF6lRBbd
r5yq3SKFapl2nvpeVCK99Pj8KwJZ3jblhkM5E4Q3OVWZ+Zeo+E3UdQBtJ2qqrKG1
98Kqty9ZNRM5W2Se2wqHBYfZMC5iMeJpwO8jiWWVJXndxgVqQOmuHpNwRiDO4rOq
SD8TB5OCzbXcLIoaNgtspJOvuDNNNYSlZQgYkVB1I5ISbP80kMn46NX58G9wz8dn
hcDI3tBNxC65DQ3Bmxlki41fa1d2wEHhBW84PO7Sts+1ggerdScCJ4VXjHMVTqWW
z3GULI02luUdT8UxX7heh8leVu2QueQXQ1d4WXfJ2goco2Q65ZiKXw/FdNfOFdKV
uaDRJpkBXqnUigG9/yPt3YhYxyKoRCW88W/uKhWFsWzANKdAr8rjK15SMg+KuKNb
PWIpD7JJXKj5Ud/TqYJWYNBRw8OHblIBxWJkcAN4Cjy/7kB+u8QRPwbKkyZmg6MF
lrNahp+mU4DZixDDH+ROWcSpNSUiHwVDVy+nz7otom27gBY7SnO3xaDDMyiuQjr4
08V9isTeYdeDT2Y2sAKhd2om63G5Vr8JeMUUgTsPDy2oE6pMgnzzdDjPKXyn7l71
Mh+nQbcC90dUQfOUhbLsC+S5QSfV8XLxxr0Y/nNM2JBGLb48MJpKz1rTAYk202Q9
u5ozUv7AblTEz9YSQQeU2fye1MF+qC42S3Qmlg0iAJTW+TNCtps6oLYZTfXgdAW7
KOXqwBVfaRsU0zoomGyOMLbXik6u2kYdNj9uuxwID7yqajgeV7ogSot9UF3Z0KZ5
NmNyowTseaeVESl2W/P5ByiO6ovK0uWcBmTKiXQ6TxOMMf7EP+H59liKvlW11Zw+
dZy/tXEAUkYa3iyquB38tqco2SC1NuGswxUnBJoPTnw1y7+ER0E83c8KYt3ZXIDj
8JZ5hp20z6Irmg5ipmAJjqlgMIzCjEieEAoeI4iwqDDhOa52M5KNtT9/9gasPukC
GZzllyC9c98mR3GkD5YN+T53OUX3ya0wp+mZpRNchU7e8+8YkCgnX4WPGPE3klRi
bOEIJV9ceK/FeEWvUcWse+Lmawlz4FTfEGBL6DY/1ljVpf0ianONsbbaJWyjXOnK
lDTaXvy42e/jNEeHWeIIfuBxvATPu7a50HOzJs3E1uoDA4+cBoy2nPZ7B8k5Q4G6
tuQyEMk5VkbqMW2qtWkmfPq53ZUrdAaIXv2p9KD0gyAiHlWwzNaM6+mPZAe47Lmk
gel+io0IgVKJTxZADorQ2ye0KqX+KL2iXyqzuhP8QsJaMJ6xbO8tHCv7pZ2EIIml
YS4TlfG8HfdxM07yEO1RILcY79+WmiUImEv4HUwLKKU8EL9FPOaAEQ5BebMO3knt
kvlf1HKEDF2YvPwwEFHxLbCDb7F24LCNZ1krPMSWS2iOQ3mphMqjFImt+YCaRKpi
hf16KpArGyDB4WGsFKibABx1QdUkYpNOUbUir4WdEL9iHyg8OAQLdssBl5GqTAmI
zGik7BLBI4w2QE+7Nj3fAtepojPS+2a9Wb/jjx9enu/5CAj1Tq1sjtCwu7m4Bd56
CGwBj7XLGg6Guwy1fQlMXjTLLh1qmPfI2u15ZdRhKEQrxzT8J9lVSUptQ3lYaBRn
t0SjYsVkEZG8zELWLxsYfwDXARYAH1PdadSOGRu+b9+ke+Sq/wD8C3ZXeiz9GQKH
tbz/B80/DZIeNXzX32QvOlMnvhfr8zYLH7Z8UrpODRdbBSfKqoR4oC/wd31GlawN
+d/jJGClchOW8GYWI7Xan0sRMVRT1o6+GNzp2IkTYLDqJtrCHb9y+gOvjUYEFyP6
DXX1ey1HhJ31s5xODovQP5PiShlKGgTcuxs8TIhu9vTqb+MEjYg41YYjPhGAD0EF
gggd7m8Rr2qsbDFDgX553gCNXgH/GebMMdMAlVZ0TvvHE5KVhESTMDFxNqIdT3kH
tqjMeSHyN0yjH2GilcDHXMV8g7FW1DxwXpNd98sk0sYSAa7lFeYS+rnRWCeRIktF
jOeH0eeuLau0tyU7YYzCwXD9nhUghhzgoImMRR+fey5ViCmMMeTe2HeL6Jr/RQ/6
fyRI/I+nT+VaG+H5zIj81R85WfTEtMoctUaprrOPs+0evcE+c4oBs/RF4r27aaGs
bGTxmHrII+3hAhi5vngRbCJO/y/JUZUVrm6VEzmDNT8TiGkaLdu7XKQ1IJik1+Zz
6iIRaw02SlZZrMayYvzqGEMtftcAfqFHZ6pcjdk0ry3UPk0oC+a0Pk0UAFyxAYLO
ssQvO0fe9A7CPok7EfRRWLsf3iVKuajxPy36xLrlRKTr7/emFgpAUHwoA9e2vxlx
gs91I4NZ76XMtJU4N39eWuXVfQJOeR9EspZ+h77g6sLRh1YiyHKamM4PZruBgIgT
+3L+WEzoDvhEO8v3roTCBPaNftwFEw78rYo+z2ztJCeti5BCcRNG3L0YFAZrb5Cj
Mxj+J9Jvwo2MgfQ8GKXQR3thcQ/D3RZFfeb0QZ1OCyi+T9lPv5X4o2+FMOTRsaGB
uyydeqZaTahQIwNJRmGDsNtRBWI2vMNooXo/XiPBQ97mVgL5h9vDgY0elnrI6DpG
kbnSahK1kemG6uP7RJPHAb7FcXsynp3f+2eDSSJ4/8Fl7mcX9+/JxiUGwbhUMcKb
RP6JrI8upGbUyHDykhCLZIK06r0D7BPy3Fpt5ee6Ed7Jrx0rV8FxWz3l7EXcewyS
eLI6q7rhNU26a13+sgzbKTuUbJ+kzZ3+BKeV/sKdtF2Y7gtorYnEZ5wpOtJIFpeu
GqVNaIMMrvW/4f9mp2ZHQFkQh9hwoGqAypNCLga146vuoWFALFuSlBQUXbf8Gi9h
zHnebPbWdaq5DrdnZR+Tvk1NFsHnvxbgj5eAaFwCj6ERXDQcSx6sPQkDsSVp7iQ5
Bq1X7meO9yDhBqRp5CzZh+4/OS1vFWU7C6RIFSMGqgOndLaAEnWhTDtltOoRGVQS
EC4Of0MThwclxrc09qxxAW4Th7C7HGk4KdbnvlxozzRFiT2EnxsDgDuW0xooVp1S
DO7ADb9iX3qXusJz66/fQ6JVt+0+LwhlBf1UJc1ujZyvD7qOnfCyChiCPhGHMh/5
UPsL4wBBtr1AQjKErPEzkPX6e+bZNkQg3dDja9owHHU3DJ1BsFjm1GwrTL0UWJht
R+9wTzEslMEwmLE+YXIN9pccyphJPJnDpA1gIKWTLZE7aGCn+QHUqXf+uIOLMPTe
BqErIYdWaVUL4HXKYoq3lXehd/w7AzMF/6XMrvjlmUs5dJuMi9prmJAWhLSgY1Bj
UDg5G7RqY2Gfbx+K4ATsF0vraX0uyp5wOMGuWk1Mt2b4eR5rVsF5HUPnzbWlFqZb
IwAVs7rMrLvCcWUe7+2NR3aH1OzntEO9VfTrnSRStWeQdS3WzixEesJ72cDUv967
stzFlo50LF4j20bOPtDO2E0y1GzIaJleS8aw/ZMfbEYivwVq3F/v1I3/fjVPZkBB
ihQyypvmjMvEjHdRYT/daq0c0Gq8sChiGH+WsI+Sii9xZJX+vlhJCniVMCG8HFi4
YT5TFjXAhcGXDXN0HKVaAPGVlfzE8zfEktFeddLnFClidDaDVnX/0ZwAQkag+1K5
+DlZYROEEHeAj8lGOL8m1oRC20ITmmDX0KKidZ57klSD0QtFwCuEWlKgs0JsWnR1
05kj78zzd3q1xSG/M8iEZ8ONZtgW7xXwDIPmwKc1k6fXd3cuaTjgbdYuPs+sMEVk
2Jw6oGFHYRnGlOjX28VnLkJ2zdPmo6/t2zMDAQ4Lb7X0iAh4pGKmho9RLZ7Nqr0y
+hW0PEtK9W38VQ/dPTeq4cXg23JQPoWsTv75pGOtA8QxD8BCc6/XVdjL49wODqgL
98TiiwByrHe+xsei5AzdjXssVJBDbn7wm+LmeIpldyRIRSVV+rJJxamyv6agZua2
SzngOy0BPyNj/iccVaCjzujdUUvmi5Tsro6NjEQ9WlyaoAdODbAGZGwhQiDabJLP
6CxchTVfV9bDRditQqrpc2CaMqlRAbtTTrcDccu70DsuGwdvSXNvlB07RYWKwQNH
DyDv2zLa+DxryN4hFslIoFbLvPAePjzn7GkzQ+cMyn4LErbR4Ng+VeRHSzU3AZHY
p46SZp7fIDOD07qg8Q3N48LUCy1aJq58rxXkfqNjmbgNCGcnhkOne4wUqlzhMllB
6QFtdJEBX2U1Qdt/S2SuzkTn9fDNyrNun1yeiIk5HxrXt5WNZMmSZb2B85v7ZDy5
3rk+0PjinnZVgC8K1q33mla2qglOYoZpoRfutWvN+uaC6aCcoR9/dtzBmMMGwasn
Wa380r5z2EGiapMYsrl81cA2YrBnZZcsFEgrp+y3MDGsbqt0W7j4hWQ+5zja/xAN
gUUh+kunGpx/aT24tVQWdWlLDgbN5a02hEC9MjCRsQRZOvRqP+Mh2UKXhKYt6dsX
a4ZO1bLiMhwVVA42djWPG9A+8TgF5+lnr1PUCq28pzcxc3bLki9AlEX9QrNCVs4o
WZfVDi3ORbJxid6z4P/5Vsoc/4TbSDMsynajEjcJ98NxiXSMFLiBogEpSCxvYzZ2
64qdVIeh7kGMF8KYs+7gQeEixQByKyaeUaJ8ZS2T9wOBPNwOv2ocboocqV5I6kUb
LxtmDbIqDzQhK+zTdMW1MqbSutJVmCUIe4+sbmnrRIJy1SAECAjPdjUvu0rHAV7V
kBqPbove0PXCd4ig3eMBB1TaxSOi3UKwv5sjOMwja8tszkTMAPzowkn8Eb5USn1c
ZHa7fvfwFt+2ymz4fXIkLbrRj+SbpAl5/ufq1hcq95pAkMAw7onzgGrBsd3BUJus
IxGEF+N6nxSCWvlhDvWfpOpg6h1Xmi3lDlv7lz6AqftJbUFIY6ash41dB1BQbSBK
KAkbxS5+dTWdIR0g7leyBU7ShFiAfKsz3g3fiHbs1K089ERTkZrcde0lnMsVkXY0
2VTBjvBcGcHGxwu6+D/SOl8wAsUyA2dnmJzKwnzuh78B/ac+VScaDmnu4IoWN2A3
4cg8HSod29Li44Ya46HwJjNB9drTq+0L9AB/ho8Q84ls+CxxBfIlt6iqtiDa/gQX
76t55WArkF35byydwbjolQU0Ly2jhSgU+2Rlcyg23kyMnGHxxSw8hr6vQw328VHm
kMMAziugdczeKnTgg0DqWEooVmIAcjILzPIs9+WxaLVXQxPmB4k0up1Lv3cezUzd
AYxztwl3tvHL6eiyiUjqiaIAgYY7juF49sXYKu5557kGKwHRXg2C+HfiAdbSm/E4
oVz7nlqnlTPU3FBhse+e/Sra/U49t/DRkWWNke8oXlPKZMFG0zazHxxFa5fq+9Hm
9KItLSER+QaBkhUh9hw9CRl9WQrpMXG0DFREZZFTpD9MpcL0dlm3GlGPN7yYCP6T
Nx7pCagPgW3mIJOfxpgUh6CkGTFwkZma2qKH8mKWoHYMQfgT5lp5VJrEIvZz7Mu1
I2mbW/BbsUjSHM0LPLxDhxTRmpl3cD9T9PYR3Td0ZzaxshvpoOJ3t4HllcqxOn56
MubJLRgoWfzNhr77y2jdBTkaGM6NL66mGjFloPRFOsKck4fAltvj9g7ZdYERWw1m
+j84wcSCF72HAmiprOr3n8rkPrX3upFpD5GR9cgGrxR/se+jgWCHW3Zn5HEBBZ6k
W38VE7za5hZjQpRXK6+vXZuWyOQUWnM5c7L8ICyYvgXCyv40vxA97RNo6Nq/VG3V
bzz3/xFLQyeAJIQTjmPfocGt/BEoFYcmylbUuRch5sey6BTzqla4FHi98s4IOjVg
M3csIjylgzOPLLRbLeqBngiB0PL3cedmwBip0HvwykPR02rfgXAa7RiCcNOeR4dw
Ah7rBhvmbL7fVvKdHU2vCW9MjZly0LXWdeYQAxZ30lZ/G/bv3V6DiQZAofVgH2rE
rD0QsXgtepxu/EeodINsf9OEremlen+hDfCVaQ0Nae5rWeC2sz7j3OVbUnDyLqGx
UhwJlb1BFHUQwwPoQgnWYQ5HQEjwTyGjwSOS/40dvw4WhFCcQ1rdfTa2VBqLRXDf
kldZrls9oJXkqVEL0+2kvstd5yuQC8tp2AB6q9r+zjULZurLN5TcdA6FC8OVEwgz
VHmlRWTiCSm6OvhMjbLwSx9/dGEqrKRQWAJX07HJSjqbCkjsnNG2neId7k4fdXYG
ZlbH5UcjXiKLuzNsWoeRG7o8oVaPELmfUPmSrXBFtOZoI1jlevj50ImSAyVOwQk6
XqTLJ3arUnuf8+yjVTtZH4nDRDGtoQIqkRJiL7F2OOOYlAwY2REKcs0D/4gMkW0E
RQkwFO5XLLBp3p2scRlOCnWCi8aBHhMdR3QFCLmS/mCTD47SNX4FY20nlK4b4O6w
9CpHizdhF/XrzzDbME2I1h+9JznlJ5NrsU2flzJkbLg5G0k8fwDQnrxmmlls9AHl
zG3gGxWT4/Q8HdBzKDo3HRaLDVRo/0C2hkFnVEp8PCcnE4qemagELFXe25ll1Eus
kN5KV1+WowuxIwOFrMAtfcEx94WUWy/h1wde8+mdG2UrGVxMyYeWcr2FR/uLXQGe
xMKegHebBxCcKCg4B62ilaAejZkA2z9KJ1uyesI0pcOSYFYFfmWo++h15rtBAFuK
Is5/HHasRwNnJ++HroWjrCrpWgQbENbPLmW0jRODi1Dsnd+VJDpq/RBGUj1w644x
VYka3o4uvra44zFw0Ysn/yg3M1CVsaSZ8UiYvKIzFo4v8Yjlzicy/iTTQRUY1ARR
T1cBTaARvViUeJH+SJ3Y5ELx2AlJA9SOg6XgGjh7q+3Jqg0aPLDNsP5mfsYlLran
OTuadpMoogb7QxxYC1L+vhhRSnfT6awF070SxEloA2k+o6bYk6RljLzNAySAQ095
YOnEgFWRtySxS/bxBWcSYdsEekcrJIe7z5yd5h0UrHbFg9CPSwOb2pQwNRSq630O
X5pZmEKsJ9qRln0ygRQfWB3M88yo+Ub2uPtjbxndD1437Zx8pIzfvlbZPU5msvbK
5fZAUkaymfWIReNQtR75vlkHVLKx8TkSLzh8AB3q2Smw02YQ/Ryh5ibz0tQB7TmF
Myz14YoHPOdlgNCWj6vDtgOeBrpIboa2sXKNnqluHeitW90mB9toWT9lV64sHK3W
WNwJGXXL8DKxighyKWSDsw2FRyxyStJHIhcddmd68kHWoh3Ym3GUgdVzqb9r9WX3
9sTr2IVrv80TC7Irr81UqM1WzuD3ruMtJeBgJZ/kPtEggq4O9smiZaVnucOcaxE4
og0oa0IqOsYVv/WxbNw4GgMBOAanofRFQB2YjrZZzyVw8g3YGXEr3cVZnRBtnj7s
uJkYMo/cVJDZUVQhru6yYDouJBMMGhxQNyqqsvlHtTCzuA6lN5KYlZ594DrTuif4
9Z5khe2y5nZVTjittRkJAFJp/fmj6dDV31SRBuQhSYzOy7fYkh6tMkHqxjnC58LA
pOVMUqUTbfqsjt291hvmbpxspKko+VEbs6IwBMLQcjPWsrkLT7FiUmF7pmnyNUA6
rN0v/R+6dZA9Bpevwk0RihgnuEKUgjmlnbydW3iIgneuU0Wc+X5GWHN0LKvleW4q
KKpF4u6T/cXW4HHJvrvIJ5mKj4lpE1otSdNV36SZtGY19GPpB+zSbI5PlEPMFs1K
yEOclwjo4priiSoZkaiHDRuEZz+j5Ohe5SnOTPgvLKU3MM0lMzdXsgGkhum/LEKF
WTv6wZYuk8MvMVzpzyqGm75cWiKVW/l7UO7mKva10xznani5E+EFHfvE7yqdxnWm
No4mHGcRTkzthudrLZDMakX9nXw/70s5mOkQ0NVPSLwMUdRnNp2vEOyQLEaq59We
oQeNWKN2a8Bead5UlVkLr/DEwBh+XRCmiykeAgakdUYCCayqen7/BdS3jUZOzb3d
Hnt0QJk4Evz8f/tzK0YcRecPBskJk/7uvMAoBxDUFGBjaDG9Zw4KY3kQD+9I0XBP
ZJo9OGc8x8IucTMCBvc0+Yt2m1GLK6pUFWkcPrSDNlu/7PwRgvo9vHXgvPW1EfcW
8HAdeOFp99Nqi3/B4Gi0qSNqCg/mjIkMoZrK4a3987j3m65bnqMGzN3+JZtjow6G
xJrCMWo18t7tQXBJ76JOr0DQm1u/DBNXT+1NeXp/gXaeXOKuGEnl9LJOUpjKWay0
caaDk0foVfdRqaj8sIaKM+1ygSwRo+0rTsJdHDtVzux9tG9GyVd5I/U/LedeAbdJ
1FgFMw/fjp9TVt18VeRDyu2OXE84Fho3ikATmFYaHSscQnkeRGUIQZvEjm96rIBc
NIjbOf/JlqclSpHJ8IqRFbh0jOwOTG3bAejtlGcZEMhb9eZ9d8EWEkuuSsT/6tvp
/kbnpRUXaOnIWURcaIhF0u4bfgjZSpQXPQEsXyi64obfIBp5eNDjswSSObuHHATD
oI7Yp41EXBD58UZTJh+SecggJZFtJpySy631OrWCisf1PQnQGZL4Q+/Ii0jV7uxl
QX4Gwts5dRHpB5oSVyyTIrpGX6uGIE9oqgTwu1BcocJCKxpKHJXga+cX3BvXxPdW
XsZQ0qz7VBHqyF7FhFMpNszSZAck6tY0aNe6iHG6Kx4hq46ZWaev92Sm/xIYmMLU
60biiEX5o/lycDL/fLEEdwJZyIA5v8VFDU0mp/G6rhk1V3+v+g/lyA8DUvWeRGZX
KMc366PIOmxXH8bMKQibfs8VHeyp5bKOkXkKd3R6RcAaDX+eRBfQ3LACem1oOPNn
esfbXyN5xlPNzR1lf79uHN4B3F6oQk5Uiqi78e2qrwSi5dwSRrfIYwJSjVP//i7G
FGRsgg5pC2qi/g8ujp/7LQ8mqcNIOs76Xw3H6jZyRuah8WN6pcmpu8l/hEbsKgQE
P9Q8oaIc7DXm8QumDkbCESm4YYR4QOb6UPtgksyfAOdc+yDMTc4tQFBI6SreWIhD
qiAkEBtUbGq5zaU7df1Fn1nUeDZfTHaHYorMhw3i6GFtvJIIcfuObblkddXIvq8M
CdIHdyafk/UjhUsMZQmdfa6hNJykcuhrgvzsM9Vu0h4okLBGYsYS6c7G63eJqVqi
PR0BlMtwF5O+wrsui8Hio8HD/+/g613xsEFIniy6e+cDfGOkAnzZZB0fljiiw96A
w2Y6Ikan50G1hsJ2JqCHervkub3KIDDDkgNY/tijAlB3j2TpxNAf16QdrL0DXr0w
vegONECCe3y6vzygi2BpwXkqw4Mo+/zoy6AG1Hc3VyCSrM7858JD1BkU4YNB7OUQ
a36l4HdFLc1o1bs7WZsgVx4RDaVVHpVMqkaWskQC+yM57S/mLxFN5DvHcAX6jT0s
k+MjuD2pAIeS/vDc8z92wSgeLd1+KhKJPYXSb0zn9XJBe2lZLO78VDyb9sTp+a/B
TUXDa3xRJhL84FWKLdr/a4qcq5wuW2wh8xZqxZgjHkKkY9PhWTrQGUHqQRG/4zD9
2/re8Z6W54ckhdi7mg39edEtargWVUqL0eP2lFibvjCaRQrJ+0QHPcrZMnZKSKcY
kAyVowr3N18glQCYt4GTrg6gbVTYIpb1IhcsHKJY3WlnwgKHawF50ELFXY8a93Zj
U+7Hjtz8o3Jbx66sYXQp1oroo0UsYi1BGtguAbIaV5mhXlE3rM0cmf2puudCAjQn
+faAPWMTR7NtkI5EDTv/2baLwoCAe9XO3e+1NBkSPcNf6boyABhQGz4UL2gp06v3
C5M78Yvlz/58om+0q+8QecalRhEIsUcoW5OXz/GUh0MQgDcAQ/NGjueeyaziW9/S
MKXeC2q/RIL+FXCYJ8B6db4BRDMBiNZCk845CJT27kS8a+ne2OkkPYiOBeCtzdwP
rhDGSjHPnrGI7RZSf9RBk+k0e65WWLlQ9+KjS3zkXcDfr/mwuhdkNUGXtnMo9m7G
y1EN9xc5PWEQGokIYS08SWMpu0SOY/ETC1fKXF4AopXkkIyR0Zd+mVaNVpyteOg2
dfukD+V6NKZvfULrteVsjqVZrXIv6iH6JJ852Eh99JesuJmnQsvhl00YcHYMVEqT
YyKJomja9f5hBr2+Y0fQdy/lGKIPYQqzEDZuSsPJhj/f2PZa6MJvXQKj8Y1wG4Uq
QxiWdERKYRl2ZFM+q+INNI4ngsQ2JgrzUIVUWi5K+WHnwgjgnZizlOdmknKc4K8/
rtJWGmX8LqSCHOBCm+503hASPbANI1o19k2v7JxZ8bk1eU2sPUj0l8/F9u1MhzBB
EssISb5KYTyDphtwo16jyyj5eDel883eJSY8KVgNeddGGXNP6otip2peUMg5+DF+
eor/HJ3su21ZoQqsA3VXWH1GP8F1WtQ4imsgqJV2g2ceCseD1Lperf2U7jOshe8Y
1xKw48i4kbEMTv5kZFuHn5qediz2TTc7uehBfLHeR2RDA4MwcGe4gwEezFI9hmud
Z+Dqunf1d/DAXZ8hVAuZ/WVMiS0VNDeF5BxqERj5cRtdGn3hJYqRVXNZ7EHohgpF
enEENtjU9ieRoXJAyOrHQhPa/sgGH9EQbIPp2KnALsLwyOJqMUgHLkb/K4WvlV6z
nd3/SdGIOiqQ82nUopOxCMEl/t7K/4dQYj5sOBMdAIqn9XEseut4DzBdfyTMfszS
AG0qOqw3fIUvZPGXIWmP/ruBs/jLc7OjYwHMq7O86MbOUSyQRIiGQ2IqQ0ojLqKU
5ZxinV+5N5sMrG+/2ZAGsUPp8zEb5STveQ/drBr90qKj1Mb4y8ROOve0lYiwjts8
XcAqJedUuOH1csHoFPSzfcMCHKOWkYhrgeIKOuhFhOnHBGCObCnOT1DVLMhRmbVy
2QqS1mTKuSV83f8QUFRtHKgjik0tsImH1twJHtmR88QsH34Iq7aGs1JjP7woX2f8
P/tLaNNoGEcnsq2V+0t+JKtUaKVcDG8GXNhcuYxT9jERKslHGtFMPQVi/s7SxFdx
guu4+ks5AM9Frpv/GqaDizu00REmT6ANy6/htzu13iuIHPttQ70bAXwyx9Ai3luX
qFv7fpU1U+1myzMG5wYiP3uFeO45NxCiUdaElzV70Wm8UIQZyLSLS1zsdtqsBR5U
6Dz0nsfBecUD3pTI081s8uwocs+wMur3Xs/o9/JJB5XzFx1fa5r0f6T+YVWJFInz
cVhF+30jh1g6AVeJ4QCsdv8XP686boUJ9/BS1r2PsdT8CNbPNVDq0BdC8fKTni9w
LdtiU4kCkfJZIhuR+pEW3VXiquLmB2uG7wAvmHp55u3cJ/RMjLOZXFu4zA2rMBov
kIIJR1HKtyl2HkL5LHm+/CQUkCzMhbZhPGLyQT5BO7ovhjEjdAXii/AtONZ36yxM
OX1yAENMk6CzK79s3keuXsyLEIvthpcoTvIXrQ2VH/OEaLggIXZJzKmvUrk+IvUC
ZnxRwYJ6fWEOz0QzTf7ZyLXfEtNzuGWLbrEvGioJRm4WPLneVjYpEQZkL7VsEbK5
g2xgxDiGfIvsWxhTXRhIi8Ln3UYwdWD7TTnDC+u26powzL6OzfKtGfN9TIFSHHDE
JmcMGBFY6D1gzt1Qpx4RVn6A660xRslC22ngmCCRybTNmktMI0ywYOilNlXAtjDT
ce0hu7bIOkTbV3//xvx0ZT7GQZbuoxMfSHK71dME0tg64SUn3XkYphx1rkBvBrTG
boOH0TckCO4oyVLm1IT9V5CRbN7qY1oV3IfsH44ymK4EBBGfKQz0EL2uMyCBSDHM
+X0VRqgQvMXRS9HwbQ4qQd6ChaSPspuk2v1bERjk/7rt2OU3q2E8dmpt67DIXlA0
c2wwdvDNJycTCnmZbSt5Z76b3/PXdBUhlGuzPX3iso/0VAgy3DECzcnfSnzThIsz
N0XnFsrdftkbNwPNP4oN+ss0SAsDjFHkttj0rDtc+Wj5fJdEJn/u7eSNcdukEGit
eLCtQj7N0d5a0I37RzqJJSK3HTWMPrYKTi22kiG1SEBjlagk1S0BUiusvtJ0xg8U
gyIzU2S/H33G0ZrHWflT/rAy8ZF4exsFy1IhJi4Xws78xtXHDNN2W0lwIGCc+6bg
gGxhw/2Ke/rXd8xMZZ8kjA8O/k/O2jhQ8wAX+KHExg3IRZgSk1E+L3I46x/nyx4D
s5ImlMymDAxY5uLl6cFPE/osah7CPsMMutM2XtIlN63zSO//ndRcTVU3H/Svmqxw
ZdmkX2knq/Ot2hcex8+0jT7JyjrqmRqQwlPPM+1XypFFvxv98Vh8PN1EiCHwtTMf
jx8r93sHX0VvKKxhM1JkZFxgM+xPG8NLPmy/YtRzRy6HlEoninImZH0VgHEyqYBU
512UGFd15cMLVovic/a6fS/4Syvk7MUjr68+rNxtVs+ppNnLMl/tnIttgu5fjpaL
aLe1usdUT6u2yEsSMx5MXc5FjMktLO6nD22DB8B/e/YJGvKJ7lwlvfMvnOmPfcZ+
lGZNpVC1MQynBks8q4VHhKuSji6fK0dluqbbF8J0bDYCLvU/1WO/JCZFtWlDYIp2
2x89Fh7V5jAeiDgy7QOoGb5HoI3cgojBGyBLQ30tDLzwMFZsQY8Ke9B3jji+lH92
Hqj/0cMlwMWSEJyXFYMJrnm7G+yjHTv8+sEL6tH0NZCv77o144WwJjSxNS+e96fG
GJhmBxQ1jNM/BnfQ7GmMNkYSV52CopN/nJm2BFy3mEI4IbdVaKv6Vzan86U++vM4
W31EYuv6FswFw4I+EnUP6HTsPukwcuhFbW/8mCAgFSvk8FiCX8wK4m8NWrx52l/V
Q2jzpj4TvzQ+PzWwnD5lFZpzO7yb+wUDNMTcmdOplbJHh0VRC6C/NqVCNb24Iv5u
RRctFzC9cJTcGkWYKQuEqsOP3WgnixZAqBaSXyUt/NbC0GfExv4qV5WcRhqZkoPl
ssuXaydYTaEDwP8VFZkKJQFjoh+uMlsPkc4XA4OZK6GGHDvU5zQbosAIjdqmYD0r
3+4pUQchWnSpY6nUcJZog/N/QUhqaCxBfM8KKo2CLlBGDP35gByOrRw5E+/TQOMd
JdjYGDOvUbzUQdv1qoMjy8uwXbkfR0esnfFgCRblkiX/7nqbsSJIzpGxK05aDubf
tmumBsAPwuvIzIXIjKBbLI0pwQzli8GIjg1+6BJ3V4aJL+Xg86r26Gl2IwXqJeYz
vpuZD7ZzIBiYuOPX8QO7DnTL6hb23L8K1vDm0P85Du3SojI4CmjAStX/r2vo4A/h
ZZgdvqYqHFOfQLbx/6qwKlJOeod/Eoek4CeuZfYlotg+YUgYWPyxCS4jY0A+fCri
w2+eozffGCVgAzZgujGQ9MLRcgpf6ZQLzqnhUDXgglDpPs/C0N2zZ8BVIBNiI/e+
6b6ktXKaElSyd49FUfCOz+CBC8urBWwRefGX35ofbwwCdcQNdR2j4qQ4EoM5fW55
RppIeP7GVRiT0nmuIQuoEiI2dMvvBbTY4KlnZq01dRASMU66TovOu8QE/1MiDPVf
SEfcd4HM5ECNAbbqioU2XELCyn+cHYPg20TD+xFm9zcFxuV3jMLwJqthsJA0Cdys
BVlV4JBoc5+b27Ro3stijGBAgpjZb5Mz9QkUsxKrmUlfNH13MGdUkwcRhILSj21p
9n5PB1N6rjQmDeOJyhknnxDGUVkjVv8pcRg4JIOOHqkwsReTTa/BLKFW5tf0dgNK
OZMKR/Xjf/myWnQ2a7y25/bw38MHl88GH/aSqSZHGc4m64KAn9G5ydNRLjMPUo45
O9ollBRPw44Ei9jMpXCGBpNgpRz4TQ5VyW/zqK/rRLMOcKK0ksZLII2u8lE/ZyZQ
0xdYklGsZxqYHue6zC46FDopN9lAm0iGc/TdNVvfFldZlKpf7o6dh0PmYJb4dLMp
MD2kLrAxoE8Gwy2YGEaQvYgkRvQdlII/nCufYPYDO/5Vyr/XYNOnGEDI6ZjCjMA+
r2lHtHR+82Ky0S6AzsgK9in4Q6SXHsHX7/Xn3L++hjTc1EYbJO3++0Sb0Xajsg4l
YbpTEviOyX26OsGiZ0yhD/8XdM5hlZPRsRcPdtmQopbos+sqoFSyjvBk5yXB1b0k
/nhGScx67kzvv709hIPCdM3g9zxUbffj0V17+YV9tMlbIbkhxpgySmJRQIzT59gd
ORHHpfiLrRhXufk8hkXJ/ySUb1AJWUD5Lil62qYMdwsYXohcRuMXNC2PRgv7e3xE
a1Hf/U1NxQ/qMM2AiAHhPd+3LseBzZZpQtxP8QcOaGCbu1DPIN3IFRl3hn3iwlN7
R2aIVWNzw9axopcOqkSa+2RKbAvP783il2DALqFa2BgdmXldSfV5PYOPV1yZHqOB
srEoKUD2Q1UQxVvxNjXFRTSmiIugtoH9lhEuGOQT0QQeyh7EtbLG/pBH76YqBNJS
Q4hO5R6qj8oiVr0LEn8f7FOde6Jd8WZjdt0fxOluHnI34LiImSv9XNDkkISRnreb
OKHSRgHRkcGJx/MPnDPM1BrDh0XBI3XsQNvKmDDS+uGuMxZ0wspgPskIQiLlzyGm
yOEfql9YoHZnF2MFDecZBzfRV7qbwFDlHL8UNrLTei42IKyxKrJfuMzun4SyRnp2
wseaE23FB1WDENW2f3TDCbg6kcx66lRW8hlEXJ4zHtEKbFSYOpoKm2L5v3zOYnEB
NySmTIHle/d/Tfrbzf0tD4vxxw3grWpSw4BV4Vj4s9aLsV2kBiwWtFkMnHtNx8kO
pD+JI16hM+CaHER+M4koFl+9poWI6f6Q5kc2vP8QR3D8pbzLhqV2qUNflpoHDpzo
xHtkrkDOpiWjgU5Vk8A1E+pwUHU+GYo0m3zv2yrMkjHJkRbby/bP0ipbILxly8Vj
i9GhXhpvu5ycEdJt6q26FGXebSWI4AsbD2FIUaDSLygAyIiYb5D+EPmqisTq2SzA
Mm0ySr2q7bgf10MpjTjrf62tt2elOtX9PD2jATHPN5pBuRpqzbUc8dEN6BfcPwLu
b9Sbo4r/LkIyoH+YofR7nBcE5enyBk9LakHdw2XwIDsDCXpOzuSvCNZ1W+XG5wXR
WeHdmXnHHGSgn/rk0/jIhDJE+eeW4VA20o95ptdZPPJ4O5lnkfWaKaJcauF9jayb
F1Hiogbaz+bnjYJ6znVpD3fG1Lr2ZlPI8+JmkIlpMbmBc6V/7QYDw3Y3njRK8yya
vqUeZBglhz08dRrJkVjyUZgVKIgVpEIPryNAhTbEknuS6ZzZ9/VniNFEiEM5fWuM
85jpAwpqKSwIz/EpDL0t/vWxGw2Aq3DMFxF3appEGZm+9h4ZuCtKzRn8rb6pspo9
sqo1twltUnstvGqoegynPG0BtsblEiSphxiz60wbBH5suRZB/zoeB21AgUEBXc9h
Y2rD9ZMRPzXmP90tFfP9k89L//kuv98qzd0cP05Yrv+JEvsM8XLcnFELXrsBm+Id
KRmicoIi7ldIo5WRBedOBSj+TFSwnPk2Dg9BVAIdEyix3wtGZ+pODbm6OZEJzi88
3vYw0+73+upU5spJc5GgJlKNYJMK8VYU+KwPQBNCqzF2IK5WlJKcz9jmO/Gjojs8
928uEZTqgE7j0o7x/NTcbQ+QVQ6sQPqu8mmAAn0euRIbI/jTqbRuIoY/02+AHXJ1
zrkK56XYCo+lszMO0P0c68r2FPHMxV7aA6Fv2dRUpHVlStSwPajpvk60Spew7gIZ
RWL7011NolFFyWbOa0Qrjn9BDhXv5pR/HkKKkZkJEhEajaANJ9TTWLKHTN5cABRx
Nac0Of71T9kRsG+kOuApF0xNsSm+S37P1voyFmiGwv0lHdVCavazAx46MY9nBGKU
FWAlcCrINtxiwEZOHQ4UH9PlsmEqKGoPjjz27JxQkjeTnOgEXBZ44yTaRsbA0W6C
sxUNkEshgsjA5SMLOYAd9Q8qKyYsl5JEB5kGZwTlzKoHxFZMUq+2JlZslNrDGIpO
9Xax7JgefIhMszT5JnxuYIM3k6vTX6wb2CTUSDX7TS1/11r5FizZAN5BzdSKQhXU
HSo+1DQYyVhANBYUpcIYVjvje4NSjBIG5xn7Yd6POMt4FKlz62QrIjzXXmxHGDcn
GAMh7FBEH+Q0ArziivcOYfLRgEe10OYNNBdO71acjQQKoLK7sG4vyXe9LCW0r8ih
WjVfucl8DOxlTjaldIZ77Cm2Cgfdfmxq9iYmRfzjSPDU0Lvr7TNACtYUUgtK3AlB
inprSoBUnzNeZl0pfXWTPBqFHewsQrjZFkIMRHRrsmV3g4MSUUjBkgKbft1QcGO3
mrMmQHoUygOPdATxPuSUKMa5Mme1cRhnS2ho6ogjTRpfXoje5zfK41bcrbdLc1bs
uLMw7GlBmgBlEKfkE4e8FqHEyMbsT+Pay87UIbZCxpF+XwJNs5YovpttQmHf+++P
glvIL/vtWbUViUqfWHrSUThLV/405yETu3QfgQLgcR+m+SRXJm8zY3sfZ21B1xzR
G/XqHWhdPCiovWVS7Prl+HZdagpq2zxD4oRfR+Dwu9IHs35aJ+duyKZ+QYvuozdb
NYWW6FttDZ7B8eyalgOT6/Kbgln2NA5eGQD8ZVWZ8L0zi11RzpYY0e1xRkKMf5Og
oApUSAIrr4Qs0uFxSuRsaGR1O3eF4AQIX98ZUeoToXQPM4IfGUvovgsyC1fhhq2x
tKeH8IBrqR/SI5vU4nG1wKdAzxnx1FSeDMf2xCvs7Nd0Q64oZrKgfeQ7kC75T5/T
LHQ0MqB7rBEDGOLFiPpTFJEwEcJq/xRPNB58EoPllg+KPVBeWgLsecW+0POtyoIz
XKqWMzzs+FnZCf7efdsyC8IW8Z76UxhhjuLCWxlsHDg4JJds6/kLJWs7MouMVnW8
YAygNbxlLRnJB4T+i5QccwlvhKpRtuVNIKMKdj8gEkuoMVAlNcZL0I+YwndVL+Sl
W9FYQKW1Y8q/TNGO9bOMxz6EgPqgd4CFKp0FFndIoIldcZU1V7d8bj2S3rWVheu+
zXXU4pzX9UHMR8W0fBjvykROx9RDCAf4iuN93UFDfyFnJEXqS4gWYn9Iy/nLXhV5
2eI8MFOW2B40L+QXj45zlv2dwnLLEMr6W9SeP0Ak58GmCmA4sBf2gRbNJi05nXQ0
OCvQ6QF6eCOizE12BrYDnZL5hApNarVwstzxul83fsiGGauiJITlKKHRIZlaaHGP
t1XgY6vvt4BOrAf/B20iKEfV/KhrzygmJKIPyRfB3C4kEtb/cxWK1q9+HINmArgg
uWZpgB7QhfgWtJx3U6q5u01MpCTlFSbgi5rQi70emA8Lbwd3ZlKBEwWIxAUtE6+D
z6i0EIZyr4xR3qO/sZeVLzVZhpyczE9VMQOsSwzXvbw7LoTpI0qHXtO7MNY6xfuH
XQw0RCu7LUQfPl3eS/SYmvtPka76iM0jE7StMF7Qd7FdK1ERekXQ/33QEwWKdivJ
MBKHZ7BgXSXqAV8dTvuvig==

`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
l8AkhYK61ayVHeteo/OFwQ2xtwTiNswruFocpanfVNQo7ij8WCRKZINu5l72t3Fw
2WXPGLkNZyOQlIugy/nw9ZsMghVGiAem9DEKBDO6wj1dllsjLFgSJxxbxC+GZ8TF
OQ/SKlo0MTsoq9hUqCQtY6N1pmavQhmqmPJcNFQ0XTI=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 14368 )
`pragma protect data_block
DDPw6/Pseumg4FK3VctbLGUArd5/RiK/I5uPDbh8fQqlVKP0xywFij5PHtplpCYk
xBsDjNhCYWb2r8/IT9rzk0RM6vFELWKreROif2LClkyHF4QvbCOM8xEQJbeY5MSc
llnPvEEqcCBJxmQHZMmVlq1DwGGmV8z2M3DlBQP0BhCQo9q+fSlcFJEcUbkkbfjJ
FGxyqMVrqQ7q1BK/DB6TO/1gjYAOaTG5bS+Y1gQY+MwnjLBYLQFz1NL1G8NVYAs7
6m6DZllFSpaGWTbj9rszeETjX+ARbJJKbxKkT4QEp1hdE6bkeNeqFfyP0kaOuFms
z7obcTGorkML95w0WybzvZVQPu9xmD2mzQf8zyFEhRxGivZS9rBIHL44lt5yrTM/
qHZfpC4izqTfRmGA1E8QH0HCMd+egnZtthTBajNu2n2ry1pe6mmHsKovK8l7HC12
VwcDrlTYKERb1MhaOGMiNdMtbbqq3VBYh9yRJ89NCoZCcvd66/8gHNLxwY611LaI
8ZNp1fvspyZBVKYXbF/KOgGXxHGfRIYp7b1+V9i4r7B2lwld/lOTozxkaVFFjPZE
MvSByVKXglhSJwiHxUDx04dGrQLLM4TPHy9HFrt3bGZMso+87KKg0uLJFLIM7RmU
pQYao3D5677Cg6rsdx8OFpZSTu34Xzpvjf23HYlK821myquML5stQqWOBwPwl5ZV
t6UV/LbD+fhhUPD8OQX+Z4fwyXKS/EapwvHpzCWhBbddP+95m0mrcVEfXsc3wBPW
KdJWIdpK2QfxQ+Pku8HaPb0cRw1XN889pRqEAJENTI4QtMyjoF6RNX4H8CCkCbhN
Gj77Fo+FjJB6ZeLJDm+a/LVf7T30MT01iGIqu3xzTnBhWAYIJ73yrExxbdSMLKVa
NNOKz+ZsrUMOyGo/hFbtH/rFAm9WQT3K5HioX6jOTsnny0zapQkPomHEQJ0u9EZ1
Xw7gxw1U1TKlPo+HzSeRJ/b45CujuK0PlR19E9jn/eiLwBtpSNYSQxinGV0xNjPa
Z+0V0fBOXUEgwNHbLzd209sYzxu4eZ8emYAZ+C4H4UOqRkt8AulzbC6tIYmBftyt
gY/rZ0+lNvHpmzSGQI9ayZcqb8/vgtzUNVeaLvLUTfOjLc+/0K3ItY395JHGLkGb
PGrARs56PS7bIuWbj87dbJ7NGUwFtg/w+snrvWFyu+vJb+HaQ7YjMGS6YpVRVEED
wbjBcrU9wIS6/67AkY/2MOVxPUintv8G7YBXdvGvTAk+R50adP3A2fRpQCIwwlZ8
FjD34TkpaayNXX+t3WI56He//Jro67YTrzr35TcbxOrK+X6TgtZ39Vntg2xD2uUw
wCW47Kuw3iGLcR5sXsIPIxl88lPZgfRVzcXqtPBql9OmD1HfTp0UwB5F6mrAOAkC
EgDQMnQ63v4bxZ280cplulH5DuaRj4c4sfqwWtMcm5Twg8NgT20qfAfeU4xWiqXR
hLG9DZowfAWhH3cARz/gvCmV7MP38lEaeTRcY4B430g3F4SnYR1U3Gr1fsMiHnw3
X3p+h6ptDYmg2ErSUoujYA4M4MfyvpHYBO6gmWGI2lmSUGhFi7elDiMPAHKkmae6
1ttVaYqyY1hdV6OILXjgZaWROpxvCTfvKdxqwLSbMSMTvJrs7OqeM4evyXfSF3yW
0rSPNAoBf8kJgF1peXTjkQwy6+SLBKxC691g3ucjk/y60Lrq7CSRALn4LFdx/GcT
YJ09HzCsHlJX5fO6SXqPR4I+naWzddjnw8o5vw5m47dTxvJPb5oJfgIWNaiKM42q
12vKroKsYa8uBNzcvwJthYS+go1ZwYTLKjOg48B3d+6vUPBTaFL6sYIMmhUko8NJ
Tz37ha21tA1YCtvcx28esOUH38Y9mZqS5YZV4q8OB4Dasp7AxsLEc6hVQ3tsXFoh
IztRbx0hxW5kEgrZOXZoLyDCl0LYsYDUhFtIfVrC2sPULIiUFCZBz6d9OEnRFTfN
Q1pTx2IFXmV2QnMQYAc6sh0TOqw8K+IV9YZkdm4s7sAeTGlGLR0f/Wm+EbOfinzp
hMBopSdp89Bn7ovX9keBI+l2pyAZcmSnJ5fAEYGbJNBi/EZBLtuwXTMWwnkyXUWB
y+qHADFI85FGav7oXRDTxLQu1nm5PPK8CgezGD7vxSzUH+v6rG5tRtGGIhhe/X9K
bq40CLI9D3p0auE51HVOd5JFiEIYImJIa2M7kp5IkBQgxM4FQ/3H+UHDemLvverK
CEuDZN+w4vQNGBvFlqnyTL5JSSq7vV3pg9d3XZgKsM9gGWasCxFIrAG5P1i2NKRA
R6OfGLFzVydLOTLGppQmVHhoKdt1tGJzcUeJhPT5sMDOAtITh8nR7B+XcgVbmOtN
M/DVdl20GpI/sTGZp++V0ZnkJgQmMeex2pKvqXCrS4peO2z/WFA4Qo57zzQCSf95
PnGxIhUp8tIRPihqNEsfdeRMwXbOSmdyu0rxzi4P7V8Ro46QugcV37k/Zb/8goqB
J1hIOkG4wtS0JXCKFiGvzN0G1yHOGpSVvfFvHTK6YhvXU09ESVbKBy2JHdPaZqHV
ZJ9k0HZq1azVPc92UkLf0RdA7FpOaj1rHX5cdCvSo3+vuWStzrKB9XvEVy24Tzuh
qeEccjUv0bva8m3j9Mx6mR1NzIoYRD6hbmH8Ay/VVb00miuf7EztFdht/jbhB00P
b/bz2kHK3yVbLML49WJDxgEWLDBR95Z50KlVOZNehLj+TKSBOHUeVoM+yAsDtSJ0
DMOXmhUZyYZadD7CdSVGOnT0RbPZlOp76zDD8ByrTwMhoCwaF4DSlzhBz1UXdb9e
xS4jLoBMXiy5TW+GTNx6bND6Lil3xFd4enlMYZ5PU0CrBUW6szYGPMPi5FbaIX85
A8e+Gf+AHEe1rGcqovazl82AMYOTj/3tbhFj/N34S42s+2memClwvFV5Pbr6T3y7
apVlItBm/2cKz2BP6TKK4yQUpbVxzxEoojFEGFZTjgyxyonjgRMH2TuGn2LFNm22
bmizL7/XPRN/Gz4co6uZfFU0rpThYvDulL4NL7DuqA/YFenUJQVPKc+oWP9kHCdc
Lr9awGzGn/1yZZKOyNFYEHIC+lix/AdtlIuDzzwYMtYjUAIUS3vCqqxiW3xruAWk
K54NbPa2mSc3JdnI3Z+u1cpjxiCytNaq8fpnh1RfWqHHv7mpPUsPaSyEmTqHrj/J
ea8dZ2aagP8JLRz/IMUj0UmADcvGZf76cemA0GMkLTxB5ffq0qjJaXq0FIQptQAM
iyRtd04Qnp5BF7QHN7fpRrB2hxLisyEzjuyzNpceXNgY8FP9Ec/JoJNQaSWM5NSa
u0cSWeA1jLSNt+fftUA0X+Jl34BXCRmicP01M50w/BUHEvbyJUUpZJz0KbBgxGFI
80DOI+BfBvSNLPSou9pOty4ILZL82HjMjo9mW9ve0KzTLCzFxxVAgXLVrGTCDJdE
cvclCCx/Fzh2zw0C/x0dtQAhIRUjnKbM4Yk4+IpkJJ+Jgdv1qEFl1ErGiCN6wc96
wF0elP9S74R8FYPMCwfyhYmVnKsRFUhuueiXsD2v2dUAbDWjC7RsD4oSsOl8cvV3
/8bjRbrsOuFR7vUBfrpiDiH/2CcWHIRoO9v0eygIXGThGxsOYi2zwZtmixKdnOfn
L2nIEV9bM4aLjMWB+QMBj/ImGRhoO9HYDdTwd709Q58DDjdkGbf8/vvRQAmWMcKR
aVqDTooAKvqxXoHQ27xk/wYDub0BqG+8OjO1heRYmQvk9TTB/mMHOopLuFQbrkWK
H6azEXW1WySk0E5EiR60A9BoCjcMVEW04AQhojmPqCAZTsTlcF/l3/I6DJpIICKt
iyfALKIeXZSPe2J27DvAOHKk8gjf59N50VZVIQjk+tRd/ctre7Oz9vMaoGFPXXBv
+c2RX5Xb86W16DL+j2lsTbCFipUIJscFpV1op10limbXxfrJ8gOgKRE2DNcQa6sH
5SOoVKHOOOwDPmLn6v0QOwk/f7MFvXJ7b0WtRaOq/j/WkFhCLY3GsTTC3AgZCWej
huBq08A6r6N9ONjLuUy3wi3BfCoIzn2t0JC+pNpMKv8Zna72hnNhQVVG4SQt+uQH
u9mXVQ0E99qbvTd7TTPQ5TdzP/ZmpwNYIZ/ShP+ja1bQIDvauJRgOStZLKTo/zp1
qP+HrsT7SsBSHbWQns0rYvC+pi6PYREfDlrrD6Mr17a9okOOPNUYtqLAgONhBLso
turfLRe4vXANqld49xorQ/VdsHxnCE7JE3eVivilfY1q0Ltj4rtiPjx+WWOjEzQb
SMDlVAjTbvOJWWDaRtVRlNalQcYhTu76lQaldz33qtYBGWuvxb3GlSI0JkB2mtaS
4MVJIhG2wMiDv01brOye9m4B0izrLVI0xIBycKMidkoc/P1BMvpwTU0/AL9/abW3
I+hu0d/C68KonIbsHBfMZTPZF8OcPUseTJKbVRmLOCbwJSqzHKuZY+3xajEZf9bz
iakA6OOW/s9XlhI6R1/OUoFKwozmX6S6GtZzEJznsOcmITIfo4Mb4NB+DgFAU2m4
6kHQ0PWBjhua/ntnxMvwAU2LYv98COALY6rF57bkZH1IBDvmp9IaL003nHVFRejb
WDMkPwznkAcSjcfwGyJT7t9yyqfMNmSWgaryM4B29D5BRbiT520WnwxUGqSgRO1t
9qPS7ZAqsFnmv606LM2TOLAj/namG3Jlah+vtQgPuv64XfjLjkKRMtPVABDGFspr
bMbRoGh4SlAud+7iCXOnrzxmkiGyRZrlISzVshntJtc5T9SsuMQMhjD3QqYt7aug
oMBWCZuLGrY81NikUhwRrJGTWXyfnbYZpzJrmtvQ3AzOmdid3snYDVV6nFGMCs3r
Nd+dKh7yODOjXi8OhDNoQ2B55MfJSCVwOra5LHRmX/xqkeCRMikGz10Z5EEiS0XW
JBng6u+CRdXitwbb+hGulAYqRKILpinpA6W1zPu7Kl8yxlFVcsFokF33YOLC7PpI
Je6QlxT2fGFPnKWhocC2Onj8pBNnKfTOVsiuYswQjNdPoKP5Qm3WwR9dQJBDaFAC
VI71Pb36yzGzCwZB8P1sPrDpWWxtU7wOpc9aMHHWZe71or+dLZvUcq9umKpJdKM6
j+wpDHi/9cPdd4usfwSwtwrijSaB7eClS0MNtcZL2DblKjU/ZvfmDyLUKpeR+6Re
/CXEIQnvXNJkEh2+eoFpeL1zUlcKGiVsSUlXbbBVRr1zuvLGRZQpMNLdykal2x8X
WPBWKazqLIspC3X50XiorcLm8ekkzySPcUL/v1a6Jrimi2FNu5Aa2I8Ow9XDc2N5
CNqX7Ns8PuALqccE6IyDHkGrIU+MLQO4B/smnKt1sH8ZBPGTzU1gfLTc1AjvxQ51
0oFG+rYuuwmQMwWyrDd3LWX0XFnuFd9JZQMK+Eh0LyCq05PNsTpL5mFLwp+nVmzL
bXKOE7tA/hmeDhxkqiv5bJ8VhoI19L4AwW7cn6aObH6/Y6DJViWvdZ/as39G4Kd/
lFnXrrWRI0B9nJ0WTJrzVRQpbk27A9wIclcpT6IH85VY8C8aX7VYa0KiqzKCsKV4
A3jSGt9HNtRAeVJOfhylcWI+9s03+1/+g/CF9HBmy0FFzehovcNM6WdvG7duhuCH
c9lgHAd5sR7vUFVWQeLLVPauN69rn2qlFPnvPAjsXaX1aP9VmYvSx09QgSlUQfA3
+EQrXBVJ9qLpLaY4WXmDuCoobmsm7vwfERqgQq3ZaXfNGWpkXTc9Qxhia6HLhBfi
J8WBmy4FzwzdHo6EEb56Xvco1a2nk7b9N4lIP95+tU3EMMKxn6oND8C4RoVL3Z5p
A+8yMeoQ3kfDVqpNF3QKcM1f0ki5kQyexkS0V975ex5/LYEPYSQ8Zx2bzO0u142l
+pdQGeu/Cm1xmJAXh8cmRMMMouNmZOkWlyJx5hXGHZq4BvzYmoP/gEpOYqvx+R+a
jDldK70eo3cui1uXXpeGhzrxhFAb6HndVvy59tm7t4yHDdFUVp2Nz133XFpnvEdp
mVyXpNiRXIDbWhTvv23/6L6jViCL+ueizVKfVc4MxIfzbMHR/j8vUhg4bfEP5m7F
b8Vz5MSdZ/W8ztPeReQmNVrxB2JuJNkH43QgDpHJ4Ej5O0DiWqtFlVR4HBIPnW85
u8UkknHqKrtXcVpl0GgUTzxbfEJRSCRtYtFFnuK4jKWjUVXu3tmvmFOeZ2w1Npem
0jDtfnI4pBcM4hOjGDLwWfVV5a0Hi5b4zbkMBhJRYs3y2I8n804al3iAtRpMoytv
S3gVsGSuznzStEOop5aXHHR7xVOeTnbnWgLqp1c7AFKOIgfKOEWihb8DOuIrW/ih
B+30tsSYk/NVEGhNQCotCIAA8lDPeWo2GZ7jAfgXrt3m60eyujXQUaHpca8TuMmN
Jm6lRH4MDA43p6i/EzKCAr5qsSb+lqVkB/XCLHRgFX48sc1ZuccB9BEj+gi4qUzB
FCh0I5AvBmFYLOLjMhpnRT+QaYjoadSKFkgszgO9PEJkmxaSD3w8AJkELMbclgj7
KPa5O7/oES2TXW89Yf6vE8NMfE5lgIu4g8hFfdKPcNlmxP+A4J6s/i6uTy/wxF3c
W8XRXFZpQswoc5+PtCLiGrsDx9H/htuLYclZRclKr+QiwcOjMnVGKEULqL/lpW6A
3UASQU13CXANu6tdCBbwcwdwJerJAMbYyYATzE5aZTqbrNLtYZaGmYqY0I6dL/eT
JJc7tME4PtAEkd8fuYgsyUn202qbmWrogHOJLpwifuBc5kESMFKWJpDtdBljhAMi
zMET3FjxGPdItOXO8dMjp06z2cmLs02gk25EdfYalXzqOQ3Ho5xJPBBrKks7vS91
+UUE+fvDM3pH2mhpZcD5TXpt8mw0JJHIW9sBkd4qMOVdBVc3dwcFrAlkgJACSaKn
D+N//YqZ+BlqMdNYgljXUwqzEOQNExxt8EBnyLu0w+dmo6K8EU9O+A+lCkgHN6Uq
rY2pPAB992pvquhPb+4zPj+BvXI7UH7J6y9eS+bjh3Dde625AV8MIDUVmM5iDuXs
X3o7hWnF9WB0DcLQfyyfKGDX65crqOYVP5dfK7E6p1Im2ZqAf3JLgSHxwBtwIZse
eVePK9D36pmthlcRdref8eb8N7vQsSqpRSwaBndru1HbyxyglaMroKSCsT5t6hm3
xt45zI3Ha+SuoTSzcAakcK7fej2cGjWgyS9f5i5OMxiO4et4KGtblWzUkKHnuq2O
eGNoaxogz62Ho3H4GSAPTgz1nN+qCBufHKiX6dW+LF5gZxBsQOAGoDFN6P6XUICe
drhTosKkfFGKsLASjuf4hko05qQRg7/4VYoTR4jl4G5tFiyWMNwb8A0jXdzngKjZ
iGKXfIjJYgJFa2/wmCVhvqEH69E1EuQf+zOcspESj9Kz/zEQH0lt3MY90Up3Gz+/
wKl7LxYP0k9H1+fsJNJed3LqU8BULCWJHWXuzz5rFw/disIZxaucxz3a/5dn6IO4
kadLnrSyNv6A1Uv3q477Bd4tvX8Xkn/f8TykMbiDbmiVzFZeTYeXU1WLaxQYlysv
I6GQE9K4O8trapT3qcZmdwcI6FfFzb8iqD+AUZXNUXDXpoXTXxWDAb8WG2S5vCVh
Ng+Vekv7eoVHZF3FRYWisV7wx54Rc454NSp7p1tqeLexYnc6ngkxUXQD1VaI/18k
+b+7gbswLONbxRuNSrdUaHPLh83rphiZQbKG+cZ9MGMgZlEDbPNj8SCZ2hPntyIg
pCSGymZ/xCRgXN68bDMzykggFp8LfimA5B4do3BZLavxqONoIvy5r7AANvXh7FHa
JN5/K7J9KEVvkzcxRNxzq16NUb8VkIUM+JdebnLLbJNgeZixBfO7rKKXwvLkPH3W
NjDOXf2yJenB5eLhXWcvc64++UiGym3lsPmnEpMAqV05DmsDXZDGFkcAQiqRvCoS
7APeS02UnSWERwrcnL7Fmm/kRjOu+Ez4ehZjWW1zI9TFkq26j2Enp4J2ONVLLKdK
Gc3xVmharkLFRtFU19yhbYaEFzaI0QHdQJIwyfxYEfFCa8WQ6YTObicWY4JFT3dA
wvc06H/PmK3GK8omI1Fmi3aA1qsZK2ZBne0dHqd0h/ibrzRdQo3Qdo7HmirWkDX7
lcfw1VcPmW/85vjFiq8ft24IlrPe7Smk0UUyiDBJisg7CfKoFgAO/bEepABlgTDB
eEZX3kM7kTEofAgzECkcyPwfnFggG+6Ds6V44aUZSdyFnb+V2LFwI+CRcOVvDjem
r7TzZlBt+qD+2b5lx40qJLdObEcaj67O4SgmxaA9y3owG8rwrvsVX8IWUbzAR7jr
M0fhG9DGTOamxCeqnewaxyzutmgMW5UVnWRG7i8heODBlJmddVfAtHiz4txpEqVf
S9dzWmDgArpQV21ANKBOMBRI+AfRDPS7RavBNkV0rik/Z3pv3h9jnaCZFomi16xo
/DsBR6OT2dOiLszhXoTXExwDsedlLA7D1RZSzZDYdoRZdqf1f7uGg6t7N7DwilbT
p9ou9800CE/mLVygN6LEh1QYfnGZssohqRDoPmeg0U9w+P3aYQ9IEGRYhkz/hDxG
k46HERH/J94t7PAlRkQlcgUPKiy9ssuswSw5k9V8xest95VRXaZb24cRtIr+tCx+
sl98NZfKeW1PWcxqlyR4Q8ZUwrSz/t6UNQYN83/qS+aUk+wBzTNsbgftiBiqDR64
7OXL+lEQdrHGfdplfM+i0lElklRFPBFMmMM2ah3ss1YepX57Wawz3lpksmunTP7U
Gp4x2dYsa4aj/Kqs9yHbak+jiTfZ8Zpg8LGN3y9mGCr3EoJMrq90LxtMcEoG1SFt
jEehDXG2qkS/4xI4dShbIlrs9wXOnFJHPgVg53TtU57R2+QsiDsDxGkVokhmLm6i
Szz0KSMimNR2W+sxQIpBJASVUtPodVplJFlN4CJDmQzwGA48iEqayM2neoOxX/as
WVgnb0pVqsHswOVECapK6MPJzRek6PsoKq/tNc9ul0MpJCcfuu6stIvFHR+Ekp/n
X38JW2tOVKO4aOssA4OQm8rPmA09G61II8lDi/GazQQACrRwqYPcncBEEMbxjORR
HyN3IaPvfW3o47HLruruwXMVW0SopkN/bA0PaXdAiMXV6s0OXRtdezKP9u/hZo04
oUSlKgIaK16/Uw0zN/PePov1sPWTF0je/bSvIOd1BE4P9OGaH3d+ZGY0xdQnnenY
BSv17ask/C0i+3ssc78i+i4Rt+5UW9WU0Wcwn7BH2hjItWn2MGw4qpT+GtKAw7bG
mtd/A9H/WTUTow4CWFxmLmIsEEcOtgoEL1Cu7ZcK9J+Px6bA2WMm1HdVnAV7tq1r
nr/00fuEmJIv1Wg6WvfnNctYQEb8Gu9FWdN0AMLglPpIZX/LhdCccqW77IomcJ1u
kubnmjYmz+V7bb2RACda9XRDAUnmv+4EKPbopvU2ETAmxAiYbjl0MF+MPSlJ2FxY
g/p/QQZNTmDXjG92FgQ7Ak0doIpNbCUEaAJRmswi0S6/s8Fe5PZ1xX3S8vh/57oz
epwwCLZGyAeUT1KRH1d1N1bVQsb2smJ2r7y5bjiOGxF5gPS/NJT9PJmdlGJOe6Ku
hsmWn6NoxgdEmptg3TpJkMRYTKCSwlDGYf3QDyhxHNFzAtnK2Q5IhUVTCn8vOWVj
CjSdAARg5mWEZao9/PyvuMDBMCh0aUOjDJiVE8Wb4BosQ5h1fZpkrLhXc7myqXBN
60k8XSrvz7q3alkHzCJo6dWDNZJX+0oVzAt8/xpaxQdt9G2z+JK9OT0nRJwz7Fnd
Bv90N7wvnHc0lglbM+TsHX/Z1v2kixFbB/VNglRCYZEbOwEFLZWzJeY2GLdfNoxF
4KQ4vs6tRoPwFEPjwDTbFWxJSWu3/U8Sd1HnwVbO74HpWTw3KS47DTOwz1sJcmCz
Idkd057zf67yUl9h5XgOYMi7niqerVrSP2o/JNOCLWLg586iFbw2H7S3GYNxPPHq
kI7u1zB4d6YpvfAR+EHzgQkm/aVTmQRM+oS96ozlfa/bWAmfrhx3/ICCDhY2PzWA
q9KUS7HUwb/joG/n6DNxOLLDWnQhXXoYEzUGQT1leIIcl6JQMUg09HoFk7MMOi6y
CG38n1m2DCpw/al/LPNWioUl6twI4/VRBZCBZf/CVwcRPqubHfrVS1kjI2qmR6WS
WUKHpKSUVb/wJAchpcdgGQ1l6bKn1JKqV3FElu6kt1lgldjVz/kKHQ8WJrawrPg5
Apnp3J1hoWOGgryFMQ2kdsRT/qV3FRkfhqo2AuzGifXWaGIDCWNrBOwIp2JSnfvB
0XXaQ2C7nlu+KT6Q1Uyv2jMg47ckAcZFk0HakT8m0aw0Fi6NdLgNjrrWh+uTnl4E
vYkzzbPeWryeQOLePO/x3xnLq1zz9olpmnre4KUdX8QqjKgap3DqL4z+sCjsw80j
wbygWLzoyYDFjywbj8R9AdgzTbh8usOBtWC6ZF/pH1Kb5+IqDaFNgm98YcSbaP1u
2Q8hZGPti8lFKOxQs2eX92Z6zPskd0gwBpz1gLrGRaronSfGzXlVc6ezC/ZbaDVd
lFWST4+kH1plI/qprnVz6jM1afj6zyzHi43rUjS2LWWglYaVZAHG9jGFkJNU8ouT
SfnolbVq93WUdqt4On4OCNDALWKkQE2/bbVYH0HozridPgvVFtdBSeTF+nlOy1xa
m/byLr69nt+HFB18JcHF2aUaykzvHbHAOKW3ch8saRXMrNIywy1lP5eZTBgp6tIo
1e7H1ODbrBKMSxqlQ/9pAi0034iaKi4ggBrpUOJ0K3UAlH4p8URg9IkAoDkEjRcI
WPGxYPXBCC+jxwh2nCxs1X+xJWkFiUz7MlWQy9nyuuazkLREGXCxSjth/ORCXEeE
blHNh5uy1wJjrivVwHBanC/zy1fF79qtznMeYnHx/OqUL2ghkCJ1hkIGWzcHnwH0
z3BJW3929XsznjFXfN1e+4E0l6PSu+bJofFozIa6MY/BNViEiZF0r2ppUfOu6jPy
XbhdA7vcUv41RaIBEWSmt0/r8nGfzJ16Cti7eqV2zlWFOvMMhm2pzsCs/Ofl7wep
LbXIUzy3KyCH/+zaFiCyRYlpy1OsnynKpIOy6mhKj0SFy4UAQDLOzw9aRb4b1fzg
ESIdLBWyjGl/h+1TL8PbanIQUk2NwG9dDlov6VMa6NlvKbg/Vrj/P63ofElDVfVe
aiufPrw+w4IECNss1IrntxqYTWRZPzRvFdZbO6wePVYA3P18Mm6NhkMp5LLCUdhl
OAGm2bxvuJ+7MQ6Fom2CwYGkIGofo2l3VWS/ntn4NkrNXObe6an6FlRQ/TXPTOZG
MnuzWm1hiJL/Fttm4mfxtsn2iFJqp9pIYNLBKSXN7RhNcte/HtrFuL5hSrc9e5oT
EvmpP5yipnl9uwlTqYMyrljJp9rAD783RSsZAKk/GhaYcWWhLA4UszylEg5zgOtI
eNOQhfpOFQojaLUm5MU9a8fEMT/XicwAR76GgVVzB4hiDjkl6PllH2gE1WkTmvDm
S/Z0EYu7pHRUIUHi8rG5pw8PUFMNZFat2ONEA1dqIexuNXHhIirzy22XDOrhV9J/
Zu9GWBfoIRkObBgLd4jOXSR3CholYMkVc9v/wsp2CbDlzicMg1AASieuGI/gOftL
1KWHxnbq6zv6PNiVWtMSujH+oe3ZZ9ww07CZzMCuZpJrrUKuUGGf4Gzr5S50sUtj
QURGa//VgBa3xuYt6ftQEskseZoNP7SpxDLsuqZsAqW4eWS+C5GufUjC3Uo4zRM+
K26FgrtY5pc8AWZHg3NknPjlBIiwV+ga3ehABTTd19lALJZjRFgxFo8rF3Ncf6K4
lDKcv9TAxur+mLgQwjynzLYrMQONJbZYP9LuWD064CVC0VFjXCHhjK+4PjeoJRsd
5xL5+ioVC6Rr2X9fqkLHlRmSEmleIwwseXvYgc/yvVUR8fVBp7Lj5+60fWAbkuoW
yG81AbMxgjZg9JjlFgAJU7cQdKvS8f2O+BIqij2nLHkaK8aJxzfCUwOutTAf1Y6K
QW84ZFsLi1gQ1ElEHsI+A9VW1Z3fBuodNtlNSFlP+yt/vOByMjxjXSMM0TBOK8Hz
Qk2Ceze3WrkWMQaVWF/K0mbhiokYY8Ajb4xB9h5NRkBEjKMDeg6woFpUWMaJVv8d
O1mOSraWRMvzIr/GSza475++NP/X5wtrRbze+uy0YtHtuWNlGeAhXEmmsvm6Ahpu
OhPnoUV23fBPoI1o6aAH2CkmLubUAJLJE3TTUa2m6jEjWscs5MBdAI17oW2gho2G
AuI3OpZk2U3CXXrFL7hdfTiAAGlsaNVyaW1bNBZ1qQe0OsCvoiwqY2d+kx1hBew7
roU9kU5eUuN93B84Fcv8hzRhePz5tcA0ZzvP/35yPJr53mXwnG8S9OOFt5teMArf
YR1H1mcdH326jVdM7GIfSQMVSx0YKL9bk4H9O3eIzL6GO2R7vppnqmzLhmVGMLTm
Y9SlQkveazCaoLinBQGNbdh1vT0/mI86b2DgQCmPYk9xu3MFpjkePZm74p7L8GZC
AtPhp887feXWgN5fVJ1cN3b1c14HtxgOwtbt3MC7DaG7HBkYBnJbhx8q9GqJAaU3
YX5jiUa4weOMZHDSN4ImWdjQNUOiuxLwt+ZNTfdw7Rs2fgg75P/+OPcwD0kSOwLw
8Q4u0/iZA4xhisWVBoEPuIjRklQN7pYaynNOWkAPI9A5a3//iKrHg6Lbv+d3g02z
1JOXk9pTsGRw5SgQxoCs1Sy1+WwdUUVELD27fhCCDr0G0RbS5Dedca1qZpkREqQg
DKwAuuz5e7nc0IxK0PvWuf1STDjJIDSC8rXy7NYKSDKyWJm9pjKjN06iViNsYL6N
Y1GpKhKMVdhHD4/7Ooe/AcgtpWbWfOQLnzX1+CodcL7ofE+Wwk3AzxddrXtgqP41
IDAaDMHdy/0TvQwagjB1g4f1rMG7co3vMWYoibf23oEa4om4x8QsPhXHz3kGEWgt
NEHB0YRhxxx0z8FcxmLlw3ekuVYSi4dSkWmkVriLjXHk8CfXZ8oVSF54TYiaGMnX
2ui3Ricdmn+VLHPUHbOSG/b5jMTuqMDl1duFf2DeQiWjFcu2lfy7CHlBFR76E6ZB
8ZBinA8ksCxY/u4RSuBtS0z4lAptRBUlMxdgRaTy1jsawvWEozXoj6hDvfYnX0j9
LAP257lVZn4yB+O+p5k5Bl2i1rk0cmImk525byQBp1zHcIi03kXsBk+kxNQcL7fQ
rHbIjxnRQKuJrFOCsq/rWQAklfuaSUlPLiw74D2EOXC26YfGxk+zKXMPQa6fju1q
HW+gh040YqkuFhMFaC36a/lpvCa8YgUgo+nhJ7bkkoXwGMwt4Zhm5BX+HXLdHW41
rkLHo+lXBZ1Di6Q1ZTIIjnCkZBehoUnnFtQtaJd1rO/14pu9p722aISBqi4ovh3R
MMxhZh9LciUo2UG1RzbENzSCwoFttCVGAH0RkHE7NUp+tz1LR0ts8Rrm75eTZQpe
aRJKLUPyzoKGejeD7YrjUX3nxzitPP/AkbcXDI1R6t64WTIeeUv4j26UkTGzCg7h
/AnOodLihnM1QhQjDNIuXYNsWym/k/3oQbsYnz+IeVkKpvNMyck9Z1tt9jX5edTk
tJwbomWjsIjGJndnfGh5Ra/VnEJV2f8tM33Mj0ms0/yu5gdxKhqvP8gxEszQuYMy
yNNoMYOVUPzXSzXEZAxczpW08gIr29Tv9rXEKNRIEMkucZLD2RvUXED52NjtsLAt
7OV/ZMnZ0EayYQntFWnOZW3JMf/2bLh5G3VY1lr1VVZM/mwVPJT89JPqHAGoivxN
Aq0mBcGiow7+hNPk70nNi4XS0b4w3SN374lLFrIXrhd4twx3n33bmDswNxqa6wTx
7sE4n8p+cxjxXIYHhZAXTX7GDDs/Am75bM8ts65DTws1OIlR8UMRajaWoD9Hfe0g
EbePe3O+vGHrSKEjkIdY21Yatbfx09kIo/hvvYrFDlnQN+cKYvgb5mr2+Cp0g76E
CHgDkWxd0NVAyElKN367+i52wqQQ14pz6pV/GEC162GmxDEhUjw7sOBCfSpjEmxN
RSdY/ta8QbXoamCMYmsZtAtIzOByv2KYDMdxTfZ2jWBM5Buy5oy3VYegJBLGJj+8
ME+f32oHzM51Gy0XIygid85lFGPElIGHhx5CT2bTAkfN7swRI8/uWUX30v/9bbsL
EQqfbKCV8ZDgfS2XlAbkxvCKwC5QObwGdG5NTv0bf4+ujRMlmp7ATNciJrbK6KYP
aCf6AELeD3zka98mF/nrG0P8Ju0ll3pZadvjHSHtEBCmO5kMAETJyu5bikubGqeF
uyDo5MHjKNfAJj6UZz2et+xgP28nCtvYfK18GKXndXUe/BayC19Cwx82ABRGaVcQ
RsN+xZey/nPGab5OkN7Cd0OhrNqBePftFY8qj3Rrq7ShYBtnME+C1xZXUWAKiPm4
D/PiEGjlhknELTyI9Z9MyBaq+QBqX9o9horg0fsc+zJvSXNGB1X/aSGo5Ll5RtM3
A9d8OlUzxjS4wiAo3JYAsP6lNLQLEQCGcfvYFO2Rjgpj+U+3zBAZX3zDzTXOqL/o
RvCqlffvkHwHr8O6tRZrzmJSPYdpDO1IYfclzXXY+iaGceh6Vqpp5Jd1E5I1JTb1
lwwTkw3YMJZtJRN7UyJWW+Ipa0prDs3a4wDT2hq/H+LIsPjE18zvH5jwVFj+YUJH
NirqDtcMTdQzVr2eub/MJ0Psah9p+Wz/88ZpZNI/0KKcaabylMEpawEFKA3IHCXu
o8pvEdlu34Fk9YKm8Xd83zzUt/MkOLaJY5O4O7Kd3JzvjuYlwLuh4YJiY+1/KwDu
pzY1BBHSboffzN96YJ4vIz4KCtqd33TJPc86MKL5jagr4ujf9/jAegpFmcxDSBu8
dHtlhU/ItYVb6yWIJTG+SVhKMWk7sAy3NnbsSm2eARF8Q0TlIe6LZKFSIpi69IFm
vYrMJr+MceHy2SXBrkupRsVUNGH9WiWis2322n8EQbQfmIUex8Fh7+WeTJBtt07n
41PjIPQwj5T2oQ4cJsDc1aRNh6AuPd2/LGYZ1Vnd5GJJ3F4qpscg6RkT8ysl1ETS
SlIZxU+7VyiOcK6U41CKur5VNvtv6m354FwikczV86ONfrPLAcKcmeJRPLTVokRE
k6ry8YvDaPNHvFMdJVnIX6ZZn8BoMQgMAuTcWtscWaYQItZabx0w1ZXh0n1rxQk5
/77vPTouJ0nuKwLDyykZAR4APyL3CML4XGcSlpzh5WGU6iH8AyMFxAiTyI2qFyJw
19lA08BE/CmkI3aR0yoEFygoHsQhsVvtNt43qkXyx56HzJfl0UB4uLI//OtRQhqN
/uxcmqoPM+TF+zPSldRptNv0jQ1H90sruNjINlyrHS2X3LA6rJNfHbg6kGQx+rvo
gsJeiY4dS8GaolWaARwbwFXrQDcwz8fTRy7VwFvuh6DcwcOQWTgEndZQe3YAVjvq
JbqUxt3R7QwzO/OduEwkjMSsu+jdO+z26SDya63nkv7vjh+ebF75TPCIOj0Npo7k
BLsPoyuzTu+ofpEvIAtpNMQvTWYXSdMDcSlrtw04wt4IYJWeEHzCsfSoh2r029f7
8ltv9m0x/FRbaWWbxSCY4UZgTpPT+/KDAsyK3d/l5V5f2cgFi6xPs+LwLxYo2RFB
8Zaii2GblsnSQWM7CT7o+VDwMWtsPi/+8YyynfRjTjUt9XK9AMDI6ykT5Z12d+Qc
ES8ocf2QUnOc16WVDHOEnd29zm9Sc9bVTmFwtZCDbhjfr+njgDGVNCnJeit3LtBd
2KoR0tPdvNu7kw2wRT2uzeCdprNDDeArdnqtID71TVRzomIlQNoPK5vxG84MV0gz
asf5/Nr6ImWwpqKZotQSFyO/fG3O52u2gwX7zUYNZzPdm6SU8/pAmhIWlk/5d1Kg
yssMt2DXYr9t52o5VLgxWYWqXm6OeDkJt/l4xL9ZxcJzJNcsLVe/gPKvxVU3TY6U
S8GmSdHiz+jLGgLWbo7qq6peUGi6scfnB+3wivuXhZoJK4TVxJJIQoxLHgSVIGfN
+IHDXuVrGotJycK1xqSAcXPTzFpg2xO/1RZgEnHQsOorS9Rq/dCTPnmGIzWEsSqE
wG/cskox4/o9CC+g+AVQZej9Xm6oqFf5kZe23NOyPUK9wI8vaiPSU4M6FLZcNkCg
gydMdhgI+JAuN2x4GlyMRqIutH9PhWzSXVvfJiDIcBPqpHHF83QVpeGzuGOHrZ9H
TK/Pc0AUVShDD/3JpMKvm73fatjuoLiZPxcPpoU7GGqUy3/bF8htRk28YgdEVDuY
f/nzWYQ9ljfCI6ARU7blROEwrZf4ZLOIG4epJofdztkJ2F+wbr29oGtJIj3by2gy
A20uIslKRvpCHTcXOgysMWRvowqIK/waJSbsrWZbTbyNJ38EX0inB5RU7nKZHHir
/KxdH6gSeSDy5J8XHpko6fe2hnqM3SgbK++F3ZMVBtQqETCG9LPusRzV0bO4RlUc
Y6HlwITEmyzQATxE0zTgmmEAO1MBfoPYNNI+6kUFYIh+2EFK3ZVJhKsVAkFNkb0P
sIHExp+Ybf4s0SeDccYtwp8scbbFYx8M9VdPODjIhP6qUkSQ+B2ctI6Bw88k/GlU
KbNjKHAiZzSLME8QrQkLJO5dPpqis+mXMkdRQ5Hijv6/onEr5Bkye7U17p5M3XVK
BuHpZ0tXTBo/ZSgrfMbODqD4H2P7YdqTqs4f1ulTBAUrR2Pc/Z9WV6nuFt54j5X+
XV0iNl2+LGrVp6SThzf73VcV3SigMfuq/MVDCr3tf8j7AKHn3p0hGxipfwEmA8v6
u4gZRe7yQswA0UWjpwBvouLl+RRusSLxZIZrTMPXyaO/mBLsIito63K8/OBS9ZUl
+R5c4Z4diiOMjQUqpKCZgrHPGGSNqetJZ9tKypYok4303o3eNSFqxeJes/CLFfg+
V5e6AND/nAxC0mpp6fm3knDNykOwF8RHZBgyLmDX8hJKHFBuD+18RAaGnj+bhgaS
w2kbsN7980J4GiZoVB7jqFMBlr1Hm3NX2ThopIrbllAibx+2Jqrc34KIzTyxTVwO
Yq6LuxqJ8tW9147CD1uDGpbK2GgqXN4xdRZjgFy3kugtKciww9gyNtTPnVxYH1nM
e858TKdUF1v0qFjNikgyySO5xep42fm8B1B2hdd8JvCLNyhv+o/XDOrxUSsFMDn2
pboNIfz50HIT0gz6XwUkW4XWndnTfxnCGtYRuTLqXR8+7431oLgzMOT7lREWPLaP
bWAmNLSvzrW2IoC2JINKWKIc3fE144+1fC1+Br2LLlL5zPoHytyqVqBxgcGxxiNS
fl9L9Mib/8N09Mog6eaLBAG/wGXD19VCeNDr9tzC1gDKbfQrksxhN9D0xh/yrAVd
Ox8AQp/4Oqm09+pPBdNZc5gbYhGDGchtF2Yc+Hb3qrGKsw0Ro3URlrmItQu+JwZG
aW9j43M0KpqG2kyQrh8ps9k9cqs2oGzB62B6fTC71e3yccknUh4RwBYGcD5+R1uQ
KkdteS62yGj6LoqQaCehGf+a3WB+uTt0GddrF4XQ41INj65XjGfIRMCE2T7Q2b8/
a2rtAksAY7oPwTrJ6UJutiI2cwJAw5ilWs2CTm7TyS46RRdZlTIpVvRtDX3bU/LQ
7qRAJKe0+qJ4AlKvhId+ZucRKtnJdSt5kxITWMlMkgyFfjGiXKKGriQMFPwh8OD4
BFqIptGmXmZbFdlEBkrxfHi/EB3ngt4f0PyTa6FlBqSIH/BoVUm6g/AK273js/bl
fBlZKPPGxPraXOGDcC8BKIQSV/m0WgDsPb5K/V0QXYF58EW+znmb0eaZTy7+4GP/
nSsUTC3/cpQ8IEbbP//VPmTZbITCwYmEEYVwpsSDzxk5EbbRIGpQxqLuAdoEzVA3
JalgAW5TwmwIUNK2tP+7gr9qQBjuFE2UBQ6lZ7IdJDGX59/x5SWKo4c/mhpHbkmw
VNla7mX8rveZnQ91uWxybqdJmt+QN/iyZKY6Kk/eWdcpD3kvorILRHgkuYjZUxvU
iemyruvA8IiDJtV7UdhMQtk6UWzFg/B8nMFCjzJNT9YNH6dM8Jp3krKcEbQH4NWb
gNBAiFLhA+eVTj6xd7v+gRzaZ2TFomNcZmzu5iE/AZ/N+nGtr17xzKf8exaLZ1DY
WPsP9wNMY1/0vnM3xwn33x/3vXcjLOVQbvXk0DtcjTCwPlFWbPggz0bMrNo598wc
H1xIpN6Nag69lpqPT0r6gpeHnhkpIF2w3KFT5wdHC41mWcW9EQebobHUtEQIb4PY
D6lYYyEHpAOsxjFGWOBNjBJQ4CJduNEoXQ8tZ/fe1Tzm6CS5xca4xFKV8M0vh/20
UF7rdTSQUuTbKBuWxjQC182uDob8fJkVi3K+65I87QdGx5/TfophgnD0lPbci7bI
+QBbFVj4qpejtny036JZhs4FQGogpgr1d3LqyffwlErC5vevvS9f6u+43lH9oa9e
URgGr1tsj/Z0EXCoSXIgxniCdcJataL63uKTGlRy3IxXJSkW2nEKQpWBxqwufl0a
jzZbnqStMalukdsfEQA6eE3Ed0gEg13p0uyyBPRKcYps1liJEoisdFk2u5oIjbAT
RxPAvM+Y8BGJGAbKHXHsHjE1XIa0h5rllsBYmJFUAccklyGThnvHBRGolJAQ0ZeN
Y1Z0ZaJ+LQ3+RbLawLhceoUpmmh0gOXy7saYTj1IpE+gywnRlT14msvqpNq6R63R
oNYj7NjaY9Nt+q4K2T0/16om1omv1iHY7kRaeP5kkeXQlLGEhTXuRyz7VtjMeJ76
EPEStcAKQvSR/vqhsHwvy6XODN5QwwWBz/9EJWWSVKLzQUSSJAFygj6HCXhjEwHo
uVYYtoEJI5p8z+GVA6p6aszsKIRawOuyqZq4qysqJUnFKne2vRGRTFg7SMb0II3M
+Lb8JxGY24w2qUYxIgxcx1NiZ5pQYjeMl5zbDgFfoKUY4Lj1tEEl9yRQNKdn3IJ8
8Rx/sv8N6WP5A7JGIZeVuC+FONVqORmKAVGQHCOYvIa1LyCOu14cU3oroRavczkJ
j61ixtWQ1y07bgsmipK55KBwbZqFmLDdCyuLWUYS9n6qe+rPpH2PhsZft5NcWwvY
B73mMwL8VI9/3E6vL5OroA==

`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
3Mq5R+F9N7AYXVc6URCedgIO1J5s19ywXk8xpmWi+wzaeVua6pu1HWm88fPJoVbn
pdFZ79Tqsz8vsW6R3gU46UqkVZxqV7SnB0ekBFY6wsrK0D7d294kUEMPNGt66oDO
GWdHTu1pEUsmqEsDhZ7TrQyaZyoie3jUoFw+OtyhzfU=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 6560 )
`pragma protect data_block
uTvGqRtS4u8p57jHprbdfH5BqF+hL4ACiX9W40xrPjvc/Jhe78zbkxxPDO20V01p
0ht3D/0MxJOips6xgjqKACdxyZEXMGzEQWjrGLsPfHYtuhFRnWL5drG6gMOTKDfJ
PZiIb+VKeeB1n2nodv/Duo0nkC+ahnKVgJU7nimopG4YARpQNmFozYcY7iNBJAyV
r8kEqlKO8cg8mPRsNqmUV7xisnUl5ftAvExLmW5BBX2AITEwnMbrHcbzeNcQG63K
ZvgICcnqMnVBKnnKAjzf2a9WPiS5wuRjPaQsUYjtyhsL3h0X5HsAjLbpYYei5ARS
/WhLDD5TeGHKzXvhgYQQjrqko9Zvs52jQ6W9XsHcTWOyrhUzIm1BMYUw/9St1xO2
A58NtAHsvWtTcZ7wa68pdif7GSXa8J4+p5/vkcnALto3lzMArISlZoWPFWYlxnYJ
Sg9SZzKh150ZVpYxzeoJpGk4Z7k/Gpt0KcFI+59/JJSMMkeOW4afDWGwVD6Qtvdc
qg81z6tirgYfRBB0GFRqKzxt/nI0av0EzA72ZAzD3cGXDw2MK4fZ+Y8AR7poltQO
N8A6F40JSI1o/BwKE6jkm4kNaC9zeEP7KJ3p4PdvyE8Jyds0MecjdnIOXiGQYx54
wOLSACsLxjYcIVqvG/cWep7ar4ryLP6PezwX5IulUJXq5KcxXBUcD2kNyhHFZUnr
Ujj1PGBuP82i4zTwGc2VL7DS1DisWJMiyf8Bw3lRr8AcvQGJ5HZN94he1FxMuGv5
KbaueJow4MfUVMmO2TGRF1LWZcFWn0oB1X0yfhzXQ8RsZwdIhAzOZIKhzRS5htwM
6hJ2LQRwa9hCkefCRjSBquuhpCXsHnlcjhnxG4cIm+qmAvOsTYpc0rhd4Xzr15Lk
H1plhoBYsff/dPEUBJQDFSqfB1lV7ruldaHDUMjqcGwTH3PPnBymg83/u9/GzIxs
6gN8cF5gGi6oQ7guFMNaEo3i0zbzAW4vSk78xhKi3It1kA5RAHzUjTgak09OHSnL
PSIwKpM9Tr82dSGmxezHtorLWiHyyQlfKc8TDs0iXfUU5zHcdlet1yFhob9uqJdh
brTAfCyGymfXjcYD0Va5ZitddvAkq7HAn6zhlCxWWfMe8pMhd7fKEpa4CVftwMiT
wMhIv5PGUyS27fj0CWJ6B9NoZzPa2qcU2/inHIl6Eh8TwCzTl1iRKnQRPp7YWgoF
SW1By7lxoysc9qRHp+0V/RZo8qNQhpwXPLnFPDcY2UwOQyH4IkxvFeOH56FZoVPU
fPOCBrPN81HODg6FDE+GBiFZBJDuA6zo04T1Om5H7yxB75QMYRyOm+MeNmxj5xR4
IUNPOeC/Jc393YjQXwn7hdkw4gZEEHIAtRzhe0hWtnoBK8ySL7oqIfZWOMNUFxy7
Z+YrIAPGtEX7KYBgmPX4w/zwK629JfmcqaYRyd4vnjeEZnku990W3EbK9i6mHvHk
bJmFxvvzf01P8a4dRnLBX3l385/hGeimYYXEEEZLI/ID7ihiEn3ODsIs6i9T+5kd
pIeBQLWRzNr95Ag3xjXsPvg3lxndSMlOf1xys74GzAZW4WPlPeBDQhSXnS0R9Oix
uSGYWFk0PvF3vimf0QLDP37dC6tVIK3aslr+pdT72Tw6GxfqE54+3VcryUnJ5rzh
KRmVmediUy6PglWTpa5U2qhoUHd1pQqKYBMsu98HPPDlV6eUbZygRXi1vFwBEeXv
ZX9UM0pPXmC2xLj23Om8jotsdhd/dyacSB0fQoi7crmT1mVk0uG23GZQHNbK2JY+
0vmBrTNFSUXJxJrYbBpK7+Zi7r6g2EoXXB91fyLy5sbwlqMgLsbkyBz1Saik6sbQ
J3/yHtnGiYcAIVk5/Lb0E422X01JhLit11Tl7uCP1s4Ti6Kh+y03g6tf03Nx9yzI
tGrnRXY/sMicf6+alpQI1iDdZ8OrvgxTb68QxH4I/Ow63NTA11cQbxiT+VcKnKZ1
obolzvM/cH9TkA2pgE5QDe8lG8wIWJlFVy7ddFlK+pbExuy5Qd5TIoVa//cIS2VS
ZfPGSfWaorQDpQx5kmHMw8TeiiNEeN2GeBQUaeUz7Y7D2XtVZcaSiAUS9UIC+Tpl
E73/wPf2uMz4FaZR82XrMQWv1yV6YONhO4R6zl/UgXRZKH+dD4JdZmT7aEplxZCx
4J8Hl4S4g07j+khjhev7vRWSp2ccjvo0mtXVwCLlZ+r3gJgg+InU8OegDspFvLiW
BznjRCqqoimQfFfW806lNNQqRG7PqrLWU+PPE5ev1Aie09bKV+EendbrNoNM3j7+
YYmBUfJzDTboyF23Vzd7vQxWvtotQ9w6NvICJa1vsEx3W1ax9HKyfNJkHvC8kLLc
akJI7sQR0Hyscz4ovlslzzns6sqfz099FbNhEJtzg6Mj7KVrt8/k+QC7BGUXyiYQ
dUMF6uY4Ysm1jI7Alm6Ua/w3OXQLLBHATZa3Af2DfCYCO8xOUUWvwdPDVVVE3STn
xtivAJv13WcPf9R37QSSvij4ytYRRIBnio8GpHUhY0B1eDoD7EYJmCdu37MLxCez
ftBjWTSr+I7B79Z0ilyN3vuCgtStluoni7qNx/nd4BAw2P3yEVILou3EBRqPabnW
ttY1mwuQeYXvQHVJtbvZMnVyTA6/sWtf/qOtomQRjFhPVzaGBrLJttSerUtxj2V5
qSV7UcjAitMoiB9JSfpgH8NuIXJyZQ+e6aHeB6Gi/NOccDm9BQ3M51TRc/afmA1h
wcDKV9VtUz3Pxp7/dn6lkksNao0JJ+TMlvGJhHqYHtHViZVcCrzQeLLFvQdOtrYk
FeMHgQzHuPZwBxBgS1oYoRyWMLlwR1R17WrKx0OkwzcUo/4ShLF6/UTQrZR5v+v7
bMW60EF7VK4TyDjiHNTRGvSHX1JlxH/PJVU1qa0+/vgtIYYR5nLRAGioQ/ac+XuY
+x7LKQZuMqqpjaGvKn9vgFjxikv0n4U3ut67ycOvzUdckIfuasEeyIjhc8KY4RwM
/kO8fRfS8wuKtd/G6a2Q6jmlswSxwJNHJ4MRXwmLQ2QYuwcPP6oGgpjJxSb7wnTU
jXHxRMk1CI0LsGkkO/Rq3v58RnPPsg/A+bSfsnRbuNa+yrCfGpRZoQdo6oHRtO2/
gsDu5Qi//Bat+/tAjkruuM19Zwmw84iU6eEzVtlxC+DToRrpwbtZNePuylyQZ+wc
Y521nb5mGZiFUtKjDQBNt6xI7BlrUUTqUVtdI8yR+fsuUPv9kRTI8r2Q2xm0BM7H
xex0dpu2YSCQzPAavULeg9eiMsFRSa6YqoU7hMsVBYkZQuTFV+rNUa72bryRHh8f
y8EunemD86aHgeIyxXdVd1iS+uC980FZHp+/SoSKplhacwpNZYJa7+dAfahQ2td/
Qad1mjotMeMtN1YaELZ69VUtmhS3Tgy6pcBwvw2efz7o1lnALdW6ngySy+OlPmsn
m6YbLPcz/qNxMbECd22qFkHhI6fky+c/HsFyjn0l4ay3tpPJkXld3kpsJ8rBDWAR
dNY4Yssg9TsKsKIINHStbXj4i7La36UiVpvJf1+/lqFqZm5z+p9LqLkgZOowxIRc
LY7lt/5gY1jCSovyYE80rg3ke/1zODlz6OY7H2QO8TeBAinV4T1VuaYg7EqArX0F
lfCvvb1q3l+Ykc/XuArw4KSuDf2JhN5AoNo47bZREuT3Z6wU24dqTCyYpidU42CS
Dajih3Ug04wt4/NVA2X/sagsdO4uEqMhinUcyR08cOLXH2O+OH99BU+PshOqcWcx
lMoPczrzCT+Kv0PIyWq2E5GkI0R4/vTdC2U8uaLCRXGqVqzFS3cNz//t2Na4aJtf
tD2VOnwnQq79m9siQiZ/vnId53excaM3nP9ke9ZYkvYCpGf18/RsJ8HZY63PJA1m
lIxOur+soRthmyFxE8vvJxwmRpLz+elUzk6cgKlW0OGq+CJ38CNqvQEgLiOZu+q7
UAC/jWYbGgDtgRt96M1qkD7R1gEeFxYbk1dxXP/1x+aVjPTvkz7gn6trchPuvYVH
IlrS45HdE5nyp/emV4Sqvx//n7Ya1EZL62Lpe0pwNgEY872TBpvJ7C58GDUkyb22
1uIiysq3Nd26kLYmms8cVowzxRdOU2zAm38hcMt832pAa3RiVaXzaDTKrLVWqqC6
odSOcTWE5v5uuJ0aZsCc9iNVWA11BuFSGgw90yWV1ox+0e37IErxrVK725UFBCZ5
hU2Z1/0MOYmokJJjJ2xEhYISm5eTfVMsgRJSvEu8wQuA0CsrJxzLjVHzMmHsNcYJ
a2wKlCr8nG7DLKifi/gH2d4Ueg83uiCxY1jkV8ZIhD/KW6BwitDOD+C6nTcL83MW
qIF4inh/y4gWJ54oFQhHmhYgR2RhgYVm4pizs3Bt9utRYpnCWZDA/E62cu8xX8xj
JAwppt/7B+BwgBjK5z0pOsPn+bC2SyvxdWjx67Jpk9mM8ffzyzDZ65EAZAGeQSqv
K5qrQTzbRxM59kQ5oxFiiBS1QC4uVBnIdVlBW+wtseWCE39NN3mOPDgTP5w1qRgp
1zI9uruhapkRpLfjU6Uje7g5a53VXOn/ykIb4eaEZfHEi8tpBI5kkBq7eyLXIb3a
6hwihMI/Nx3SzibIqFOGo9+bKpS9/WZ4qG2eLX9uslYlwF1gxLNLrAAv17Z/3j++
+Fm2Ovq/t34qmeK2PKDdOK3zgMUpORpjPTRgJKvnUTlMtbRR9XCHBxc8IwMDcJ3i
y2iYn3AI28Au30d6DnPil40tR2Pwx9+sMUO/ZD6ude8ggsaV+sXWXf4QBbA/bajX
eJBzR6ONn6XO72Tu9+cRgS8Zu0oFNhgzg6aSlQGziOtJ2dYV0tbXHs3d5p53uyJE
XmcEKj/h2o6hmJF0dsKmHwR4L51jUZipnloAemULlNVmLVnqb4O090O1ERkjNp99
qAuZlJf+wfefIQL7KsHq8vD8PHlzP+0N/GsgaLwzjBViQtSCXmqG9vzL10ZyxqP2
sGDevbPIVPo9nPeAigx47cS4a9dYqFbIDei53VE2KFAmnjq8PEK88kMkPiCYIRzg
1iMrSHD0fkTKkaEzqMr8TauZyfb6ohHJ/m1uhAmMiVkKA31EKwoOBE9IYc6+/Iyd
RqYDdl1CeCO8tKLeEvbMJdaQF0VP4qmahUB4sOiHiVMKcvtFiAnbsIOYz7M9NLa4
VM66HAMflXaUmf6Pdl3IYw//m4JnMWFlOwb076VkWkfw9+il2cws72ipeJ35Gm34
Cp3XcJ8O5XIJucMHKlLvCOazWcluh0cVx1tIRuVamFcaJpJIEYt4RhT9cNIjcNBu
OElSQdUQL0yRNxWIx2YaaoTHsI04jqd4NGKWbCV1ZjC4fuCXaEyqgpLZti4s4DhR
3XU8cJc/pEHLtoR04lkfxYp+dT0ufpeRpus/GivQt3tNtfBFalmvmAFRF2cHqo9B
SfC23zr+G3sKfusE6Jqu0awcxMHokCPSGfj5mV9HiiMxxifOvwOZhqjzZb8o/lPB
bQr7v0/DDMNGX+QE9CtaxC9rq9fOh86FwNi+E2N6XnpYrYrqKsRy/CJ5JYC3H803
qDg6exy1YDsyQOfsvcOa+UZoSmsuj163oBfMp1t1y861SnOw7u+l2cyq6yR7pkT6
4+tzppqlk+1W7oPS8Gc5K4qFQ+VkIyWpffcMlJMh+EUS195EI4dwOQ2lCY0hWJum
q6j5kWvHGCpCXtyPKIh3Z+7j70CiFMgx7wFSpJxpops2epNw2/H3H2DwZnKoafZ6
naiN9w5gKq6SgRMZ9HeguJUZ6iFXsOt7Dtl6pAFGxLadEFnjwgNhuiAPI3X96iYX
Ode15vn3vsdCxcCcmYudxYOsR7p/g4pt512R3LWmtoqyyelL7TbFhfSsJHWszrZ+
xAYn1kVA4u7kaMdg4zScHxMskX9wqe58YtDI0jzvx9C9mjYGrjEAWk3mDGBplPeY
ouO/4oaIdEhoa4ekXcg4OEJKq7b7DsAMYQusYwnVt8LNjlbeqxZTVnernDteXe4j
yIcng/dkwDrO9yleIh9WRc3t7fc6IbIOUjpAARFjIakj9Yc+pWLdniBe3rYSlzZy
3JZBQW8BeCSI0RT2HqAt7Xr8xRe+G9rWIcLry5woyPCjcz0LQVUPEoW3hHc1xuKW
fLY4rnoKGM0tpVUqcrv1ylr54zkszrhqUMy6MXFD/22wmT/URjQchmZ9Zz3vrwGE
bIFP7BEXmGt2YgZ9oIL8t86KrXURccAtTPhf51U1h+GuKTX/NH2sJ/d4X0CG2whh
Q3gETwvhySchQxmrVzSAX7+gIuFnDRZ5SGm5Hy2klsx8aeHFj/3et20Rqt0YjRna
olLOUjPz9kijcimmjQjbN5MRF5xttpctuGUcZb3qZ65JwQlaMbKexI1a2vNR5z/H
aIwWw69EhRxa76cpUBzSnLqzwNVlsZqL18JQcbW6O58UNe0gyx4OO28hvoRIB8bQ
KthHN8bBca9eurdto743/SzOsN5l/tzorqhz4fz9jPFZ59gzodfXkxGq3c0Fni6F
cqiBXjXLiOEW0cv1bIAFUnbSQUx4319UeKtkzZt/yu65rpcoauI1OifYJSOYMPaw
kQXm1h7KjdffFmhEu+2tMUBCM9tjHHparzB+MvcOl2rjYfTthMBCD4gOu1/+tQJd
Ci997MsNAk0dKGUMnC6WGTlxEgHwQ4Hj5MgWtSK8rdjo45dV4RoMc4sCrfnQqr7W
n0Qlwn99hnXam0WNAEbJTwXwE/QYdJTL6ZUDha3ruOsNOom3lTvSlfCm9eOYub7R
B3kWls9A3aye4KvIfcYz3xts7zHRsgOGeCxrkRij4VKTp9he9RSnsddKPgDYCIvT
+1b0I2WNKjmZ8tbsWQJze1O5N2yRvkCT+upFTfXFK2/QjqEDs7vFkB5EzweodRkq
DF9EsTqa/GBpWk0XPVCI2gGBotrt988t0oAA9K2BJL1VqcFag2VKtQEroWqJMtkN
p7j9mbaGfx1M08mQH6t8F2leuhqDjUok5SAa0sUmpfZlk60G8W8Q0isHQ1ux4nB7
tbda0jbYG02h4w/PnqbIs059Pgr+7yG/hILPEqo5qIRU8fj+jW4Oka/dN7oJFIDj
eB9L1fmvG7nw7yNMFr7dAbFIhH2VavwsCDXS1yIMzNPM4WnT0jwHosy6SME1mWIm
HocFAUahBYLSIvAa4sSPPYUKLbxo9Qfi3hl/XMQgXQvbHPPOexy0/WA2unIk52A8
0GKApLr5Z8GQExqiqiFm/HsBc9zeU+UnqcCo5PN4yegZfwd9WJFdkxdLbUFrFolU
/UsrplTLxYP0sVpPYT/KPupMujHw2ULxOcJZAxfpfwP+WCzAMDculaQXz1JscxuW
HzVs3WfYywacwmgr+vyTwPrI2DG1NiVD/3TXGGMyucjRAmCS4Rv1Ns4xPnefNpgP
lZYA4ji5EODmilq93rfVC0mRgHwVUN8oSDG1O9ZZVKp+Fn25BYdXQR1eoRNW3qOs
75bmUHcpQbp0UcuMpas62DHJIipJyTeHKlGjPumVNYasTHUHVlsKhyOtdC7ddWrw
pJoehEGCbxWIm7r6WkUH/Cm6IsWdrYDxhB/yD3Z07JaQSF7wv6XTPnk3e2iR21fJ
zNlf5XgzT9xDAglZzw1+utHFHn1t/Q2hCLNNQE9nhvLeq5j6W8dVRd7KM+xmX8ar
iwkk7eA8rW/AgVcK5oy+62RID/RtgUM9yPkF5zb7ClTZeuSNR+Y6hTGCGHbKi0Il
sOmB3KR26xR2B0CR4tWK1U+8WXxXLE1TVIsXd3qWWXyd1FV+y2ph4LMNXyIBVsX/
BQYFj1Q0It2U3HSRDqGW4wFEW2Xf5h+ltW4BUEfpctrTxO8UaBKUXzrTQsw8HmrT
BOsIPkP/rc6CbPxLkMK2KEPh855l3Aml8qnLteJzVc+PcbqiEAw7ixXrmS05AH6P
apz0MkevpELYlszxzgfseFxxzyWeS4/xpFsl5hVK02SbIRmc3Xf1ObWk1ztw+Zln
i3WRkhewgXxTek/80s1YUoQQ9tV+Kr103W2eyXd4FnhYxxTgifKxyUID1BEvCu/b
idbuixjZSp5wkxHLpVwO398wqSqiTka/Gu1FC6qzDInA0NAFEYhDpkZI/ZTpmBHP
5J4UurKEslLF4HWeUkb+zDUAchgagn4+KvwjqoV6Awfk3H1hnBdTN1CJZd1SpN2x
kcNKnfpkEnepQgvDR4YZf4I74Efflw0el66coGskL/K2urlIVMAFcfuluGM/fpmr
KhM1rz4Igvx5AcHKuRZyCztn5k+rBd8tfFyOaOV5RDHATxXXohpOoYBZzA8m54E/
+sMxVUsk+3zdXD/fgG4LI5+f9jscM9Vp3r+ExpnUHxeE7BqwqQKUDlAHOc6DzROT
x2AfwLAn2LThe0ZGB2XhCIpQE63oDVNeix0eb0waxq3/5yrJAP7Dp1ZjsHuONrja
CAE5By3cBNzyKj45V5r9kAp88vNFTjsQ0YKKGhidlUutLe49r7b3pLqpd6z2cci0
X4hkyfVFFM13IkIOCtd1Xzr0TwYwNs00zPT+msjZ3HM2vUQunJAIMpHvJoWBh6oW
vZPY4lmtlhwrJR9AsSVwZ3uvT86cm6k1a9K9iK9VzR11nnOxVbnR2vX1WnbV35Bd
om86ysajf/lThEo+z16H1v/JtmepyBPSmwnHs1PwN7SeNrJKXqZUHWI2k700qITj
EuqcaAkGPXNXGp5j/GI6UZdmATkRRHKwRPqg/uva8M0=

`pragma protect end_protected

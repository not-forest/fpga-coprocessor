`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
EiONMIL9RPgWHlQECOJ0nGxoA/1/9wzJVt5bvZz3Wipxu3zw5H5VC144WN3yCaha
jMojW04O1G3MvVRGz7EgNX67apaZAdNJ/iFt91M+CYxSHLsR8zvIh8GBtMV8vnHZ
HeiDOODl3VtotG1xO+nhAv+CcGjxZwZ3swILkNz1vxM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5072)
TxX83eJJPtxRCsdLwjDItZvoWsaYw7cVOozzmmfMT/dXGXkAeznfvQdG4ZTL9nsN
6n9jy3883j3IS9IK4VznsQvgm5a/t+UW6YzNGWfWijHXlMcTnOOdyuolevCVeyuO
Y8OvM1XJB/L0+ip+mJT+CjiGqEvtWtEX7DVISAT1IoGV4aw1XXjgApI9yCTCwKSq
FDqzSvzUs/Nu4Qylj36/VzIlkJTYQMOV42oDEsos1qxsXjxx1z2CdUR7TAPN16nu
lB/xLnbR62e28Bjkqm92Oo+jZInIC6YF1JpIVuhfrDVrWAdslY0hgwD9wZi1/7H/
d9eORBzvmF/fhQbwte5rs0JgACflV73R57cIhmdRWT9Kj01Z+6oTX78NYh+N4qLF
QjTxNC78rbRc85Vlv017q/Vs7WDn9EC0pzYBmkjM1Stsh/qRZj+MjFBI5ti+Sh8i
xH4Qtk51HaRHGXT0e2AXDMgzy7xr2q5PXwrxM1k1LU+Lc/3c83PtU00s+l4aheiW
Ao43jlJz8DwjCPIEWyjI3Wbe3lcOXKl5FP/h7JUj6oAUzxFzi3awL/f8/aiEyhiq
STZs+dvjd4bkq2r0yCBPhUUP3LikeQHEToqKt+yIEQ7dKg3ykxHI/7aoHuNBnhG2
NLkC57ZjGIfNHzhFvGLY5WaT4XiIO8nZBN3xGCLy1d1pLhT7+UA0uDROFFnMF0Oh
FOoeblXzrXDoIjJz8NG4ZQfox0IqWUGduQ3YyEKBU4UxPzN067OgvaXaG0ca6y16
f3OnKhfZBXCjJ4ar1izjAQ8cqXeOi/iqm1H3TikUvonv4RheK351yKPOYdDwvPBM
14VhtZFRhY12GIybw983Up8QxqZpdTeW7v78lMxeUaS+iqE09vA+7yFuy1et6rpY
JNxMROkLWPEug0DSN98R0uB7vxpwh+T/rd1eT1gpbo1ADab28CzcAuC0VivjvQb+
u+GA77+Aj+dizZpoPBTsZtG5OqGZa8ZrkLzOUYmY5LHrbjgE56AyUGHB1zoE4/GL
LqThjjwHtSoiea0RG+VovCaxfTaG+8yYgh4NCxVpl84DrPcuSkRu/J6m29A9bXhV
6/DhvrtEHfm6HDKAgtOFruDSWSWrq16oRG2t+XGirhI/bhtymefLA9zLDiwjZUDf
PTc4NZDpdlFtubPTe6IfcvL2r3L2bYWeVE+wl3G+v3oJekJrmY3W9fN0M8R6XqWY
Z4FQcTMBCWp73+VRcb0ZxZXKQRuunRuakghQG7j7R1P1h1/I2K5xGcUfJ7bgkwZj
fC/fuaAyBTMoPZVmM6Ho0o04wcq8OBX6PJU4ao2sGdjr7cU+xRwNKhJPU6KfFNPA
DqjVtIpqKa/9yEqOHDZAkAAQqEmIGmW3bj8nuJ4RFtefXR7jHasDMqeYNbBDLx43
3E3My3tvNi2wz1Z96FXe3FsPCRDbBlKM/2eZYR5wroKi3gYrQM0UEfLCA5lCBhmk
mCgGpxVteFSpMoKMCTFBdDqqOFDq52dIiHxr4j32fKrnL+CttljSfWGhKtCxSfMD
aK6q9rfZyZbJnoYgT2VZ9FUdweG1uxJWGXLhmkAMLQiq/gEeF/4TMRFS/iAi7/1v
+9o7qMMXRBy3+IWtzjERuU7B6qhRjslGMB20LOK64tQEvsjJf3+3o7O7IZSe79g4
EemG3bZAgV7v+hUIt5GHzwi+zJpjp/Z50lIhwri6uRSm6UEd07/qK7JcfEz3oXTb
uybAz7OhPyXD5H7Kzvw8giFurebDCl/0N6Y1wrGMGK/yMIWy5VSbKwSORCfKrArT
1/jPDR56fDnZrp+lC3TcVwu25YIG8zmrBJLHYxR4LHObphAGC041W2tW3rGlraBF
fWr+kzAm04JpmgAbd02Y5UWMhFQvdLejbKkKOb7Yx5duM3J+uftv6joJV5qFexQc
20uK0HC7Q8nH2UdOLIMRDRn38XmA8p54dqN+3b4etGSDBPR3ZIp9qu5P0yBtiuQl
eHfpcPekBWh/ezgUdckcWFb2ZKJIR90HIK3iJ5QmRXDpsllWFIsmdxOWUfU3M5XI
eG52hzifdXqZ88UXW91lZ5G26zjaMZZvs2vbkULdO7tHAhWNQafgOUsYTPCJcttB
OX0I76blVZg1jFdqegaXhtuMu+5R5lI/i4i7XMcyRTnxmxBX5hylU9leZC55rebD
75cAYH5hcw7Kvsr7bS7o80pxU5JAOCKbB/vqM8x+tEx2WoET9qJZuTT32FJRK0rU
F1mrlMFcaOsZCw1pbQvCAcU8klRupCZpKOBK2jWniSwkI+iFYuFNE5Pl1LFyFj7h
Ihk3lVuU3JAK997w5AjTlgcv/0AONDRU4dWR0EIA5R684YV0GY+RjkASvLsVz9D8
0+nxmsEozzXvm+VQNeONFof/PqML1m/ATkhy522G8Z73QGEGFopeLaGg65rjRKLq
Cxbe8tJttENSPkTAdjmw0BDic6ikkS6vOUdd0dxVCwK+q8aI/n5BITyrHYMR8Iwe
92VAQyXATbFyw/FoY8WHSia9UE9JuA8M8qo2Gl0lUpG2iwBsyLkLXJs5Hri0fCRR
5W2HTrGWfipd4wrbrmqp3+lKaCU5azOLyonvdDayu2PmDxJYYEy/WS6baq8M4nwy
UabQJ0IgDhg4AJjGszIH/ZfObSLceQdA9GGaM3UAHeDkli+jb16E5epd7bjDbZtg
m/2cr7vWbU9Wph6Eiap9Z9yh2k/UxR42hg5Vx/7neNnkRTa90MA6AL8C+EUomYZT
S68N4zFnshB13R9QB57Va5O1RHrjncRqZBJjUF33V26qtc243pzKNVyJEvlvJGQV
BWVzmRUxaPkAZTyQDAUpHeBqGD9/yTmEDYTlCTaB54d3SjtTdN0WbZFv+sl7afYW
/kzep15qxI2B0m4L2lpsdBO5RnWu6DFMDhNo8GSmAeb/LZBZXvCtKr4rPda1XHd2
DV0/WRqKL/PDUVjFOqgmxABUTkSD6iwA0YMxjL2wsP4cS85rILEIyPH1Ry4V8Dqo
aq1txacn06UKeGw/AUBECnvHMN0sDUuqwRsTXarwCBqX1CeH5hNLaAIHJRzji3e3
PqQFmSqvCJNcIhh0JDHau8gO3S5+LK3HHCj2lbnH6eB55V28V/RAQIaePUbbxF3R
rneBApS64nnC7TlhVpxkCNiMy/zx2EeOCXKL0upJfn/+gMZqPerbXUejGBSnaXXg
+dD/hycNJ8RaW9vE8fIOIPz2/rDLIJSSAp2cI5jaVkmkQus5HpKt4qngNY6boMbO
ra73rLJw/S52Z9KlhqnyosSaiNd/vPyduSW62yr8VlEBQEtiXZ6BgATyIr8ZCZQX
HtYsxjZZXMXeibv+vg1sD3nZt+tBWmYbgEvI+DzVWDTD2L/3nhVGgaU3dpiJsNtj
RcOJ7bwVLNb3NC7gLuqi8dLtcQaIn4m1eHAMA6BWZFREO+JyPI1NqAvUbNbl+VDz
Ce4rD6twBptyBeagyy+E/SRLGRPoesme8F2r0Ws07NwcczAi/4cOLtfJA1PymoD0
TcJIqt1lkVW+9V1rg9h3s3i16lplDnWRVfRTRmkrsQUudtiwWJM1xUbvutkfM6fn
X1QaJvknbAudAN3flZnTYTDozRrPZ28Wsg3UBv32Dc3g+Ic1ocjQkLAwhcdxQgV5
muyKIdFq3DQN/uFxYRzdP4qhqSZWBqeiv58zO3xUA2eB3ehbbhDj9nSfeHhibW3n
o3ev5oDqYhL72ElED3CGaDmiC1fxqL87mEKWnN7X/opNFtoZYpX+ZBm3mPLWM2LR
VJJw/Fdus/dTCCU/YoBqXj+QlSF2+j4eWMmlxePVdVEJ7AQnZq77bZPYLEngd8ED
A89M2qjjdO/GnIR1hXBjrRPQKkvcs17ejw9EjsiKTlPpfGbMHZmYsD22zgzJYIbO
Y4UCRN1e7NCnfuLTu+X6SH8bUYQITowjQROUxQ6XgFSpqDdLf7QEgP7GdjveSSeN
v5CVsz6ECA9TENwka2pZ0GzXblmA3uO4NlZbzxHoEZpToXuL/cSatTpQcdgTAq8u
7vNmjOwY7wZAl1nbh5JqLnGmAycCvdHc7NegioY3ZXE+3ukBJmcvH8Q9OE5uvp7J
j4pyhBBooPRIptHdM07zVizRmRwsGzW74ZteidgfYbGBLC3vsJJG4RJX71TWxrfy
j9v8FVeUHWnCuE1/ineM4n1R/lGZJB+q8ljqRABfzgnlJipoDblG2GWai3HklNZd
pkSPVYacxbcaPZzloxYzOBlC4Xalw4WNdush/2wbuIwUSVvp34SCPmFo33fPuJZV
hCFr9s3sBNBk/FzKk7I0Bb9VAqhclmpYx8csKElzJUoQVJQH/00svGRlbe/ysmmB
jma5OGnCtjk+ke/Q/TArCs2AelEu1cKJVXw/q2jKrYci649BGI73kiMdez1eWD3J
HPL+RaJjfz0Is4AtAqLbUg4qnP35SUVq90WuNSX4x5uZtFf+EXYMrZXzXtypBW7L
sXEccL/pAGQSqusDsnLcVnPyc765BO+k99i11uiRqmmxxhATWL1FHYPai0MXGjjr
gH7KZanlA7ecMRNMUDo5N6zIRVniKZKqYOT/feX/df8iBOWZXkoB+bS0XkF5bGFQ
uLKoucC1V90vPg1gpmB49PMWc049lUeEgYZfJzrgKt7wllJfo2kAiwhnfiTF0W69
id5Sl7pzRxN+TdIZXfPGCtoQ5MPkc4plEAsuK48egHuDPhBf7uTMW1PWaKx7ZS9L
NV4YkrSJM7j4gk8EWBm7L5novMXVMuBO7ffq3TwxdvlLPrAlB7T057EyUeR1JMdp
g98DyJWfniMZ8eHgaHI8rZR/jFX2lX/zuGAb6zuq8LGuagC3VdRveG+lAT6t/jJ3
rbT4kSxKDf4RO3dfD9mKQOnoNKD4ASNDnTiw5nZiDCxvb3L1SNAsMQSSA/iUPQK5
sdl2VOTRdtme/NwKnU7Qv8olRsSWGIdhrokI0H/NDuQjW71vOITVn02+VqweWVdF
oqPswStQm2uhMH4siGEmy4Wmy1EOD5DF6IrLqsWj5BNP9mjyBLMxSKZv6bS77Kdm
36QsV9nkNVOHH+SOTj2aoZ08Aft51xXRpKj+U2/1/tO/gApRaPM49aJ6LUfw9XaP
77DoASMUYQJCehqfOLvEumOGz7WbRwaPrnKoXPeNGQwZnEKssAgnNAJmgJ/T5Vcf
ETdiPF/CvbP8Hb0esOYTKPl1PkYxSeuXr01RfltdFNA5mS/kRL64dTPwpQsuuR6y
TRUmeR8pmxcqInn5MaHQm4cgExQj6mA0umqxNw+PXu6NDdGgCtkm5esNbHUyneVh
mJLyvV1H3xoNpgEX2xwoUZ8fMf/vQBz2zkks8w0XS6ouSSSQ9vIkofXrQnvExIEb
604lOL9AR/NAJbFrO9PUQ7L4Q/5iaOsP3QD3zvPvvIFrvNE6SCz2cCuVmKo6EK4e
12odjK9+F6+694yg3Kw+czYIbJuPXaEt+riU06Fml4A2jpc7Wp38OYmqlOvkMTp2
pJyYXdaUA76za2D1WziR+5e28nRqKLf9FywCq4z7QkyXqWxUvDQHftnc3tPGfm/c
Dp5TDfl40ZAwZJoUvfcBgz+csgsb4CtMp86SO7vpSmD59n1sL4ltk/MzAisi19Va
RnrOrpKzMtbWLeVgSfI1t53fdp1XepmtK3brjbgHqAq709cbu1hWplpsJosZ03t2
ueH19cegVehN6ljlZ8Iz+1Zck1vJ2Jt1B1lig57KkjkWY92+lq3ok6gyImCp1o8/
49fjCBWkfuaiOwPmsk1VV90x9QA87KvJu2P9R/srIuu4iyod2naMPowgGiZWUmdy
bNO4yd1f5rXM+2UbEeepATzLKKGJMbBmPLcOypictnoFKZrZoLi2jMheeDbob2UB
u6AUW0TnjRF1ZiAVAuwwWpdI8XcwsqqLveyoI7+8cN4AvK86u97HA6mxlY4Di93r
GWiohOKgoShy27KPQvvKHuK/FcYZrRAoCUaEmtfXqfkT4QFta44bOyLl2JVrSxu7
EAbF2UXLg1W3QZhKbu7/GpOLVQ2Lv9j3tgFnokrMLU64n4dsdq/mZIkT210V0JBq
0KnA0NVXA7aZfhSfMfecTioqDyuUTmHY8hiXuv6mN4ebi47dGVsDc9cWgExYFGCt
cY0DMfbfPHtm/arrT/X76oDwwufRaetpKZtEuORVyjIQcYbg82VSLJUOKl0hUD0C
Kjnb/37Vfl4Xl6Mau7twh/2s9wmLmrfDO/8jb1h0MDLAYvEE7aXPbxsS1ksE3xkF
3FfElFR4RODcPp8ClggGmuQu+WXq0QMBgeKo+q0Ahbby2YzSrwRJtpkQy/UqMW1V
XemE6usfab94Vs9E+Af//CQBN+lE3dFdXd7b1KIA2TRN3KYWO4VvujqeCNWNp8S9
muRNHS0njh8WqWrb7iwyV2a+T+9tapHpvHQGTI6K1gSA/LqcrQQZZQK+Pv0XM/KY
X4Er7MWD9Seai/8MVb3G9OsrCzSzr4c43oUnZuJ+O1uleWKpFHEQltcor17YvDah
izewy9XtdenXXtgow8mqbswCm2HS9ROwh6Pc4gv3sXcw634loWQA1CeSquQdhTkn
oYjozZWKjS2cCO8muvBTiHf6ro1boqv8RTJzaLbthlXhVK2337IMbMljBZKzxNEl
Hnpv0BCVYVo3nawVcwok+GqO5zRjSs3Myb8Rv/1+Je04Hj2CKWHbf/O6IKqOVGpi
Wc53bSwBha1CJsYGKZMeQff8ZaEA0c7CG37e84rshpo=
`pragma protect end_protected

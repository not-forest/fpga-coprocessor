// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
BpsqmU1KeYMnBC9yjyPnx5V1UhU/W3CZHZ0XkvRQLpi1dgzKAlPPzvhsTxZ4AQhU
eWJnV+ZYiEDnT9XsbI9sKc/k8SEgeCepXITZ52wKoexaBSRSNHlb+Rju14nUBb3V
gmFBxwDTw00yftF/VfrCiULcJvqe2BqpwKDDGiWQTRBjsyBp8SVnnAmoQKoeO0+y
RCQFYj0yT0bzOK2uE2Jko79Tip4nZEeTQTRjVqGjr8l9lmQeyypMn19i+L9AazUK
fNQsXt9/fxBPbtAxE4VZoNpaYVEqsrIEmxz9BqcfzbEuEPBuIOJ8dTBBoeC2pdte
8mLIqyAQGbqyv5TToE8+oA==
//pragma protect end_key_block
//pragma protect digest_block
wtRqgFwrIXt+o2fcNi3oCh9QA2U=
//pragma protect end_digest_block
//pragma protect data_block
ms+JP3BgQC16c4Y3Ep1V6ZxjQNfJVO4ytsxEoXyejb+c1ppcGHu7/QyRAlo7kl1s
XQXYPObVq08AvXix2VgO1BU/VP/0ZIt+obnMMnaTts6J5TTd42O64uVmZYmkw/Tj
JOvWh9+7rh7X+sQ5YtpinM8Oc/Y3lHpdsxBJoB6EtrL/WKTf9loyP3QtdoaK5/Vp
5vI/xJoLeOW/SOHEp8zQm/VHNIVd9nZmJN2GlNqU0v8yXM0XGWzsyZoQl8nrwaMI
Z5Jw1Nw/mCodLWo9HQPGvbHxDCGTo+XP8/KLuBw1GASUM7v0GSFr7V7qHr3TLJQe
32MqjnZ7/LzwE4JI/TRbYbwyNwQ+haE2PjWvqxlYIsQcnJxmbJgfczUzRjZiDrS7
L6QqsP8Ys9/odr70YoCb1ka8waLVe+PHK7rmJPADCYIz3AeFOm+4D4S+1cOyySGy
hl/3hhHYBVdrF1Ozt/N57Akmwu5JF1+qh9Jkc34+hltItxGWA7BH7sFGseZb4iIG
5Ds09vUDdkxEu/H1JeD2RepyopOJXx5yzbN7Mt806HPaui9CFg77BdGoovb2+Kzv
reRrQXjVuBm5J8l6XyjxGuu17jaVVDm9wp9uV6evjrj13U/vFa72Oui+D8X7v490
aQsRpBI5eZapay+8pLDqdfpExaaQzY2hUCaGJ1yld2zE5oqK3F5MpwK4R1AhgPx8
AIZ7FVS152Oma1Ps4VtnkhPkK/j+I+dhLN7mx9p/60T2NfkEDqvGcahSy25G6arp
ywhSBB3iQkwVhDfu1LipWGsp378ySTQJL9MzbV6ERaP3MAyk9kzSwyvNEn75M3T0
uLvS2Bgjbl2PM4Cox6YQivG5RfrfqHQyLjSet0ufLiz8YfSUL4+9MehMXWsvM8vW
7XT9n3159hq7SPLLh7WhRx6FZ4//zoRpQeT8BcXhNoVM5Zej3TLpo39mM56zFRN6
oYsGFmf5S96IqCbhUTiZzPPhLHkAh72czuKhrLKMD4r2KJj2HtNpQkYjxhnbppE7
dWCLfM9j8J/TCcK+bOhwbeFOsPACIiwiuzbfntOZkXeW90ILEGfuvP0lJq3sLYTu
cG6bKLG3p5BXAOOXomHF/ncESd173JGgNINWuZ/3XtWBLDHI6XSMO45hgNJIKtQo
/iUQbSYrKSBZLJH6CVJ2UFbpULTzHeMFFGBiswN2fa4q7axYPRUf7lOkhUQ3ONRI
XPDZhiLy893iWQbYBjLA5VKXRSLgWH093kN3BkPbpUR37uTY/fEaxQVpWZwFxLri
dASPL8EC5PhEfo8Z0QX8ovbIuuy7kBWe7iXxYCNo1lGfzuCaMYtZhSKMdf6fC5zf
Bl6LtZpKRCsR6AbeWbRPdCa/m0Fw6GkR0bzkx0ZOoG9OdW9UJE85arwHK4YjUmHu
tejSPDsyaikwWgsx81BdnaEJg7k4XCmu/y4l5z2eVbpYzlkWaAPcAzW5w2zw+dZn
c/SMrNx/LZnD01ybl1mjKdnegV5QowTwvswTF5vQskpYQVLA2eJaWMv5IJuMl2KS
ne2Gs99JCmEC8Za49BqNWf+m93siMk9QDAESZYvNWhR/KvjuDavHTGsw9kYLp0l3
EAFe5usXT68/KeNIcynghUyh1lrFdPKGECmU5f6bqOkz3IldgDb0BcaF7rfJO3z7
QjBUzTKmWromBJGZz3aBFOlHo+pAsFS1KGEVPtGr7vYBnsPNjMjl01SyEA7D0pRF
WIOBgjffoBePEv4rz30ptxaQbZ5CAAvIE/Ld64zGFL+KUxVu4IFkN67OgZvsqIhU
OsPleC+vLGEw1APqkbTSEQKpzoefntWqXtyWwZIu4WYZDcyhg1EG6HYrM4iVP+l+
FDuRAMWakFKn+X/iGQLuWY8k55RV7YQHOLs7P898oYUIdjsVbp5mQmuRGKRO38tI
dob9N+eWlIoeD7wxsOCPWyWmvX5xbhUfZ4tVn3ul3+cnq8VtImANB9xJLoBnKL0m
xU+r0L4ae48SmcAzyA1MGpFJ4RCeesCtxwEMcg4dQSZZadmmfoGuBwWqsjdwWJTj
RKAHEE8jNUj3T5eF0ThXebjPdDUeNhni0AY/BQioZPxLQ5NR7aeEsxGbkLTAHYQ+
unuO+tbssV65qacf0o/NsCcIYGmTT5TfjYED6JxTmxDk4nAiV4dMs6LkylW3kG5g
Fky71QjenuPe7CEi3Ryb2rEWH8d7bLOUJ40hbvsq8bAI9NpCfzTnOlu45/+HISk2
v3TubeYjP7RDJVft/H/7cB9jCyvKVjz0jhVRCr5d7Xe14A/iLbbCXYZHv/FJIOsO
HpuqmVpZDJccekjCXt3hTznS6hARSxYU7VKT8+R+rGSXmnYQOI639ZFa5Gmb7egn
PNXcW3Dop8NntnHx7tC/HGmXT3CKhON66T2b5EVKS0xdNcv3iAx+iSAKxvoT2G01
7/sNVth8OeAcHytLcQ3Dh3pyN9RicfoDX+Vkp2HJdUDylXRgkXH7tfJmtpAJPauG
Ip3cNoStn27KHxYFMnYJEwqb433PMee/7a2ESBV1ZTpb2jmRefLPjkvlYFVu8A82
QCAIjJNsd6TTchNZMPO/1OX1+e19lq9NbcJRnilxIk//HHvMkLXast+GVhki24iE
vTxD2PjdcTeLetsE/judjI1xktaNFokpvilDuQdXljkfRCgaTNqMh8QD1ytNO2FE
+tZcs/WljyPS2tysxstOaKyUqwsV2MU1P8EOGANmYPprIa/CnuQ0uwzjAUbuuHeK
9bGrumlI+q5Z/a1FLQ9lxrPhn4zGiYg2MEn6W3YwJ5tL3nYTcHC/0o+xHhHGJ2+P
mYCchKy+WwURuSO2JzjIN2dl+umK2TAWPXA5CcJQ4cKG5HavPIDz8goP+WvZ/SLr
Cn24L4Qww3UyNe9KDRUOeWcuXoVMWiNswSGIhew5/U3tejPctXMd5WNkuFbK58Iq
QXZofabCgsMFWqlbBw5a6qVEagd+D66yN38BLASfide3tdt0OHnogJFOuIph72Xy
YdQtTbnK0fN7O8JQu5wi2iPJsZmX2w8GuKCEcLVdm6Vi8vp0bfGWnyQWsIILO8dJ
XhlCULWgLganGcKOK34VhcP2Hjgit+3KvLbeUYzmu36lKQ7ifAg9B1Zn85ZuoX4e
7L3uOdR8R0vD7+Qg50vumNRCXDLFCjOFyOJ484q9eHVpG+xVdjLHEqMzID+jMu8G
PFY7gPVwvMIuMsYFs2fas2O2wb00t4+HQoWGzFMgsraSQBqpz5uovA6IZGeHQGIq
J6ZPAUeG1SCFH6jD+gdqyWqAUV1ZvUOarXJkDZwgbbyemLukkWj+n//ugPFsqrp1
duMYcVRIXji/v36Hb9XlGMKHn7k0ry0/hUF2WuXgfRmtDgRu1WJSNa88QaUL/auW
NBxoPPRbL6d7LiRc8rq1Udly3Oj/BS+C/OI+5tMoGue+2lDb/Yh0+EwVJDrkcHWr
3Q/VJYQTvbjljnaizzE98g45KS68bJdkR1qWWdDVnsiLh7z+OMsE271XS4U41SkE
do+tqCA9nErDWqdJzqVpQFRUKqrNKFR000dWzToK3FKOxNVe+Kv+pliaP3qGgYwd
W+5YHBtkZ25fuxf1dSBhp422yN4u/5AKRkEiPOa/dG2z/K3b9LFnqdixtkBfR4l6
oCr9jwBr6tuGUywEh8d0+HheS1IUJ3a0Sok86bDbKFTA84FQKdoFpb+pp9KtgmPS
WUWn6TNWtTm2NlXNO3hQmjunshdw56qFdUksR4TKLghrl5bBIBqG3Z0g4x34XQci
YLbYCU25g3URjSbKdD5oM8Dt7Wb7GKzvQiSKZ18WhEFHLH0bdhPCUeXIE7M4+Vof
0KFx3LxXWgfgx+41QFZfX3Nazj6PzIJvZv8bcVLyH826bID0lFx52Eee/CTDyTeD
LRkKNDLGt0C3z6zA7qhg/kU9gMU7HB9T3Zh1Ilalwz9dLRnFusyO8NLcfDpAnlfl
2E64kozVk7qSdBRBwvXuhTeS4niLAdshO36+b5PqvyxYA+BD8yrb4Qf9PKgLuVtF
TtVnwc0pXegHPy3Pp1insENqqccvdE550mZZGDK1D1LiqAqIvcWtIz4px1xlgthN
H9KS0ym8td9FOMZtRxjAA85+R8lBe2qCugnDiUfkfT96Artoh8IH4tQXqfYc93dw
2tTFf70TD73IHRHqo8p7MK4PI2RRQFmT58f+tbgYXS8H8Q24GdA4e9GkwY29vjW5
oSbTbhTGuFJKNmn00TMa2+kMtNfH7nt7bklhtDGSbuo+fPV/je1kWvYmUvur9/Wj
zrLHVckIE2hzUb4jZS9m1gJxQWx5FliuPPiIq6m98m5xQmxsoTiI9aFPmPxu0FeM
oYx5S32FQoSi9nptbTCoYVp09SHPD+IyY5QWOYVBDKdM0pRSh/8j3rxvTSLI+7+S
Xcq9pjf4uIoScsasky85/Dx3UA45Mu7E9YAOsuIEkmJ+EMFamDu8/cEZaY5DCb8C
dGu7ZkPowTcUEEaC3Df+fGSvU5l5BM7HytD6Keu+MEmzYEc9FJPatH6oCZga01II
dOWxQ2b7gbBxn0umMIT/NDYxI4AD4azmzy0clG5U2oBmG1bfMOhUbnYgQupj0QU7
dhuT7K5hPI6F9BhbYxo1yEHviAN2D6yUJT6efpZpx+7r1avyReVozSSYrEgykpSu
LbjbZVaVgjihC/LpGTTr6OnW/xOVe6V04VDn54XwJzLRJfq+NgroJfg8S0u443Va
9D6qFTERefd2k64eiPpZR9mD9HOvemBK195CRlaJaA7CasAG8v3nn8BR9WaXAx2Y
IuPbAbxfjATbC+I6Qe3wUNhsjcCi9QaVi5Qo2lmLNNWqCrMpcDQQt9ywjzBeJqzx
6BTNPl37bXLCjjC7GTVrw+/vT2rKaq605Cm4UujRLNut0Gt6u/fXT3B95UBL2nnt
JnNDrrNeaoLvPO+7Ns9CAifS0jNN/Fben4mycG3wsqKmlAkW33QJt1o4/gZ1ZL72
L5AXI8wZTqsU3/gadLV1F/Cl174ujKvRXejWzqP0b4Pf58lLJlTqHk4QM54IUoK5
P3YXWP2LGLw51Qa3kbQm2+4F4281dmChBk0pzhXfvI62Vp3NflCU5YMIq3/Alinj
DhBHyl6BF5T8AoTURYr6NYiXlxy7c+aZYKQ7iL83OY1yFSg2HvL74dLpiSbjhNxW
xO6tIlk4Ckbm1iRz3r5as+IxU0hzXH0/D034mLP2cMO2Om/4bdKEF8xtosGE8Qzy
gzEZPs6af+gsujSN3WhTXj8NaBi5Z6FBcyfCkszNMeTOaptTYWNQMzlm9ety58Tv
CB8+ueQ30B4Z5KELebLQ103VNy3EnuEUf2du/cE3mZ8+uKGqTX5DCDc9CdJgJ9tq
QyWMybsTVYM1kMq7EAZ7vZUPuPscpT17rK+mDlOOQk/nc0Rxoodsiyh/XwMVdTkc
HSchvLJgXq70b/vCee7ODyhTzVFovm7h24rnxGvBlOlkgNk7B42d6E5LpDhjktgW
b/bqy9NgbRmUJ6qKAZSLjf0V5iX/meWUC5970Lenb9Uq8gdcFG/L3cPRHcptYg9X
IkQZJalUzz3PFvExEVqhw1l+nCvk3GQzTATYjdaRKkLLN8ECbhcjEeAZziR6aXrm
LtGmqufSmvgTDvcoT5u29Rsv2mNk/TnarrJ3YHO1Ut7OjbCzZ+qEZ7R3MWYTVIJc
f5iRHTxSU814J3Lp8tmmDVLGeOS5ta7SHopRb8r+7QwoKlTB2ZHQtbUb+L1zYoxw
sJ4IhJVD9I/ww9iDZiyuzmOFbg1jO4R9xgbxgDnxCXA1JJpWwy+1WONCP2wiMlen
xvYPulfQkggWCR9AQ1DDZ2mzy5K2CjJGc81D2yWX+SW7OjRONSyrcb67o3lQBUKQ
EPGG6umq1A8NalNM8PGbvBNWEMpS+9PgNnSSukoAWsU45qP2Yy7zEJG6mrA9SaZ7
ZLN+h+GHpe6SCx0VPTTlsErkShmZnrKTlVGV/fABN59j9RTfwKGrI79cIfGudbU5
siiy92pdxu6hNadN7takI5u62NNdGyyv+Hq+U8IBnBhulQvtv8SrXhI/930KVU/p
nvrPnnN/8YXVzz/oLVwj6Eeri8TPX4Avry6C5CqtQmU2rg22F+F3ywbH3U1EdYqg
dW+En4vf4L+xj5h3nJvs5+1i1dllhIihTBdQoJGGkQ8kaiduhmyGnHFkm9ZjT5iu
Eisl1Hba2AQfIV+lD3+qZ0VLHRAHQpMBbF6KSdb+caqXpHsV8eVtl5UOR++cJvMh
stD865IWIkCLxlodBVRQ2RCzVdI9QlxEH5gm1KRBNlq8HD22JbnTsUkL1MfUCitQ
2AbbDIx/lQ7uOGJSvEXkI1UiB8pCWkJI3ouw42c8NdLNBALSWW5wPMLkivlupCXe
jZYSpz5bw7VLQ9XbRmf8j6FOBnauCtLKr16LcKielugLpRsE7qHkxMDPaq161ooR
t5zm06qhBNlyFUrrYQrpOe96pVs0CFwHBW3hf6Jbx/vWO/hoYvE31Cqg8Ocr1Z+8
P9NVvccmZPGaQVpLCIX8VnH8/gdjsRI7vgYD4C3s9eT7NRQ8H6axSv5Pgg6OJpq0
LlJ/I/YJPnqU+5hh90QPzYSvsCYSIuJ9rmXwp3u9rDtipq3ovFfsBARi4tIqN+QI
3H060WaUMpDU0fn6Cv6ccHx6nCjE4508PLH7itAofumBoP3089bqX3kLJRG7zuNO
TIILsEIwtQ4vrbBSX7ohKeIwNTzivqr/JXvAEYggcOaMY3zLiWY44Y6WdiENyM+p
SVIgWHMha2HqFdvMXZz/MKjFMOzeyACHcXahAEJhFXfCf1J3L8pNIB9HLqx+EolO
hP7witdJTjGnZ14Ihsbs7YycjaA71XDmtRYxiUeZQ2D8ahhcrAxyVCYnOBFKmmyy
BeojROTY5+bkBAtNL8k13P8K3skD5gTfPsZp3PMRwht++ar3sRHX1PPRlgt/OCUr
ds/3tx75Mbxoqqn+yppVmmwbCK48+hKg/BVks8IPCMabUfbyUyi0beECwkOPhcE+
4+7tJuHTpu5sCuF23XukWuXX4DyN9N4XTqRvmKJjAFFFimRmI/Q54HdUvHzBD+W9
bvdzmbpZxwbHuTfbd+T0aKn2TXjgvJJ4J4KF1Q7sMaIq7HlFYQerZ2VBe8oFDXaw
69xZ/X6WjP4zADtoYkVPrYcIgK2eM7ISnMV8SZwk6En2xv5CyklEq/mRbibKsTQI
oYG9ZgWm/G5IX5s+iB2XyDQsapTTZ4uS+fgrW390e7l+XV1PWKYbAtbWr5iqReTt
znKqRn5FouAZZ6rJ4IaKbMJKwWN3DAioxcT19kfBNAGtuBy0LaPvwaqcwcuDDt2K
slUmlliosSp+Kp7OyZejwaqxX9OGv+/TriPa8Qz4GJyqd1H4XMVmi+2KcsKScM1k
lyfPeonzYfCs+cEITt6rZRxh2lVXx4rj2Xn7L5/+phdfD009jHD3dBkxcRfeqsth
hAj84K4bo2qfVv9qiG7Vk/pBvMJmLDHZpK5bLHxrwJDeZLrv5CtfuUrHh8XMLrGN
c4bYMdFC+mwvVbmgGH8Co3et87cW7v0myiik1S2bh4oMfJRXSruU/Th4BF546xy4
TcZDvC16kIg4BFszy4rE7HJatqzsb0wVGVInR/81mNWpcK8eDbhFrFRiLzoHC4tf
DKAvHjj1gJ9wR3c6259bnATWnkn4xmplEj8y7WZ/UTxJxwDG8/xoEM75TQy6XHFt
JL5MMZuinrnCQfL5W59zxJktDgzs9rzcAwr/5NraOmL1Jqz9GPfZfGD4WDsczATM
/j3kDNzBvItZJ4VAsjq2VI4x0WBNckudt85oI3Id9XHuff20vJ09R3YOE/ukFr3j
cAPuxriGSTeamoGRDW+HKndfLSwu1wEUdPb/nfdM34LtUC2OAJw9MI/CQw1D5dv5
LT5ITEvRTdJpilxxwnF1kW1ZQRJGeAuE78f+Vm7Y5ndRSgOzPEneAxrMyMVhc1Uv
YVXqzNd6JhzOwfmzui0iUXuQnmwPJocTgTCLjONYLgJoSLSM+W35j0YuDzcqC1LS
RUQcnFv/d0rpwQAicctcClMwjAVlUoUpFGthXwKwGevX0ZowB0AGiHaXF/18+ZHS
hUSF/TOfohpgnwp1wAnSuqXOtBlNZeudKqouQM6L++r3lp7DKjifhrEX/NkTa6LA
Ka9g9dLaYkKu+TkfCWEutinXVOcG/Rx+/c4b91c6BLXXmY+Z8UFGR9Mardki6IRT
oXU0zaw7BDIbIJOpguIJL1+aDfVc9mlGIY0DwZ0p90/WQeP545O89gA+9Iz3HumY
EqMl4qiZsxN73phIpRP0VmND9FN/vPeIWhddToln9wk1Qb3PixBPOceBisLSpkUC
wbwmpBIrfv3N93GgQ9od5QVRefxmkxebXyRy6frN/m5CdC5qloImAyx03kvRbwWo
vptAWvyBaMEcsV0e66ybG+xUnwCU8zX9nd36KASeJX6bt+nvDMykIm4p4RSwzZk0
nlOjjah8vm5DNhSJtBjoioSReUOolMhaCmGHCtGA/9Z3RkYk8X4GWgxC8yZwpbMZ
h6zsfJwEwmoDXS3se3md8QtBKDEIZoaI6tjGqszgl54yPxb25sKZpHeP6zCnNS5g
R+agLx/YXyVBObhjUfFlI4wxlqy6KikC7h767RjwnajzkBvRTeGSKI4IrNYnXFdJ
z4skTAvGsWNVwRrU2DKg8ek2iIPV13wTZj2xzl4qtj2RE6BAIOK9tPi/GF7gqBk4
GJvZL88a/5tlmY4KLJWIYIlfZEXrYcovJGb5G0LQJf9ekVp082Tlq3BXJYWAShxz
AU+7si26Zdjo577ecjl50TCmO7KJRg2kIgQHN7SJKHr0pIP4Tqo+Nw8CFCzpomtD
BtytxsGLorWZrKq9cp+dMN9w8GOuGU7QvNhKZNvvknREbZmxiODxV7SmMIcWr8j5
6z7Jj/7FJGuH6aUcHtWzNDqgeUjiL5HvBQkHvWKUIlL4uCDKMQkrZKYd3Nj0N6Ib
BC6NvdbIY+lnG+x1wjn2tUjET/9vaO+N9p+QeVQQQYUSSyVsc5w7LOUDmS36HMkV
CQybDDMQqH9gYb+9rQG5fsX7G4vZuYoOQV+vNlKcZQJlnolySCsvg7NcJfGV3m/c
B8m8Rsydi21jV/FE9ilsBRkhC2e/FVxoBvknomBylfmJFh4oEvr5fymjxDWDCmOj
gZk9H6Eab47SImyx45ghFsEroPKiLkDkZi7wiI5sjDH/CKY0aCJt1wbz9gZfQ2Hb
8Vq/DnTMMqQJ8TXxv7Vue+LnKIE7cRzhGykO8WthTltyyx9utw4aFviU3ugD8/vz
SFP/CIfSAh0Z9AXm+uTmwUNv+DciiVFvXrGPrc8Z0JeqL7aB9bj+SyCbVZS0dowq
WSY+epTp9EY4+SSJRTlzTzx+BzCO6Gn3Ep6QnGK93gS+k0T973ElmegxBL15/Amw
emthRTgOrItMvsplR1ZjLB3HghCI1n76bk1P5S+EG4pEix3Ug1vyqeqgE6G9Vrw/
+LassdJujVvZaXuMhtoGye1tgEoZ+CjW8CMmL/6iugVACi4AQwgSwG3FYfqQKF3a
xvda5H2DnXJ737pHY67mgpumnuXxqIaYvfh16BhqLF08ZH+amwPBooGa5Qe68fIp
lulDD0zHtr9+AnBDv9gM+xwwXMq0JJAgFMk77F27VIULElhsXyXRYJwOX9D9GGpf
KTnBKkoOrJxznrXIa0O29Yxj3J437IUQnZauSl2aRF4Y30GjGb4Zw5V/o8wNNue5
NrKRuIUJ6FllSxrQVN4cik+X9UiyZ7GjD8ZraggclcvRPu0M0sSCP+IVJ9ElKkDq
bYsDQnlXrz2bCBnJ57KZQwioobQuNuHMwOkxrotRo0Np2V1PGAFTRtcdkHrv8VRt
Ag15apQQ8pwVTlTbCzsUqX82i73J5ivg9mB8uztN1Ch4hoQ9gadN8xRwSPxLpFrv
2AXV9nOSDR0bf5j5tgAn/DBZv49KdkOEo4Qi6+lnENQUB7kPeDLWCn7bbJPRVYG9
7QUUbW3AgtahbNgwCQBXWnTHTxGblYPIdznW6sVLkFeFRriMTg0EzBp26lZ+qiYT
CYXKfGbdOpoZ6jg1GaE+HdIGn+Cmoc96JUjh4YGAPHwsCE/WYUE9Y9S9HJ3sTcUQ
yqDGlK+uYLGDYBKI3znmX0d/8522Fwui/fHEt7NvYRPov2Y7pO4OprftvZiA0eVK
ZgSeY92QIX/7FeAE45y4Yscmc2BdpfzojtIs39ZNV1/3Vxv639NtBloWlImJOlly
l/x9gV/uFQ6mpVSWjWSR4aiifR+nq6VgQn4Y1rtBD11nYEseEOYwgy3eP6YCT9iC
z7MzM1w3MXl/uJva0Q937RLiKfLHfMfbg+KIpWbVkChJIQQQVS/WBOMi1/5QvrJi
dZxB7E4CFuz85vTh/HGLIYZw0QbVajSsrs5L8Fk/c8Q5bSPLA4J4kV0ePAoSjfoB
YrqW2ut0CfL202Je7HjnwohzQNMvmIa6NBlewCNmrOEwn0Sh6FdN4RO2A+FTfHnc
KaGisPHJRRVr6ZvwesWqbPVAlc088GBiI4+9x2AdmzVluboMwkjZ1gAPU8k5tbzT
pZcriaY7sMpGziHKD6JnCRtzAVdORnHXOvmOgbvBMjCVaG0lDNBsCsdBQPLde3L/
DAs9cvnY1b8Dc4JpZ6kgjD5evSeIKyY4nqte2tyUOqCMSxuh3jkRUiJuaFtLA16J
x6O9BIAXadR3MqRe4DsLqVcotjGAiaQ/pkGpslDcqf3KAhBbUtVQOsth0BoqrjHm
xBDbiQdOkC6TjCxnVTNzqEKqBNAVtrk3m32rlTrDNLT0dO475ptNk6W4C6Ta0y1H
VbmPHBwjtCkYoEfDK4wzy04gia0F+pwQXP+oXUldIy6gAOBITAxmo9CmOZ/HLsRa
iaLb5AGDYs9vAnknxjaCB1IFJuwvMDG2E1jUmubGstnNwl/u0B6NK3C5fuYnp3Fw
JhapMWUi+6KCruMeHCtYjskaxaDc0rxjEfvui9maS3OkHUfwa60itrOBKOOr6LKJ
67br/EhrC1HBrGn5/uBbtnDSyzg0CvggYCJFl9FTWV8zvtIauu0l6oPMGuwaZ2yx
XuF1L0LxFuLF4ass/ISgLnRwuo8TPiOf0SaanYimajSKx+/tU/xVIJpQHFj02OaU
LRhNJyvv8FHCI3SthNaZ0zsK39FF8vjnh0zorHZEQJRCaEs/3Pa7z9P4nYm0d7Az
kxsR/7cM6R9y29Y+8yiSIF3kJ29upHbqkaZtbr3fWvkK+TWVIGSMN70n9RIV/JP/
CgiZLmoGUR59JNxw3Oqy7wEkgzKivLXV93GS0nm7ccye3jLttS3xspcD8UZ46qVR
EZdRkqK/biu685bj3RyT/O6E2JnDR97CU+y2SFqmExS96Pu3Q1mUOLoWNUhwc/AG
PfbLsXTFp8rhyWEWy2WAied+CZp8WaKFBBf6yuJgb23/bBqWsRcV4qv7PT7UjQO9
4bFJQfKfpyVEoT/vjta/f6jvuDEYwjhsFASU0Lh6zfjUM88LxkUDKvF9VagfXM+C
fmHcLD1BPUY6V+Q4aPc8TSceLVHIZLykC8/lUxDTTL/Tvaw3HMxxRy7lWVybkPjA
GoGp0e/WFF6+9manoBq97SELeTBVDG5KcubhtWGlr1k3uO7BKlawJVnQ3WK/r3IJ
a1r8fXXKJ5T8n9FFO47vHEovcmSsY2Mg/Yn//USjRQSRCTXDHA3229+9FJP+nKrB
wvI2bnSKl8EE8aQwccuXxIRp+PC9fO80alQB8WmyaFOcAyrMIh6xQTY0ec5ZKL5z
a1+Jjilr1ViZm8V2RP24DP/8NaysvZra29lT5RSI555wZzqKDvMipb2+sio/t8vZ
cEcUik+v5WGvICuNjdRdPDfspZEODfNEO2aXgEHcZRdeINAZEhCCbaHaLyIIFtVq
nk0WZQGJ4TbT5PRcgwskfVgSKYqIt9Axv8PNC3RetGDBbyglvekS9wcI1NtD4Y6s
xSHLNCBplFsX7P5gOrrIChbrPCpqpraRNWojR3xwoood/5XXMMNinA0NFyLWLqiv
hEp6A2IJ+GM2bcyZSiRa0qu1cuCCUdNqUKxwnQRKF78yVgr1UCJykDGse0SpaRZD
Uv3NZFXr77uePIPAy3Y+wX8HHSymxdqoGn7U7LGo3v4yrvCFZVU+mHTfgZ1nJzRl
zFQceh0/LJtYtL+kIob3UzdQdIw+gsD6l6AJZ3MQq2rOIZzhoaKOk5pSC2luPonH
3VeTT2MaV305GqNG1LtTlUQWO5EpxQrGxCDFZfYal7oQVAygSWBkupMWw6VIvI2N
3QEHl3vY6BHoJt+8Sb2bcUCXNhDtNjZpA9NKX4QbM18Y0RUjHZolT3xZB6duRpcK
/bSKhwsmA4rqm1kkQXqxUw46POyZwG/GaV/BYqxx0wRETnb9uK+vtxrM53cFhavk
JkqyNDAG555+NM/a7Vad/EA/5G/+9jWF2WXEPgEKo/EsKrblV7GWCVSV60R/0Wuk
hpAru8bzzjpW+ARENT5ylhX///yAAmIQBIBuZpv9RdM9JwGW2bF22yJbIvZjwuRf
nqZY6lNTPYGrlKUmLo92UIW3F0Jgzew5rNRdfYEWK07L51m6X3VjUGpwVh4i1+rY
W+Va+cuEtlL5x4/Elt+Uo7B4Uud0GCW9A9MWnHUwYuaj8gIXRcnH+lZShMBvGCBN
Ske+f0qsJuCfLIOQN7Z7XgTn85tF66aoXFXp3pmLuqXEdvI6y1u1IiV+waDM3aL9
fYse4eqxGDIULlsp8lISqmlWwr8zyy/t7P6tOZF/v/ae0t3+j3qSpjHhvhOR617c
IlCUgjmpHJy3jxy7zfRw5GVzZXOCXOISCPxcyIlyG8GV5n0h34iSIYeOCopcMkFj
E6muR9/MwY8g1P0RSUK44O7/B56UcsZddSvc0YhHgwBLV1ANpPfFI+1M7gkrO6Z2
5dSTsdaLn+mVqu4iz8EHuoiQnDNi/9VQ8KoKwoDjzxWNgLW0Oa6SSbJJlX9r0TJy
vGqvRjTy0f2fIqnDDD8MzHK8yLJto6HZzixBnBhekAAD+uO4zPxWzeghmZ7Pqtk/
2Ao3qfhqt/eQLXehlY43gDfO2BvpmMGWmQf5UxPeQYfgiNHZeQDCx1vxbg6X9Grg
VTThMOOtW6KdpVgynDZ3En1zuJbcIbLjJu8+bpl1/RWxUUARHDVD1UFPZ5hZYy5S
CUg4ariNHSd97B5LsCizCtoNkCIUk5MpnEgbQ80sSBhCOFyrHjMuuONqVrDPUp4s
SLem9H4cCHkTtG6YSlV5Oix/LZ3dGgpcm905BQKswS6WA/wtCds7HuhunXL4IrTW
AhgQt4QQ4tyTbgyfSRfrEBt/uLWoqbgzPR6DgrP+tK6DPZnXiHJnoT0QEajxPvpM
60/offjvdZlNwzS/VhvLtV6uDN16zYFRln7BCR/OWu4iDKTsB2XEjC+UnT6xgReE
sjPqBoq7Yty9cig0nKyDr2/gK9jT2W04kndMjIHhW1u2KpOBHnTUyBeM6KrKiuOs
ZM2ERXGbmqqoAvbmgUvvhUmZYf9eb5kTdgPsofBf/txmeOlB64rhkrptZI9rGFqq
zMTmJx1ewcEEmAeV7FdVDbrfpcCDMySJADTLAFjr0aitMSGqa5sRjZnaSbbeWtwU
ZrrIsZUizoQ4PnzBJB3Rx8hCeB2Wwk2nor0qy9zlecY5dRSAmQy3p3YWXxBW2N9g
nq5/tadY67S+N7DnDjEaBu2e0k6vYSsL/HCfL0KUWBNoP+0k3eMRrRl1OAchVOev
Ytue6/vab1V+z5FiTIhTmY5t0BJb4UD91YsPhPvCmz0FOtxc+o2KIBPogXx/65mB
xwiy7mkAp8VVwPk+vva5/3xvuAp/VEZ9kaJTgZ1FDHwqhA/UC1JK9sFsWs9E+88s
jOasg8UeSFzeD8yipXdjq1TjtZTAsmN0Y6QsAGKuZ52GfHJB0frZuEGNaG6wOVWr
1A8bJ21eOFbGefth2CndSSiqDVFarFpRqivDVm8RXBB63wdj6FSdi8oOA78EL3fJ
PeS9Q4R12VLEQy3/iyW4jxLa3AMi7mJDHHBk6yCpPLecfc/URCAmSWCm8vGabucP
EFAjObb5oYZ8YPVTqsfEQ/Odi4Yc0ey6CG5YBsj4AOburZ6T10Rfkfu8K0rdNPGe
yqbRqVAoHCTlV1/mgQnnUzKx6M96lCzxvr9kKlESYXIiTeZjzcYvGHRYPk7PzmKm
3tdbXR8qvW150F85afb4O/h1aIIVBdphOdfyDnk+1YfDYdpBiuPl0K0BneAdPXIO
8stv98ziy5LQRGWxZFZAh7WQRvPaMEedAcPw/YH5Dk/gGJZ1GNq6ILAJmHTwcJWF
07Ybv+RN5lefV7uWeI/sBkGMpvXaDhiCsj8boUVfEGsEb0lSYZK0jYWYgFbH349J
NykbGlm7wDbWkxiNoECOdmEl1/tnpXzfdikOA+fo+xqASgGFo+R//FP7tw0DDd/z
yHRQ1y8oKtwn1vyB3md8Pe3PBZw4ZxBQXMoQ3x8JJU5JRsi7wcOpCVlQV2VB5hVf
dFjkw2LM5U9s1CNLV+bk9wFkFn/3PNEtJ56+8x5c1HHNjM0o5AXztKB/lVEuZaF+
Y5NCnnKFwzsmncLI4Xu8iIDEHIP/grgshMOSmBsAZT8089BcMuWv0WrkmZXzrdRp
lclBnK0/f1woOCJ9mtffM4VMvbZbfnn52YN+wKdnL1UyXhiYCimIif5TQGZlBzHg
tXF6p7xh9e9me88c4htPk1xbwibt1/f766gk9bwgK+zmmFfsnBij0RK84F5GHVOG
sx6QimYcdq1uoy8TZDVkaB/0+l9/QO9aS+ZqDOwzTRD2esBnQZlz7DToOwXV9dC2
1prWXBrpM5m+9qEU+J28HEYhn9bcB5p4OIxZzZSQFXHpm2PiaOAOd3ohzAcwR3pI
kIOwfNhDWyl70nAsk1szc/cx9Ivv1qAMlUjw/lErLciJIL3DFFTxQBTy80+951y3
4BaH9TgRbC/gwwkf/kEWf3rwK2QoDupClQiUK6ERgM3Sqdnjx+peQU9WLgbAwB0C
At6LcZWT/qQRFi/E6oc6CjxqyIza3HzQghNNF2ouK/Yyny5kIVLq86Y6UaaK8WXd
UmQFvZO1xybbxAjeKICIYFZggHRTGHNHGaEX0TRxcN5AZkTQxpEnPC921to7OEUg
kWiW+Z1LYqbD0yaIsb3pRRhYf/nFWbIRO6XclZ2FjV+PsehNlH60Qgb+qXWgyI9R
ma6I3t618UeyEComjMO/6m323rjBvygJVopfuFj/U31ME8sUq60QgCiR8Y0wo8gr
JkyvUTXI45dTeApt7fpFq07AAF0zcVskUdzIy86rJfk3cXV9mk9zwUK+BvTxWsPJ
eLRaOc4vI/KQPXZdDe+Tc3k2QvBY9oL1fZFG5aJ5qYwr0HHhY71eaCQwyp488HeJ
V0FEHjnMh95qSUVTVSpkl8A2cF2LhvlBaps3grH7FLn2Ujq0mdhy6obt7Znhwm3P
8c0Iqt//ylfbg0BrTBrBUH4wNEIMNYQfbME4Nt5dg1wirMEuTti4o/8dHiksRcQc
KY/nSs+pcECBmEzkmm/vG3mu8Zownbl/7Asc0HbZpEHZ5/PO8l0HSKnKN2eTwM79
N033gW+FzuzL2gy6jpEWr77RMhI1CUuaAmaxS97Ia+YEwDw1VMGe3yW3lNmNtblk
g6p2pUXVxNqi+O8ya1rIRyHDqN5kJzh1sofGHPEwOpK2Z41SxA1z9mQj3TYGeu7U
W2/BTseKZoPTPIAUgFwaLf8x/ZNfaMJUe5nKCW4mbjBJ0n1IqdVL14CrWX7EGziF
X72WIZ84GCpNtfbYRvRhzhmuisCT0WpGt9Eu7C9An5Z4mcvHjMYyJdrZ0Dr/XmSV
9WntznY2o1x6lAYfGKfK7BJZ4fjTp0cNpqsf4eexDXGxc41C69Rpms1QCdccDDfN
WVVb9vku1l8c0PYPnpHfG5Zcb4boyDlyYJ6s9bBzAoLzLV38/cga6lXBsXdQhPRQ
l6bG05gG7CUjC3C1pzpi4ek8q1D54gkrsG2BMTSmE/fW0CjI+8y96PbrubGDVTRa
vNh7PyyJdtIiIyZjpxuQwVHOQ17sC4xKnx+YLqvcTn2nwm92jbmXbtinPStPDNZJ
lrLRqmC6s/1ioNnArbxC4CbguaH1OfF3y+T+uqAJ7W6GhPiOAaBwzjDupU7oEO11
c37m8RNip+v0xWr4YyH/pXGWbs8kzairQYUgRc9KLTzGPz8CcUrMpOWXIvFTtEMW
BT0WBFmgHNOERU5/CzrkWFvwy0NqsEtuWsdAD+ylU7tRTPy+uK0di/CIvGfEhMTH
SCwWfyK+BX47NWnMZpGYwlB6pMj5n+fIm6wW1z+vXKk0zpk8o6RTCBeENmqPbgw+
IHFmmFn0EhBsco9ihWsVFj4Kyc5QTr+MzUrNx7K9yeo+ZD8oMTDqDVcgu1k4m3UL
JpoGjXFLn3bxXC6V869ANEifYy8j61tJgr9txkHPa4U5Z21e6RxMGnx05GEzd0Yn
SUSjFwiY2z8OVqf37eVMqyIrDknPTRYUBLMXYrqcJH4wX7XUI9/tfDaAjV8vMb2x
DyvbYUPKGp3myc3dWsDoIvg6YTHewx+Mww4Uc8nX1yiMDt8P2sB8aOnHyVkFmsIj
4tXLQwmw+tq30vh6dbBLojarPcfBGMvAUOZ0vZdLCYk8HI5nwDMx1lYIZP7oWG92
Y9ij9Y3DOCG9gVju78IdmUu9VYlkBJUIBfe7TK/u6bYqG34arxn2rM9uF/ebznrJ
x+Z1GkwiixUUL6L+fopJeWfv2RNMbOILJ0+cAqK1h4HDtncaudV4O3aPE8e4p4GP
1xajDAnexH7KOBwBBA56Dka4cTRbKiGHiElaM+f1zM1ZbSAt+BxjqGfhpIzAlyek
mz8UEjCTZyfxuAzoVEfyTXLTt0cdX68NDykM1roEexJR1jYw16P+S2+wFME5MeUS
ENHaAoYsRJo1LYim96niUuHEiUbWe0hlyA/0GPKg8Ap5a+flFiAPDUVLaO6iXg/P
8ruerc6dnxM5l5wY+eZhweZ6nbS0jpn5ODpOmz1WBpl4kCs7iCntkuoRqq9mTk5v
HW6txXev7OeoXkDxqg1kSJ+faCqIQHzxi82SjKvWoq+bQoZH42HxZlk/nG+vRuaS
FF3P1bOs94G9AqJ4XJrg7/YQx0+wKZYk+QLgEwx1MJO/h5FUM1maBKkAD5n+d2Nr
l/Lu1pB1LJ3kJHQkCJnYKObBLg/kMadzc0wKye1lxujnOt6+fVVbA6cmhoEaESEC
WhFgAvisrnBbllKjCe2zlDIkVzgJVIXS9plfRxy5SjKRK4ohp4xv7KsEDDdhikrj
vTnajHiM5gmqKkaZfbAf9/jEWVcethDV2Kfje15KtJalpeoMJHNQKY5mkDrSlTbC
kNfEtzbViixFp18Zp80hmdLLGkKY0SW7Mw05q80iRB6UuDyFc06u3Op2CDHwn9Dy
QkID1qRHX02s8+ubQi4mNrdj8QP5THuB7N7l4ax09GDZuDvTXu+aEUDbtKMExcSa
m9/Gf8hpNKak+uJsbXY5map2KbqxplzRrJnlb4DdbmBxOXXtodx0Kt6mRtKXyI6c
zijnxC5iwcVXwXJquCLMEhnGhG80JnLxSmdP3eP8QN05qdIXQT4sLSVT0TJ+HxFF
i+yuVIrQO3HCtz1MxW/ozKja/bIAKKiD75uLQinUTKSoBlVLNKsRRY1+kwTvMijQ
hLk1EdjkUPciPmnC2xMSjwLPAwgQoSiRtz2Ha0AbXp0ZW3NBty2LfK/XFjKfFIiE
rxUjG5v/SQe2q2guEgXiGz3RQXCU3DIEdkf17JQ6wLgdvsISxc5lXvVSHfmyOpUz
tKhLlEpaKvKzBJhK+IQPcwiGOODBlf6QOTkvXOlieV2zj6YiQSe0dkLVs9xA5VmT
Rm88y8yeNHWpPU1sA1M6+vxmOuMtPqdP3KisornJSmtFzSEzmRloHN0rYnhNlymq
NGSHy1tX9hHD6x+0CJd500A1vRLFbMJAehh9VbZq41JscMtuGuQHf5fHpviJ/h0N
j9hQl1w1HiR0x5iUA+sTs7+VSnFCMVFgDLDQp5cyDT98D4D9Ota87HsxhIcS9/Mf
usz+KppYpcx1anrMg24ym9wvwEbViTgeizUrEgliPyCUjQNq2kbxI4Jo4TPWrZhm
BMnITxFuj3hhcc/UBttp7NjmRpNtcEb7vmPb1wUV2boyS2Kh62yceeTIkO1OR/3L
uCVhUANFK3t4df0ud9QFyn8vvHYBWK712np5Sg+1IXlzxbzsZ+Q5U0qFVEswoRef
0yQBKQsqAywB+5sm44X4aRy+TV3goM3H9cJMHOjDpzWQnfJ/Xhg/fDnx57PbnGPW
jA6ZPcAtdWge/3nOPDbeOs5ndgUoIU8NtQybHN1q6SpYFpnEsWiGTjzzjM6xzVfJ
1bDkBKM+KyVtErGR4xyMwAtq3sbdGryfVJBO5c2IxGhzkhxlVckaFtP5GPGE6ZAV
FNk9FvwGkFVYx+FIHUG+Vwg1+7124lI7JNedpthbDzE2aFcjRdHWyANlNCfPoQzi
swVwMFedRIKiKrp0QP3L6JhDBIjPAUEyR/kGyIQuQL5UEYYmgIsGHYbzajoSTTt6
fol6Y6p5HuZc5+I0/bg9HW+M0xuhcJUFLzKkKFT2S9jcwK/tmJPT23tlC16+7enO
sdbIcaYPo/80xS1bg3uTzUDZ+hCWmBiStenilKKnEntD2+fb3/OE+T5lytP4cz9I
WoNmFAjQfikAk4+qoSrtNNkwcLrPkaB+9RmdmzHMymyJ1s2+qoWjzLLfmA1Ty+ie
BkexN/xDz0fs92IzbDg9nTdjjnIdzTgh4Tx6TFtgVBc80n5hXR+tHlmlsSp36QpZ
qA3dT9uScvxhb5rqnLq3LGQFdhTqGkaBv1q1iKR9cCNjfOwQEeoCtdooC9YD3ifG
A0hFTC3z5igG4Gcl8E5maj5G2LVrrbOfy5xbsaiA8C33dfZJGv3JwkyToprs576d
6IL7Ax51V4Ayt5PnA17OkjGopfJ8aL4SCE7fBUQs3K1qisNiLLf0AbdrP7jSPWS1
+mLzxqwW6yOpA63VoM7ne1mY21ANFuy7nqlWtaK9lYRqT8u24tJU58wgIjHDZakR
QQWDd6qATSFnbgL2LPfS8tgIoPFVdmJp1aMB7NyDtgwnEmqrZyOBeQ0QCDIU7vQU
7HiL7tGMC9BvNMZTMc2mCg164x7s3Mq8uYLtYsd2b3BeN6+BdrNrn926K4kHKM3W
zXi3QXX3HIQ/8k1IezL17lqjVdqqBsuJ8e1W8QuuYN+Sfrz3zt6CD4YFufpC4z+Z
G2dbIPdnGysjReNs+kbdJE6s4f4kz8hKhDgSqC8hAqVGw0l+CEpMogMhPmEoEqkC
hhH7Hy8WmBI5gIxMeRI/HqdA/dI0Wze86nrgs+dKY+41FChSGQQ8EIlvzx2USA4Y
ey+5+lqh+Fymf2n/JrYp9uGqlNGVK7rGvttL+laqqU8DKJLU3MB7xtCjJOc5Xiec
AJjsJfovD0xqwiQUnsY87d0nimPdCi+kELP4f985xkT3ZAqOEbcoYLU9Rs/+syHO
6UqtczWoiK11cgseJ8EVnNK2rTzgeGfj3+UXEnk2WBLzkyEktJriMqEHzfW2gjnj
Gt2KkH6YHTRB7GT7Di9HyCy87Ncd+JXcoA08lc1IAD8kjqGUydBwX+3ZPsgfz70z
Wp+7QiQq5n/oDIoH1nlRyZaS7Sxed1PkW2K2zZzUep9Uiksixe3/kobPdE+IbvR8
kO36BqhV+JMzUG0VnPyjNRSp/vDnWlRogTs5l1noatFy1xbK1dSNj8yo6+W5WT/c
rSpS7ycqnjGelUkMQwsz/GNePbWK6pMplFibx+ByFabdTr+K9xKexGgO2n5t6jxT
dTBkPalG8qhUTJvPA9+nGyxIQLbh7cOd3XgqU14ISPIsfSk8CwZI9x8pTZAMXDnn
Xo18vMNfD5sZr5aSOrJTXpFU0qFxhHnbYrm9H7trEQsfii/YvGMyKfYuwaJV/u7X
NHTe4DldsfpmyZG8z/jGSoEqJzC5p1xbRhvbIxvXYtAotMM5lLbtMfRyiSsuHL28
n+Gvx0Er8CoVq210DolGbqF9sr5zhaNWLJ6dXPggnTRowvDy22EgZVXf79S3/32/
rQMtxk4kF76P6aq/J8gquZN3Wg+rcJVtnyrvWVBCC7HfB1xeVeoalcBb//C4m8N4
NuJluAGye60IXLLLYnHlaP/178gxuKnqGRI16Ub5rY+VqCqp1dJiQahJhvCzcWP/
h+IjNYwsZcoYU825QCO1BrXJWWtRr4dqlEAwqoqC533ZrdYZpSZ8oo2pB5YxL4sd
DmZrNRGeUnjvqOZ1u8nhi9RixqY2uKJNmz/EiWgQl1B445+vFLP/0i/oY6XNRWke
vW0NNtwdlC0Lewb6TlA3sIg3q46MpJYWsnjH27Ry9kRRdqkbKeP22JzsI9JllHhB
sXEzaLVKZMYN9aJGj5mV6j7pt1sr1jNiJ2l/chJhrVNxz5EsoBgTBTEm9d761e4k
vk0OJ+CwfJa5sIz3qGSbhx0zEnUTRH4we+X5W/fkRCp0O4bPXICpMPO2V66PHn5q
vFJytJ9H2p58IY5/FxhTn0/6KPtURCwtVFsM+764SqPyZH/thxy4qC1g20obdXee
RaKFKyCfG3cwFqYeTi2m/3N4igwoLVzFzOj/e18XEjODeuGM0BbwtoyrszxGQaNA
Zr1IVYCXpFT8LNshWoqVio3H98B535OOp4P17HmT85UwBPKtuRtAM1hkxY9entwQ
asJ9hIrCG0NMWS+4CLa/EUUu489jL7AfPcEVKfLtXgdqGB4EayKI5W6eF6bQ+r09
AG6tIlxe+wy8nNJX+3uYZ1uCEEsQY2sJqxzTFWRUxO26LFs37djfNop5Bw3k086y
k8kjD4JMvLFQQKCcYw2d9znU1hknsSz+DWJz9zOTJn+IBWhPe4QC+8xVSAE/HmPB
C0UK4JzxitV8YYuht3fHLB2Y/piqqmhZKatIqbADh8fuhWoBap5i7ml1ZdcYBXBy
MNWePKiP7niDQZKM1+u2IvjfXXkPC++cYCswPBShWpzAva5v6JG0mSCTViiDC1Pi
WCV6C4GNyJ8+DoFXjzojsvRLq/QMLYXFOsBaQYfxRUMi2tpE7lGfoY0dksxvTprZ
ZwSoaNqnahVE5OYnd9aozTW8lIAmwghc8NGG0yyfRkwJs1m5cJeDPcWJYycL+0EE
1gpNQHfa4f7+6LBO9DCMmotnDBhwezWYRToHs+uiNRClM9R3FJilHLOsGunjFSsn
mtY5sZcJWZCrvsxn2cKQMEao4k6V24zGwChpchVTtJ/ANsHuJiyKg3l99J/84vYh
I9Riui0vYeW+GzaLs1zpbD8f/+HC4Pp9I6soDfR/ihvPPWBLTBAmO3+tCgvb3Amt
xLLArp9gOzXaqWEgwcGvUEwSPQe3r0jeuc14tKVKrH0JYamAjvgxUyqXHd/q7PBC
PEMdYEySLQ/UjUNjaRD0sRzSuLEsPNSMwaskYNOdn+QBD+/Do2IbcZTN033oKvDT
/NU+xuH3KeOlDzicvdYoQU9663ZkHp9GDYUgHP8Jolnp/6ncGbkw/OUtIYnq+/M1
fs9b/jbdzBW/tWp/FmAYSoTGwZDoTtQGf3Udmk8MEmIadVHbpGyS01FbjepOWtkh
Ck9RpuRn7rjjfrNnoJD9JNPWYMjxb5Le6jkkc05624KEuD6JkXWLgzvtkXAoKcly
CZ3WH6SG9i1kEs1ArK4ZRsQvEaQUigkQFvrwn6Sieoo+tbYjjl2r4KP7nHrbuVe1
6ZEuxMnZY6ME/N+/NkU9+Av5XmjGWmLAG6oragpS2UpvhoRaE2pM9kP5tCypWMxF
KRa0h/yPKZwymh8NMkxf2t/Z6g25gBtFGJfT+wV8YpEo30Dpb6aEmJKF5iNr9nYH
aQdz5Joj0By7FGJncmrc1la35G6eovNdYp2dMdGFnMnkhh7jPw6aLCcflHvdevBW
dCuH1HdRtWd9d6wMxjFQJP5vRh+vFnuxzzp6RcRMnjrM4cftoFcvuWVJxKEzk7NN
aJUrwFlOiag4RlWWLNko972hJwV61/18fPF/XZ6uh9mnL5H+WcKw7qG9O2ceUC8g
V7dnreLmWuj8zdr2XBPowzGE4wbRVkqdFzRO/8mJLiddPNTQaSCA+7nZVh+aRSvj
is+XeRb8sMq3+uxsuu0GrFPUqlhLsJ0o7fzEO0sBGJ6oTeH5XbajXsLfp51/HiZV
/CHPmAi1CMh7IQtT6SO6ZjXNIvLZ9mPG73cOolfMELAfURfRjnx6mn/hiL9eWOYI
Jv6j+hqtbm4MGOn1jqoI7MKlrzXMzNbTx8P/y4css6f5JJc6+8DzQjBjjmnACNvN
1Nuiz6QrYGQTsGCI5bL4Q0dagzPem6+UPdAUeTTYusloCno5Wup1MFIu9Oo3U/rk
CY2kfzlmjwrpjL64PAvukbjOmyBy2a3hhcP9g3dbCA9WiHiASJ4EGFshSkXKQtJ1
bm86i/HPGOZBG72OQxJHou83CooXN2y+fWu/XtVMgWwNYn9PoFqwyqwK7Hzby6mT
jfQE+jAJ7fzFy1lzd8Y7eCC7t4N/KT8nB0Ji7O0iWAMGydP2JAP/dzm17HAuhexb
Fpjc34LrUOE6QOfMIhu0/zJ9szdsUSoSwEykCOnTZlZAyY8er2QxMOp9xvUYrlgh
J2o4U7NS7E/2v0p5N/U/q99zx9RwWw5yOwvoOqrsu02HiDZjsBSYHcEDC4w3XoG5
pLLvZ26xV/x1iB/5hNQ+Bf/IPJOY9DeAc7CUZ9zRAljJxEppLzRQ0tE4s7oPWfCb
+VQfy2qNgL4DsYCfkYEGcXSHJ19kEQ0C90q3POnPZfMLQRkI2geZhkGYTl/QnBoH
auu/jb9/HZAYQcQOr1tfb1M5+YsZe/6BKAGXf2HC5aTWjRVEn92n+8+ro7hrurW4
CPsnq7pVgRCUV/KaBQGtel9DDzywVboKITm4tjzeX6kTjyEipFu4/+e81X88gyy2
o9CbgbEUMZTLewFkFMqK/ONeLNjr49vu1ST0U/qsJfCool67VYVBz72YQYQGdhBV
8riJ7Gqc4RGNEFuH2sFw5N2UUvyohquz26PlWG4ZSG5WeksQ5vUn7W0mtIGujDvp
/+Gd5xHsWPIS4NHxHJvmdO4bJQb9pjdc6EdfOMwG6HXwXJ+mIflzEwz0M8U6oNu+
C01+/VU9hNDawhL45G+TReSKgHMOfoaOjK52MP0xmtm0BKmTCQL4D8/S4q9KQVLz
a+rnQi7WHv5ceN7F7dNjkjZmoHYLRN1zx7yjZl45zefSc0N3+7YOs626e7cgx87B
bXel5GIXPeCfcMel2ODHXOjYfujQZQ6/0geG16qbi/xAidA3mIEoibe5RTwnbh9u
73oAF53QkVHi/G52MnEITwX/yFK7B3q9euOlUbuN5weHHln8LFPSWUNFR1uelrAL
FzYYnhE5uGEfPV9RxXpL+3NoUEG69yA7o5sAnZLPoIRRr9FBJxJig/WxFUbdelUh
JGMUUxh+sSNWm8sqx7a7eCtcdn0GkvcgCcgUawayD6v2m0irOtXvJEu/KkpwvY5B
eaugZSVIeAd6TzeUDvOsGCp1DHhi//JxM0Igs+F+0omv1ZfA4NskSnvD8gQwEsw5
Nhr1k1EbTlzefO6zFGfxVzFU2KBLRJBEwtq3ztfuCfX280TUfQnfd7UYljuv3KKg
x2OFND7UUxs+w9QiAbt6BIY6eDzO1hkZsL6CRkZ2huPXhA8y45Yyi2MuyDxeV8v1
SiWU/SxpaYWkspnwGtZpP/dGN8SJWPWK3yogKHNuNslaKOZB+ItpyIod3uZvt+vx
U3Gh0Q78z+1wbPl+YvFJ/S8KtJng1o4i4UnlKVPUmshg3BODa18IWwC7a40nzX8N
+qJK69iZtomH3gVmd97wsO42lJP6RLaincAUr4pxNOGmnLFzwkIWLtaLqeOvcUvV
ilqUoNWjN6UbFjmbtDfG/G/lLP2pPBRmh2VQXXzphd3awxfXgUwf0FeM073tRGoD
LCs7DStFM26a04rZeNHk/EGfQaQ/DQw4/NxEC75biZUyffSF4a1jogsBoD1NyWQ7
u2PbOWbDKTjaG6/FiWsHp8asL1ypu7H9roriEg05aYTfir1BPgW2+mQ/D/xdUL3o
hBIzoziSydRzZ2iiGwNyzNYbf+luKR/mfN1+jchpZI8/CdKh/czlzCIMJE2Idpql
slZdggElcyXgNuWJAHmMdox9MDJ66sVRb2x+YRYIPrpTqPBLhdDHr2fUa+ug1Oyj
WvQOkqsFCodFIV5PYyWh2pc9sFUmKKuT30b4MXTRBqrfUWlugJG+Np3KFjTTQLwI
LSZJcUOD7XomR2hQ9KmZYQErfanNTVbRwSmtwZzFG5mhoDOAvnidMAmaFwwBKMxY
PBz1xSU94XpxsWlup4S3rMT4r6K86Ly847yEgAQz3+y+GOUMB583y0W+riO2MG5U
oEXgMfaNpSnR03YfHgkjnAIWqRyiZbYx4HOuYd0xFlLL80AddU/TW6WIXflHycqN
nxuNzO+NF0IXQvjZLX8uj5NwS0Zf0uLrUqIqSN7azKPOs0pBBq9wC6zSiQW9JUVT
6AT7/P9JsvdEhxJ6Lttf8hSdjX2Younh9GtKjFZuCYeKoKo4t7REezAn6nMMwxKw
kVAtgH+mSyBPQlv8h6eUy/7zpUZhVxRGfwTTGbDk1nrSYF+Pf0LbsoApAYtywZfD
l1WjYQkkDwmS+T7oYfK7oys95KeSMSC5bvmAOytEKsGrrDSFXBfqSv3N5Xu5pKtA
8tr1hRu/82rYICgWo2TG5+ihQoFcKmBqNQDaijBUgBuLG2k+oc/bR/7tSd6N/iHe
x6Q/9T+iDbnukAn10lR7j0HrtbfIsJkOMiAKEGn1mjHkFrQOHWghB+nc2xKE9Jgx
XJR39heyXNhxMKzBl7uqc4JwD+2QLggAYrtkD63ahGfCWcz+uSD1PcHz6sVQOEN9
YMA6NRdbbKuhIJIDLm1r8WZq2K+MYrneBAIs1npMypxdlDlrklZxRJ78lNlW7k7T
jypgclUJa11Gpj+znI81mThJSlYUi2Z3mkEBhDjjcAERbHfoV88OziK9+4pr5ims
hoD5NS9RvQSbzUL3r4n4W1BB53lbbSVAT/MbcF/qMFt8mrciemBWAwWsUwBdafhe
vu2P5hlxsmb2lnlM7AzYXrzW8oub7q+N6mxkfZEXNzIlVTnxjiEfluFLxYMlmIPT
vaxlPJelFDsqnwoSvCtxBTnf2iCdVwlRxum3iov2i96zjz1YGX5Yv5emsbBhv4TV
AbClx+0UVxvBhbyyuz1fOLh2i5jo5Nd0f5b+wjcYnB7S8dePqddWNOwTos9Jb0Ve
dSdfdK7chJ678VboqvsurQjc46plpgIp3sDDTTNFTPa+bo03zvCuG1r49Y0QcIBa
SGiJj7l4fCN/eOqu3V623TyqQL67ueOREI94i8fWGhnPsgJmwhzv/tETpQN62jGf
etZPluMBZ5IAuGJUpUm+dbf04sBFoOc1Y2Ey6C/HaFSFZoGOEE6ZhdaQUlCdM5YO
tlrNQN8lS6uKVNsQqb2NRezBMNvqLsboWVijmCnNuf2kqUjNB40xDL49cuoFBVr6
Iw8Rx9BwbqnYV7IRlE2yaZYxtBYceOek5G29C6MT/vjoLjSUodL5JkqoIxLUpXlA
RUVUX22nJ7euyf51/H0fVbvXLYzOqq+7t6C4UH/FWO2A4Rz/ylAfrt1+7HVEcWnQ
9FVxsVTQjHpfJTcoDgXxOkZXXtd1qk3A4Hc12N1co4A8ST7VuRHP0nw3mBnrEJtX
Y+IQNTx+Oy+yWBdTxU/7GsXy65+/Kp9eJN5Ij1ctM1yfvUhZQyu+AmaZzzVV3AZb
0enLAxhkBS5CKqUnofbeUfBLmzz+KbWlcluSewaZYX2MW4GcsEL1wjiYq08/5yxl
j+SMOVjNGmdJqHnJJ0ECKEfvzTtD52LEIIoyR3cAlTamVDX8ayza1U5Rb3uhxUKK
yEPKGoA5v2E4VpO+aiRKL3lEJGA+O8FJac4N0DqKIqEW3E7jfGDh4G4ztRkTAoir
SVURB9r5YxTc6d3OpeBhp5NdtbSvpj+dDO6AtifepeuLqnLraIX1kM10YkwPDl3K
Daexv5iwQCN37hv0CF9J1qqqfBCs0rY9Zzlet3LMnPgdYzIjH4tD84UZIs5IinIF
6hRhR2QCVj+IcDaW6h/E4D385TEzpBDEaSRV7RBlR4BzIWk2nAVrewYk6P24tP1O
p4gyqizfTyAbgIgVlSSFBe08XRppn0pClDVTEBPT1wwz8/EMSutNo76N5Qkk+SHg
FCL2gjOmcAzyZd+RtCEQwsmgqBWntQocKwg3kLl7XKuh0WPjHbZ4Z25Mtx8v0I+g
EhN+d1ilmIyNJrUT8qbSIL+Us4X1c7xud10HMM/Zqe1G/fv8dzxqCmeJ0dvo8eYA
S7L3QCGnWd5tK8dE1LkKRuJY0jMhBiQVTD7utTQFBCSHFT1nm4PpD9SPIorApkY0
tqx3JI7xy/Rbt7boxHyGyeJwE4zd46OKKQMIzruf61XsgPpz0oyVhkXYRMg7Zfey
rCpURx1YSnteaE3lZ6z/pW0xMi5XnmtR263NSob8t5EYYYL/vHDZ2ebSBDMXqX3k
6Le7aEEZzURclZimCMa7g8/Yh6yqWFa1qwF4gvD5GS3HxC4Uyze8guay7xrzXjw3
nQZRir6qV1xr/KHozuVSbFioAgDyQy9bXyaQbpJ3YkoYPfM0qzaV2HHHnzE9iqKs
jskfykXBIBiC/vl+YpxHNi2RY+5NU1h2AFmhe5zHHPw/XP3+UPLvvolj82Zz77Ue
Tl9ldzOcjaM3wt0Xy39vTJUA2jwVcbLObMzNXi6Kw/ro2u7FGVYtkWwFkTslzMAq
xWTwj74Y+bOH6mBdS/7yjI1hekNyrQfdshQtzjMcsvZjdeRxGDOGcrMnJ661vOrt
0ivco8XMxAhBX2hC2FEqTbgp/sncRU0nhE38wXHTXivGNqj6XZlPCbypYnGl+BgF
kzppnyD+UHcMoXMe7jVRCOG3lF130vYcI6cCQiWP6annmfj6jUFRp5AmkudO7zWQ
MsdWmon5DbksNP6yoK9sjZHK1v20AW7HTFwa95AXhwdZ1SgqRa2D1mfk3U+Fpor1
3GtnBa9uvL5Nc3qsfybzGeK5QEYOdRVg6cC6U/q8U5U/inQmgS5xAUfflCE1JdiO
86InRWwgbuI42pI5eHD518gZdld7qpu4HlaGykhH3IyC3a0ccz2ez91f8RLxhy/T
jSLuyIY64q0I6FBOli3PMgZKMo86n4rK81MLmskt2anPHb93TKtjYN8AlMsNyWyo
6L+3L07W/6tYdoOgD89GnHhnbj0GoD/vDsTit4qnboqivl/EfgS0dPfxDUlBHrcL
nH9t5/+2d23b0lq4FATup0Tyoi7r/Kso49FlxvY3ql5qQaChJudc25NAXFtp1rMm
2sj6Yol3ZHaPONvTUL79Jk2tDWIst2oDs00ZzrJICA5QvyL/9HlWmh4p0sPKbgQa
hVt6fFRxBM1DNHaOh22oBxT/v8EElo3DXYTu4np+m2RL9Yt2l19nY2+q7xbNjDWM
X2cfMQZN1/hwExNNh9P+soRTE+XExpjoaYJed2cCyg8U8+8KWhfoRrMxVvO1h3xE
jiQVD442dskGbThAPUoizxfAHldAbFKAjPJIslgYIHjLgBvkbDA7bR40mD4iCrUV
nBbeC6pVf4DTgpkKKoyiX9OkHsWX2f46J6vzGC9i+z953CiPKy0d+OBLiZHIRzOz
gF/oGG+1qHK42g8y0Q2AF2JfziBfHFUEfHcwuVu6B3+gzTviAeU8Rnlpri1Qru0o
qavPpMmpMP687bVZZci/L0BPy4pgyWZpwuBekZ1vpu095ZHhDqDcagKjgIoxsPhX
W3kdhb8uTFfhVq+hJ4KFvH+ZtLisa5w5aGG0FIh95SLmvxbI/ex/6aq0BPy8YvYC
lA+AuI/+aAUIFWXCpMql+Gy0MTG+6E6YGOUNVny5MuiRWO5iQZXcdODJ6R/3dPyV
eR6xIL9wZ80JGZMXjDd+Tg9o3ig3+MPZfJvx2snEY/u57tXCdtXoGgkpkDmvIWEh
Rd0rSejYgfLf2iq2YMKAU61Y9+k2rFKIrjQy6BrJ0xt0vWugpl586Arr1VQuSjPZ
p8ipGKCDV//jkEJLk6A1ZeFmC96Stkhx80T651w7iNdgQ7ufP+2g54DA3Symrklw
ObdIBwoO6RfO54S1lRUhPzds/dZnEP/HJf+T6eSdNYx7QEwZd5P1ZpVmkOk7ubp3
3LMuIR/hcHbVuYSU1UcspitActWl77ikyb+Jq9+lqIBnfvJiFxP2ACt2UGZhjoiw
aEC6jT6IkR8d75QaJlKlyNaBU4Zt4WgpJEkie0lZ63JfBqQgpP4EpL41uspMLveB
WADbnY3frc2roilPUqGCGUVlujhwBJJJAlTJMeJ3tSaI9n0tpzazmWAktJNqrOj+
uAIlrNbP21hmJnJz+M4/uvCYOJvZlG7vMWqabQihGesUfeulefnOMyoGoC/AUjXW
WKcrQ3dJr4ajQTcuXIquZHVRrcvsza+zNgpQDZHjWW9Ab7k/wgJWZ5kHbFbgYjzi
pOabSmgtQbrK1WzO6r9Zk7l+7gB/AorfGgzovfer0FqBZVRFtoh+JsW/N1/6Jbyi
wKP18h+szO189Sr96FPP8Ni1cdIP0yT/A/rYM1mVW+rHuDdXHKomj+stANhmMmHw
LaG/uyTVSUNqqsag6nEdqnPopfh4DaRUd4p3+qPWl/hPa3Uq/VrYZ8rGKHKsubyy
S5seymPhlhcWixROmzRPHaVgFRK2QcpMwowsl/tiEKKivDZRZuiPYFdbKbqXottD
TOvZWrDii/dsdNyNbjj7/1RMnNDuYmtzkyp3ih6rxtkuel5mbe4pMN4nh7zlhR23
Gt9q9pHLR8CFzltgp5962ou/MMgWtuRL666l0Z2zLggB81UlNtljLSVdGjv3KC/g
IIGHc9m+5e6MLDjHDwTaXVKUiNSQd4UW6vWN+Y8fXEDDjYm4Kt7ZPlhQPeZBPfJ8
iH9KzxrXPAL0nfkz9dJbTfpSVyIsUUzmBs7A+3KoWJaO4v2ThC6J/76DPEB91P6R
ARjTuavm9DxOoZvmD6yJqAE7HtkzaVsy2i+bn0erLBErIpDGPdPcrP2XPBp/gQ3p
9P/MkoRSsJblg+/TJIC+A2f5wOyFN4WZCi/FOYStH+V/VRS+NDcQMKY2oYRwIAnP
MfP2vNvhOZlCH9izuQ+N9dgSvMcC0V/rlMLdzagT2xaLDci5h9+hJs+XbcSNeoLk
5GyRioCK1YvY01n2gHZqmBIxw2qJ400s3h7wFB2uC8Vg1niKcN1+xXMgGlGaMZPQ
0EbjH0IDys7sktbyEDBnYqHqC55opwv+g2QngIotoC+BMn44/86EoINIMb9rUPfm
rDpmzBP1uuxzs33ohXik8A5E0NrQTj4jiz4+4ab6IVMdntYFXV1ttk3rm/1qrx4S
Ni5q7QA7sBvYDPaBZZfEYDn/cY7SuNY5Sc5VpCSyr0tyZmy9tCFvCK6KWmaBluRQ
hSo5MZFZzZWxAtZOn4gwfnrsA2+rLxONPbmfpAaoXt4dW3oTI3//JE2T3CQ0KKRy
UWnIgC3IsRhAZHMv7012rGLvdHD0PzH2U39G8ZNJaE2Rh1EmCMR94S5weNYo5ib4
Gh1Cg+O7z1+Ce1QrIWzu0tS/N5gSblPd6Lvr4zch1A63OmNogJUKPzeeIdZGI/Oe
/kInBuJVGufxhXyz0Uyc7pGRxPAYGzLb2qlQHJYZdiqgV7w8cdsUwJLDXiuGOkva
mYGomsYpD9+uo5uU74zDO+fikEp8lGnkmcCkTU5XHC8ljdufoLDAn4Cr0Zh4Hdd9
8ZRhIiVRW8EAP3amTnuRBEhlKxOIgl9YBTnCqD01SB50m5GkwwFozYELNaKIDt/s
XI4VCx1X5VNni8+T8cMxVYBmW48rwPbXDxf04IrNL5G82AR6RjDj9G8jQkKsahHq
zXbks1D/QSvvPRa+7j/7gpdnDT72VGgdxImhUn9UqWWMWcRsQHZ30+1yDAT9+vfA
h5KzCp/fVQcLD9TXxFFlINtf0wqjzedARGGHt7FSOFYRX7CZfyuQ4q/ISyBu0Eno
nIeOThzlpeTOT3MCvDOWIOjpME0NalrOf08D5Q0aMJ8swTgM2SjEZttugrPQX5Q0
r7271N5fkERwfvBN9evV+ixiaxUXA0ATbZKaZCYX5mX/y/cSe+5kkFYiwsXfB4T/
uOtF/RzRkyE0G0JDHfoS21m8ToSCry4hnM95czRXsNjpLlVeMjEBLjoZW7f0RAmO
2z94ai6oMeYg3q7d+hgAtSV7F1qTkb8h2kZDSxslNiWzgWi7WDtbv5csAvb+aCKf
M440/LySs5OyFaaZpeIGPYxVcVE5POfzanFtJR1bvk/UdS8SfFXyjc0l+yidq1E+
2LCfY68NtYCeKXu4wa8qwldck7X7cRurRLQx6SwpM3WmnzTQiFnvvqmz0mfCsxwO
aWn5SGjty5V1srdk4RR1kbWYyFVnoeUMjIhDNNOgog4wx5ewrTBGY9kzmxxGPVZx
3Kqu98vYwKTiQb3adJt4wW14g6g4eGlxNRll94RtqP7SqQCaWaRCNN3hBgjT1Hgj
WLuUZUUvWzRpVqQBgVnhfEkmO15Tp03styFlx9jAJL6QAkUj+Ka1dSOopj6aiBxa
2TzGXMp9XoPnOmDJVrIJYQXVw6+YcE747V6VaiGVCAi2Lt/JFfzxd4a8rSwIOy2n
jNDFz6IqHLkbzFWf81tj9578vPOKRIR6SfFNrz0IhCl5sKbbc3rW9e58Dx1SwiiA
bTJHe0UkmZi1N+9TQy+2TSc8CUbInzGIIyCJfdBnWsPoReYWkSNmKR1QqboAq8QE
3OzATpLJahEy1Adalp5bL7PPBVVX7HWxTlUgRU1mBlvgF0WedJlAVOvvwZeLYLmz
jToJ14ely+5D9U2UdmHa1DyxfqRrRZvyj/f29Q/7b31SFp2/VTc+mGxHnJKINoQV
+b0kRfJZNueZzp1u4AXWwdQRsniEA2BqiByF0FYaiRI0yvui2muQ8tX2EVrE6oSe
tmV7Z0Tb5g87yVT55G8VgA0PqUiiVYtLppbTA1QeYga8EkRfIngspiCO28lXzYKv
8wL2S/KkoeqbAUtsRxoryxpl/nqBCa0mTAJcIBltfYa6y62TMJQOH1AOprFGqHto
BKCPU0CiS1a84tt1s4Aa4nZRBnBPSKchn0iLPwPkG4GKjVTKaOZ24GzpYS8uz/Cy
0oLz7OggQnYmsAfQHRG8t3QlNQjlbX2j/n3Gq5CqCH+PssreFp6ZYMGYue8kejJr
HwTcD3SKoPJINB8XCf4p/CzJivfrXJ2PNI2RDYwqqplo4jMJ7JLSiY+Fgvd/xnsI
+fn43LF4eeHN9IoEOPIiFYtpGjUazfU8XGKgvyMr4oVl0EAkGYfTRBDTD29iV5vs
2qWYHmhD4y2OaUbfwvcwcOzC5Rfn/8DyAz4rAd9ilDqjekkM/SKMT3Fdx93nZGiV
NM5OfzsF6ys1YioJyYeIvoOtsAxp84NwNE3x2hAKQR39m4wMpfSTn8iU5WSaH5DX
W0RHB6wz7Z2Q+KOJm/Ne6oxbapZmeoOSSkxUGTMYoxNopOKxPpgwb/mnw+pCJ7Lj
3GyYNa7qapBlup0HryObcNoojIhLJJ62OIQPDPFCc++4NJPId0lTf4RlrBaBMiNN
Ha3i7px69OZXMgMrWx7mchsGrpOrlnKtYjzSnklUeKAG7HHmbeyiIdTsY04idqyd
pL9AtlWt1VJRQG6Id1dSGmTjcYiEnO+xWM1ThHXeLXYHlmnpyh7WJbNWHYcv7lB3
BaVCFTdE5aIYvXDkUMzKK3Whnnn8Nb2OTT0MEDKpsRLVKLZIEQqLzY3k2dRMthJq
O54C9jptOCG4N7ekdXPP+5O83GfOzo11v2SZUhxEUNiKIUlLgmwR2EI3YGXJFq00
DA7UnYkhqoR0CkDy5pPBHlP1te7hPM2WVKKyFiPxyo7I3rUUjkZ3ijRKio61Cc4E
LNEBa9jrIo+ahIf6TjKxPsyZ1cO8OSJ8XhZJCrtJ250+m166Yfb8PECSIIr77Gtf
g1WmayQBJQ9BAcYGIDzL8masr4c9OUsuBZ7i3g2uQ7vRFvdvXWwTpIyM7HS5n4xp
LKP5Ttlc+MHvpnF3gJ4n0k+XrnpNk+2Qw4p++Nm/KuDkvwyjk4yYGGwef7s4JwEE
Dn7l0Vrpo/2ubdUAhQohEw+tWSemnfX0E0cP3SvjmLvuCjXbR55RN/gvwmHJvo0S
UlOpSqdhtAHGLG9ljEK88xO7T4ae9/yoYb1F+F55RyHpTKD3ERP8lCr8jmMkyXYn
48Gq474tQ3MI7HvZK1lAcokk6c6FjZyfSy1hoKCrKVs0Qv9GcKnHfnSsr5D2bRVR
xwGtkWKDpjyl8o5cljJVPrUUjyAkZJwrGvXZGmYAVHc/n8pBHWOmZaDmCIkprHFh
BENQ0qwGhqauVIW9wdU9HXRUfYvEzk+3FvCODq4a1y9VhQ/l6nOyu3fJglVEK/85
i/bOM2owHLkm5JnE3JhOvKUOnIjQtbYaEUBiYZCGjDyxj9VxJvS+98LDOfFEkluu
ajFxEDkuPVIKc7hXwtw3uzIfxalqzXRU+5uWgW/x+QaA+9o6XGxoTvLI3BUKJctn
r5uKAQnDJCF1tLCv81oNwOAsq7CqVE1svzUuuCmPRsjuWOPQx4Otp0QojzLHu0xn
HpAukm5EmKVfza5EpBh/MPO/BZS5YpnZRPPDz4X+dxMZALJ0qFwZW8CiEnjpqHt1
zf3SSAiJeJQMGFqNN1WkWrC5CdRgiVnkKwKi+XusMvCfsCgXCbz14i5ga/tRyg2R
daWVzWc2W2cnVe2iJe+Tc7ICIxHBB0L3odbG2+1jNW8OVLWwtG9fSWK+WxBse4Kv
KVzUQj0kgJEMV2kfMHyHgz9917JPt7KqSH9dCH5wgKegQhngjkeXS5XxBNG6ZFGb
VL9rw8Q5KqxuuMF8+rMuhHyhsAYmSEjXzay332HYQzafxFRArIoT7AC98FaGPq01
y86XcUhyhF9WymiWHvbtGZfti2s7GrDNOENsyjsbuLHhC98WU/Rs4FIAW6rieD0h
4SE+IyK0AcA6U6dtLf1YZcgJVjzauv8i23gUnLBLe/fuvRx3o7R3B3kOEyxvDC/K
ZPhfgLm7ZVk0xIODJD7LvGbwtZYY+1PB6/BnZY2btc4COfNtEgliKnGSNc0svktb
OUkuSVZa+UMSfE7UjYdr5ICTr9lUgOQZCGZHCF64HPrMLXOS6eQ5KWbqsgxYJBbU
+zHCP/3oLCWtyAf+Lht5c4178kCHeuvFKNb/wgDJo8IfVYD99b8x6H/WarW690Ku
jSR5Jscm+xffDAym+KWebJaO3ozxe0D4iRKZe4UsQ4CwM8u6+LkLME7aU7QKeVCo
PqmADgZ9eN1goC62pIdKV/BykqI8aGMAssPuR7Cru+BFuqBHeBHG9oDU2jbtveZK
pKjcttTJX2AtshrISMtVAN8i/IiOdWhmnTeuOQg4pLOQbGWvz621HYWjd+GyzWkX
FpGG22i68/tNBQELS3QO5pYcSvXi2nHfEpdJGlyDBu3ynHFokr9HASS7xYsSTKDr
6BlBvtV/Qqq8MejiknvFyYTgIL2NBMB4LNMNFN6VkHpTR3wBMhRxjOu7A3fmERNI
wiB5vR9eL1bmR5bdOg4cd3DAD4NdQpJPmIThksp+gic4Txqgx1+jjId4Gjydu+7K
CRQIYgqDn9+G1AWI6RcUkJwmDqrxBM9R6LU3bBJakZvxjSxG3w03ahVCnJgtoMZ6
p0c05j0v9eZMLql1D/mxgt7tfSPIG/NwHcVUH4xTdHAOnBPm9qBx1HFi7O5P4N6x
1LochkTE5u+tEhflB6oZAt+7ABIfy7uUqK89xu+7RW4Is08WpyYaMXFbN87+Jpsv
aROyk2I40MLJopK1dg9QFfKP9dH5QTGcMxgPZt5/W2JflLmVEsctWuMNY1A5zKPi
xjcy4DGkQYY5YaZHO0NZrZuuI3Qwt7KI7iE88lyLbKM44Gt2tnRJMvIn5GYQ13Dx
3OExmNNYERVZozJn+wQ8jD8CSBkg9o6h85HRNVc79+O3J5K55JTDJZZM0Tk90xrR
hlauo/YKUQXZTOOGUQ/6SVxqnx7NEpO8yeWVOZcx3RnpW4YbDvATc4mYZpyoLKFp
Bd4plslwT3zqiakNm6TFe8Qwkyh4Nwqd+9YO72DCReDeb17x5uLS8Y12H1/IAlCV
zrtX8WxCQtoJ15kPUlVabXVruaOxaiWFc8gIYlCq78CNDA7BrnQwFZzmJI5RD98t
aFNZoKFgoHk/tFIjc2UxiIh/hM7qbOMb5GurMvuRSA70nzuEpINKaVdX7gmo1QAH
fT/mm7b08UyVd25fzRTF+UMG2vW8Jt44tXIl590VnkcJkMLj8/cg5oqrlmxLW8ai
pR4yiUHbavU4yHlaafWf/oGiF0p1TEXOPcsAZ1w7ZpVpAm47UEgn1O0f9Ivh1j0e
qXEdlVU2AaMAusxq89TqACf5CdRwLNzFSlGe5GLhpMXtzh9ZpJPQJ/lB1tj0og/r
04PtPWAqAreZVIhGerFWIMDaZhXW/RD/RLKVQga2fJ/D3k1COhRI9/+g98ALumL/
1LFmMwaJmfa/cb3zVuaq5F3fS4T66wYDi6YG6k9GJVPds/9lPKyfEACxHGdTbPpI
UjksF70F6RzsF0My6Bd/wO9Krx67Kdxv+tcje2wdsG96l3wL0mkD8g6JoV4smkFO
MUs1pH6Nq/jfOru48xqFAMakv0rcFoIQZnVgosXbNGlnfppGdg+sv2g6if9oiXPL
Amx7UA1TJp499mhCPZBuSdS7xVbBQvqXhTckei83rXelWBU8SfkzArZL+SflyBj7
4eEi896RtgK9MCDcHO5CWoZxy6kNBoFK8iinHewqyLUVQb5sw4U/noPssHaJiXFz
ZNbq00uDWMR60dq9WYRsfq7tbWRulgaNnl80v47sx+wtge6E7Dug1XkSAjCmmCvo
Sgz2CYs/PkOgJID7npEwlSiTCv8BdQoJOtZJWloUqCKaAV/EaRVRgX88gnYIVYKt
SgrWbvvSlYKHUPLGLATyFDOZTs90akSsnbyLqZZW8JREPwpKBIXqbMwvvyfviOs8
kgAG1jjPCICQMF5GHz6FS1Iyz7ac3nC3ZCLEL7+mxwzCwlmh0L+P0yR44tHfx+AJ
3+wK6QZ4tlkqBzPS6zSRqMHqSQfL19NmD1uEfkWte0DuCMwIfyMWdT4XcCIdtaFt
294Qb6CC7FGf38Di51KqTT1QyYBWMsIGkO7kBGi2wz8t+jtLOS+oa3Xnc5pLei0a
9blVMqG8xTdQKselBU2vrTiSHJb1DPf2eSxglhvpthdhcU+CDBZjJTKkM6CzTdH5
1/zP7UkVZlC1uh4ScvlkTgZMXNVrRwhjwvQMRRkPqkLB46Aab3g/K8cmbBihYhtR
yUXHVHpUHTbv22b7/4qnPdIcDsVSwKSFdjsvquWG5AqaGl6Vky7MCp9XGVGdmiJt
9HziVTxNvwQUmylwV6WawB5P+Dl1Etj07tB/oyhECng8wfCm2l2PUHOaNM8ULFfp
54O3P8FE/963x2IqRkVv6jDJl0zkOpUe6D/90V5WsZJnQZjuVfMmH/gmB9lFH//P
7Pf+dws06nBeAeV/5mDQUNnGk0NNIJpYbuwCslxZ87dOgoJNwz1x576hyQhC195k
+NPMHqsKwLr4tCpTUdPPhN7UnCLsATqi0N2TAD0/k08/sJjECF6XwMUCsLIjOVby
Ays1fWHVyGosGNqt0x3rwmpI+Ydk+DPpc2a6ETLTMq4EDRtuzks+BzC/RIuXzZIt
trmggnpzLAmpsrUzVowCaSnqOlNmX3npvTlnW3y9t9Qdpsvg47rwXkzXlphoo98M
g6ABJG49n2ksqXB8HTbkKh0/ArtRD9EwA2dEjCTGYubH0+4Es+IYiwr1fzt1SgZr
gmwVPcbN4QWJokVB+OIzQKAGyLlX7BXGyFnY8bMpgkNo4jPMeR3hDwjeBDpnbNuJ
CWuxBqinhofBS3uuX+UrC5OIZ4xZrLPD/pCSirQIJs4M4Fs2TsCuTHFYFMQNuBHD
uBKpHhF3GyNkx0VOug8TxI4PRL9af15Nbl1+pQfZzGDulullJN1RC4oUdv98diVj
bJd7QEMAnof7SfdG+o+pN2pkfILhmomQUHQ+gOcsa80sFFy2eyZXaUT45cInnX0u
RWFo8zmC2OxVGYSBuRKSn4vtAoSQMhv3kgzug1Z1w7JR395ockMNGxVkxQzWxEcV
6ecGV7r/b02Vv3ATq/5usss9ARfqJfqOY0qRe2Zt04RUdX4trVjItdZi+j9fUI/Y
kxtHNe7z0jS1i7Act3/0DiVyw+9ekf5wexV0dtoD+OeFz84irz0L11DLXTKTRXSH
oxhWEMvyWCrMSCdJZAGu+1OXuFVtrpFwCaQwL2/kflLHe1IYpXs1L6w5ZfoYgvHh
LB7WGgrCvJopokNltfiTcZochbi0VhfN75bd7Ek36YDU75yzovto645U1KGDSZOQ
pVNQ/YgZwzJ+aR8eEaYvLjo1B6gC0YKfTzgBaPDOjUz5jbYv4dGFbJlpW2SbHPGM
dKbGeWm7VUPGsTf6xuFri4TuqVGbdPyaYr0lFcMY5zHGWB0nUs6k1WQr8IyeMZRj
NeB+dzj0Ht1W9tDjZPX4HXxIw8Uh7n6Up6v6GqIkx2TgwQ2CiH398Ipg6nzow86L
30Tre1WNDI/Wj8Qs/bNDeB4uPxVDK6xWKw60gaYzzmIbLorE3g0XQQv8LMGeZru7
JHjLhF2bt1rI2X8Er7TRjeTNvTox7UcJmorNwTkB4WDfCRduaGXbAFS7SWm8nrg/
w0wsVP4qMzGH14oE3cAg91AjJGfz3IWcTTTpWq9nHOkHHWJJMtuc56SKRd7i+ugc
UlPExxwVHi03QAFWR710/+5HnQ4+nR92hd092iuCKhpoR4feMPcvVZFNvc7TLPqS
2yc34K5CieT7HZgLbfNRutqkCY7FrQX5Ju5VpHxGrdOgh6HC3/j5Wnmj8feShpTW
H/7edNFWDclb2xWZQxeaUkT8Y681BPK1quOoEwz73YLeAxCiu6T5iV6W3MllzyRA
1Smyci9DqFTMbeGThM6rqAoYER9ZQWcJ8eklegt128/TiOtlB3WYxEIzS4yzoNDV
/2TBUhnzxmtCEYhYPO61xoLlVsNQcuX77svR+k7vBK+IQN9XHhwgBmsWepdJC9Nx
z3chm3jVvnLBRV2ufaO0Upvyz/ovlf3GvoqbccQJyp/eN6h8Y0f1c/TFpndBOdX0
H7/0IHXVMqxXmJtSIrMndki1FFH2UHYYmF6z8BzX6n/utOTjA1/M7tQzVf9vKrL2
t6XB6k6Xkx9Jw0mlBnY4iFO8tZenausiyNmRVdpwWnGKMFKxCHjnGKbaAC0v/VHg
gztqijukgWMOYksAXlqomPrWodwHtbHjdPYUrBl6hPrF7uVKTzengtRge6s4Dyjd
QSyDerH3fP5BqGhrLX2urNCvQP5VTFT3FHMOw8u4cAd4rLABC9v3Yf3X0EboYyG0
AL55P+u+LIhXdV7c+4v+j2GH8o6zxEKl52MapmON+x8RCgtyTsRJkPUhj/Kf2wM+
AK/l6smCueCPlZRybcxp6xaSHxZh33rCI8aLKEH8rLL++HG5uZ6imU6671+/A/EA
cZHb+k7/0rig/j2/Gr7KEFk+6I9pL5Cey4x+rbDAlQprPXhdhkFyvEvpys0yDy0K
aMOvNdEq2e8LNyJo0EX9MQDGnjdN62dlHFytXB77vc+UxS+c9Kp1yeQtpzC2KXO3
ux3NHz83Fg7hSBa72n/Ia7nBd6KiPVeR8f7dMhX/9UEYQTSNt73eyKg+9GqztuQh
LMw+d23rJOp71kLCovaPPUzaD3wqOn/4qJuYotFvaXew3xXAA4SUT2wvKHMBrwVq
S3iM80019vEwcdXEwCDUSddlUWVAmwSXcLyJ0N3nCNKbXK/tgW6/RS2MfqJ5oRjC
m/EQ3p+aUfLz9uYS75T5PTgujU9e4xwKyxvJqpgyduLzv5qJ0qMRB0roTBRutWe+
XVHTEwWGOfGyIgz9m3IxLzAoiPUBn5YIKSAndyuDR3J5Wsz9tZLfBIGFdz4OlBBD
qJoca5rHELfsIUKthZqX6Toj18jmmGrOZm3e/89iFiOT3nU1qE+Q1dmh1WGkGGA6
OmY5zWja5JHEfSsBjIp9e5QAD40xfUOZ8p0rti68LoMvN6zp1zSqBD3fci4oTYm3
FXE4eXxEPAp4n9zmoQyfr22wHwDQ49Y3T+76zZm3Mz2wvHhqauGlR76J45YKZciD
ZFvV7U1GhMPubnJxQdmFl3Lg9bdyRBS+LMebNK2SVfy8dmji1ywCCvzgcUD9SCMY
HtEkFnEtEUuqLHmVRu4Fp3CwB0nPZLVJvCEbHi8ZbGEj5VVnZ5SjoC6nchuP6UPK
cEYs7owBi1yby2p6UVGSdo6+sf4B4V+s+EApM6z1Z2g/TJQD4Nd3bZHQbM7+hsm3
efuEsbMd62BKm0f++79IeqbqLlNbnTJwuVqoEIF0MxES7iCO15Pqda2RMKIU4nnB
m81wUSZukabChXMXza+giIoOIP/nwZys2JydvTaBoJUPtTMolY87wJRnxrqNge+O
KXt45C77et1p6HZ+uufUNyV3nl/hMc1uky8cp/AKe1UmYok52URcV2y+G+LwdLsT
5hAc/Y269YiwPIlNEPvRJjU5vn6MUjXAkd6HUaf8/JZn9o+gpXqRb3PDVSPUCUFp
DU0bTPLbrUBJbTP0yw7WNzH3Io84nBTrXOrHb9/kJz6HZ8tnoBPkMwqAAtXiN+Xo
SncQtziGi9DDl4IZlX5pYz6aBg78X59+O/asQ6yS95wEozl7HrLU00yAdHu37I1F
PpiOazAen88MaDaukyJhm3gldcpbRxdPP4eVMsbdar/fmdmfGKLDuz0A+8/FijVc
UnBNNUAgDFJf5MP00j5NhyVcTrtMyO1oXbvBZrKcra+LgCvwlkVzHqIqxNP3p+L4
3dwYtcmPR7mWaofgm9HhiO7lytjYNsczlJaYifZfiONgvED6QYIKI5psbYdjyOUa
1sUl8xgx87M9PSajVlZYPDFB8mstmDWMWSj/OqPOT6Qf5v/srQUxPinXdjRKa9YR
QfebbFt6A33bq7M1FShBj+6cCGFcgrgs68pvMDWD6t/tGcQkBLg6JmcFdN308uV3
rpPb8Sz+2jN5gc3dSMZSt4RTJvuyLY+3m6foLXRVOXGvZxpxQZs5j90E3VdSauXc
1JQYZ7+OSUkpPzl4fweYEij1hh90v6cIytY8gZ5vdGgK1/zW1iPXPx6M9DpkMINr
0NZjIbT1IghCArcwAp2aL1VBcoVNqksStAnNScRbGWt+oBvTE1ZAIy/Ou9SRukG/
6hTQ1DEL1fZq/mAUWq4u1PG2DivKKzUYzLZ3LJSecWMaXvYFi5v32p81IuCRY7w0
H8xnRlnFDZAQBZ6O1aEyb0pkEcALWVMMpqd4iHzUdIKNfq4ayZsnr331OrDNlNhM
tmkaYza0OVNVUU+Co8eh6yaOmxz28zrC+a+MD0oaaHulHQKmtQ3F1scROQh3CS1E
qhwsd42IMFe5/CNkKrVEii3kh4h1irmXuMwVQWbXHdOVvSKBvTCVjpHoxX0f+6MI
rbP0gFX82oMYYWHdJdDvgjsCRvD+4xt4kAA4WqFRywXQfmnE7yTtXFoM5agvYFsD
h/t7i+jR+pjaYlTQ2yGJmzEUZUvr2+HsAYMiohrOkc92fIxkVyLtmIoy3/CuiUf6
s24IZksrRQdSp4egMMpv7Xylm4fdxfYJ21rNa9Y4aYIEA/tdybAT88G0HApAd42G
vBhtfhmmDucBtPlKcqkieM3GjdKflsMRH3cgWaclDlpLlfltvAoAS4Z0A5acByeG
BUaFSRb/eN2uIIa5imlnIY/jfVMRKxU3tC5fILAjf8JcrrG/BQBMzRlKFqiilpRC
Fe0bKVdRa4by+pOJxQvQzh/EocwzPvks4uU3W9h4kVSXU6LOhABBklxutIXWmidM
ZjDNsD9HO/jiJpHuVwzZzVWfqg2xM18dMiTm/LKcOLhiyMGaEqwj2n74pvZ4pQOA
MVjOArw4SiQQsfOsZE3/MrmnAy2Uclnxl/qv6JpONm5jO3XWBdfeuAzW43lkHrxM
/VUmM2yiVAdoFLKA0Dqt5N8nWmrfwMSznOCWnd6hvA7m4J4ETu6E4qwjdZZ2YQiS
kMlTFym5HCNeCb6FEeuQ/SH73udm6d7A/DJLPzxUS2ZOt9FNKikZ8p0sSPe2MAPo
Nej2FrP+RTSXKkYwuDdmGywusyogfb1zZ38+uEz2LMMVvBp5+j4yWuXW0UJ1q2HO
QTImfdJeA+QpGtRV3pXV0sZFc48Zg5PFFzgLDJ6Bj852Zs/jWZibQltTalB5mdLG
RCujP37ujAJsbX/P5sBscCPSeJ3/y8wcoRD0FrQNbKHc1ofxpG2n7kb/79pWa6Sz
qqJ+DjDZS+iePcFfxrBIBdPlIT4XjRkmxfbdPFPUZcE3R3s9V+TH6I+4LmbNF8/J
V/6PBMpELKns18/qGX9pRDlE0VMhg+tuz4fbXjuSkBZskn1uPkXr5THltWK7HwIu
23olXL69CeWPOH2VdEgUqWIFwUdJpYSxT1Gg4Y13VSoy0Jy4aCfmD81Pq2N9GnZS
QCatz6nLlviAh7X3UGXnzE/Am7KiIwTrelsvVkGZXKP+AXD3niKF32A1ZOLFx1p0
OXUbnHiDus8/aojHzts9Yd0Mw38QU3NrYIlFgX72gzxEiU6g3RhHcFu8rxdo+MkZ
E49bN9LjYA+tiW61lv9Nb0fMA7q/hN6DrcevXdvkhUAavY80YypYDq6shyc0ipda
ObbnDj4KMnf6wUHik3TpvLqmzqtIxlIMRuTtzkG47UB/mawuj2Wh+BazVWbducF0
E0UewpMUZ4FBSLthjjY0mWqNeejg3v2+vZ/3Kx9LsTrKmODHBbF+1kTI61JCWYDF
HCU/YgfdUQru5S9aRGc5EeLwaMJPEHCFfDZhEPXNlUEF4UGB+8NHdZNMlR9D/itu
U8ig+scLusTqyfk1sFMZF/XKp3MrSM73BtBMb4Af3S7lRUySo+eOVhLs3C/c/Ev4
2h0xXQknaSkCCTKkFk69A5vsuT9tHkzI2UpHpxPRgl+oj819+yLEQoki3pizG9mB
KFwDf1J6/sMactwmsWhAfHy2iiMPABuNAmUys9Lel7w1jaP0gfxy3lS14TqE9sL5
mPMZWTNDWfFpSNjuQMmJmuetcbNip+cuYKHBI1FbbqSmDZ+WEzAUZolWcB7p5bG8
W9tIrr8qG4GH8KCegZzRn+PtAcdw8bRBh3YziKu4muecQ4Ptvq5hFsARDCGysbgu
EPTfdXxSTEz4gF28A25sEDwEbKSTSrMol6ajXu7AIGym2lee1oNlaEWrIMeeE7DB
472nJZL5epEiUQuRD1Q4ZRLJuxjYUEt1s6nG+wZK9K9ZRy8evt7LDPznKGUMJcX2
wlw6C6W9zDOvsPnh4N+OntUEa1hM5v7ya5p/bVcgTi008WMysbHBsShiJM1XX62p
l9Tppn4C5o8DjjC7l5DUrBt/6bdLwz0o3kUnz6g3r70xRqZBEjPy9wWZLb8EW0K4
AJCF061G1fIHk8vWCaSYW1jsBfK7q1bDfkIZT+4+5Nmo1WZHjUZtq7hy8IO/miE0
yFpJG5taJ7ACxwp/kcaUSrNZevVFg2p52PMulVXp2JTT0UUYo40gDtIIUprqhav4
+VkKzTFuC+GWjnCemlJzYH/eFOQyKXiCjoRH6hqSwTgnFrYGjF+mf5b/lk7GVO2o
NKawnlg3NHhKhv4djouKVPD+OIGIVpUdcqecuEZi7GCw9TTCjWFAltIaiFy/2ep0
IinYhOlMF6wPEp4Nd7Ufq7IQ/mlOLN7UmQrD6+gjNhayfEOej99V1mf/q3f5bFTZ
6Nn5lshqeW7co7eCB2ZXZ6wyY5LTZMdFB9reC4cdhNMWMysAJvDMKKQf0L+G4E0z
pKOWi4QX8XZH4ljIRCe0gJps1LzggBHThkzdEJ6aZam0mS+Dn/egiOb8oFGgzxox
lZWkFMcuvxa+daB1/TE9eMvoBEYTVnQsMYOaZmqG5woi2l1tJFAqlOkZ2ZPWVDZ3
pgx1f6NELrTScidYZmsYDSqUOTPVnrH/4UswRdfovplxRPxNOz+n1Um8s+qOXTWw
WQvkHFIjuAZAPmKVacpfq6EiyKy8X87UtJGT1dg+PAehYhw5BwkDoAjaO23TtCLk
3MBoG1Z1Cc+cF0S5+m9WCYE8wrTCkjH5vo3tTI+FjTVLoD7D9iCYD+U0KQ0K8qpH
90ATg4z7unEHyehjAcGtecQsc0santaHTD/E/NJHsPp8Z9xkOBgSLJCPHGwkBfBg
J8jHqXMVT241lkEnpCqNfu6/0KuuIAAMHNnRJ2541nl7tt0BOOIbz/jS7mGxIbIx
X8wv+5MqYl2rNYL8J1A9fea1+4Hdmvy8b8A/D6yOXraqbitx9OHDRVYbgdRqq5Jt
NuHSF10HSqtOx2HNYKMtjPij6DdVxFNEgpa0+BObgmWZZhEWZbqwN+dwtYZFNFib
8engIRXipZF2xhnA+QGJUkKys2WXzmmSP0ZPXJIkoXM1R1AF9bc5riuXgXIpCF/C
lFe3chmi7k5De6MC9I3X8ZUjsJk1wZEJKGoIb1vhMl69hCRYFuiAJh8gowMRAM/L
HeFro2LeRos1tnaEOlJOKCY+SHdApMHsoV6LdqSchrjomPr1EGDYlzPjClaA2ig4
G2k7tJbSGuAEAYaw0BrJcYjp4J7YoF/iGiYib+YqODvaSJLupy1ssq1AgKznLGXS
nkx1/Feyj3WbGG/6tKTn6WUnjWmf2nYUG7bl5IUL2bD/rEFVyHVr/tX/fuCk8hGN
LeTpmE5KkqmNreZxVd2hu+XlfDiJ47MqtPD9f/1EnH3Xuy1xJF1Z5oLFxxXUwpIv
SsCfUDgh9L2IGTGW9A+X+WtsWCemca7CyvYb3A6YJBHup/VkeOoOAuo3128flqU4
NXDppQHeYYxBb0OgBlbjnBdr34l5OMB2zKLQmydhxQIKkzoIxIhQhHD7FFKvko3G
2vIYiZQ8HNaEKCSTY55fjBlwnjjDZwTOY7dtuH1cQg+z21vSlbjehFVYhCSt8EJa
tFL5+cbJ+kmTjbTSO1BH2aTnUN7i+kgyODA1tFrdp2MCdNwbWNFGb7nVi/clymgm
rfSYC1r7/kcjmlixnIbBpaqDOcEcy1CeX7E6RpAFu17Sf8FAXE6Eq+AhDamJov91
mfEVXTJPSiH9oKeKj8JWcHDM6IRn4ZT3OSjQNTO1HaItzb0SxF+WBh8A7q9/x1PM
tAb6qrGB4J0jskG38/NVjIAFZkHbV5xqSEPbiIxG+2h79INZAf4z8FyGJ+TyxqSx
wtatlGtRAiHz6sZyslcwL3obFnuMyZfH6KiMyWOMl6SkYQXPc4PHRpVElfcgcusm
y1zCbIeOwCU7EpWzlFmTrKQIvOXZI2SHGe9g82z/Z9NlFA7cVhI/9fF3GDJS+0My
bmbUAmBC6kiDh4E79QWb+90GiSCUJmHxu7kSIqbi48mM5J6CNl0TNxhTSkhOt2Wm
ASQ7Qg7sKdEZqLfyR1GPphyL7ZbZ5R4MY+1bWs1zoS122C0N5ycOysCBYDw5thn4
x16zZZbrABPOHxxuMhVZYE7qdMDKTozrvdF9Zi+WSEmXPqBGHEX4P71PG/y+rEGM
NtX5upZbEMhphJWGdvQJbbdjipBWTKlZysajzv9OoqsdzVsbMD/GSATLfA5T8ksX
o7/jAkO0DR7JMeNGHj6r9GKp9s6l/HKrwrLmPXsv3u8c7PehNpGXO0MlBagprg6g
BoEc1B1a4AYWdpZNjBH2AZOvUwoyTK937MSOViEXhhjyRS4JuZ8yesVbc6OtCQfx
j3JB1V4CT1wYlmM0N8MHPacTAPd7LY5JSevZW83rKAqgfkTiXWUFwI9ca6Q2z+fn
IwVPAgW52mUPt4JhzdJITIoOqccd4+wr2dmWkne9gFfB+7+XwaU01bPu2Hk6ZjJs
NdPL6SI4Q8dt7wa7J7+PcaqjRfVW0CZvYg6SmHx0xRoBdccnnHumaYZzKxcdC7/R
y5sz7URq3HkBQQNqGOWDh1Q8Q8afs9Y+QPawrAxTnC7xulGJ3QFcnhcAoHtwBl6N
EGKlTrueZX9WyuPHiPomKBmmP8vh8Ix/9MRYROB0lztVvsrbhZhQZfEZDOz0SIuV
iS10OuYngDl80emeRsuKt2O4GUVKbWahPqa98sRrWTvU/CAthCJGsaXtAn42SpVW
8k1aGSyKD+gcTRjJfg9Ryp+F/3K61wr975waHkx1CCZGqmJU1m+hEgXvsEoZvPEA
buS2EQvUTq0AkLESlEXxmfDfucy21/PulV/RnSNrAFZcZWTfat0yvl1PD+oR782l
AmnFLOx95SeFlfjeXrtxv34bYjOI8D2Mh6w17yB+2nYWabKPexAkLEy+DM17638m
KzycIwRyeZ/jHMbSrYQCz+3t+dzy0Pf+u/NDAvuWD9F89GXBvny/+i11H1z/R2Lz
+eDBO3VAigAzewldHwjwFgQJakUGYA2SPjblB4X49ou9TaoKQrDrPTYXoG1c06ay
E13oEgt60xlJRoEc8bF+kez6e9Qwp4KNY9iK1KNfYbr8Z5IabtscVMt9WvsnXydx
d9zlORFPFR0uTU/CsVfxq7E9Ko2IgPZkYVCJf/urLZEQSRq48NQdAEWgqVgmjjDl
siXtNL2WfKrdr2gSRorxWCpo6ABzlBp3Oy31cETjLb8FxGwIG0AaTqpIZdtPWJTd
sasz6Oq9EShlWlPWz1LE7FCu3QAIR4D5aQcvLO242ME1jWfTzJnuHNT565NYfInH
ibAhYmGWlkxRq9PLyNqqy+nRwWDZ6cwsyJxie0gS+rf+5eK2ap7ZhDn8LXQiwJ5P
8Y/EolN/SvwE2QlYOCVI9VTiM+GFQgMPiXrnj3nFasx5y2jUBe8p0t/6al1G3Z0J
ZOCZcjB5SKTkdkAk/45MgC8syaAv4zMulL363RZIDaydaX9Ta3whKj+G9rTHwx8j
GMu2373r7kTg3w/SJVoTOVsItk9NTiN8JxM9IpViCMD+puhNLRoL/DUEdnOooPw5
6FN/ljznxS0VMBZ6aDo8k5yGy0jHFvwKmvNsWgpZAHAH6ZKlwNxgrO81a6IBzKNx
Nn9IKI+5tKNh2Wdj68ZL7p5SBHJ0FsK3zCfSKQBVSeWlAGSbqPa+jFWWD5CxmtT0
1tt9a0+fFgaXYWHoCzQ3muwOGQwwR3Py+mK8ZeNuF4QT3FEPpjvjZ/JV52zowkjZ
zTO4TuXoNVSu4wgD4DmXsNLUfeLosIr3b4xSENQWc69Ggs5kpCZVJLEDqSzwjdA3
MLjjultCvEzZpKfrSkqM3GXEh44yVSqsatIAzfuX/S95BagIy4wI7YVzoPf6mksX
46sSM01roiomPnFKv4gmv83f944JzBC4nRd13sHfqnm/QO5MrhXplqe3gQi+awrF
V0OZ8GWfkJ6PYelMYNc4CQZrVmiBPtcEQeZYhOSPSL624iQJ8i2nQDJeB0M/tibq
QFrUfJ5/tY6N+1KmcUOqRivRrIy6iEBkVrT+zNhtAxiuQ6bNMjJss01cZP1CiO70
OT7TUNG/q1WToPc8DYwbgWowujqISXPfe6fSd2vISVe1jASW/g/l82InZjvpJP6H
0U8/A9rYlNIwGf32G0qxP6hWzZmgQDZAM5UlrOLFvbui4KO7540bX7Rziotzym6o
A/b+k0YYKXL6U3DF5cyZVIc90t2mRUQ3WqTg82rOk2moNBFiWC4vVx5PobJ2q02t
KaSxSEpOtKo62bmsmnYP6Et9Lzay++OXZvDVBBzVXkOD2K9NGfEOfbtGlSODylA4
2tGpfutgmXKLlC/6DcvdlOqHT5w0GgvQ6Vj6lpmhsVBQAbvXHo3FoQHMZGS+qvOg
wizhswWGdI7vk3YYAIhPUfi2N11g6huKyja/E1cB+UTxUka1PD2j58KP4bf/eMab
B1vlRi2UpiYTsg6UMHzF64c3z03Wi9hX51hCdGcWejo8E5X8ywxWE7UtZSfyzHCL
AH2SY46Us3ESSDATTGbf4m5MVvTEaUakJgAEcQaJPLdcN3PIzMYy2H4wDCSU+GbZ
RhCP245allguXXO7diWYtR9aKPorb6pk347F2Sc4RDz8Jzo9FJ8Q+JBW1S3PfJE2
NLSfb9yYgG/GobH9/LOmfTf6sBEBkI5/sPNzXmsxd9ww1Y8qMxXECnYnndFdpi4+
Gjwdzxv3fgP7SoBNHkw0i9ciSdVIjBK4Fpa/0gzI/jWoBJXfYUsSB+PgLyw4WFGj
K0Zzu7TUvHWmsx08xgh672ySlVPF9jmgeWhGmo2RhJGKuWy+wZY2wzyx8Ym7j4fV
RNiA7yz+Yp0DKPqzrI+2Ldw5+4vMb80S/b+pUId27KlNvr+u0M1FCY6XqppFSXMn
APk7WhYG5ji1400f6NyWcboXNCOQVb4DZO90Wh51GjaxAZOoLYMKprE54wiSfwZ5
G2NHQYjtNgkYgAHGRq3XcelREHCkdntkYksb+NAf6YkToKESyuo0gxPvFt5Bxmwo
WThyMOFx3aWNGargeyfeWK5v/BrsFnjbEnLhCWOtYkVrh6aabXD5MJsnEHppViEl
RDCViiTxblK2/X7CloItqI5vMHXTUl9HgMxTkJ0Qfo1qIY8WhTtcSYgK+kUFk4lj
vs6B+wPJh/vGx9Zo5nzJ/d1iumInPKTBVpDviPyfazJvOU5Vao5Xv9OIw3V0bRvj
5k65YGOhiopY2Zvvkrekkjyi63QVYYjJpUym8x8JBAF6AcRXtMk5EeYOgKFCFwt1
Vw8SnYLXWfV0jZhVavjfpiL/HtEYgXYbA8cgVGCM24peWNs/KKnCwMiOICUpuSVc
3ZlT7zb9i5jLGBtTrt/t0S8X4B/OFYyg4bA/hA8I39kj+nMHhXBvlPf6Ni5IJobW
/XQIH9X77haS8S/ef/BM8FDlXGyFQg5kwCgvHAc26HEvNW9w1rNhbijjeKoozkjx
lQRnKSu5jUhHNULyXKo/5NQ00s66S4q7wALVLAk7pZcerGjKaWP6juN32JEPz0ve
G8IxTtmAM6Vs2/QSjurJMadWTMdr5FuY4aRwm+2uRsmL/zofckGTsrjA0xB37RSd
2IyGjGYFiXpp/jpiIcRYCdrcfu0sdcxzqMLMEQcmxaXNit4Bt9hb6ddeufnT9tLv
uj0oWPs2o7O5kSzFkuC0uKNpkhOvhptAKwO3aG9mlAxSzEv3fIwtesVMhwxrPk2T
a6HoO/bUqQJbpOCtG56MEIfGb0RHcCARb4VAhW0EIk4HJOhq6KEi/yVFfLvq7lHI
iO5DKyTSNgQUHcpqfAmr8d2fuKq80Rqbi8G9tbiH+0DKt5P97qw0vfC3huWBJzQP
fREEAgw6EYDMC0yoPKBGphc7QxmjIWv2e28EyUofoVfSJ4LTWEixC1nxtgL8cjkQ
043hixl/e3yNBDeiXCaP+ACSBVxyJdd7mNqrE+er16ldmKaqR3GEgOigwZX7t/Na
SAaU/1ibYChpJwb5l1MzXcbRQ1LsDo71GJ1Ulh9DTAwePopCxVmb++TObXEtvpKB
KYWSI7NS1Gke6iXeGnqbGeuR30q3vnpjQhVQcLSuvtcsCww2ucVX9ydF2L0xcEOk
3YJ1tUo6CFi/kenkPeDQAzmIeTrBJF338Sb7pwx6OD06pAhiD+jDroBdyyiELfik
b6asoMriGm8Yl4A3W7mQEWtF2D2OFJYP/2pDfi15SxolipQ2L0mzyXvuGgQeABTX
st7VYda30mYJfGTVtLnDq49Gn/nDN7PM8zFckZ+W+V2I9ajrS5xxohw70VcAJ3Az
Isl41zsdsLn2a0zpXLu6o1mkHfQy1T2XN51401Ar5SSW3riP27UYtj9PN3OmjeaN
V6tiVqEyH4oaNFTLHQC9Emw+CGd3E93rqalR0mVyeN7+1nW6VrRC2wK3VnybDcNG
R78rG9vb8M+GMOSwmFUer9cNgZILQYIjCbZZiO2FpSpUJVGzUOMjMToJgUmf0Tmv
CIdNlFYp12BdxGR4WdIQ+IW1FCdRn90ikN0ft8K6lC4SqWjLsK/x19mU1hv80VVZ
nma3/BohqJjh+ybAqmyjB/ikEU++yurnbD5qumB1mAl0yoH42PNV26p2W+/xULCP
GVJTYJw1eLwl2A8hDHUBbMu6+R0vOxiRecOWUrFiDgTcoKVxk78yy6MQB2RIDY7q
j+5Et4nDN1WGnGmxEMONLm2ppffAf//1fkZojoZkTAO89UYb7qeveE4pYfI+k9im
ga0gH4fk4LXVCrakbdGSfO2OiIr+VHjBwfaDoahlA7ay7G7zhySNVjqTf+EMkY3t
HF0POG0QMPq5YCtEdiKK6xdunRSoWl2FkOxqX9YHE2EUOuN0ILCzQF/i38+pXEcr
BUsysdLoss0p627ehFaHlEJnEPXU9mTOjf8QPyJnDW90VGaGbuAFG+CAJJXAdFUa
4369PYUP+KCyF3qrNQBGzV6mfQHUoUX4FOQQzWM7XnqtpIDDs+6IDxI71Hyy4mkL
fw0I1KGubr6EtNKh20CdhuCCMoBLK8JAFlE0lL1/8IVmgT+7Sk1y7BWblxyaFwyQ
829MSg1kdoWqmE1A8Bs21t9hsJTP7KuJIiKC5b3M/o0lZoRo4M/6XskmXKi5UsF4
4Xv9Lcfu7iY49v4XeBfWWPhbyT2jXAaq/QROLWSXkC5rHeZSfdM4kobdvZVZxgDK
sTfsb82EgTRhzQfCbYoCtgN8TbRwOdnSCxQ96L0/UEspDWqMYCsJmpGH+mhheC5z
eiLk1EcHSYv2AoWMRQbDR0yMOu6EIjdgnnM4aobMjFABVra7qk2738cZfTAWHodp
+rt5FjQIDIYm58MMk32oTXvoWQjkazHif3CStt/9W6AeyTqzaR+cLdtmGCXCEkhT
wZ21QcZ2LegVCWUfl6EN8iaE5WIIup6ndR530ieHl4EghL9WeUzORWrDZJBdvkfQ
B61d+4UOklIGI2nT5A6ysmgg3Kt36hyVWdJmn1tl2HC0Kc/7H6YV03+4XQqwxnMD
mnSE9/XdyqTyV0Kxvyv4uZHKJUs2xg5blHY4VIpUKrtl1gP6TvleIBvjaJMTWqe2
KOKjRjyuqwpiJeSvhdxmW94IlEGF1tc2EpIu2Fg9oAq6sgnH7jrVN6QurOc2inWD
kJBOxJPB5vwsR+t211r8NnfZX1h7QOxBt4jolmgOqBAKdtxKOJ5PFjBWrv29nEUU
23MoFveuYtnIQdHp+jtZc7FG58wOaD1GskO0XJnmUvtGQIwcBFUtoHFe84EUdq03
XDWL9IHg3Z6emmBf3EsBJlCLYM88Wjo9yNXaT+Ch6ZMO47icTg3wJIIu3zjWZjvO
PYVk00lA/jqCpciVPm7/csHk02+CeBHvWsnDYSymaSsHEg9aw5rU1dlSeLt5L9Lv
21Sf9oLi5+NkmYRew+uvXUXNUhIkEQCqjVOm+p1u0fy9B6bEZdpcLgz5qtqG/Nzl
fTQy6sKIqUdG3n4deravA5CXKqx41n+bcMjLIqZpYbZlqFVqJ3YFQhalQuHLitSO
dndqKhBMJzMMd5G1kljppe4RMPT/FWGrSViOa+E+fbVz31PlOrSQCDm6iZsCePYJ
+ZANYUD/Uk8syGcN4ufexKduV/EcqAzpPTRMs2NP1zXUAn68A590ZKqQz3yWj9og
ZtxstMRg54qwvyBC3iJHSokM63xK+vLd3Yf+JgbzeBym5Gmb/s7y29RTHLESgd4a
eG/1HGjqcXonMonVO4z1+ch9SRDByB6N3noAT9cNnun0qKbD2M2trdLgY08NZsFh
7Hx1QZ2gX1tMEEmKr79E6aADawKsyOWvIl3xDUl+k5v8n5xRB1t4JYZXqFR82gem
Hs/GZ9fnOtRzU1KJivZK+7Z5jXdmuH0lSWU1CGgtSXJjFWxzU9aKT4J0BVgu5XU3
EjB3O/uF4lJj2QfMxveVWzDCTqKJ23ttSyBvbQC09JYr1cKWvzHsy0swlzx6QSfy
tpzLCDlWMmdrPupkjNnFqE6c1yTesv50w/Ha0fWsRXLrsTD99i7/s/IRDIUBrfvI
8iSvrq7UAGF58FJSVWwvYp6+/sUsJqvh7woHOGRP5Tqhqv2LN0HdWi2fbDFYksvA
MjMv6kFmFzi24CLRdrEg7r5G92TvVyfXbzIvuAypA/Mvq/iin+ZDEiyPdF2raQ94
07wZ4SDZ2GBGAysyZJ1i+cB86nUcTirjAgq4vBjm3APO6LLZoOUDX0D3opotuBbp
VA9JRSRve+P3zJmsF8ioKGN503XTcSHDQQFtsfhPbC0xqQQGH4qvei5irdFqlUV0
OS6HP5wtiEwuz0LabS/YtEBarxOW6PVWqWXX3PgbQcV8XkIesPQRrocZnT3MkmLB
1ozigAv+6e1/QvpIwQzrqBwcsxzTUG2HAULNhGdBGZb/ysd5v5naRo7zb3mweh78
qhjq8UzePPOg8ZrbguEbpkyRsR6M2SaP7U/gA+tn1L4CYYgOSwXa6I83yIawPM+v
TRrcTIcZcth6eL5yvj6g2od8079Fx2HHpdcFTfxoNv3w97/4qa6BYvRBKyKtmIW6
EHsIf1UffjlBxB26b6m2didi0+ihnOmBcv4kIJeibGXOmUCGwqgZwayFKU0vnR6z
D4kewgknxBBh7UfCq3JSrEM9EFPn6EQwRN86BOjbwy/p7rT12XAhCWle7YPzNJ+1
1xNcf/Tb6Bq7f5W3UAn85hhatbQfDLdP6cePs4r9EGqN+1GyPy1Kxdp5PhNEgKRr
IBpcRckEgJcpp3W5NMSEr7Qci1CYhgferKbqMgQrIJ3c86ZRQqjTE6qpoHmp0yxf
OUxDx9BHMIDSGucB/KLXHmCXBHCwaywV9cpqF40bbLYJrWHB+9PWfUQCEPbtDgqn
yLUQb+KmvU9uyMD6PHJpvaC279Th6DtffSrq672SX5ucpYhN1uObBfwSVFjBI894
7Kl2VFMI17X3PZqwPdLGGxc9ZLbfy8ulSGzsGp3vaaNrcSBLP6crYlxO1eXCpyd4
c0KDnLGNLzAqKwcfQfyPrOJKHnmdzBg9aWoPEJHkUVy4MlCAfUeMR3TtN2WDqb1y
1GeSp/Y8+gagZ8sbIKIGxudfEdlTO5OP7xVO7MjdDS+jV2yDR2ybpOY5bA8adyVC
2lQ/aHIGjSx7lIsD8ehk6m2DPQvK3tC+DA8KjXfb00KP1hhtHZrLtIH1ovaGZWUm
h27BYQnC9YfPuOXUzNCmedgQtMWJQCvLYcxZXFv3Dq3C12dZzvxW1GF2U+yeouT7
gBsjKcLotYPHLDXJMOxJ6FU5EwQ1iITuDxLilaBP4crYM46P3iij8S69nsg/bZVe
29Or6PHSE1NMWKRgxDGXpO0nMyMI+INhcnWHE5xcJKoFjTLFut7q6mqXwZ4upFiI
5T4zFTJD5SE0mU3IfYqtmRVE3AzAStk5dJCa5FDoUE4uGUKkv9NUwk/24jFgqz6x
zuGpeGsU+R7p3dxeszwKVRJKqFvO8F+04wwvx3z4HZTwuo952cszILiWN+oy7YnO
XYV7Ktz2x1Iv/fIb3xLKEs/F4r4M8k1MUi++70gUNX7KbXqRN4IiJOmvbbiaGZDx
suEF955qSAbetQ6GJHF3zlMUKTi9or8cKpGxA9ssTKNWMweLRkiszC1VVem6hZCt
uz2wre1z6l3PttIXeXlQ2ZyZwa8b9jfVDIwIkWl6K7W5K7+c1iJCvPEAKv3XhQXZ
SCYHQirc0i9opP4nyoThU8f6v2lbcTISS5iWnVLk2zv9lHIXo0Y3yHb+Xuji/0gO
ax+yiGtDs1G+q+pwLfOBSlR2ZHCW/fP+M1saWW0eYxHS7/FWZyIwniMV+198Q7OE
P8II7raikMvo36xCg6jLgK98MwE3C/kkR3hrHht5iaQRLpJsoZFZM70noiJdRi2m
rES917KjEaBRGI3pwnySQCCsGryhZkYAEeTctHAH2Xv2JUeoViDXt+welU1KQeEc
ombjwxz1v2Gfcr6Ym1/0e7IuVjdUwmdtpzKK9EgdHMFi0YLkoQrlNyR1aJV8VHVh
vBPc7+C/U8NSMPvzlC5fji4OOhLlpDcsyVGcX1oFZvh+70ftMx6MX3jAQU3eEskm
gKsBRk01BLfddeY++yvnSCGxQNMVFug+7neLQgh25culQpOciRqT5EzEMVEmrO9w
NTqw0wUr8y6wX4+W2wCHqBB5wJ+2o225NXSt+CNFsICrC9ro2GrdclLuZzF/gk+C
bT5RwA9XLGc7oK6pUmAfY3YkwjD6OIZX2uCGY0DRcJjLUAguI6z9ll8QiGelLT0z
c7LrqVPCExoxxiiHGAxR4eqy8CBzbIuYhNVXE9wZ2F3uFIpp7/RdrEE2h0U5c5Z+
AnYm8otTo49fP5x5POLFjWMLO+PHPK6OmMZDNldEasS7pjcTHNqVSnAeMotCdAu5
Ke9/8Tzl3AQ3nTGm3ydu1+wNp8S1rG3pssXETJ5v7HRa5jZb6mrEWus1epSYq0OR
a/Fdu7dHUcDRL1V/FoP45+eSGTx+xUmYqflcdgva268+3vI0X0/TsNBBP2UAnaS+
lTH/fydx03JEA2S1IyBunV9+yUjz61uT4t9zDTbUsHlLqIgCyz8YAav8n2sxqH9X
LcknI0I/z3XUVQFRwaUDiYeDIX3yKt4yshf9LGO6rURdD4bfwd3ibc0YkqOysSy+
yd2vbxMjvJfZ3ePBComLF4dAXWK2RKy+b/t3rfv1v5jHpiX0MD/JtB6YjQ6jV/F5
fJHV/E+rs/iUuUvcRn/iiIfm9toxw3wRPk+C9+s+Ui+n0ShNQhdBes/cympgqOa+
rQn+Uxg8QSWCvbgOZnATYuOWyQrM+o/nOYzVGbBEQGuYJLBT6/L7Nm8KZl8YPc1D
srvB7VZlX3FjnzxFEaz6kgFKTg2fjmfV6GJo1ap0E5ZENkaWkYRqLuIAQCSritCi
c6CeHy5izwrCpanxWB2uLFEs0dCfOxrcu0UcnCAIlfC0B4+ZBvL7ppmw4zpVBQjk
7qS0JC/YjN7A8qybTRY3mHDvTr3unOOE36RPttItQRt45bDEZj11DPoHEb2x56Ep
Czz5Fz+MjaZZYpDlaBsAXOlLLlN7HL2GxeZN3ewlqiT37w4QOVZof0cXtg05vspf
VvfhewLnhLAYwKrGNq22MFqllKjMGxceV1DPBL3etoVrBMjiu4JPxHXJhOKt7z90
XE2hhWT5xn1B89LFK1swGO1cgJKIl6QAl9OJMS9FW1QWxjwAGnNQln9xJA3NH8ch
aO84H97oGwwbdDleYywVWS7urBk0hSTQaV49gjjkclGByNxzgJmvLzYudQAOi5VX
ny3VyPfz64y7LJYktBZYlds7WG4xt6jeRyP/SHjm5viTgyVaQt2aTq3eB6+5bjTY
VvxHR9FCWBVlkD/nBpZ95RcWcbJKueKMRl4qMJoERmpdALvWxK/VzNyYafkIzMda
exaTaokhy59IkBMiveaojsbUrt/ETV5pdwC2Q5Cou1IjuagFNDISYeI29+GEMkf2
4XM66fKN8dWmGK5omskRxd8QcKY6fXPMkZj63dxaGxGljMIj5KRDrda/4wW0nwdI
aOuEn4sUa0scZ6mEsNaOJTMhmTGyN7PHJbfqCYvop5C71EI8N4F9ji8+4OPhegtU
+v/VDNQ6Zx6pn5mozOopyg9ERbOSSeGd2eM5V2/sSHNrUb5p7/p/rdJvy7YuL7Dk
cZ6oLefnbzvohgKj0spgACVjN7oQJRp8p8OVyRYAu/NH+MXU3w+G7vQGEmvhkJQw
WQ6dAzDsXmKa6BPLgI8UtSgO14z+LAxrBdCLFgvKFTDqa0DXmCgKQ/G8xwFjAaZu
4daS486Ggwzwfs5sMBwF9S4q0cSVwK9sB+x7v9NVGT1f61BDhKz5rLAI0Xc3OTcz
s0V1AabunQyDQJs1ErNC6H5V/qikzeojKgpz0mNuBWhobiv3qvHctypb8E/5mvav
M8R1aGwg2FnLINtADlmZhncvu+dzy8EU7XOR0AmA1svfQk5rsxHFlqZ6+dQmPcEh
ndpMggYnkksJA4oZUx/t1RC3wuOCuHmIgY0/2I3L4b7yDWDb0N9iTNFCB8DlN2OO
aIyTTuw9SVz2/bEDfwwld1TbJRxeBfRSV/nFT8UVbgHPKicIbe21n88nyLeRzhfR
YiSkinfQ+yQEk6kMgsiiMcGG2U/Te8dhh2Qxv+nk+5OHdl3wFKGbc3gADMILC4CG
LnjjWAGcVlaJMsGu3jSItxnFAa0Gtn+eF+nv8fjMW4wjgi5WrLhT77jLOfvKsBSW
LAClv4s1ZAF04XcO4VK/fiq2mzAna7086FRcPlSG+mkUrMWu+xoT5hVeX4cK6vWS
yMSd/J6/7kn+5T2f43QUWD9HhrdgrcOzg82GlBZzRDLAuz7jTWWJ/PoeMzXZnhIA
WKA2EO/YCHJx3fxkPSOwAQkkhnJroOLbl/n1xpgsOGzWYpKuax+fgcLXmYDhtWjZ
xyYsjQN6BVbU5tYJ6PnythNAy1h4I0fWNz5lP95vGXIHO+Mmb9Ewfqig1ozK4Eyp
XpJ8KaPfidCEwiwc2LYLfroYHTPvKncD+eaDgAgR1DIT3SC9a0XrgUExyYKiVa+l
IYoo5lwN5/e8zWuBubSdwxyZIogJsk9uy3XGjekW3ZcA7mUrgCZCC+7q5WDl90Jc
0pEuatezgZUR7myVY8CDhzjGtDcFX6CCVIHH9JdjHuq93vfHNf8yECw0VvPEdoQF
12jSgPad2qGQRuH+QiEnGC+/uTn43DZCccLNrqaNiNzxjUbqgNucGUlBRn0Cf+05
ZdW/ejiEemLcH9VIqs1eMllPw8+W8Z/yOqTOMFBW0msiPAKEStSYogTJq8zSPqhj
TQiXrlJR5PgGSCbss+7zzXVwLpTZ0kvXUxWjDxv/3PTJJ6Be7pWqHWkszcEDxT+7
tTDqCOU4O2sIybPRiQAVrfaxC09sjSwiVEW0PKPDUxdsqkozQUaKYwsvh7C3vtoM
u9zY9gDb61RYuFdXB+ZnKrA3ECkENy5HtDoZelUU1Q99vKEHRiY7oQ/rmUAKX29R
VdGUXVkmbuzBtogASmAYe7sIJqmGCXaFlhtl6FS5XHlJIHCVM+B9Uh0/XOFgHsuG
JwdoKxJD/7Za+uYzWfex7/VURiOKZZobNJ+xr+7BAG6s8I+LvPip9zKFTWeVL5DK
I4bQq8+YO0WwD7XoqLfA4ngkj32SLkk5BiH4jnisK89FRAEsgrFI+zPyqizZTrK6
UQyhcJ+B22D8Fwop3UxC2RbfEL6rKfJdE3GFsNkc8zsFxZk/R8RPd3L6+J62aohB
aCa5m51c43mvvJmtRCmkXTpdEGIblgBTwmct1tONe+Mf+6zjcpl5NEOn34iLeBvt
D956J01j9096Mg/miWTvDtyPlirWL4SYkOeB7VSs3r0/+TFEZqbvYHsobx6WhNV2
sl0mGS/xQEhY+TaeT4sBZP7JNmvsi644tmkpQqVWVTwSwoiV3e4D6JZ6Z3TUnHGk
vdBPDjYOeAC8eL0UkkfUCqMVfxd54r4RfRSwovB5K34CHcSKPdElRFNDFZuE+NfI
wVecyZfI6VnXi0gKJzQw/9Dtyrlll1cc0UkplZMtjvl1S7auBdshR8SIJSdiP3O+
KOX1OBZAbzzNSBKpv4fV27VLz/kn7VG5zLCNpivHGyjZzLjjr0gvwsI08kJ/ZHJT
ddrAJuK/Z8RA8yCUZUXgk4xM1AgHD2tgpMNeigNkSZF6j5lHYxQWWq8q4QjzSW4c
FQLEy4QLUMJi6fFANKzxubkLqMVZw3orAHo3TXf8QHg7pdDacfmvMf6jvo4SLJwZ
UX8fprGFlF58s6eV6UQMGZcX4FUyFNPqX6b9Se1vw0TNMQI7L6ixY0ub40yeGIfB
FWj0/byPaqgNIcdt1Wt4To/jZSGc3w58f1vKJOWHy5p6FM5kRI68d6wOqjUN8a9b
pZJuOGSQvlNP5+vl78cn/VXQVnlZCFd9YxIKZZLFczBJWwOT6oGo8KPdPXMmHpqI
bIv8brsWBPt48NQMSoJbyvTa7tqz/qvS/4BYnY+t19zXycBA+j+244TqrGe9bZVl
NmPBn+Z+aOy2L66UHdKFPLZv/6GXzEDjov2Nq4BGaYIKCXegIvDtio3k2ZGMexOc
nKDyJ6kC6eV+v1nqmuI4AJT5UJEOo577C6WNGMyZUttr6+ZJi/rmjpIedIhdDS1o
baR1AUEH03fWyG2U/P8Lhts0GHkdg8IGwk2ZBCg7od/IsulCcTRorrdy1VVruMls
9O1T+NlaOv5+JCKFZcTn5/7pP9P4zveKMVan6p6NnmpJ8qHiUSuWjUBi5C569pKY
AyKZKDiO+26KUf39MOdheEtuGzyKjoNttfCwojpqjEumlehmMqivMkora01tO4qs
TVL6IjNzIOrrUtMrFkYGwoIw9ShYsQIJLKgf+CvNIAPp4z3tDy8c347ah5gdg14s
zxct8d5fv2BNiedv7d4zqt5XeDWaSD6j/EQobGpMseEiVi8aeKXFeRehCJVOrk5m
8GVjRKMFTs3Xg9TzhevKBkrLbt9QaA8h523IdxALHjdpnhyTvj0xemWQg7PIBg5S
S0Zb9dF73bKmHngz64zneJDyOMOnCujKWK2HQPpgJqowDdIUCNLMHO3VWbf6laVw
2RpPTrhNOuKbL6s9K0Z7LnkNUDtXPMacJJTZ0+znhWJQOQAoRNtIh68mRtX6AiaY
FJau2Lb3J8eAqY+ijZqzBFhIQiRndHJvk+Is8KAmbvtwmAsfGq12FhSuLNmST+V3
zHKDbLxZ1CwFlR3D/L0gYVNlepS74ObNggZ/eWAvGFMEtqTYsrmhoYkOt7UVr+nn
+TiYEZcd9gVm7WwkBvS7J9ImuXr3rlhahgs7S9A2pf5fPfLG4unw4dog6wplAcgN
v+z/CrIr2V50f8H+PV54Yr3laLZXvgmyFzslVU/TAGMbK6otZw+kVPjAhLpcu8Mq
y926rVhHIIzIyZzRhGWSuiEqYd6D93R/EfqdSPBCnUbcctY5x4My/Le+ptzgdgDt
/SLnac3KZwdKqftbYDgnl2Uya/T91QG6ZBUdty0qZIxllWdbfqEVnxNCKiHyecu/
b4LYBz48weSuDgxwfyF7lZDee/lfEvPUwhZGRxmVrRLpp6oO2zpDV5FM9G/7561l
a/c1AJwZ3IF5HNBWoeedaoNsCfcZCGP06A0XGkwnZ0KNqABHnFYrHEjByZl7iuVL
yO77X1i7u3vVmhaM/RInMpF1Yy0zWGEBoLrn2VE9SF7ixM33h8iQ5393Cud/9Qtn
ia+6LmXyfEcS4QDMnyQmbHTSXZ3zfaO/zXZE/6jvT3K+WeZiT3RMba4VUPlB3zCU
J6KZsJIXA8t88vhzN7P48Bnost+ZXgef908IminlXBC18Zr/+2MkYaNxRpoJqQ/V
YfTBEbkMNSGMpQozcWPBHl6FdReRWIIttfqDHUXu82w9rJJsMXMcdvP2GVoniHem
8cCFZqY0vt4vO2D6o7IICH6HN4JOuj7Ty4pA2c9dT5uvKmIW+Fng03jRL6UF4y8y
MMm4C0A9zAUx04IMyLUMIdCTgHUeB4c16UUYkx8fZn9SLjVUcW52rd+kqwlU/0Br
uHvRtOKK4Z/RibUED/9EujhaGIJFWRp2jazgTLR0Vz/bhBJpZLI6tI37GI+Dj3U7
HnqdvSjwtoKuTXp1AFtQmVNnaolK5O5IJRXKiThGPVf6KSp1AMfYeTdr98Jc6oXZ
ORHhvFbxfpdWW2VfyAFE4MWOJszU7kTupMHZUgciNwpJNn7hH5QVf/Kj+qZQGjhc
D9hRL+P7xusbeGRfWm1icpm8/kspaS97eUG19mvjKq88vcF+0Mlg8w4jWROBeOLE
QdCfnhBOXlLDf2JELvozBm8aMZPHjrkAt9bUor4vsvB8rRnVp6m6NOMBYx9s9fgd
wzvw/i/heBKnvtsyVfN184oXUL+la1SJc1aW3XlIGEpjptEkUZ2tDjFHdXMulC4h
PzTneqibbQYJMlOeaLG4WIqaGcpww9ozO/2XCiVlY7gHrI47vuZQhPE95oc1fxdu
iWeSgaya8TMvRelaH4+UccQj/57WPF8qGoxycElAFdkzTa+izVXSjy+mTwFUNdKb
d3QNy8jrxWd4ezTnZK4Q684Ny3w2ga4pcArHs4Ds/nXJqzXXZN6ddy0v5lmPhCv1
5xKTEViC4kysbOGhyalX3ZxEoTeo/8snjhMOys4xVjRXBKCWCcLbEY+f9yCOuwIM
gdlNpMqTJPqsjeX3DbPVubNxUGt05xqVuTBb0QEbZzdJGL6/ubUcgs5z0C9m86dl
9zY60gjbMsb24QYHNNIqNdT4ga2jpa/M6SvJDSktNNSduZrCuTaFHvLGxjufAnBW
qsf/AJSCR5xLWU3OK4fTNxvptb7JVZ2r7TbOSknG4cRxZUROidzgjQxDktax1/wP
P2SWodIFT0vAwaXDv/2nJOEXC+3vBnLgR3uQxH8W+LN0sHlhxHYX4tdBcQ+DZQVD
Y6PBNAUrprGdrCq53WaXStnDWcoOsJ+PShvjkG3lCNy5vZaOPzWaVbqrZ5zTxis0
hFBofOOKW6/UAoDzfVCzDUVy6r46mq4+xqdZOLtfuz56QLmoEe8C81iMQ70kJW2a
LCTLgoh475pVBHUq6DnyxVhqeUxZ/VVzgcc9Ks2Q+2yif+9//hCC972FUMjlMCsN
2fP9WchXYNKNyK5AXJZ3g+AxBKI2VcqKA8MQx/xL8Qjq0cpIqhx4XhzOR2I4aS7l
WU7BtPnE0gGjkzIc3+2HOY7vNS8QAKcDzkY64aQjnZE7HdzNtMDolI6dy4Pywnro
CjBlpimnf4WJmEONcKDaprS24jmWfxjO3oDTYHPdD1y/OtNh+/PMxGRZ7iVDpOQ0
WxhbDujG/u8Y1NuDt5IPVsg/gRspphC8wlT9ibh+CxxbivtmBupB7Sx/sXPAPdze
Aki3lRStDgU/yO53ewa+0Ua7VSbqFNNis8W2lQdAFhoptNuNI7ZCrtlYY8qgcmsx
fgq+bN2FrUvLvJPhuOxNUZCzoek89xS3vxqIUuoLy0LwIRitnREv6ZUrdMeLXEcN
iNzYR0SAFOt9NzTIrMN2gKf2JtK3RrbzzTgda9+L3Eg6OhkyITTp8zjq7+unF6Og
a6FfY3C+8tYcF9g4bau1IIJnMWWwSb6rbuUTZnAG4jnUKJ2XWklhAYYCWoEHwjye
8CcoxJGIYo5c5K2NlMoGiAC+luMfzFNjj/XsQpVO5xhwU8Xr9nMtLJ9+IX3/bLe1
NKI141aW3x2CnjnSwnetaeCmxlfOP/UqCmNf8VzbNui0gZtJziZhBxNdV3yxNHwI
/hwUV/TRDlZ7pVk75zHFwibg6JNiPrK5pwt9wNJ+drdc56QYeKS+jdS8ndQ1FhmX
Qvg0p1XZog21jkHONM10F0+tdBSkyz71m6sYZO78GL16PzIUPS2rYsP3FihtxkJb
0ieoLT7mZxnaocLp/MARyLWDde6DvsNqYdlXSekzSkTtlp8PIwGeRkPjn/lbxr+Y
PxVBbszH77c/bfhbpp6zdtJPytidk7yl36jOQQRgjz0ckHaYP0Z35qYKhZemPLLS
WRTMHTw1SaIYIkzIqrRwWgJqI6ThQ0j5k/UIslmP71fNtf94QjrvnKLOzQOFJy5y
0ic3+VdaLykEULfbKaLxuQ9XUTtk+PEDVljTBv05VDJtpjkDBzUsTEy0mkU8wB0A
eqXHuSJ6d+TACZ5AZV/mYC9omiWryZEHeV0ua++NKWiqq8ZOGyS1faNe3ZwtpsEH
JudYq3WD35SKlNJtpImPvslwqyWbetBQoR1lIslRRzz3n6ZhbX+XbjO+OUy6osgf
psyihQ1z4iMdL48iPJ8V8x4EBPruIdZirDnilLxeCR6WPqc8kamVSK9sTUwMi9KW
KHdEa0ZnBRpsCg35i43Mr7IXFBu4mrME5jqX0vNG+GQz9jpn9wum5nxUWLTGFzR3
B2j/m0TMd4yCw39j+N5uQpTW0BKMbVSye+dNXP5U2YuMBvI8egk01TYehVjWjMVf
rjCSsqV0Qa36U2SWPKKUm8HNmCgur/giUc1aHhO4u4s6nzLRg4p44ew2x96P3Nmj
BjeJKW6LRY6EJNYQIDQJT0NJjQfr3b57AfQcTQVCvcV0m74fQRAs9tpDMhpxu/wj
nMwgxPo6nIQfq0lJHuBFZVc+50f9ndWQ4in9g2gbmWmYX9wULXWG5A1jjVTz1z0A
wQ8GlmLbT/nR076zK9boqeSJwo4P6Igq+FpybopD+fMGw/GLJ1nLlaj+xVzsB6Pn
eALxId4nG8WaDDVb+/6tjAL1i96aHJiuIQ/i2kQlSu+OkPpucwQ3T4QKZnu2Zj2o
uS+FEoZx/zwe4VJUfusAZ68A+uOqFUOCNQSI7FaVwn9Yh2/0l0hAfN43+X/MJ7Cf
wpA122RKi3xMZsmH0X+mPeSJrCg1+v7F6QfmX1/tmBVqNRXojbe0t5lqIEMIQfG5
bhJzSj4wpEvutWDbPxZzmWlDW7SLiTU5RjVGelcP5dnTGYHhw6FZfw65xo9ISLeH
042WNbZNQXPDz2v1mROHIU4ICpdFus/4XrkCf8QwQdsHWd+k3jMD1ifxirkFg4c4
meRfForYp2fXvOFrWoEgBweqf/f2cJG1BCcFsMfBFHMD+5ksGQZvRHD/E8Scpq8R
AFf0W+s0tWoljhwmNyM3Q229DpmNEz6dl8ga6rs6w0F+yyVfsQq5SF5SFHIs4CpX
zX0h7ljEX8eaAB1zP42VNgDZLybZptRPyYyCFBT8WMBcgT0LiyFCUnZlts/vPx27
rxWX3NvOyAZXQmzSbBNL7KYb4pJQXnn9cHhJZ16dJkHxT76yGZX42bIztJWFWpgx
FqEgk2ajiUoDaw91XNLsTZS7ugEzIeSnPBaHZzGWvAmjVpj5+2Hg5QmaFp0cb4oq
o4oT62oZya+c8Cag0lToiBfqHAqA9j3Q++AbBVsbLaNrV1F4muD+KtUGCyBehK4n
eWPnXp9ZwxbkXGX5+ly6VEjOL0yeb47CUXxK604Pvnt3EI3rRIH3yPNxLGuSi3kM
1WPMa9AnaLXHzosD/M1cUFrA21HsQ5VWvnTVN4DmENX1RFNN0oePdlZzlyjw4Ilo
uNPDTGrTISuE0JF+yWdKmwqX7wcVMxKsMmFo4xq/QLZ1FRwvMt5JTBLafPyjfu8n
m8qO6xacLcqXT2GZaLejXkrbhbk9klB9xvwbXGhDHvRHjHPOUvDLvgrqePwq+Jj4
wpTC4Zzks60YHVuhxXy9+OMQ6kp4WTCMoEA1HIGxhaiX5Jw6ZJN04EgWaY8/l2OS
HO2UkpnDWRnJDGEq+KebbMgVkCjxUxB9phWnCgTxLa5Fzlr10YoWi8+8K+HNrgBG
Nb3erw9o2KOLx7hl6rTVHw3o4os/yT3+m7brWR3Zon0X9578z0cUI+oPOaDnRNY3
oUYnr1MfyGQ6IoIdp9MxB/DDRAVvr7kN1nMz7QDUujf9K2eaYrG34embJGwXtC3m
6MQoCNH/E06hziNFJ8Umxo4/FjLzc2uh2vaRSnlBesbxttRz25cMW2XEowjIh9u2
yrWqqztGbLoNCxV5zkOknsKbYAyd3yaYzeBJ/WbkABYDD6spSCgd062x4t6razhp
FUAxzhpO0HvVUfG9iOmCTGns25UrP7rpbBCsr0Dc7TfeJ+XlDxV1GS1jw17Lns8R
scoM6kjCiEbmWwrvvaTTep9DXJo+YUX32E4M9xQPPgiZV0WZyPglIUzS6oflNQxA
EsXdug2CgxDj7Fk+DOiOxrebIyAGYsbagU/vM2jLFJLRVrKt44Q+YG+RrBI1XAII
H8Qseq0w5OpsT7/+vF7UBI3u4I5HaqQzYgRD+Jnvdkn2zbFMGYk+RL4iQBkYlbXi
mmFoUnBpGbRrzVNnYSWJpOQmapalBoPYbpxAQr1WpBh5VsENoYAmViVdkKhAuhPP
SSOxgESJMb8B0iNtdBkr1jvF+ogXZjl7Y2kZKM7fveIloQMViJlf1mAVOa7SkI8m
+0lwtV6lpSAZ+J+1vDcIIqRua/yPndYGqf1SDS/VtIRzSTRD9yiiQB+k9ZKiJkNh
93DosV2VmThF1UgEE932guxiaec2MzluA2AjyTY8K0LuXD0yjS00s3KcKDRCTzAV
+JkAhwXtLFeBK2nHGLFtvlYxfM15SKow7LFeyS7y75UHY+Sy2+RvZsqlz+b7YT/2
sDPmdQASdpFaSgLo/enuxGH4eAp66dN6bXfW/zoIjG3P4HVD2vRLBKjWjF67XKIh
Fq4N2i1sFX/j0O+kqLsG2B0UXIcyfGhWkE9GPVLdQHtPTfDFmzYIkqzsVZFqQdxm
R7hgI7c0W3WQ0toneXEVrO+18yPjxUfnMEEbdQd85nZOjB307ldKxu3FAHMHc0tR
f550eb6SYABXZX+AfNZ3c2SSWACnBMY1MEtO5yOJYD7CmO/CYxoD/Ud7SwAq80PL
wZwKTYMsMVKV08sOKl5edEPmKKXwpkH/FJnAQmf1e8/iymVpy+p6czdQBYZZX77t
/7SnVihV1rF9Yfh6TtTIohjGnGp1WVPsJqD4OsAKFiYQrVwR6ScThzlm7ja3hyWz
2dWJkr2jZam5cUK2yQHWc8Gx1Gy5y1vbni4qW6SbEvJoFWAzYOLCDBvNbyoJwn9l
QAV0GlP91S2dOFmta8vFp6uYvZDP4B7DCX6ul24nfhn344q/aEAlUuXlckBh4mYn
P+4Ef3TyXVi0F9BRw46pizGPvEK2H6D9GBHwVlhUigony0rX9a48TXwed0316Qn6
i7contmoddDcmHwAIg8tisseX1KJ5i3mtn2zWwNCRF0sbHgmyacOcbe7dvCMpePX
T2lS0DusxZ8GH/yMecFbZqrwCypef2UoeDxWzWtjTz0fGot4rlZNWFi6I13rno9w
MckF67f1JpN1dHXZm72K4Akz6OwfyzoXPrFi/LUWkmqLOQRU/g5T4l0uaRv4euz1
kUyTcGEtFojQgB1kTlITqBY1kBXUstZ2zO0dAAtlNeRnYIX7gBJM2W4tF+QgAJph
6BnX6BPOZoeiBDL76V2bU+iuX2+s8tWfhtJyO147oa23W5XzRmE3PE6DVkGGCvWD
qvWxmuiXS+9WxgBo4nHjX9QguHDbFpF/rXbxZS+OP85d1b0A+tqSVDSLRI4o9geI
QFTib3QhXeZXrEyqh7p6bb+5i2ZiTuDF+9D8AiV8xzE3wcVScuDMexgkTNUTAWxZ
UaNyEquR6npbPDqyBfRv7R3ym08VAh3MHsAxrzowb3vN+4sll+5XSg8fvJVkL2Ii
Xs1ha2nOgLl6tpsejTX7/TpCcEYA9kvsNdkwxjCG050sPM/TYVNP1Y/zehSmeaFP
T4m7i4DCp+jaYvFN/Tqq77D5rx5hSvBEcnqUoJNJ8HhpzBXLrkycreiihPpozGvb
FMLYwqzYIzSV6DhPXPaKJ+u3GWYubKYG37qffYkT+QAjy+FU6xZCLVHaPboUqlbG
+KkYxP7tbFBE3pZrB0KBbmNtUYlT+NFtv5erJQ8NUB+bqvPxXa8cGX2l0sTb3c/8
I0Fp0pZY9zj13Ops5dfyS/gb8flSJhBIiy1Nf5UK1ckIZFshImZY/fUl+a+mOny+
BCSFjmXxHlkCm+xPtSG19VLwyCU6F/Z/rQurt7fyrsdHiQ+2ri+/DztMcGluzrt8
MD6r88DaL8mTir+8v3KD5tIsjyC9n/36AbBz3dXg7kyOS80StM70oIItuU3OPhCI
0V7MnMrLuIcU2wCeTPSKI+qE8FoTJJLtBed/mBTsAHxvFce0Z3ZN4x+depAEGJpG
vNA6aAROOSPw0RaZmoBLmkiAMd/t//R64+BNohVVt0P8C0IUorUTgt5Vo5rdSz7W
FTMlKe/EJZ1s9pkfgqv2suMJpnbdB+1CmjW6fHwhpfztAFO8F9YoMZcGRB1A8aV1
St3057vwKefaD7NP61CdVD8Of22xKXl3lESiav2bAfFFiEvVF1F1ZeCPOoEY1oTq
Qs/N+CdYVX6kecSYxWkQA/ZDCnWbDGHBk7uwbhYnTgitge646eth/3SheZCKIfhb
67CXJjjeOMIsNYxCZ+5h4YYtOQskvcQk/x7E82H3PA0mznJbrLW9sjAUyPCG409l
BkvbQVWGyRG6VSjvT5h5snPwBQZNTk+iE2McvyVEcTLeGpkp5EOmw1LvbwilP9Do
1jdS3+STXZXN0QRy8B+tBe1JmSzEvZobiGiAN3fhKIQjtzd3WZyoYX5QHhJN8Hzz
VSGL/Mr2XfL6dtw7BT4dCYspdQk5hZw2gTobZCFXt0j7jV3/gVqDLn5IdIrHZxUk
gew/yU3sDEPvIeE37ROUA4uEewLATv2NM2F2NgrQUwWTsmuBUoxu6EOuvHHWfWub
ra5ouBsndfNI4u94zEob7mZQNa2FZY6yfWP9lW0NnUYfOpJ1usLx6dqND4fg45Up
/c7J3ulYqrnKf83NkueGDk5snUsO6/TJNo9kJwMQBo8bxPAANmTfNzrj0iPHDCEa
XUJQ3EzvOleKhUCwvo1RFjRxP+c4lgl0RHXJCMyLJb1pZrMnFINImMyxEb9sh51e
ViUHCZT3rHY0CtBkvA533Kw4pO575i0U6xCo91KL62ipBZ6XhCIGab0+KURFmtIR
13QGN3GWDtWhHj+ymRl+ZHIZ0OijxlYg5rPIbHaSB56bPlsrt4A1avR5JbcdRZrK
hVp69D5AFx3SEU7S0uutExCG+7dyRXMTKCxvtcHXpdrrg4swa0FNLB3LSAOgVnUR
WpiXbSU32TBERPeHCb7K5Ly9FR3T7LMPOEtRqBVG445/bJsF3kYrg3uTm6CEU2bz
l5FQsKcNOPYa6Y7zUJAsnvqLnWJCH7Y2PAD2430CVLNEzsVIaHoC1ldGZLRXIyjN
MHjLPj6WQ0qbL1MClzjNs4kqB6N8rbBLxw+sjZIMdUlg/G+PpIKRBe/CVn+7Wu24
3pFv+p9Q3BP5R8ceswkNpvjUBkYpwbASwswWN0nVrnXUO7SHNjXCLIY3q3dk0MTb
7+ThiL/kU9U26fuaGI84Fc+jWAnZpKMfVLyMLJccasS37+aFrBFOISrqsJHA0VFV
mpMAuCu5WFTiiunOEseXFyx2VVBrT7sKep0djZtGGFVv7xLtzDXslt5+IyFmnMO3
w1Fv6+EpPag1BiktiFWnvDazROdVqHhHVwCMcWYZIkarvIoDTTRih+29t1DSJQ/I
f7pKQ5c+0DUuU0JIZKThvchlxMo8B7qONgte9COvSmsyFYskrKseN7Eul9aBH3FW
XeYa6nw0JaT6XXqNKl+9YfvARKrSJy8JfBSYss84e/F2UTt3IymqYdmN0JpDxYTS
ATVjEGyxQ9mBdtdJe2NFdR4FG+qRsyETNhL/6JnAkOt41w5BzLfCueNnGjM+dB6A
ohYybKvXCU7ddSMasUng4AG+Hu0qeseLoPcBKb7+0jaMgRtOOfrydae/pZRCEInK
E6txytbfRNRqKgWmBi2i/lg5k2R/ZHJxecJkJIsGzuwhNXkuL3x/e9aMNlQs44c9
ryhEHZoRqxAG+iooMJpxkXXiJLi/8gTT5Z+cjPa3fHVdcqK9J99U7VQrqSb8lPMF
VMC9QqVggZWIc5rLgSWSE9ObJKHNMsGVMnYj5e76fBOirlwCFLCpcosLQHzsRmkh
Ch4FbvoVjkoxlAYEn3eCfcOTPcryak9Wl/Sqvcl2gg9Wj4DBo8UMZ5Y4zn7DcUb6
4sX3w+sVClhaxCjUols0EWOsDd4UeyRE80ZXASDuFUG2nWr8bl6L0qSqTq7Nr7It
D19NCLNQKSSzVqaUKDjeiyQBTPs3H8pzVqgZbs3dpFlZxu7R6nASv8uPZvXx7xO4
SKwJh5azO/ltdFkryX060vb5CTcWsUVh4rn91OYTBTUHHSCZ7+ujdLW/5jYKxfaw
RML+348S10i59njomut1eVWeoP8ShRqWifwLBT4EJ6OavbqvgLWr99nJh8esTHq0
C+6VS1Kq4S2roVYE+vVSu7i4Ug1wMW07s3bwgLbF8zE1w3jGvOien+SMkSi624om
pmhqJRw2z8QxrasVtkQ3F1fjKPuGQ2d8eGEQidXOfrfs5JCMKb7Qeetf2orhpDNM
vZWpDLrIrd7TEcN7Ob6Jpx6Z6ZQEf1oo/L10SUutUVY1PnbcIjYglpAopc4OG9w2
T+14TxYcaw8ULS9aicGKSUjjOo+jz+bsqxmUEk8mi5hNknyH3ZeXxqmiVjlkL4KP
o0NFxZvowNjz6I9yBnk/2YiP4caadRmqnepP57rtje86BGTViljIJEKWEtaVpIYE
nEsxiRjGwwFK8NeIPsTCJHt+OTrrlieNZmoNGr4WrmKtXAuQftDX6obfpXSgK1ao
CyUwFCaHKLw6NJU2vHxJZoPHb/5TtGtST9Lx6UsLqyu4u9avdRTQK6nH7fd2QJMR
4bJWF5O7Ye9YXW1yQKWElKe1HLCn2lZ44Vhrtvz4T3G2pukeIc6cHP0V1Sxwe16n
iQnMsGDugM4jBfwOzo5YOWLPwbDcSolfla4zV/CCuGeRNVKaHKc6OWtIliuGpA8m
AZjIEnkvCNQW2SYl8ghPW/d7fUPWyDO1KjS/B0UgJIR9LGXqD2Eb3UrFaoVse05w
HrL4Vm519r04RCDgpKThXFza3Q+TAvE9wSSD11Kn8nsbNwHQXMlXLSNw5V2/uwVp
S05ym5cYJtGRh/F7QrizXIiwsFKUIypEJkNYa09r1BqLO9bwKrjYhIYqJyI8BOKy
YVYaIIvk5a8ShfR5IEaIMcjpDBbTWoewZ72enWf3IiNmjoLjooh/RGyF+jW+105Y
s/9vR/BGeJukc3TXCxu7ZEUUUQ0DYs+r49M/YCFL6Or/Bw4Jea6xkqhXmdWvtOQu
40UaYfA6bpe91hlbXhTZd0vxjYNiycocgpeMsTnW7aXODfpzCRiwa/3/viVyMqA8
WhhmfR0i7AV4I/v8Ughnr0BRyyC4vuF4z8Sw+S0poyuMadJN2Oubq90pT0tKG+Tz
2aYWkB20UuCAamUc4Zeg4zuUDO1QxaWjJ5M1MB4aIdXoiHxR39N3hDy1pKb7s8sy
WdF0psiJ11g6NWC/kEQEawyd6LbX4Dl2xhYhvrNuikWwqKafAAe+4yKIZE6hjxpG
w76Frbj3JgPSx+m91EECM8bQU1/GmTd0oVz/6AXwHPHOQ6EUTM3j4GjtJNinTeUg
b+7n9nyb5++NoqTAUMX1mc3R0k/OF+zGnO1zGirDw3WM3ztBFEqwn8ot9e4leA6R
2W1y4l2GFy5Y4BHxe9boNvNha1XHwuoBwXQIq8P88r8H6KzFP0tyZLwzu9joq+7N
z5ecPvCJKBMcTXDvfnPUoEWPyKZif+rDeGv9tC0bahJ9GvH+L7UGueag5YnfRHPC
ScBJO4dXlrLbzuAvami/lgwV+D0jdKk7SyQguM6QLrqNuSQsU2R2q122kAtROCzg
soxlziqeY5gfGKZhAe+Zf5Nm1ZQjA4/UjhDlCHwsu0yD+l4Mj6Go3vOBCnUPZE5a
FlNRNNOMa6anAlxxdJ08xbcZuysgkNr6v0HuzAc7i7WRs7mmUfdIbP5nvvS68Tqa
vEmpNysAkP5iSqRjWCtcwPFN78Fr9EVlIU1dZakc+DCbxa6n0fyLkjBzmI+2W8tD
5kx+jlfRm/iXNxf+IS/aGlIXHKip/bURQagVABSGqrClKCUxYBCkagCM2LOQ8o0o
nQae9FSEvD6kiQUGMP9i76GS2IC6RpI/c5ulTnnyzVm9JHB+/tdYoWxUKz+ZnoY3
rQeP6asZIKgCum4RGzq2qzRhGJKeSiRiZJkrwouNxxLB7HLAJm8XGYpdtOdrmttI
Cg/Dgf6b3o8YgYLCsG/ZPjtmtnKTbDbEorjz66R0Mm5wbIYSuKuw7EOIctQ1AiS7
6UcLGs2dpckNdX/naNMCn7eaLsJ08hhlWmoBqzK1RprLTSCqU+KmaX/c+LwuUfV1
qD0Z8CGTsRAFCeNXeYI7eLgMY9ajPzKoPjfaBu5NeZvvsfZgdLSuC9uFH1qJsn83
Zrp/1nCCCcbrrI1hzi5AhqobZc2/f+424jAUu/Xjvxyl3gueTNyMCazj4Dkg4bkV
aCDnPpbuH937WObxUKlmH4az1nguOmr8GpFG4gq5pJu03SszOkBPF4W/RiW91/R3
K0B8baros6C1ARZzZwVlShJIVVTrdKnqa88Fw5lzUA6SCP1Wpa0504h0TS3p4Vfm
OWmkhdwvv+Rt5vNnucBH1xN+96KS03ut40WzYWRyL+weeSTGHL3hsyEF4AIvJiJU
AR1YzvETNtvmPnUbrcgxajZ3R/nQjmbeLf8DlzxwzeiF0KsIa/cKNgECnr9hWnJv
r6+aCHa1RHD1Wu1/PZaDXqOzssRSIr21KpPvrtygLdXPoCJgsc6yK0htPyvCAj7X
tLS7d6VrMMk3eFVuLJq2G0Lf5saIgF4pUCR0rixILyhPkJqM2loM+6XIO51V3Obl
fLaNqJaDzQbHM0bqEHQBm/AQqntQRnEgY1pKWe0BZTi/QISKQFmhyzssZumd4j+8
CzmSn6GYAKFD88NUI9tDGoDWJAiywVi4bXoAflH424Te2RC+unbllQB2S/UP3sHB
vBdKtJhzdbSZ1LYKq4UXhBxKtGzkpnhofzG+KnJ1ls/e4nh3bF3U3uWG2JK2AUj+
qsXESW8YgHD3iRzyEr//6pdRqyoDSKJ4Hv0/rVj19V0/HLLPQaIQu2OjKyzg5GZn
doQT6w+CirLt0VQmI9bI8IJMFiwW95zmd3B5nsoMcL4btnGMHp+gCMpv2NDZSPrh
lburiS3PaHJheJk+1qwnUfFAKTbu+VUhk8H5ou4i3cM10DSq5xTLi5hYhLUUVl1/
su8XWLmmLMd+dfHBVqs0n9LeHU0qcXXaL685TuH7Aun9jH37rz0m2ZWuAMERjs5/
bXsH4jsi6qxs3/dbEVlxHMuDA/1BzjPlt7EFViH3lF0QEvWh2OegP+jOidlXsmwD
El3n9WS9bdU7TbZkqgXLkV9M4DckkcsU4fBvhgKm0+hOvWUarOtqiDzFFdH9riwW
xtNmk82cG2urfjB6XonMxpRobJjgBraqaWUT5sOmhLrd2V+vxjj9/YEm7J5hLwk+
hLjxmZ3bIXJpi5aSOURtObbF5VO1l8mAuXxY64XKH8zkHxmhBYzfcmMCkXHZw5Ln
3m3c8WgnrwOgo31Hq5LyjprdEUYUZELnhVu++EaRdWW4a2FupEsehz/guC2Ic8Tt
C5dNSATkPReZwaU8w3+mcH1ig/mOPsysarvgEzFImJvFvpQfP7z+rZCAsevxdq/a
ORv+CHCaM1l64ub81ubABpVMZJAP19RXNM1n5fJqfgZR0ojqnJbr4rAFlWI3SkwW
HxOQQmcwNpwhx9CNXL0sR2gnn2ZrfgQoMnRL6wF1ZJIjBDyGsKq/I/xP+K1C15qp
NWg5UVqAGktpfla+cXbfIxbu+qim0xgHOelGDrgnoLlZmTWSx+c43vvxwVthypKg
sazOHlOLQ43QgIInnWvmS/PrBnieErCEMRzGmOflgSUao8uFr+qSP9nA8mRhUD40
KUB+LWxHWjYtN0+RiNixmZgZ1usCPMwpTr83mf+NKkT4Wcixv9VrrBOeb6Abzkcs
oq6G6+URvcWjTmoGCroek2gs1KVTwQ0CETgFMTaCkDDf3kZlaMHXx1WDs8sNLBif
KaHEVfvQvpZrJn+rhdIvWESDDSeo1CAIgdt03Q5p776s+hnzAb2r1+Re3SFLe9lG
tBja8ys1+L4iOsKPAnQzpA==
//pragma protect end_data_block
//pragma protect digest_block
ZmNnPvKPxTc2FrBy+gQYRcLrpZk=
//pragma protect end_digest_block
//pragma protect end_protected

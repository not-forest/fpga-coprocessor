// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
oyEr+IEm7VqJEITbFI1uThBn0GpxsrZjpFnv6ZMWRfAOO9eyZk2M+/kJ4vfbAtzd
d+c5fkGvftZI8g14IonDh0RQQjcXhdIixOZeQqYZe2nYuMJjIXSCjnr0NW4YSmcR
O2ZfHG5YHBIIinVUP/5z2zjg2WfMycXCrZGZr6nkD7I=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 11616 )
`pragma protect data_block
9KRGiNHYcOPmvac2R3fLnBEHT0EUZLLCLs2ie3IJPgWuWYr7dwKwkFkDKKRe5Q/J
aF4KtuNd6MjPOjedHsCYwlM5M9NHDeFMjWv60sq1dMp7pk21Q5soAzibwnHZDUtd
GF5dqze0EXlvV2YcVD9M4PigfvdsIVp4hljKv2kUcNE6kK8hHcQeDnViMV9ZUq8r
4nSgtY3orcxaMQwPu1x3XWaYACQBPgrW07SJKpeDz/7QAxp6Klc+WBwDJRVHIJwf
Ttf9yNXEvs7UzQY2NUypupcg+kLt1mrMz5PHKSfckcl4yoBJzW7c/m2G4NFiboQp
G5ZIqrjBeJD4ktPAparGEYrvMeJM4MCb3/neCIkDViAh2w6d4C56RXanXdfJ/4wn
W4tTt8Dqkxr1/nALk2DIyHkmDcXsYNnR6Bnvx7sYiTYoNeu5O/oktUeJ0if6A4fQ
lTjMqagbwjq7iP9IbWyya0zmwtp6rbxY0fx6Bhui6BOQ2pFy+Ll2/OgRkpik+iOe
JSAo4ZY3F2rHgL2Viy6CXNrdngxsZhUyvJjE+POk4c6CSZvHsRWjh6tk5hogfHWl
3bB0egTqy/mw0jzQwcGckL32d4W+pgiQ7HMD0wMHDnZUvXYp+H0hihCefmPk08AH
G7IOiuJSsUJtG0GArRVP+Zw7B2M3BSKv4pmfllRaRpvjNN2AOUk3gT1U/dhsbSS2
rzEgWdRJfKOS/JbzijVXrZJejHg37I0OyafhMZ9Ne85CVILb4BXVwHUfCXT8Uyhg
w2y7GUuXn7m8jmbE0/Wn03dMUQ0bbomkGh4njBE4+ROQ7BXs+ecf2EzJRIenV94p
PYKunjAkQXiSqFbBDB1BySRtdg5avpsntskRIUZWwu2zQ5tcTEdEAuEdUVtCS0LZ
ORB78rULD9W3/eiImiludzQqatndDPC+/MB2uaUaadihg5hUTroGEV/szoUx+QEp
piDQk2q58SqBxn8LERhIhGJSS2gVWmZeAIpOqm5SspFQXeyJby43sDkBQyEgJj8T
q42ePPFWa7Ux3iGxOHi4NLUONGLt0c1B2N1f99vi19Y+PLuWv0OlT9Qe/qikNVdg
secay8USiHgahn9EK34Yu0KdMoLTvIdu3Sbb4tKXw9Eyxp3a1z7r1GwL2iKaRmqY
vwb9OuORUXBVGZJsD5M8SVLfQZQZku+FLMRKMuS6hZGiomiK6lNXS4B/ehyoZMqv
cxZgx6gloP8w+nGvSLyab6kQ53PwZT7SSW+daMzKtVy2i2vOuxrs6kw9Oyf3E1aP
dzpjHr864+8dWQPDttlBSSQtB0RCNFDM6Tx/N3sg3JhYwgMv3AJgEU+bh9xY4DNR
Ri63TOSBPM42EDbnXETvHXyfffxPVhVDCHnoD/yHx3+mNMPl+Wg3rarAcJnfA/Tk
+4LuVer0Y+PJjUqys5GxPZ1cCU/ypLIRKhWTa1h2iN49lZ+v+kmSClhWoT1Hr0f+
mayqgfb381h1iDxjss9DYKIjqrm27r2NQj5cLVytgelAu5Y+2mm4V7mjpGxVvLgf
eya77lCOYyWbntpxLdenxNBWFjk0oqg3uja8L4X/P08MxrZU26eGadR8MPnuIzS2
avA7+gYFLuIKM17OTNmz83Swie04qYww6MaOA54qDbImrf3WPtMd2gChZqI+UaPs
AnDkhpIgSW7TRyAZ8VYE3AZfWCT1M8JvlyvQ1lTfE4+ZnbgaezRADa2+UOZLRIzz
p9xPOA3I/ybGVAH6mc+Hyg3RpwriYokZZzb9rTHGs4IrWhhopsbD8jh21pKk+LJm
DM8eHPkVs/hpbYRl6nVRJJjlD5Cpi4EIIs4qpZOp3y8t194vJQVTlANw82Td8yQs
G4fI7O0pEx7g/VbWPMcvVyso5iLBSymQM56DBXsf/tKJiaUabvRJb5WVAfdwGxEO
JNystiaEb6eJXmDs9TRNuZWxd2Qzlg+GGBukzC6z3Og/rRMisCGmjMy+3jOwUeJ4
QfuSrBvHl7v7YMOr9u83DLyXaAhBlPjVBEpOx5429iUsyJL6y4FGb/o/3G4Te+DP
6rqvNLrJLBDUv3OA+zL4Vvnrk/6Wpz7af35GNpl2Pud9FeiMowiKtU/h084aJ8sf
nryjUgB6Ulh7EP0NImLNSzp90ScvDBZOghU6nG/ICOeWslP2cbBynuAInbwZZJLU
vyjnA3PlNXVHV/V8lqKNvUzE+f/xymKlkCwk0CLBpKXvBSCdcjtfxAVAf0p8se+t
mhbsJSg99/D4QvzYTpoC99B24sv3Zp0eNCdlsSgp0aN4fKCUdXu4Rhh77zMV5byB
pcfSAiLEOp21VDrP+KT91aawjDVHRdU0W1rqExfLlyGgY5YTsMpkwx9Y817My3Zi
RSVyR8cl7cR+zSNo61fZ3AT+/1J5ydkPQ3+sZk+Aelx6fm+4Smpf1F6YlhvULXOp
qUsfTyUbu85NmXbzA7HnFFfADOhlZ97uky1Q1SjsagFbYgQSWCh2xQ/DiR0IJBJP
HldWpDj31XWF1q3XIupVwT2AKT7po57a9LGoBpBNloE6f991hoc+D0BMj7qGlz9I
muBfrfLPrU48r2/k3deE3LHCTqp8Y8iokqjvEKIHy8q+Yy++iJh1JX6FEaReGI5V
oSiQn1i8hg6aMsKGy6+NBkXCURurOcBK+hUgyXvIyhUUbUBtn4vifBUocJTg2Uqw
JNHAAvQ7nJxs0h/qCECbQxc15g6E4TGOUpkHKe0fMNEDLGVPBYc0JdnGxTbBireq
hlLJk+qwfXsunpa4mRbnMsmMiwn336r7nNtyHgtphP9A+a52Es8MnAUi3sL6XCBb
nlrJvuYFhM4e8axTEho1gbyFkzKEX2OYikeJFkZ1WQKvb84zCSxIpt/1EDWGrl+R
ayhXUWmyfQeuoV6N1dbaKVygT7RQG0isp4g1hrkcNKta2ulsDKJTKsOBht3q9p10
kUWzYx0r5W0hC5yxqELJqaxh2OZDd3Erq7SiXgcwHV4QW90H7XascOPk91n7i95Z
mZAKo2CsuQoVPAUDNChkHLyNtXDL90aN58qOpSVmOdHOfS88s/MCP8Qve4y7ufgf
sYqH9+HaYMTJ+8CBXbphi3/0u9/cOiziC8d8HeOdinEC6hDlRpyfK8MA5Mpii67y
MPDi2elGgOW9d5VRUR/8LB9oO11bLvC/EsmlCWgwAXA0F7XgQKv4N6nHMTDNMp8s
iPV18GjcTkmOP+QaP8G9Kgg72zJuqYv+iqZTSGP66FbnK7Dhs/mmDofLRF6CqfF6
XL8FnBlX9rnJD5ChfHuBbpiAIihC3Bewwu784NJOnDtGpB2JHlUlJluIE5HrLiRl
hCKtaTvR92LfS0XlO9TQtcXsiqHnn4mR56KLnvtbQ8M080qvDNoZ6s72ilhgzLyK
9eyJT7fuqya6phwjjJDOJfThz29xHCeEP41smUy1jzJrT9GdpbE4a2jCZn0t8eeN
9cNSpkeso7naVQTfgrKpnvuFo5IZ9hbajWIBAUZgkpwjcQO3inHwcLbxT5RHEn4p
WVWPuno+9YPrws4r4WUlRVGLFN3z3le6ux8m8t0/D1lfoQWW1Tx5ppWbXgUT2Opk
uMYqc5oTkEMz9GsYvvpQdzc0BvdFBhi9wsIdunx0wsnO/FIUnFt5itKITlE+DMBK
mMJSAztXJe4djXbe6DcCGZApbBCGkPEv6OLaRy9pxj7Wjs+yzVzlRgZzvNGl84yA
Q2QvwYRGwDqHe2egCZiDgfIBcrSQHWA+fTJzxqrtp1qd2JjIiK3x1L4Dq0uNE4xe
3SPWnG7vi51vYp2QPkDsBnb1vRUBavh4ISrkaaJpPcgO3IPCg2/SaMRGEjrgbZ0o
BTQLMhVvcISLRHu3oSlFJfa5IU8vUhyQseooVshfMZ3mFBH98Ga5CyUg1Yv/COzt
syxzEhVLUg+a3eT9DcAjReIk8/92SyF5heW5EVAcsYhX7be46NinBEWtO8H/PJwW
V/FB0eENrek9+6FscG3Ee3u+AM0gETwrrLPxf8k4/DQhPxcS//YWV0YiwbxGbIqH
IYulGcpIdwdU8lW4F9FJUm48zi6tr7OmIL1RlQceZ8eu7ByzCFMYL62fVkQhAZyg
dLQ4o8BBKjIbPJZ1sd7ugSVgRY+avUgy5NrY8neOoswQ/NpDYS1Br5hua/eCbdrn
pecTeb3b/sN2Kzp74C+uoF/lYsFmZmSYKz5THayOntGogikeMN1ngASasJpxgNgb
7pemHhoZXevepCr7mXtEk1Pcvu0veRn6qbOQAFevJeOJs/Pd2KtyfAxQ7QF0lXlj
/b7f5cf2QDVKELFARh17sPA1y5ZntC8C1m1bU0j4r9vw93tgtLTxHwyOIVBRglF9
AtvBrQLQft1O1Gw3H9v5jNumL8R4/oOfvYfbUzTXiDSdvEPmialqKkIE7ngwRFFd
Zw141KpicYzKftPgsOrkSXddt9SoQmo/+U6ZTvq6UdU4oYYibkbVIOAHlKUMEr5S
9PbQ77UDdakgwVPJ/EaNW3R1Fv8ZDl98i+Qw7NRuDWVzAkm1i5dMVyL3UaqmZMCL
MCNkcgwOD04cldn7slPHO9m7qqlvDXBVOKPEdqS7UQUGcwGYDcayOvKCyvmwSd1K
wWNGiDqyVXyY/zXc6v2yVzR26ykxQL6dtp0m57agcg0vBGxqZp4hxpOj1LJtuhke
YPVz9wRCs63V5MKUW1ccCsdQNmMgdz0V3Ps/PY6ZaKMRp1qUWhW5wIx8+fm+BIXl
JU20aGjilXCofD8OIUHnRP1Ryf612tm26/b3BL2NO6maQSADjuSgtPWj6GqAzMwT
ciFsrX+P9ClzHpHXwAkkUyho1SMZ11xO2ssCZBKes58BS1gfe7k5zvxYSo9uDGeH
rl0xKS2UnwLe/TKW4x2gATTpiSSNs9ThGExF5GqZjE3+HtBu/Sk5+wek+kSQoqd/
6Nq5XB6FAa9JLnb4w2uTd4gky4nxXNLcw9LfGrZABmQjOBaKqs6GlRxorORgVm4z
5g1/hWgPF3C3mVbe3pXDRl23Q8pb3+ORNDrTGkPAoPlaj28kz1l/WgexpfaOEtjg
+yue89FzW9jWtNKDKBM/tex0fL0Nizorau/O2N66ajkfKgkcD7C5UiK13Q2rC/0T
Mb50Jsln+2vshs8rpheQbvsziHy3wQeEM4tL5U2DT6nSCpADn15cv+jbi5vGsV+O
4XnURMzh2ShmeCwcxN686kgxjwWHsiF1dnBj0HeAndizSGALP8PrmlFb8YOETovX
ZOJhWpJhunkqlWCtNaanSCACnLqktiKPSYxOEtLhNp3rMGEPSIIKZ4HvkJRb7Ob8
EAmT3kfIuFfQ+fwB1RbABEN4gzdxW+VEzQH15mUzUzue+el4MFTP6Bti4Vs/NVib
baGYwNtD42TwY5SdEm326uhKCOUyqmtWGV4hkMPDMX4EMwYHQZe6eGd6xOfNmW7D
mDD5fT0oShmW+u1zZPip7gqv4Y4QHbeicW/ycyLot5icMUAgVjOQK+I+va1h5aqV
gSdL4RrYxAMHGQNDP98sym2m8GznMBqYIGe2s8L4sWlRrHyt4WnDLVpbVT+7+HKk
xOxm4JKAxw2monQC1wlCcRJsFJiplSHCkZZXtCiTyi4wByusx1c/bEOlkLCCF+xa
WOqQFdGSK0cPuHW07DaPRv5cgRjoYS5Nvo4r6OmHb/sGiVWd8uVX2/nXXI+3vV0o
+6VVntYLOTF41Lwoxa4eWw3063hdVI9uAI8IRi76qtsvemvh7TgV3EfzGCF1FLho
d5+cNR39OgpLtGdrglCyNLW816Mjp6wyBqtQCXCe+uPzUvSwAS0UEko4xGuy9CBS
XRXEDCiSJxbTGfv8ZyrK2bpMnXRX7bRgsjTJAFl0f1fDA2i+wog4VKscEeKNChCQ
YQmq1Ch0fJMTiqpPzF4ff8v+t1nzSo8FFWju5BX5BHDJqa3wYeNNGQwFzU7xIO6/
0PUNAcMmVe6eH9+WC8qUO5Eg8wXSXut1oXMsQsn1IG6wXdatTzggZpA2B9CXIg/a
a4fh2eLO1kgUAvjzDyGlYdtuKiQ2gVXA20bmx8LQ9rwIsOOqjsnVciT5Yn2pjD1V
aylfd51orO461WRAdDjQ1KlK8z1kL8/D+/U8ohZ+zZcoeXd4Lebh0bQ2rZG1QTua
lYEsq7BV9BuQ4G9Qd4GgVOMbG0mS3xK7LS4tlfFeO1Es0AxEpZjFEhwa9jCj8K/f
7Wf3jO2m/mpmhWkTFz65RDmonPya8a+LsRs4oJ0EaV+HHuBPIpNZ53fMEvJk9hLA
XKFoCAp0CzRlH8R+ieK2MptSyidbdMlOR0nSF/EhpVs3pyH2Hk+uYZdl/1jldU9L
pMrn+nYEQZWC9a/HTcL6WW7wBQ4PFq1WHTNCCpkhrH77tt6VHxOhxtTJiEkRMakd
K7x9kaMmDMs0BKZUvw9ebTvm7FpJLZUbRtKz+8DRdX2bTgJyoWZfF7nlbFc0fk/q
PLKwUUGX0Ms/Z0oGf9ayd0CIy29lw/molPTriYKxGdw7Rpsx8luE53KGxrhX0Feb
4dvwJmS/VftL++er0RNmADXftTfE2bwbUoBqXkAf1nvh+0nQsYDpf6oYt2n2LX97
cwyZ+fkECe7/dkDh3HQ2Yywi78yNpht9+B+yvJn9q+Nr/cab+i3jEnm7fNZUe+fH
4GSHReU9NZ68dVfg72j7fdGSoyaaWF1TTjCd8GEKZNeadvpu8aXxIvuGNl1X+wbf
CLSZpHWi0NdaH9cY5+3zrTQJu5luqGa3BYeLc+c484LV7pcKtnvddyC2FIGkaJsY
T43BiVluVKaGzr9ABX7vI2l9E93i5++3cPOpC9yVgDA/zByFPpJ9V0d5VcN816LL
CmDmXLp26hsJYfSSuZevBPWBGlSPr08xheGpMbdsQ6ChzzxiydNGHh0xIBmh2tGF
4zcUW5PD16OwCPfHMnJD/ugPZ21NtpkGut0rXtjZ0GhS+iVr5zmIOGdFjTLFtMIT
kfKX26ZJ2VhKR+xiNLcU1PiDaq2Ut86Lo1ciljjeKpMwdcFwz/bakziaCHbJIMfm
kMfulACpsZYnEqgQ5MkbI7dGX+a2/ksNQjaSgaYN72+398lH5UhVI2MkNxpKbWK9
SnaZJ3DM9w/nMm75H5J6E2j1CS5C5CApCsLV42Iadx/3jvM2DRTrPo1QbxXW/qLu
3FpwZmKy+r5fThTLl18/3HgsWa661p5XVFMX6vYAu+j8wUnSYGBz1feuV+D0Y42O
HXYFPvDBvi7981oD62E7dy5xQUo6hxpOIPBUAYx8S823Q/seVnKueHtcaV5zQSPm
xuumPG/wHHq5X3BUZZYXkOv5gm4NL9lAZfLQIRjLbS1D4fbdfVS7hqFrJnwn9dkN
HFEiNgsbPD0KLYEYtaFh/UXCi9ageEsDmBiKHVBoz07SS8vCMNVT/BBKbR8CUv+b
U1IRA4dEpMjE2aOaXTueG2vJ2uJCFF9HI6H+HxQ7nW31WFhVv2mCGh14fH45ugi2
DHYccuEgHJ3qTE4Y25fbzZAqoEDVZQZ/91JLVoHts7/Nnh7esm746oCt0ywYPEsz
SOGm4+fQjvRW4QEDpnK5K34wGPGJ1Lz2MyFOKbIWbK8EcJ+oPIxdwchg1E5Sbp4L
QDBal7OQi1PmMtXG6726pNASHk0F15rIImdgWCWYGwXvARaRmVSo/9eGsffDQYeU
oXXMD54kYsP8T3qYtU/Eu48dJUtyohmyA+uqxHcriaWPivDnsbygZ4Y4B5FC5+PZ
bb8kHtUP1VFSagKj62373XsywHyQaE/BHxhmuf5XYBG2yoJ2sqMqtlhSkJzR//PD
GBBSD5xwkXryLsjHS1Fa9IrZa/f8xJAzzE5EIThrMgYg3irCfGmtZklTLsq0sQLZ
8Q1ge4X+gNFajoK/UVxebQiKyf8ISChmuiD58dQpQlNqqpE5mrcrCY5lVx45Xc2q
W3Rx/AzqGpUCL65OWdMNRp0F/YMn/urIqdYg/j2YFewNXKG5zU9pO2wK6azyaxk/
KGVwh9Q7LH7Et34HnHzj+ORMlCc+ZwUBU951wuemfZujiTQUlCSs0WHJAaYAoOFK
maDUqeT9/rqmPL5L9tJbVmsU3sPtTw8+WLQS8KF3jLqYtebiEDDy+e+oywGomC+h
5pAnLcTOuHgB4kI9h3cZxN7oWwA31er4e+gOVMCQLmHHNxJdiKVBijyx6ex7yDAA
jl1OFPOHQEAT2wd0VdGVxQhVAMV9RZSRA2mDC0MgTE3ID9qLwngukA8Zq8zMGmEV
iOATC4guSptwHXgBzvxseH17Q9+tNhMOjr/s44hlbKm0557p9N23LMFj0BFJNPaA
RZil7pFoFZQf1CfIvy2uyeuKUdyUIXzeRE0hj5c00zfEQSlnzqAySDeoy79Rddh5
Lgvg81+QXskz6oqia5p2eEvp4SbwRTO3b1+QsJEv5JSxQoT9E93Migh6Qd6BGy7H
MkFzjfjiTj8f9lUqeHviFFIaOOo2N/61Ft6LgyZvdMT9qfYvLgmJkF/kfvlcqAsN
tCP9gblMmjxTWBmaECqcRNB5L6C0Yak3Y+0+omKUAuwiVRBoV3cd0tZ8GFIUe0RK
XELNrn/34KQ1AtcB4lh891gCRAS/fI4z2YMi3Mow18e8/7az1RXxG2f7rz/wLGzj
y7sUffqvoQxXWUa/YJ8ZHtAWIphz7Vcfe0BHvONXV99je+q5F8/L8TeECF7n/k9I
4eu2vfWVOmFdGtoC3HJdxNRxdoU7+ySGoHmklkFlJ/Jgl+a2yvulXf6IPxvrVSec
KK/0ZEs+8J5U2aMMyGrdo5PSGv313X8yEmQ0RM/s+zZUtAoZZlGOZHczYnLckgWI
Rq7wnujH2ppr9YQUbMZXIw3+EwosGBaJXe5LMuNuB5Og4E+15qJjybCfc0bDGdl/
NFeLqkmQTz9UOVqcjuPULwK4OEe45V75a96ckzC75UfJdtoijmJGtpaWIxIdFWZC
mCaYJhLc+KktOgHCYBxh6yQzbkit9FXo7O5+91/aYy9tFYW9hIaGP/PgxEQ1dip9
jZWNFSxMsk1N4+B96ZGXoPZ5PcscMn2RvhJ4K5BnDrZWNuryBB0kqnsPJPj/riQS
iIfOxhdBhGcx3/J26/1JGiYHlPGvtKJhSTqVfiBHY5953THiYxGBb78Vqr+Jm705
7SwkkBlmtNX1GjZ/xq2uIX2hVd6C6i6NN8S+1dhq2QVo9DCMH3rmh5+qKQqslo9l
u2LsmYF1k3JpWimoKxJjTEwnwrG+ogPCnWCmaoyDBFDg+9IkhaTsONa3a2a58UUN
V1Dl/VyQqL20JsGsr+z5H449xQw+bEdN1i64LdN9TlE92vTYY/zUdnnjz0wDE3xe
shLEPB1Ro8gRvE0/9jUjIo6K8t/8qoFjgU/2oc0OFOQ7JqlB+ghK7R6vQZA09z+0
5HbAUMpeGp2JHWa/HcEZR2znvjd4dCtNXAX/U8tCYxD/jwUcS/gMuZ0GqJTTCV+I
qV+TXo+n/06IQBi4f6279xB/lM9hB3Un4xuesfE8GCdWXwgRyQsxhoCJ5sNeO7dZ
Z1wbgLwck/ZT72OXO4jYs9Fk647s+Hr3Ap1vO9hv5T1EqmGIeOBHSv7B3XAONwfe
2v5Hca+nb0UUGbjOo+3qUx2RXypAGutie9N9aMhXhvHNPLlZpwEX3IDIT1tp5S6a
fxTdozrQe1SBXpW473zq6dVL0mPaguiABKkGzkEUX/YrvDihjJZf0TSJh0/Mic+/
Gz67MQ2carGtO16XKDNQpXTkk+1KXbXWpDd8E2vtxTNhBLbT2u41D4GTLCm/f+FR
He3goSRjI30QmMiS1Uts9aEVFQrIyH2nIr2YIGihkMyVDUnAoRibsMcC1v/+qKom
o0YaKI9ALkUaLYLSUI3AU96/x6D+p8C4u4STSl9pvd5C36kUoebgae2tzouNhn0U
/t+on8G0nD8EsC4+5ryrdfhg/GTKQ4AkTDHFLXnzJ5NaSZYqlvXE33LrZVnrJKnN
yW227rDOWbd5QBFivX0FCFPW117YNImy7r4fKnzd2tpjWNpvmWqkq5Kj5/+uuJ96
MGDmuYrqwvZuuavG5TOQrfbNVoNYvIs2FXJAFPYfXmPPAFXRsaeFzR2SEVc7h+Hl
0vcg2K7NSJIuL275VGCTx6ALW0KNEPb82wSJN4kpB3BKwydlcMpBFjWr5ASk8ntY
0Yh2bOvLLXZg69JNOgNMbjYxofoDvRXx0K4zzZCgbjsva1yTuHqLE4iuf96ccA/1
a6JKCiIX1AibFO/BMcNW52zSGj949tHDyMGJdj4np2kaZ369QOM0pAWqTyNybNOZ
aTY21ei793biXndXabALAtZMT2tjGmZJHeYBDtecMVTCNVqRuwugGG9kFokRupil
6vD9LPZsEUfCekxsbSn22NY3wSAEadN3VTR1au+sHoqb6ZD7BHKUVj8+oEUFKzWn
U8NmN1vfZOL//DFur2YIj+vEAWzivsjvpj6B8mxqVZ8X4vJlb2icQbBoxnQhkkMo
3wlP8IjPmDKhTCUO5sUS9UsQYcS0Gxncruz6JydP3F9yfZhNA76/uJkzpIfI0tdd
+14KmxGfYlmADKM7EIhEIt5MVD8SmONxlmHtzCT0Rw7pRvB0RYoKlNDXfH1o6Bmu
lihjRdXNbYy9CJ44FvGvkiPmoNAZBzHko2kOJbYwkgsDEMtTQ9Mkb8nJj5798bYN
Xu6eBtLtwugwtt5DPjvpAsnTgpsm3UE5YsGnQADIzfT8Hqls/ZItpshwFGWnjYGe
iDF6Fhn5w5f1/+W1+MrslcHFnQvjRk5cNhLPo3fs2/vslF2OmaLKuUpkhkKGwIxI
Us08YmiXoI8wuMpleVRS7qu0/48IixwkwA0gBpKgWI16Coe2XWeucQNc7DY0uaFI
V8nWJ33vt740UCW8TvPjYoulIE2UcvL03kv96rzNyT0WPMjVI8D1VPNHwnIIGOpn
bPYSklV05uys1wX+SAy5D/4EL6y9UZomLDCS7wsvZMOsCKO3/EuoSq1h75lre+tc
fUjq2La1eheKyuPWqR1RhyRyjF2hR6pgy2v7vv9ANbrsAr5o3mjyw5qLLsPnAPaR
rNFIdi1ZvfoFM8kB/RfL4KUhy4jVYxrYy2C/S20NTmqXmsgsDOPOMcUpDu2UE+vz
0ba/v3lpdNXP7bSxFbb02YZvWdpO+X/7bpfHNrwE/1AdtqqPkb6zXtCWPAPjAJSp
yAA9pu6qBeGSmodz//nN2pJEHG/AWcJVVZWpkNFNEE9xf7Zl1VU07O9qeuJY8aVT
wBo6Hp6VEE6nsDUW2vl8jNiJXn6PXi7zfShkuWGKWphWZUj853JnLQd8iMY5Lvy5
KIT26VQtjd4PIws8Uq4uwhPRBdOHPzjZ8ixsULUvMKt1teRQXVWQeYXmouO28xv6
nFS431TR4HWEm6vMN74z5FBKpcdNOuEb5lPiq2TcJWHRGCrjIuByxAokUZZmSgHf
RiXAIkIjA15Gp6m0s1uiO72BiYAqNV12nSxVgCtfQlttepZvGXMp8L6KdNvJTK0l
3DxW2p8v3PAjM/FoYjkaLHm03AlW+ZiQq9MOGZk1J/xcl8oGRDf3lA7vuxVFj949
sXOMCwEiA0NMrqrzSALhtA76lxbIUd707pnKpxzvZxvY/sOIcnfsMxV+txC/I1aF
me4twEpgOXWUhKSweK1oVkkF3Uvc6fmdTFWy/D4p7k4YztZg2zIzlEcf5mqL+hBq
B7DK2jR/BCf/eTsvtkS1aO3UkM+2kh8WsNse2oJz/siZm7BxDA/0PCm9LHBl/Z5z
RQEq2illT7Wh28kyelytU/WDKulFJCVdm0pWs5K+Ix9rTeaMJWU1Wp6AsbZwLynw
7JlK+m3x0hpdEI6dzUU0CoeSd19dgZAeZrcyALU7e+6naZxHsYKlKzZ1b7z6G24A
4tDvT3pnEF3AVU+rc0upEXn55z9Gpvng3P64YwB1NfsdMOk9fcJfEe5Ye3F1bX6w
G2YoXPEv+CPSA2wj1cudQzK6HlSVfHoDbPaEVoenlCxuDKNveC9reZee5vvx6E0X
atCBhjtsQOlHcohidEy9J60E/zt7sH6uqXlqd+OFa1f1dBmgXk2/wfIqoCrRiCHm
wGag6UCr35EUDcr1xOALGC37XdT/bdgzG8SZ6LtXnooGYkRLFjSuWHUahDiOcww9
bw3zWjTo+tjUXXkSY8bcVZBKrOrCufpMUeGQI4EvcC4DcUKHGpPIIUc3XU8FqUL/
6SjPPS+/RwyLkli7VRHkj7n3ASjLQ7NW9T27cDwKb+bH3TW26pzD9tu6cbDBznOB
cSbjRQvg/xQr114MCQgl3S7DzLO5d1BrRUsA78TNVS9zjY2NIEg4xPwgA+RGq1HW
c73N6PA/PR06WCyi4IYTk9YfGsNRSze20vxBkzAmV26qRXpcUQmLwY1jZIQdFrGW
fYCY9JM6hMmksUD0zm52TBUFN8+4SrHfI6Am+DbP8KsrGMJSds4eckKOxAP/Sztn
NTBFKsoPVgE67ADlLu4GsUOshmqiAxAw2kXg4f24plL8ci4YOiZ6n8G3cP2LZzHO
hyiz2WEQEBm4Ak1y4gA2LCCo3jyZuNlfRH3trY/evR05UqUW96KKE4RPYgK0vJ5b
gSXqIknBoczbELjvLPSul8ZB7rS6ZnFFI/RJU/KB0QikMDNlQ2yW3Bb/lTOzRQz1
i1XYLMWrnFIE+0mtY/j5BNnnXRsHTHHwBqHEUIlw4iRF5CHu/0i/MU3P0W5GR1Jf
HG03VhMQ+TxXsAlLsrPde0LAdjXREEBioCWSXPOY1DUO9L4yQUdI7+XnKo0F/+J0
kpM8awIlrV1azTEaAuaK396wpYvakH4duhMe3aWkm0DJD9o3Ll5IryML2PNBWGFG
3LdwyBgwykPX+oFwVmT2BvgrdM31hTyfOtyNH1zOxYI5brPtHWlD3tDGiqlrJIMO
+vfCd2s5kCjxOYUQy7RIrKFHSIXqtnfqWws8rZ0BU37ZNQOyuxF9mff14kxYSMng
Lp5uDbViBvuYwONzAz9WUXPWem6JnPs39gJYjglusIx+Wp9f5K/ztysESEf7v9qn
Ez+rU69f1L7NQzfFTTI6N/6mKzCwM9mmzjeCiXZHPN0R8IBOd4LOCx/B1BxZLH4X
NclvgfV6JAcFA/BxGQONJH0HjsuK5CfoVOgMmlOEktlu+SmnWxgwLXyOo/NRZ9wo
olp3BrQbESXFRuP6+E+0OJGHMpuXJe0N08VcYb5EUzsaTAA8OFwhnEbRed3ou+xB
Kg4iKpMZme1frf+/985F5WCUbcAAqAcpArX6cGqioLTpEJdJq9bDu4Twr7l60L7h
bL1L54C1N8MCrfkBy5u+ZveKPDm85e6gDsSzMGhlbK3MCXT9jFeLWecdvT9ODAZv
fHQlVmO1pL/bx1pOdYd1kuMD2j24fdFq1uyfyxWSGUDelVHnJgk/YpZjQ8ig4Ij3
iJ+J7hf4bhLaZlL6GdhYvGQg8UQ8qJ1jX2UACzG7nIlMPXfVqVMCY/DdxQa3aiWI
N1LwtI2cXy0ktveWUz0+kB/zzZMV0CY0EFN/9RtyO9GPDO61DEVnNh+vnMIWjDi5
ktQeD43yjUbaJLV2GeivKdW15hpnHxrl5lrSTa4uxgl81VLO7bORNs01g2bJDQ7n
P5oUur9gc84h4lsFBShWIcdsD56mdmNq99Q6639G64wKMt79mQalgWJMpxKfqc5o
zLurjhz3X/8aVZaFocgvVRQbwqQslLhg7oeenSi7W+0s11a3segO0F80ZbxcLegq
jlGKNMN/skMAMAlRuI00oSJo12jduP8RSSFLSogM+gOg5AUYrVSYMHK24h42KSFl
ysB/pTbFTfQjQV59UW562FPnjCvVQA56SJxiZvU01Vp5Nw0Xrw1r9/EVrQ7AhNhZ
x7fua67AjkDOojrWOs5hPBhKN9gGT8oQqE4G5I5wOr3wkLct44vEaStyL/Wq25Mj
7b5yIOSpTUXHLlhZioPNNFDGPmM+m7UciOcBt2EU/vP/wKVWk8Qxn8msEA1Xhfkb
7m/Y8/yplp6PGo5hytJ+g2hK5lTqeYKu5xKnivr0lYnMm6FPLLvXVphQAka3XxTs
I0pqCDgFhfMB+MGWlHv/JovXO/6yy8ubAwBfTnoWlhqUBdGVfcutz6aFJfxoBPRF
F1Dj1c+zU7vhis5aRdrFnUVOzPKZ/jpzyAdr/HKO2RLNvaicA2kWwot2drDuFYHp
BteWJyrPlNwbOEgafoaCoHx1eUtBnKPCG03DXzLC7BLuRT7XnImRSFAOcD2x7Npe
pxNwNmWcQXTXMGouUbVW62w1C67Yw0u3ZyqqfWJ1w0CWTUj6+yrQnj1+V3INogZ6
yyCvOqku0k5C+HbyzzmNyqDQ2d60jJUZn88+UUAXSQ2ZWT7GnqmLGPzsfj1yFkFb
Pt9yTF9/fBtlTrxxdMwzmyjSQvyWR4dZjHmA2PvT0fa3t5g6kDjLaZcQjKikvI88
SrFmaXRzxN+mlQS2BMeK9IMIYlFvOBwJ3wtJwp1mFmMevuqGCjLPwGp4FwRnkYBW
LlL1M1OQuHdMEAJQ/Uqo3HCfCv5tWGJ//xvx0vJVoHAU6d7TdV8k292HzNngPVwY
8ry903JAuaocxMfjP0YG3gFD24g8MKs3Z35Bm6KpRCTAa2QetNCIUTd9TwULokxp
SiK02TyBYCCyhrY+qfQxMrlKqhW545kr7rfiOwLQSPZeAEUkluC7xjj4Md5qet+X
a/cUuJvwzfauZymsemUuQwDML5ArkxEc3mWfZz6VouIsBJufZPyDfRVjwZnRHh4Y
9m6kNU5DXZGpxW2LH2O9W1Gq9/f9HrKdeXQAEQlX5QDbMZvUIKkUSVHOmHP4trfL
oD0a1XtEEci399ek+AP98lUGNHToxJkMrCMe28dPkYkmgb/w/ddzD1yC7wXByjqo
Hv1FcedEfj2+AQu1esGm//qiAFmaPzk8VU6R1tcbIhGUKWpxyk9jwmL/4Ercj562
+Q020ZwXM8coIg/DahBMM4VlXMSjEnMM2VN5Hh4gqI/EZDNrqUdyjSYMshymHDYj
vykgqbNfcFdgNpSHsXxA5BedZuOwWys2EZB9t1OxiXlAmUSnvFttT/Z4aqVT5/m9
/XZWqJioNR56SReFcMDIN0qUYVnV9w2tRGE/i+8srNi7ANTvGnF7Nd5ht4wDkqZy
Od4g22jRS3gJmy+/0CCif/IA98upWTlO05DCL+//wDipO5UBf9Wr+4wYNXRKIe60
h0T+DCywdSYTuhCFBV6cqQk7CZRr/81dtuilbHHI8iFcCyX945FxJmlZ0G1wpLgS
qZgT7C80BdYOiExOiaRgSYFfB7fn8122DQ5elyexKGSMQ3VQgf1Sako5RJZLFBum
E89/fz0LBOQmIFToBMjaFWdutQdl0CR1f8XmyEv9E+FmFkFJzZyCqazasYNDl20f
mHnj0u88Ewmt5p2HEPT+Q6UXMITVnBF7Gdp36bZN6+wtoGjtHqjfU9dnSj0sjWsa

`pragma protect end_protected

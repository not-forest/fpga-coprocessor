// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
oNFNZlS3kA3qnnCS2bOHNMgTFwmTjLH74LtIA66AyWAA7f0mPQn+LBrLvmZKkMZS
6bBD7cDHnZJ23TlHOovXJ3wmYP3ryUQM3v5j5QXhaas4hk+N6G2vomz8uUFy04UK
4zl6sKSK/PT/ytmtpSVy1JVsuLzBeiCIVcelQ9UFcu0Hd0R6dSNyKphU/XSwau57
DFg0VkpDwecySqPUiwt27I5f10K94gdM/vQpR8Ga/lKHkWpgs3UAw8GOhOcJ6KN1
7Cc9GFebyv8bQ6Woy5dORuKIbnn9jyaLZQ2pm+UO56fO2yFAwxIcpDKAfJZrHUC1
UYY2dj+chx4BRYRqfOMomQ==
//pragma protect end_key_block
//pragma protect digest_block
+nC/sTSrCBmxQh7G7kRKA/tThHA=
//pragma protect end_digest_block
//pragma protect data_block
u/unaUOSxCUafFj1vlqbBm0ZU5Z03eYrrmBaK3BSwAEpH+U1j8TlDwLBMmvlQGb5
ypJV/pB9apnemsMPf+KgkmwYHeks3RBPv8JVKg1/Bhqgy6W7+Eew7z8BUkF+I0K+
2WcNZXs32Uf4NL7IxMPacgTJKVjW/7M3h/KgNfCQpx1rdro/zwaQy9dWJbeSwvJ5
0X8kLaDmXrCQ4Zv6Y87Ijz/6zRT0ayYFIaiUHdhc9ws4kKKJ+V/T5mx2mPYSgiOK
AgBkDIcnuWc82/c4wJsZsZrPOFl8mM2JCPHf993kszdz3XWIRtUncJ/wHBre4WVU
muNkV6sk6+eY9tQP8T91iRRVMqeAtfGnX94HrJWppdMlaLBwSKIs88J8wNyur85w
0WacxLhDSEOwIHn5HgJgLI6FdoJISD1vSH+6qNX2a82J/XKPTWzG8My1uNxq+2IK
ARo7QYocwXUoE+eor7HsfphNKywCTv0x8C0GU18nywAs08440HILpZcOPnx3XZQu
V+f10TQW1xRoA/5g6q349/zGyuXNgVfN9sjT0rALf+8jrN3mA8eIeBWlryMzQSnw
7OYCdv7HOOczOBOYV0OOSkNlN0pSewKUn1JsiRxJeA8iz5hAZkKxwQDa5E4dPy8c
9GcNNKx6w7W4ydKpQ9GeCY4u1Q9NYHcC5boqIRlqDA6/XYnK5Eha1jQFD11Owjif
O2R6Y3fR63WPIvBmSrbhZbd5Vfm9pgf/rO8iiP0du5Cn/oU8el68KF6FbXVA9OsY
fdOREyD03x8ovp9qWv+at+XYlHS7xwgEeKFyNxoCxFU22hYPrqv222UWBGi1qCjI
9DLt8goSk+//PVcD0ZxDe1rhktsBXkkub/09v+N1AXzV2gvPe4V9qRQVi1xAUFnQ
902/I1Ji79qayMnlk/qx/JG0m0LSWzPdSvzcLvyEfVYfD8UdXf5jWslfut6CbX+k
qUbhmnhy//P0eJ8aNSy4NiXa5rjF7a14PnVYFGZ4eu5SEw6oajr43tsmeUq1SkLo
wdHM/H1d5mNxteQsYmF1Sgyznt3DpNL/g1w4ecF5OfXYYvhGhEOrWpCV2e3kJXV+
InB/M6sHcbWbB+fDI4+5KU5MAPb49STs6zuD0MTmwbrlY2DE64gWwoao5sU4koPa
1qljtOSHzUSuZsIIHEC5cPB1cNAxqNbV6fb4GX0S7TQlOitN0q8VcOHoSvFzzZEm
TQsasFldPNnXZ9D/lSD1vwv1nlcPo98GgeZ5HWnVzRirVuWHXoiO6FTHgFAH7q6n
x0/7eL9trUGXhmtmWlsBBu0jipdlVRuyG9+F072jE3O9T7EcmDzpyTeOVqxO0f6F
L4CKyULTGTx0Fq/6GX+L44XuOLZqfCqJdIkdkzl0ARsdm/5wRRDLk4IkX/hYy/0S
nZ4BZJFBYfdFivXUV66BGL8zVX2RkjJu1En5Je6lKJayP3wIgs3x+WCNhlZHGZ+/
ZS3On71Unfujbwe8NEFOZydocRcC3iACz2NRTw/F0orXVOFKZhLLmiO1+a1QVSmA
ERNlCuhddiCa7wmVi7L244WNUSLkpkBDexrabwL3hcE3UYfsaKIo06SwpuXkOpRk
GiW+rfOCMYwcQQnHpS3Q32SygPFZYs5Dzh8iY8t7ttmQQm6OHL5F2tYJpB/+DEA3
KH8NmgfWpu5EOUETpTKKAXATORdDkEfntqCNqCpyDD1jN7Zy2FEWeeFWF7FBuOro
TDHj7iVHs07aqxJOj37skt+r4+qmYSQjRAj4n2OuvAglsB3RfPaewEz6XSRGt48H
nCENgC/r5BsfC9O9ji2WtSyvbzGHDlf4YUpsZhSxd2eunG9yR+MSUiozySmctYyP
TF8QQZfuJ7HI62sdtQky6uILBAUMDvyticiGRynmEMd1E7Z9lbGh/1RjARUclxif
uyZzj2tFB4xien3nzgJlAdXi0RimOQsItcc5kwA+nNiukvA58/4UV5s0xqJsoThz
4hfFoeE+UrLYZ9FEOG0pnXBKrezrTAxE6oOT8mp3sCMsDSjMVyDYEgjGrw28V7EZ
6kH2dmmVrrAzU12V2skIJ49RBwOxZPIaMaVTgcIYnexjDYSHcejWHTEgnl9iTP2A
9Mx1s581PZSWbVI3VfSa72iDj/FKe7hiA+i6XlcmHq1/n4JneF1K5xA/ScctNuCK
v6AxP3bg5wlSlRdWki4WSUBoWlD1vwr0pXxWyXUQkGjU4NmjUeYgtb2fvbw1X6eH
y2js5did5Dp6IvC1zrGBqlLZheKdkNVJZtH3/rujcQ5gbVHk2nd/0/bDKCiNGbXr
LfxBwregEoDgDt+6Dz0qjMqSLvUuIZSOrZB/zQsUcjayH7LOaJUS8g54Jd9T3o5N
ZFXD0+e3UJIVj0Z6zay9pEuKdqQBnTB94s0pgwqZWZbma+WF1ywq3AqCCwGw2DJz
RAdDfsXTZE8TYd6HcblINuiFNsiVQx+10M/wSEBNYwp0qTY4gy4eEYsGTgi5jRhA
g8m+NmujqRbPtxcWHJSI3yqkspR2XZ9J9Tn9iXfrEOQ9TzhqyqxsXv62hd9dXoVw
p9W/XpSdLsHoCsBOKZPkMtdvPv2PaGMO+SxWVfWmFw0Hda+S4XtYHPA3lAzhL2i7
Cl9E9XYcBauRmrSxKqbJzPUQ75iI2kuvygCyqKAYQZ9iWrRcVHsCdUBAAK9x9ARN
WxFiscLq8toHxHkynyDqFUvxzA6BIximyxekLjgTyb5aM6CbJdgFjnyM6uhgq03V
5GsEBvtFZ/KM1NkEmyz9eJGJ/j85ZxNCSO1/5kl5amypjgmlZJjK80R0R3G2SXkf
G+mfXAsXf+GviX/Vg12sM3x8AEZM8etwEV7NtwRCxZakMxwcdaGIZgf1eAOVPVcm
fiLNF9HtUKIl0Ky+boLO7P6ehAtgNuklQuMhuxrj7y0aX3jLFJYa2C0lqlpjJxGb
fKdw5kpb29QlXJi+q4g06UFqYgrq6iQkmdCUatGpf6M0PIarkP6cCJ9htbVrzw2P
Z+S9vIAwEoK1HdbrE+TLSGjxa3dqtMMhfdrrh5w1SfzdIAcwXNGorzxtfYX3d+zf
5Djk8pp9aUgo5EivC8rXMh+5U5VeFP0Gw0d9pu9g8oFDo0uz2GeG8+B6lLsYQg7V
XPxUW0sPGe+3XPOWTj589hZxcvn5cnYx0O8l0cx4hicMYRIibWentEsd4+YFTA3A
E/UW55rmx+HbR+qiAAsVrO1tgrv4uRZovyohsWH1AiNZQnbCMvmPcc8oOqvLGGjF
ABlJpCL3/vlBL4jD3/KxRiUit/9XSfd/elLngtpJ0PzgtN2Ogi4bUE9/q6NCGckS
PBkmQXZCkBLzWzviCW2s9gVyj+d2K+kn3/RkZbJH2ycQ90uWHefJhxrXSwutskkK
EJXj0F4PrZsdGRDSxk/I6nbcG0qQ78MaDKqiDN2nQV+JTQYieB9hI0qcQmJAREPn
z6syGO3FVyAOwtNU8n1VxAo6TRsjUz6gF26Cp1sZ3V/keZEhbwsDvP1Ta0HIdG/V
RAAxFwj+/7pewbEYSBmspeo1r3hAxEBliJwpjVDWEixccMxqHKDY6IvzsIr5+25N
TzuzathmXbtqTqvniKDGa3VY5kPHbAHm606Z/4cPJdNyTlYh1Jxn3T55sm6LRrDb
AcMuYvnKkGwu7hckyOClVJkK0IoWeu8ZlJ25yHrtyREtEz7p3vrV+VFlkHwTriA1
LPnb9hSqRlIb/E0Zo5gGVKm01HnZj/w4PpEWKhuDp3Z3rnaUSWmekmRX11dH9TWL
z+3BaVoYzLptB/BPXs8XizH/bUFSR5CDvqBvJdWINeN47uS+a6bCEwoyq8StG5F3
j7uW1SAnQ4rnGHim9EVagqmSa+q1k+HsKyQ0RWA2aZzTvKopPIaLYy3IojBd37WG
R9P8sQjBqxtE9YGlnu7n0x/y6g6f9EPbhqIcjF/ZkakSJeKCQ05PbEsqpbkVZNq9
SFgR/PU7b4IHwN7aIpsxoe0Tle731Li2fkSMV6fGre0lXDEG3XDCraVau6MF/9/S
nXGQvYiIC4umvO09jgvAsh9xtOHORFOvZ2CqpuzybPhkBRuK8O7qzO3tBkZvERp8
fc9jSLfK8mKlXM8gBo4F8OAmXcSyoi2ow6JcFRjb7xRcd3kYvRFKVaTJt6OckW+y
gE5fKnR0scvfEIcmYgn8Vm1WQUHpQ0XLpvMbb2onAvglTT1s3AoXaS/Pn+vMCVqh
6SxH09hQpbVqGNOJpNaManDlyNixUUgFnAoyh1OizxoDzbbzxFPQ2eacwLt8v35u
DzpJjHOvSEFyRjfrYcPJSY+L5cqlX5zEoxEN09JfCYmX1J4iSSB00nuQSBfIBg/F
Dz98jEPwb2ePj7EihmpTeNYZ9ZngDGxpkztghy4sCrGiok1WLrAqFKawpHxHA+GZ
OOZnMz0q30nKclc0G3K1LD6VMDYtlaeBqa2axnSJBrgjRKHIX8junrLNAYxlGtS2
ClVN5+HkE9Vx0I/bAbg0BaDP5BAFiF2Ov9nOJbfwO+kBioMIA95o+rhRHw7rAT1R
cLpS14yov8cnX+BF62P2pj1C3y4DgW2tQ9Clc/SvwnqiNuC7IvYoDFl5ieIsqgKf
mjv5JFLPow+Tebkg20Pge1/yJBpCL+3uJWVRfpjGVi5ByibAcYD6ClQtX0wDjN3I
Vi0Zyvs117KxSJxJ4Uq+VW+Q19pZcMUD+bJqbppEIgWfo9l5oonl/oH1MEI02O8I
23GAWDseDBe3Ed/J80lSeOfM2P2/mBSpXcI1M0ytwODhY5KswTxwuEIa0tzFdVdb
+n+bfMXAviPzhQiMnhyIxxV3CN5LJ4StyJ9+UkIMIy5muQ66FeQ5PNXYyut8ilRq
ELRo0VO79w/WEm4v0EnYBRMQ0uYWDL3X5KKtkMlooZHeug2+FhR3PpelBkGzWDmd
QaPaLJRPUF8uaJr+2MRq4rQGwArVXffAYWxJRJH65jFJL2M05C+PmtH08FmI1d9F
1Jje9O+Q/5Z7yPCRQrLtxOgoJgOq858ousVm6dn5wdQz4EHaxXAxVgBnw7iL3wIq
9SsHGjd6gzZkSfDdna3ct1uCLdYP2/al4eMCZ5ao5vZPReIR/C49lT7BG0jgzIC4
vHldz8VFW1DLIlmEF6M1bC4R0H2g7UmFEpfJV+G2IJ1Qu9TU74vZ+3YymPRRMbfV
sjYD8V7z6FBVNhmijzlwA0+NILezq2fm7A9Gepp/uJrDBc95Xf+A4QQOkhUEDQrS
BYrkTEvJt5dVPrq5aBGRv17OH9oOqsCyOtvpfID3B2TdAJYG7MnPksGMWZzeAN7P
8qkCpSfiTU6rxsGAGK3ErBAuzelAjc4E4F9oi1quIzSj7yypgXgTEqZJ+DfcK0ZB
04A0Yzk1Y00Hrvw/IWHDb7N446aPbvgqgljgUK8BnNcRhLgtJMZfnaWXNQjyi4aV
cI6vr+3depzJ7c0XEvyutN/pD4PNarr9wFE26Y49ypaXBIqJ7te8j5czKwl3cqPf
KQsd72iiQTvzfGerWiFCpu3YNYNv9wixb86P8tpZ+FmJ1kZp22ZF02GsjgJQrBUG
MMdZuPCkELF/mpAU840ySfI7Yv6QmpiDQip1oVwQxskDdVbQ2ndlKfkykAqyRQ8i
uA6sYmQFkPxtWj9j9Y/tG1xqRNG9eRpchhB/3x/UYuEnrtsPq01oE+EFswR1J0TA
cTDeioELRR8ToGOuMmM+2GDXgUS3V56BFOhMthhQL87hs8VVWXood9+rUT1WoFGL
7+zx12oBctQXq1uf0Z2B4uFiJaZgwcRL6Kbtz70XTEkUnpaPSk/7w8Y3s7Q3qpsf
CHHLJ+ru/Mdl1V3Va3dK7zeDIb3CulxQGk0dHr4giRfm6syJVj2/OIAhS2wbMQXf
8lx9xgfkjGOr3KpgfZmqklfeRlOw9yjgtMp1+1+C6qx/KXlqP7kEmU0N0Y9c+XYk
iys0sIGY6xvDXfc9DprFexUnLdq/lHguZ7etJBGFxOBnDH9aHjQZAQzhSMEKz3F3
nziJtdlQjIH8sqvf7Nvjn7IoK0KfLrM/7QsJppcxKX2H9ccJPS+46HbXNhGwq4Mw
0548/naWLJmf3x+eC5SIT1//7P5EALN74IonM/gRF9cG/XKY9OvGUDGYjeF7LYIk
6OScI/DTOWBN+VKqrBaaLY5SAdyCAzFraJuc9+s1YaFFHALJJ8ebKKK1ZHu2/CA3
e7kwylNgM4YmiOocgWC71LAw8TAmawujILV+BQCQFnYm08mXQpQPieQrd2uI6HN7
jiKWcTcSmoUvgDLPqp6zqAfcEqAYhJXNdQiFxicb6a0TJ8n0+lAw/QuXE/Yf6njJ
ND7UY3W0UKzhnNazSoyHcSDZ81U7qJgyrBMhezbqWjFV7zhsZt1KvC2Lg+Ci4en0
WeoI0juLKx73AqjntzfbaD5Zxba7Dz7G8oJ7oNulm9yls0U4o50mJcDuFbSplTiG
hGNK2piFytLVrzC6rHCcav+PSJl46C3z0jRHfj5rbuHivEYvFK+TNEl4iw0brouP
B3zYFGTmhu3D2X+904yUdqax6fhfGxPbXzxF62Q+Y7EJIfYVKDKj6Ek/g9Jt4LmB
B/8rdnbO6JZmwrhCj4tvVDR5TeJcVJN0KYfrokWLrCbBqZuie/dVmuOj5LF7gzka
6j4ckAW8SjySeEDnkIF+kR9PB6KSfzwBiRh+VS1deq1smsAVbu9p8EMv1d4cTCff
+gYCn/CEJQIJkuvuOdtV5gQKfHiy2keJz71e/UlMukpW1g12hRCjGOkOLhty1n/6
uPq1TfRAFKEfCGIoqwkxdbVAc8NAtQXkEvKuwRXoO5IbB+VyF8xdgkHBeMhBRxy6
46Sq3UH7OctTfJqqFMcFZNrscXTuNRa/SCcP0JNR4dbxHiJlydCbLJjJGuDkjGm6
JeKBStI4JMk1YEWAqLvajse1XEQm01Zs/Dl5tKJ6p5vcWy/ZFAiEHMR2Uzd8uH9a
HtkttEBcGU9OQkuCFDVZn0r+x+ZQ1GtSR6DmyrAE7IBMJt4PBnIJ968U7/8V7pX3
ijw2IEqy/5Sl0aFI1BR6xp8d/ak865/0+aXTJ1HPF4Pn8hV7sPpz+2gTntJcDpzg
gYAwRIA8/K8/DzMS36uAUPMmlBNafGs8AbCHNiyz5qZihATgCaxrViEFEiUXbFhQ
CTm2OiiiqX8tRkJQPsTrKdo0oO1e+CrUz4vrJOV8y04SWbEXa5i2fRhdy8BF9C4n
M37LwHFijYAz1ujfmyvcv1EUDF38US1ma2hmmvguk8w6b3HeBTzZhTB7zQZT9QZ6
BWCTRKx6orqFU17XAxUeS3OAQV6naIddHMl8xoM7v9oR55RowQo58rXq/sQDQYnD
Rhh5CmgwxrqnBV5ojCJ4FUdLghQWUS5DdRHdYJ0j66rnHB7gKYbyzrVsms7QzCyN
JPDtAMTqOc7FFFTiIcVMoF2ZshmnH5DsDuTkm6WLYB9ouIWhk61ZtFxLZ5ChE2zq
xP8Yz1ttFrijjFLUO6ma+UGR2cDEFpFplaMH3kQPd5kSV1KKvhebBXq+A5fR2xG7
pJkUsf4LbEHHKiTuQdBTvi/V1H7f0I+4tRG71+YpcAIc+XP7QUOr7fmzQAIg/3lv
+/z0ZUx8mIeIniZAKBr1sncZK0OgAJb/JusxHIKXS1ZQvxlAme8Rd0CQtmrgTPZv
vM5shCzPlBE/km5RXzepJjUUaVDCIr/iJATFqUAqHIVqPp7VAm/Uuzi4IOqiaxy/
ZzDymvL3hbIw8QFczlnIYlQXVgQ3W82r3tMqe54r8Aqgar9YekWrehMLbmROFu0L
xJ1gDYX6DiQ35IIlKuYRgTulPNg3p9HxwKhjHKVU7O1XzlShEH/Lwndhw2tZCfXW
Rkkk2Xvh2TYczNFfKTwZpFg514zehEZJAsLwFowCuE1UBjWpmXN0kJIzuYMCBFGj
E/XjkAtuU3KwnjBGKTiFXhZiDII1rF72C3mMel7UghiA5VYU+K7E1ULrxYZn1AzC
fxREKBkq/GLu407yABRd8N9aISjBt5dyEk9WNUi6KVAwCtRNrLN+bsnAYMSVMYx1
vQyuyzwDQo+UCryocEQraA5m5+h9QJcDIClPB3Da3+pUHriWKxuNjdBaK3uKsS1p
4r9adweuaZJwa/F1xeqwp7dX6Vnnt1mQ3UeMMSdGaZFqYUXty3bbb+S3J2QnVwB6
Wka2HXSQFD50WELwCRG1C5QzGK8bF8yJpEyGkqK4+WeE40NSWnbn2kioGvpAQrZK
uBy1ovtwhNfydwyU/9/7D7DQgJpx4KAsg7obuu4/3U/TQ18WVpkDmODpH25p+bB7
0+FQYCkQ77A4RK0t+xjvvJJ7VjrE5Tl9LGCvSp2XlQNzNaJuUomiiH+QBXfK39RX
ehZojC/UYzyw2E0Cq1XvIEXaO3kTwVFLylAa/EF+B1lPdJyc+RNiULhTDlcKJdZU
4IL6i8stk9jUcXE7D0lSk9J0hXzsV+Q0HLj/exTgNuh3ZFKQZOHXpAtE11/cKisy
aBxxvz5QURBiwpSoM8OnDKvZF5+8JScYWY9ezf79GFvI/vbTnsBYx5thXmneZ8+r
fdWm1V8F6cRfgw01qALwt5FQiLpPt3/hmwtnt8w+9emTAPcvs656kQ+AqWbjald8
f/42rm5zaW+CirURcKR2ifQeZthK4XF/S1omM6VED1qrhX0xSqVbrF8yltUsaqQF
4CjxuGDrD0a1rGnhJXNESgQz+/S9A7IFhZpcd1/6P4ScN/bRU2aql+q6K4zNO/FQ
IHVjBh3tufV1HJdwY3ZJUH6f3RL8n422K+fKidgSzT+t3fZWKP0eig1F7davckfW
n8/RC53ramB1pLI2Wf1aIJy/dsrGm7SuqVKPFLPG5bM/c1H4lFVQY5rYJh3m0ezw
+tj0u4StKUH4Vk4bGIxb3Hy54OcHFQAchbDZPvDWKagemqSQT6Q6ujGWaKwpoGng
NeXipeflARKlricosE23LakafP77nkEsX6RcJ4dB4HN5MSQqpKxul5ywICLV7Vmg
iEZIUAznhQrjwEJwZsy61OJYi/reMJwIXj08XrC+e4u11AJRPN1tCZ8fjIJgU5q1
GyQayegAbZ78h378Se7/q4cw1XgeJBNhSc9a3KcYYVl04iM8GAxU/eArQikMKSSu
OckvDghlBeJ1BsPxwLyVlGFt/1uTwRwAvrOOgs2amXimXWltrvAwUuhDWKsySXLS
KBXETrtiSza0wZx944UxHTGKnNzVLq6cWc8bRlzBgCrTQyuN00MQ4z73FvgIbCZQ
CbjKPVSozsVgB2ouI3abmxY1YSLvnI0pbns6KytJA4e97VRiPb2q+r1ySN9Xj0dZ
qroMXQaAHnB2jjos4eVcS5We/c1aQztxQglk++Lr6LZbgUe1TJxxYT260Tvo8c1U
Ybe6uVq0V4jLqNEwbMQnYI53R3Q5uWgFyjS501BhfkgiOQeFbWeAxSwJ9HAQhuhe
y8j4N4VKlhOd6vOYlryG0jAxtZQPkdsPEGq7Dl3o+BSE9+PgdmBuJeR8xoy5u89l
4TVkqSfBQg/d4+H1Kwblhbu1UVWdueZOE/J3o+8RafjC5+lKkji/Vu5UCs3VtCYY
k1gSQ6UY2Guaqm3a4T9V8ew/CEdAcR2uOOT9u701VTNBXoqqA8OP2CfEnhMRw4AE
djvwB2FgBB0gMuHQ85ujves2QwKBqLsUv6bSRMvVOwQ/DHlFUfCSFHUJQVg82dnD
T73paDzOuhXavMvpNgWJexJKubmBLWSbmrgsJn7FFzC31VlQJEwDuOvCofk9kMVO
s2ZKCmgo6NCUUazPniVKVCtyLOuGlF/8neTK3FChbn5NHOFEH42lwZovSEzM2XYW
yMZYFHUt8ZnlCJUBcTXmVwwrKNWgrWmpoDdkMU55m7PX3OQH4SJFLT1pC8hmWYHG
3xeEhCHXSMrLattR21B2tkX9SGql7zXo3hJL1k0SHOlWAk6tOnOfpv3IFBlzlEJr
y1RD/xIbOZQa4/bHJTdbMKLXKFZ0FiQ4dmF0EtLnVwIYxmoxgSN+b/RQS+gxG/jU
ZTm03D07U5PTVz6OtO3mzgLi6qI0GvAmKwNr8h9roA/Gbhyw8BxZlDE1YMhEcRP8
XWIliBLt7AxH5PhmithjLhdTu1FW1sAYEfwNIw1WI8cdXHo8Ym1bipqSnGU/5StX
sBgjDOG0nJ4PK2sDdUopV1nSRhrjrKhqDcuNCT9ADsS+vJtVwKv3YOiHPRTa0Kym
N7d0oe/S5D28cCb6JeHol7egDh8HrVAXODIc5SQ8oZiRBvWh/JmPlhuDrVMqQAQw
WaRFkvkdtC3nhHGxWFbmQhgAzUUTUOJ98ZmggVdeQkv4S/sU1mQXrhuqN/Olgg/s
lgXPcNXVwZoSAONCPyv2ANgYySrSFt665fhwXe07TEbtuN1/LZV5RqLv41Ip7oiz
XF8ohjicgPgf+uY++eZ+uZDtUk7lsiepKNBr6BP2wv+TlcHQkxIU6l/tsSGybgls
rUkLAuWi6RcPlcARh/eMmCpVejrgj1C0VJIySZ8LhGFo7utZHsHtcI4hNWzFN56L
RTUp2FhaKfvA24uVOcnUi441rpZErzJU4aY/wyDl+cjlDdUXvH3UP1qzOVtEBJ/P
quMkj+AGTiPd9NdlH+uW/nC3zqXCrP6w2ExkPWLTkbfJE4fTUTDi5rubWEc38tzY
Shb84Fezi5gHefPO907Q4gwwAq8Q6OBgVSFA8f9VtR2FpFuy2jBDPC0zGOiklI+1
6jAwOsdSefiJyhgnzV7EV29I8LFyuHZO93BbbCOgXc2cylp4+AE6osA/xnMkCsjT
9Rxj49bEktz3HnTs/jSBpstBo7ZLeWYLNSotnbRB7jedSnbSezP+NX5qsQz7UP3A
4sCGk3IpWs1IpmehF1cbUpQFY1xMtiSqSweChA3OzVA2EI1/nmUtmTPbDWriMrOH
DM+AsjwvJw0DwAVmBqsU8af2jDMcWV961LnvtGNlDJ6tFJTm+XFiDKo2Qn65fw4F
AJXT5e6I4ZnFT+oBfye2VjgeiAD1BRvO3tMreanzBnihF2EIuUpWOoQDIK1ut2Yp
SG3zMju5qAk1AyKAJI//fjz0xTdnT6rI702CMDcWMgE4ERBAO/pnYUUNpopz3DjE
KRvg85S0Q0JpGa2aZUK9SDaZ1desVDDi3mFKbTXqcAtrPnqs/7vr1ezA5j5eaTzf
b/Wrdw+oTHcI+9KHuSqeVWtaG2yBKnxRzoUmpxC+J8HkHEdEed7SLBGhz9jM5X2F
uFWrhI3bseaFNHI2jVnaxg4N9NF+ftGNPK4hx84vr2sOIVwcOE5caJRgPfjKians
fsJvmslEmcYBs4kA3uN5YGuoiLSxRphdYk6/fLmIA5Bng7TRrGD1BXzTK88dB0yH
c8Q58JLGCSBXf5OAeu12+6S9yxo0tPVv5wqnDTH06TnyHq2/LRoVQi2lxEY2r9tk
TIT2x0wpKzL2+nZnzrbFvuSD2d54ToSjNrXFbTVe3UpibCLHT0k4x++kw+15OhHE
EnPtdfAOYD13EgNLFq5lFZKylZ6ZqCz5ty6wcozVvhpQwQrPZ+YWY9tXxinT/ATL
j9nPa2LJaa2oUtpQ6I7Qd701KglqD26+Kg6IBfVpOSbJ+CP59L8C1+Yd4eq7XhYJ
RJhAO4AVL68OdXMlq+YoJP+mJF0+Mopfk02YORa9cD6YFxRFK6WSEiMZ8K3uKnol
/z2CFl1U8N1QNKYKsYKi6li2n1tO8MjD7jkbLQc30l6ykSxs6SWWygsAI6TLff7A
nlni4K0jjM6VOXVdhWA2Jg5BGLrACAKfiJVZ+EcIKfAHwi9Axr7Z70LoWkrABizY
H9anDyPcN73gwJMguOr1oXPfXstnVA5rsPZ93berQ5bpfFAyI6AOTAqE5eRAhTNR
KRAG5BBzutyv1/XLkUO3YLEN+B0+Q6WpGkyb2FkADNMxUX07WeITivhubnEr9k+b
iQFNDsW7/OOwpwVlo7NsuUpOU0f+CvVHlGqu9GnZH7h9LauOePqlGPEuzsv30eBi
BaZoUvAzHUbxDPeNRMxG0rRegwJ4bLLz2mgKaeJz3iaURtVpiFsuduhMX0VAMtRm
uhUrbblj7Dj7c9PCGBlTY2oM76pptGP4nQd6I7NqJA3MR7yeDwLiBXqzJbyzgRvF
UA9vWqnhcvPNmGsRZKfqWOM23NmRowUF6lmT1/zAWYnhDydNCbi3Zs+d4xEOrcTU
nDf1H/qKmTUiB/aIC4NSy5lu+B7wWGFoSOyXEK3Z6Dxib3Zd3iR3mgXTWJP7MAsL
/4KJboVCcafRG78D02eNOTyeo6PS2iILWQ5ApEEywiRviyk6Ztgh9oG0ntIwlGjA
T80wDqoPgW5fvcBX5TPTeMhbwM/rA0aBgILzmnI0yf7VsETKx0BlwOlH600XUOk1
BNx2uRaMNi2Y1xNT7xo/F5Is3CMqkbzUI6xLczqojhUgn+p9BxwWXehM7sAVof4f
KifmkhiTMcPOg4oXHI3hXJPII4IgQq83QGT0GeW3nHsn3+hpk7svg3Shu+T435Yr
JWUBrcdZ8zoEu1M6R4u7idMoXA+Ac1hVukW1eEN2mbg=
//pragma protect end_data_block
//pragma protect digest_block
IyYxPo7Ju35BuS0/bev+sQo055k=
//pragma protect end_digest_block
//pragma protect end_protected

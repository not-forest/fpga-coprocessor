// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
u6ToXiZl+/42mlfeYAeaNeT9LNYr4w4lpU/H0AoCcRrPHOdkJlnZn18yLjnj/+cqhMwKOokg33qY
1eY4Inb8nayO/sRoeitLPXleR/4JbWTUyOrpDGFnJ+e33e9aQzTnZkkJlSBYuWMX8YfeK6kqRonB
tH5hEoo0aJ0GvRfJqgaewPoPtZTyoQ1BvE5B2AJNK56hBraTrl5vebNQJavMTRSaP9X7aFbNWyw6
DCUcvckBQmiP4RFpSPq133BIr48QCmzWm0aUGoiFyJznwfXjFDoOSP6lLFto1HmtrqVI7x1UiR7J
cc/mNIgC1Q0F1ZzYjMi+IVgbmK7DaOm/3E102w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 7472)
cmw1J55jxL+nB8rW8wOBKzTu/xOa0Yk3YZBz0CKClALvtoMVz9EekvI+SmeJipkSlYkH+2doCPyi
O9G4UnxSc8muTRo/4YdetHEwyPSXe2fKjGSoi3bF5V7U7drANH7mHS0aj5XnlM+fgVCTCDvkMJTu
SjF40jTvNZOsqeE70CYnLH8/bxXHpBYFC+JCuHvuQ9fJ4HDsmvjuxoJ4q811pzhCN79BIlgpuM9i
MYB80Zp6UocSw2F/sj4nX/ZW517WFv47NvDAa8BEN2gVyZW2JHCfs0EeY0VEBOyrDsM05rja5/Ik
UvhwVis5Tj9JyDFo+hZ8LkEBuKnCglg7sk2IzAXa9kWTEHYWjIc9Gg+IxpdNpdQho2y82RhbuAVf
PPI71M3UbQRLH5m0qhui3vaUGY+QwvX9hig+JrtZX3k+xXSkt2kYxLNDm5Ybk6T8513zpGNO4Tx8
+LiQtyCL5Hc3Q6N1MxOGf2YZYCLtsvqmvM3SWpE3aF2U9V628V2n+Z/C4NOerD/W0ZMNswoQM/D0
0LwBP6cBqYFby1MBAI6X1NTsWAbzQKOq9v6zdi043oCeuWDjtth1/SoSA7Cg6DI16LLl9Yp9T1r9
mz1F5gSUyg7vzUBfU9OPgqY1NQKupo8OsOsqcK2e9C7EvSHmM2ie3zKCPUuZW50YCaAm+45Ol+V5
u5WaB2TTPBSt5hAbnUavpw1qtsmsHNSRo6C7xPkUm7kq5Zn/Fo7WPsA9RCL+OF51eY+wZMolvoCs
lSYtL9mZe9y0oBEBUX7c3uolZJv9nHHnPpJqYaxnGh7yZkAThWzI0kZFWxL/+4YSJiXh+TwBN+7B
BEJSQAUqS89EXSwQn/QAGrnlNibIBPjLu/wQfhvqcpcT7hc8SLBO7sqqXMy8rXixYGTOr8POacXi
DU4CaypYdK051VYsVZPHBveelu54m0FcOwk1CVbDKhSmbkEYQz1n+z+MdOvkOOxmH1mb7YkmNts6
11B4xUhdGTaCJwfnl3gdiZrylUps11aUj7/vds7xv2fE77VvQlxF/6+7RCxtMCeIs3Fh2DSXBNyr
3WWiIOJR8V5K6wYt0gf49l7k/n1hQEnt45Lt5W0tNREDD4+YpjhZmv+1NN6+0MgDwLNJn1P3AkLE
hxwbl8dwf3qWm93s0eWVK29m+Gaw4hSXY4c/dQKPUrqhdo59s8/2x1ySeOijEfDdobEAdEeLQHw9
lgbMcSAwsbBCfaIQMEu/kb+/4bmnDZA+XDB4eOX2z/ztaHi7oJZWsSiE1CDbPc8TIdyfkm0/QlQp
KTilMnEDM7NKksAj5gfpTisY5RTEeb6Iz5tjwZCBQsadepIfHry6FF+/3Zc08B87tRO386zlp9ho
0dasRljRUiqvenrLwLP9FoloJORBn1t4xcrtnhkej9yhZpF7sjkfqK/8H+cYAPIZbwfaFzxLAH7f
RK7r9pV4VBKy0IpHlS4vknJJZaTtdDVtNFUTR6tcf4szsUSWvnLFjA+OcX0leEjhj6gSJTWmHc9t
VcH/wGtkbMSEooQouTVSSDXVUNvmC/zSnjakK0UU6N/ph/+NU9dYOxEGCf4ZHq6ET80QE+ltiXED
hV1AzHRkVxDZZaehw/ScZAoZ9fHB4lSUXYaFPwqIiu55D3ZAh0xMd+vIqz5go/UrBdmfdJ3W5jkA
7sb/SaE6O8Jz1n/h4d5pYlLzse/zW+yh4zgdZmumLYXm6sfyIAs/HYcql7pYVsD6TZbqEWUle8jO
oP6edSdZrsSegKygYF54ohnNvSfQYdJ/pC9uQ0B5EEamig0iKrfRNEsMHWf/jJfTsqnopUCSsnOH
yrBmRoXMbe4TAOs2WSqfUhPR9xyqU52aZv0RMb4VOWvHADMT9oUm4SNdJFeQMVPcHWyaM0oZmEXK
tDylGEvfFRzQb/WmhNLDk32P94xCjApskyrpR1o9SOqlOCN64E/rQiiUfRd8t7csDynXF7FlY4vP
RuQ6886E5lgy3zLBVsYfoy/vfmfZyL88QFev+KQIwTUeBpsLw2p59gZdob5ekIIghO5nH71ksChN
u2DW44wkt3Dvy0/T70MKxwpxmt4kFKrkp2QPsAAHoSYF84qoPeuMFYXrzabsu9qMutGV+yGiY8jZ
w/By+LT0dNuYLsVLCUn6OUv0iJvCcDS0TMUQnuLoTsZJPeATUtCZuE3Lcg5zt4ZrT0M9xGaD9DX5
prWPB1MkAr4pCwLUFQEdHvHYdtL7B5ekTioB9u9oJuJJroFG6/MCu+bmrXQrEtRSUSQgFxAKvVvm
ToCs89QiMPpECvajJZwdcigIHU1V9C9V0jWSre216YPbmhtWPOqBuZcptXB33qVT7h+OrpqEyTWU
UVkj/LI24VQBxPcn4KGesDHCSPbPJDMEI+lgMA1eU6ENPhQP/1CauqAMuP/TbMxPwyCsjeCiGg2l
3EsEuKllyq1LkyW1Ff3UQzy1AIGngpBbCTUYQQuuVQHTY+AlmhW8NeT2MmVnNmb7omrRmklpCJrt
WNV6Nld0/7E67igewfmFj8nbdV2JQeu+YmXpDObMegQdSBCtdPj3OC32EYPGRcPEWo+MpGKDfrZx
oE1zEOPJYuZ0IdjALEwbnRLBTCRMMegDn85FaH+O0WJJkEb+X3cj0r101lzhHVgVVQc9XjitlQpG
v0SjXBmtDFJQB7apK7776kXPQFl5qEJyRXnedopsAvW7Cd0rKIMMQnPobSuX4U0pjFDYQaaNNitF
sexBgZ6g/PnkFK1VQUs6SOhZsL+eOaaiUMwJ3eDbmgzWtq2pAJoZ96VkAAf/qThKvnHTDuiJxJus
h0uhGuqq4qmVeBKoo349S2rZPV54ZVxf5Pdt3vZnGPTx+xpPm/LikRVtoAmn6meRMOLX4YErxDQa
bqi/Utu8R0XQZ4kFs/pHnF7WDjDyznNNZ+aKT1CfIzGqDI6vSGVKegX1cZZxdjvq+qMhf70jgkZc
b9O2AKy+l2EMOzPwxBccQPttUDjTdU8mIC/TkrdncA1KW0vn5SIUZPHtFDFbUF6d8YB2FnMCdqst
pYZIoIS2ATIIsRr1HuxLNT/X1fAd7rxKZYpxIpvIvXKuGoVMnaQe5DIsGEri9uGQ9jzSlCbKZITO
KS+gyvxZB7Tb7sg+fz1pOZxkoAEtf5ur+2JXnzDZdVCI3YwpUnn0BX3pLscG1sbQMeLHGdF8hZNt
3/De/Qkl5d43QW7xVugb4Tz4Gvezsn+iA8VSfzotk93UTPYfR8DN/RhZFVusSLTTGuDO8y9rvCVc
DI2uh6raMhhjh52K0EsYzMYg7mGKtPiygCSUtkkfJ2AcUZKGXKXgN4NUnzVIZooiYkGqNo90AFsn
URnQzvxSuvp6oOlTzB4KQO6sYn1vWUT8f74Jyu1SH0O8pmaeKRRXBHZhclNUAC45373N7RwJFBWU
/w3kAS6n8aNfmYhgiUl0fpdxGKtK0jk7jWkSU8CiYFL9GjK96dAki//u2qk662TRc20Zz5yZ4+ic
XxrTXbeCIV7muqfBcCxcdzEiuYyAB8qmpIHWXvg9idbyjcZAKDX4lVq4Xq5TFW3PR3Pn64kHDZll
Fv60gLlupk5jK656VtxL5N/2voD0fnT4qeIbqHv7C7zw/mI3nrWQ96Dy3Z0Mo/Cjd1TM7Z54nh7d
6e6tOyBLsUyuT+rbunwZAkAFi4KKKxFluISnblOALG/rdf70upfc4TlRHB4EJhbJP6HUhNvyVYaw
E8B2GwBMm6+0hzdF+nJX1Hof1N+BYo11ZphaN0MVKOZNbam+FWbo8MYxfNYffLnQImlrYjkj+Jtf
b1fj+QuTA89poM18IaT+YRkV0Y2HKMS7P94QjMsmtnmhOno4Nrn5RFXIcWQbHt0aTjUY65NOKhmg
VFI9wqYcaAhNAYqH0G+9tXaslodXVe8o1OSachIdWyxEnrD3B/gKh7KymBjOW4fG4mcwvy/UN49P
vKoejM9SPZ77h0CJKBMclbMELIJUYNlO3G2cAhLKpaWNmUgtgnJp2BDAUhAWPpfQTGJXbbSpfLYu
TTVtx8gUX/Z8a9QftyhA90QuziqO+AP/snQ4E5LdTUV/CkIupeKgR8WVPw3Q7xEcKf/bIu4zHI2x
rmmnhIiKWgl6GLDdV4zfuFAN2yNZeA+93sVb8EliykxPWx5gbiTcGxii1+Vu2GB7z9yF7VbyRWz2
MyRGvNIdIzF5Q27GFtichDcKx67wttdWa12j/HMubUHDER/u00Xp4LkPdhGkCY32i+XBv2ayB6fP
N+L+AhqQDGoypBhB9gKHW6ZufqkAYYQRfq0APF5iT7KS7N4fIhrOUIQfMxOoNoDxaCmovauBsGbo
AxTNLecHh2QVE7ZZxEl/eWPSOqy2brKlfsdg0zho6/Tod9wdUV/EOVrTqdxNn/7BGxwsTn3rDUAx
mU3zmfvIvtR4pxVWgo5uqKCJ9LMPWNZBZo/OxmeYlDkfCd7T1LWUTf8MMJpvJMoPj94uypmzPPa4
Xc83z7NCYKUrS+IRs6w41JaQUr6Yu8bzOABhJ7BvEiiRQexzcWBHsfb+hBmkV2AxO21kBYddUV4w
tmtasqqPuzXrILBTQtPVU++gjETfr5jiWvt6/tGRBJFv1Wgi3bOWLZiv0fBoFqD9lj5a3LajNXTJ
diuZLQWGY/rRbZRPQOgQqRsG2k5Gt0fmRnT5th/PT9TBrXcKRwIMd9CXGWb5JnKS9DVXvm0YocIv
9UDq5sndnPk5ZI+79I+UQvCJjU9I+vBVstxE+xPmOVQuYHrWq0ap/fO125brOYEW1iwUL8x9R5OT
eIRhwKfn3S0i5mf7gvvwl8nIIaXBLeRqkYIPbBRWwiezLmUrWsn//Au9ulAgHnlFiqxjAgjkQMFb
qqtXCWMvuuvk0MGd/EXdl5xqSdEeKgnHErh2JNgPEAiPuBFG0ghBSSAIxp//3dDzQyF4qOS7w76e
3MNn2yuNNjIycSGUL76djO+QoiPctXNJXIpz4J9/IyRwhog3qBRDTu8T0fuJn5OOivgvLv8Z29Qb
jJvfMv9VUOmb3W0DvVEU4WOmTZg4OThiFAMP2gxTq5IJ1saWovQxh75IRQAXgvmQMoVVVCJJcETc
91uzmS209e+XAYshUsTZ3/ci4YZ4i4NFPSWeKvmsPuyuz8ScOFCuFs+T4Kizn087lF236l3t6swe
jIE3jQLSYpJ6DO2gOnnpNTVAiGz3ePps0uuUpCms81PozIV1PVVRRBmw+gtPlz8RUTNAv7zJ2ig5
44bJPbUnBJdKJyDM5EhBNNZPClrhxTyARMD3EHdqqAc+MFyDpptbsFOGYChMHQ66oc/cFKqtkOds
25gXsaDqY1kQCdW3LNxuYgJiZgLBybyGxulNrioxUPUQ8X/W1T6EbfPUu9t2keNd3d+aTiATq4v9
Qvp7ewRul+qYLQrCZYuHJpxPmfWtN/HqTb+KEpqv1AcWEWD4ibBDgowNgltANhr/INUUXtHhbXKx
SAYCxPLjav5Q5qyZmmfpC89mJSWHpXf7dW+nMbjlqXWHXeTJSy9lMGKZv5t4ip6J+51LIgu9p7vI
q+MAHUDBghlNB/h5R9wHXeV7LBwhIA8ftaDeRr/kwS6V4N6mnv10+RnXyNBbS9eanRUnJHr3NorT
B43Phhb1oHeYyBgmATIYmo3oODLnN27TCfRbdyoqc0XAeTccFqoVete7eK9qP177x0PHyCFFcdjR
SNSPEXaaxyoDtT55wKAlG+PFUxbMlv6Aag6JUqVTuJ2ZhGAlftf17g5I5VgKPHHXY7zFdgWi8ssC
Vb8+wHwvVEVZrWpq/Qt4j1ZUrnSyzX2w1h7OVhkFit0B/S8qJ6VrDMRUNsjO4dMjAGXAswPKdf0R
V79vSk7imG6IgH5Injg3BNpRuYwWi+SbizKGQSWMI4SyXn1SEoT8i+MgQ0Q+++IXlK2IrY3GC3KO
jTySZbN+BzBhYh0zdqYx4hW/+V2Q/3ueD0LlKlTaGe8010hpRKhW4lfSjaE+u4a/pLQX6VmcinUZ
uiKi+/eaTuWMgfEQstE3MwmWzOWNsNcnOkVwgkzV7TggJFJwF8Uj/8kKZ/tUItqSSqYP+4aoV71s
TIQOj+y5q5VVYbBJucRWxNtR8BCrR4KBV+BpUuGju5IfwtTw1K1HgY+iPorbZurXSv7NjwoZkiUG
DBR5zmwtVZGFKoE2oF/xLAaUgm3U+Hlh9Ft29kVOD85hfU3FTRNSQTGFT+DDdhEugVPNsd/8XaEH
c/DQflaFZf5E3fxm01U23mOS8DEG4esDEWreOirEb/796OrFpp3tQdzYHG9rC07gZkyJFn3UDlmY
QfikxGndtF8Jf3x7wFVAoZINgbKRC4OrfnGyRBDQFqMHHlOPHP0UeBixJKWGVqXWsbfCaAVwGyHS
0KMxqu2NKfG9dovVqIlma8jU8sgzkd2ZBhK7h5/yqH+Q2SXCR7i1Tm9l5pOWtlqEFNCQq32bzSvm
US8GBiUQXs2a7HtyKqFi7gKYpn+LguUWIyrm7R1C56SN9veoOXdN1kAntKWTehpx+VpFvW43JtDU
wstJZUxgm2aGuiXFKIdyOAlwz6V7Iz8axrjZyLsbjYCeHBYAQK6fg6tGFIoSwdhLIqrluLWLBLmB
QbhU4M2izqr+PPyuvdUQraDiVEFqZUO9P44EvYBhUXV2/wLZD9GvXpAsFYjRfBsXKKd3M6/yRD2U
T5+SMiKHsIK+e31RPGmPNmGHztlMIPardg/HqC0j8ho7ENVLV1jFZvlPKL8bC9SnBqULK4nRJCJj
X8xjw0PtkxGukrF6Q38uxI0MTP2K41hQ6eXxp/KdCAZbSjPbWKX9aTlgHZBETi3pUb1L5L+CtMEO
4tzQ0rCfeA2l77yoSu8kPrJAVkG/ERwnnw8wWuuH5BRg6Y/vtB9YDyQn/10Tluk3XU2eWTDqQcjP
Gk7uYYwqCttbJe21aTl0Vk5JxsCknS3VMYRYjUnCxw1xNd7fvus2DTqJjH6jRY+vz/ZB0yJzuJAD
hdG/b/e5NxkD/zPiiHQomBIm3U/g2ZrG05y7d6z/xryqSIX+JAI+I2t+YmqsnUsaI+AjuDv4i404
iIOrHY/dG4vAQHnXaptWQpCa/Qepne+CmSSr3vVj33cxQUsee1UIoPRM0WAB4WUyH+d4TPu6Uzk7
GQ/kbRNcxQxnnM5ofY82iIDwDwKx03FWpc/iuhQ3QXffQnDSVStpKT2e1/ae3Z9SyjRIhnU+szQ9
Dq0Pcs80HT6DSLOFv0q5+Tw+2CpalA6Ls/H1EzqX0ofbI01PMorUZW3VBLO70LYFZdpK4SrZkmg3
lbeU+lTOtAYsjtfm/d6dW/UR5Z9wiGGxArDKR4wVBkYs/S7+2mUsCoVPFwysUQBNXm4iwNiOaGex
Z4UVdKy2PkO0PszAjUmkV25Jrm6AlmDJNSESqeZiarpTiDCtID/ypuZI1ZqXUT9kxevkPPA03eyC
9ypNTk70J0XQ62QfhHfGO143AswyFgYcXZFI1NWLfSUJd0O1E8iNtyuy1U5yAKjlQ4tkKcEby3qe
UneX4TLjv3VfdqPXLk5uxR5fReoJTZkqsV/1LtxpmWjV9LQ8t9PKiDMzLubrtVqDfUHlDbHrg3EK
rUClkAfRb3Vymbjn3RGUCdDcXkPZ2OW9AyCzZdVew/Tgal4rROqfZQVyAQHhZzYxjib2hTjIJZdt
axhuFPTzWLsOMUCaEFxo2JrPmWLxJVCcRriuq97nLYZrNH8pM5EP9yG8n7S/WJcy4kGJC9pkg6R5
wVdxbh6m82qGJVl6n4nLRv5wxbM+EE5+BApef6+LOJDU2St24PocGridqyGZ6rIYYqks+bY0mktq
ZInTkXBTXIKM2JUfpp7WnToeiaqo+8m/m8FaX0ABunw1peWZiYtqe60L7Y3zvS+rCt6szBX4wCG1
4e1Ab8bi/ka3CeC0S1KTAvauSKVqJKKn58ajVQhJkw7CAnARmRH64IKkkK6OeK9ZPRcEyRndCOOD
GZj2J9qz75BB8wCNAp2wfi3B9boD2E9ywd1ZzZJ5UXjsE6WJqYxTp09cEfILrWgaWbiksbRA9+Ed
h1KfOM4qojcomOvR+Tv5LK4LNG1NN0SF0J4ixHy90fTaUR/Xy7cP4fv31A66V3064lqXyamUPYUf
kMxsUwJKD9jlSanfBW9428NhacMnOyN6MKB0b36W6xWaK7zEZ6lGn0huZCk8zKVPActYuHMXoqub
Nw2Bu+dOa+nUSSyVfbYufQQfk29leHaQHelTJqcfiZtvEd6RsyNIBgfyoErq6G4PbwxCq0bzE1fE
/ISc6MWzEvtadrCGqR9axU16c8ADHz+uXJCZ+P/gq9AEhXK6v5mi3SONmVmT3JY0riS33Ofo/xHp
A6poniHRoGViUmsy/xaG5tvH04DmbqYLo4z0wJUe3z3fELfTOjLYujVQtdiDJj2UBZEbgbVEYB51
ZZ8xsS3mamM0ZMMQKViT0DtEW8OECNMKwSDYsrZK2yQzgS2qBFvRVD5KOwU81l6tXvvgtxE4e5iX
VDeKR3BUtzIRI5VwK3PCV7uumTUIs8FHrRIYNuQslfBl0nyB5ccOl3kh1D5/loz766K/1E+qDW4z
kbSU1BaVZaKF+tMU+81mRtrYYdp8sPbv/2Tgahf+1v3zvVWPK50V1iRLibo+J6U+GkQj4RNd1gHg
anJPRggoN/4zs3b+I6fTbsOZ7xheQWUNF8bgEHfJpx0uNJt73InMA/e5b1eBgVFYutCVpVjoVsvq
E+jMuQl4pkmRe2vOJVuwx+sHRgm6S9Rzv6BEx85nlgTIQ3dTgWSGlCWfPs3VyK/GlwiApvc19LNl
skZ9iuAeV+AN8ZiOWnd7QZLDw3O65qEMLoIxa89C8GjWgp/eXzT826oCw8JguE0C74xHKmjfGwtj
6twqn5QGZZ2hQrc1B+E8+bbCv+BUnzJjs1k/JIT89C9o+xh4Ni7XwAkPNwJ/GtgbWl1PiZdOKXIY
OYGmkf4TjrZIJoafnV8JsOua+ku8mdzwKt+FzvV33sVEp5dKK97Pj6Yh1l6UGO9z13ZyVMvBk3Ff
p5ai1hHOmH2wxFDf8RHl5yGz9XpHmXxKJ2F3v0KTDWgKyQZbwUHtjnaWAzBNh/D6Y3YLDuAaZOEQ
VD971X+EGKj7woKeoXrs76QStTu6gXJf6PyO+FDvFUrLGGbHNPCgRdChXvWuhYG3yf7yIaYqHGR2
ogAmar+Id3Eub74Np+c++pjyfG0HTguM9VhaClBrc9+8pb/mjbsowlZAPYZJHyM6jHkq5smfK8GD
+VE02039yK+dY3S1dfZBSnu+tohGBn4tQgxgi++WmqEbza4M0CDs9PQNlCNHsTv11inpj7tLcOuU
gOsQgQ0l/8r0U6Xs4HU30VFibADJ6YFdjJp90Xc4e5uSixd7+UUeUlWBdn7IFUkh7rXxFdgjazWe
6MLnmdwtgl8oTlUvgZ+X5jG9cpntpPO9z/4EJ3xM7fj7OEI9bDivSQfjfSZf5lnFBn+woGxiwaFX
YytPfcIdSFEkvNbGE/LB82jlUebPpX/utqlnZNLmbFgK19TtIPuvP4A0birUn3F0Z7havsYbpbjf
iXAxX2Nq1+H3eVrTThbmuq/fJmDtkYAedRHw0r3cVjCdZKEV3BkJlMgqncrYRlagqU4tzx+AOyrB
/gE+a/Jx8gR3eMM+x76MUPZQoilqw0YAqf4RmZGIsUT+UV5vDtQDjaMzL5RVGZjGnCi16tKuYSgn
S42I0rzuAEsRmCKmTIUMXuiT9GaMPsz6h+T/XdFkU+1Bu6jIKxukZhGCuPBooJdnEOnQGCoq09Ys
dLMktcFEP8xKGgz93kLUvhTsuXDcV5xxej6QkGLsDhoYEtRQKtm9Ex2exe1bwARTJV0OYov0DRi+
YioRh795fUdRAIWAiaL5HNB/x5d/YnHIUbKDmPNFb8Vw8FeCgUn1DTpZMFMWdfC2augE8gzh/x//
2RtGcp0=
`pragma protect end_protected

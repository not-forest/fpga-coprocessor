// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
o7c3vBz2ow1ajclqyiIlZnOoYckihq0Io8/ryljReKrczrq7CsIUvCJELpscu9np
0+JBjB7E+UHHgvOjIbzzm7KkOeSyk4Z4WpBgQS+IGBzZ4Q+Zq3HtU+b8FN+LL9wV
xQjtaCsAEL0aNXehdN8LwTkob6u8jUsri1l180byrzhgBMozFQZePoyGJiHw7U1D
eu61I1djsJwphMSV3oHButDPoi08GA36t2teBTqwfEabOtzyt3NzYrTIXkjRYwYN
LrG2InYK7Hsf71AJ/lriyEG0DsvwEvBCC5i8EoPL7HRzMa5sR4Kmx6B1WqvPzLb6
aho0rxryGnZlQR8D7DJZzQ==
//pragma protect end_key_block
//pragma protect digest_block
QEMY5TE63rT6aLBSC/iMPieyu1A=
//pragma protect end_digest_block
//pragma protect data_block
EMZopa8D7WEdfeTCaIL+fgHwRXByWd4jcrc7NxjaClXe5MLWBaPdPnHxDkA5yOq5
72n1no4AOVJn18+GWOaj5naoC5taWKfUlXmwqgCYWWhRwiNhqP3tRokdISBanLZF
OPxqFO5t1bJVi9VHFUGUBYEG+7bo16CBwObJiwwWvAQall++vs8XJjGZT4QD01jB
a7U6+hxBZ0nmqqKF15QngoFofPD+QSBGxBq82vl1b4bgTRyOJCcZltCo/r/DiKUP
NZ4p1JJddl+1ZkU825Kde9yWkBeT7jzNIandnvyTR47PtdierAp+MuEIaKnwuhzC
bJoUT4s+2wba0cB9ItI98I7+8Jhv0KpACZIkozRJBkxoKTLFQE7Eu73TczOeZQnX
b5WSTiRpXWlKKbIiWiUD6URf8/oOS0XGWNGyRurUhvWLJ1Voe0Hg4L2sb4XZIFTN
4KdT/E2qA4+0FHyZvbut3QomeZV9u4ohHCB7orFGckeB3Z/WF/dFu0z9PaAPlfFc
rdCxLhl8gm7JnYSqY2Ii24v85viOHAVSBh4JKM14z4zl24HtI/vrAmse9HWZH7r+
WiiOotRvMXLZiVou/t1VMZec2FAuSVdhMnWNyDQb83MklPfMglY0qJ3uAJAtC43T
yPHH19yN9pAlRgj7hYUBplLRby1koJpL3WWgviIvC1Lqsew0QC2UdZgNPnBtodlt
a6ZY2bc8G+/CZ2gcg27ITlPYt3xxGOA3ZA/XnPd8zkZSvd6mfuvB58n90V5M0nGF
YV/Yrk6JaYi3+8BfrWd7Rj8ZmoZ5hAR5QVB1JyPoQpg6KzisAAj/9DUnlTDcz2ud
K6RH+PV4KgEnevZnk0U+njyc4SuohP0cljEjc44K2HfUfJxqb0y/kvNNN9ZQG3ed
GZil7hKX3vaBKFkHNHKq8p2x4r4PiLLu9nl+Dmfg66uXBLduaYyD7X7qlDpKBqQt
NHOHVUE39EmdgenkvkTC+87uAYBPoyLqeKOXlg7kRfvx1zT/N8nIVqWDbYxIdvuH
6IXKYg5ptCjAd7rMFUYcoLI9FtpOoW4wqZ8Yb9R0Plt860i/oVH9NIbZQlp76ezN
6A4J2I4RbqAT/Sp3HsOVoarW3Iwo9VUFrfcSU3GChKMhlKNwaw8UH1ZaXovSsGSF
Uutofnwk8IbZ80pParTHlYorRS1ULzrh0ODliVi7LK4nW8kRrZhK6u0D8Pl20u3Y
Lv0Dvjms6KMPEF22kUBUxWkc8P2DtpJ41g4eeZ/CKlLTBb+tw7Yo53yIh3KmqeCF
jxZAQ0OAmnum6fjuZWJWtn6DKpMs19g5nCTHdq59mkZ32IP4+jkDB0cYTT9JXyzH
0YiSsg0P3X9THvM00DBBq5jWI9ubLIZMncoWfCoNKt6FR696xk3MLVDzF/8DiSsP
4x5i5FO3t5SLKGA9YkAAVuqFQC54BUl7ggVarukGdcReXI4Iu1pg0ABHuWLfQXBk
gQolmbVhYWZqfR+IIqtVtOVPnwxjkhxpj+QMWYY9ziSt2UOfnLQf00+txYBcmAq5
u2ejsJCGd5rdHZ3tLzKfCym3vuPWLr08sumhjqnBuTdbUNlr8/pZdJNX1YEW8qk4
YFWLkjaP0HpQUY2OfczMrj+kCNm8mMOEtDUCgQOvuvlehKhL2H2Xz3+NoBlOOqtG
hL4HLnKuo8neu8kW7NoS6/2QFVbxT5zhkjF92V8Wykc+wxl1RNPtp+3ygyHV9Kkd
JNd+d6NfxuW8zWhgmwt+pkcukP2Es+dqRBeNsQQohcZ+E50mkMiIyHOsybjRVhNj
PAbPLqe5SyvF70shfs/6MJHGZilMJqILru5XRHpiMhloYrh3X1g/p0oIXkLY/mvb
1IxF6ODHo6EYRjD1TVbpd8A5Qeey/ih5B7o5UdM9QhSb9ZbnSDU0Hdijyfc1NXrY
LZZzsyKrgVgJRTVDznInG0UjYy2AJ9mPAAqpgp14glQU0RozGwAWrSZTPa0T1NvJ
SIwZTWCIzyVDtlRNCfpIVKVMTDv2E+0wTuUH4dmNH7K1Zr7m3UjWX+gY3HL+/XvT
hnhCAGDGDupwKZmeFJcAvl6QEgwUw5iaE02h/87O/hPkjSLmGUmhHhlmDj4KVoZw
v24wIU8f+Ci7jIg7PetnxMvIecgmeR/XoteHQPZtg+GOvG4wGwOlwpSxc17XTd1E
pV7iC+/ScfJQNLxx0JssnGmCRkUkAJ00nH/PflJND2HyMAefaTA8RWlxDgmVa3C/
nFVObcTtLoU0ayBQ2mqycAgrw3h8WUhE/IMFUoiOBQmNVg+44ecYmTnJzdlV5q1q
aLuNmnXwuwVp3Gky4qFuh4M4RadBnyCwwONowLgekocwZXUnOdHOaubTqlsOlr9G
aCDnuaG5+b8XQ9elRVHUJdmaiZp9sp7U7tBmaTeATjJE/8i0MX64ijX9cZhpVqPN
7JcRBuV6QLrVVekyTIjrxNOQnX3ksAOrdrfIGcLH3AK1ywpbnZTjS/sD3OupkA4f
x/stlJdB5t27yyTbghS2YkwKi964MqeKPtJSGI3ctM6M6J+GuPUDp003I+IqNyBg
+BOOt+E5TX0mW1/TXfFDoEJ2D5elw9hX4tkswv8LumNb2a2NEESDpz0of4Or20gH
gS+Rt7aW2JHt+/D8gd+vVghMcRpNxgwGYYeZd4q13SUg/rHPpSbuCDbDzsrUENbS
EtubKnL+ihOPJZ9h9sdG12GUbfyCwJNiL2ISRd9RA3XWFPpcmL2qYZDxc4ZKpgQQ
gqBylUN/9kSGCox680j9McN566yiWpYrjWzqmYM7Qpg+UjRY5D1oG06ekCgXQtF5
joyDcR08HRKyA6cIqjZ0XU/abTSgYRWLj2WrCPQQnQMivMzVOr16g/OzoyJhdLzh
jy73td03Z9HTpLtH/wTy8mnoJv3XlQtyaAs8b/CJD9qgPxrg+5ZANnh4f0hJHJJf
0TbmJ4XmNyBVsDKu/HGnAh0TxoucolNei5juwxwN6c0d91TArtqJmZE3D1rluSAC
sstazgPjS02EWyuYlLIiKSGf6BsIetLay1bQMszIxb9nN+RYdbJoQESvI34SnNlD
24LRL7eBbyyIBLEEk39YBJhtqldg5xc3ePN/LYJ1JOKx3r6OwX8ygHTDQE1cKYJ5
N1MJEfRRoGvAveogLj6vTg5+m/QygMH99p5YHpv+9pY1PQHB3Oe85RDYJHt04AF0
uC2eU+pCdzbhFHmvLFFAYW2DDf9CJHSoAU+GWe6DB6FW0pNHCN4EQoMU+gq29OHD
krlmd2KwAeRDgz6Wrf73YMjH2d3rhmuApa3Kr0m820+A4myoMtKH0IBzvtj2HFlo
c6XxVrCrfETuaPBdNRkqs9bkV+qUuDtBmQVvxHuPAQ5hQYT38aWQhrnVNnoSbdhZ
xPvtFQTdVGrniVyxlBCZQJrGgwChLbb9T5MBlaU0+C68rZY87gzrifhrq6VMFzg6
pW8n1GvQV38Zj7Kw2ifaS0WlAKRxHwHd1PpGCE01TlJhbC39NtIJuvWqW+FSavcO
bAyK6X+VZ/Z5Y1/1ONsbA+jitqlnmz9cOkVSNzAOlMGs107Ccno86+p6T3zqWuZm
uDBFDxP041FtFy/vRxIlWwx8rdR4+0l/afo7OUj+pNYkX+NpUWsxPfKbryQH/0/u
Tc3oMIferdNQIirXr1S+sRy5gpTG0LZNr8o+OJa+bcW0v0lZhn9eyKTD9WYqyVQu
eCL6KYpGL0Ckq3axlyupHpe9HNaPmI/AtbEn2KHn3G2qpo48DaquCBKJixu02g9f
bnHrQGE8s1vD+aSJfY02DB8eWDwdPAN6y2KUX4iS9SIibhuKAuZCWLX3DjvcSRMm
jOyn9+fiiPVgNs9eohN82RgMX52elS2b40AfNdOQFm2soSOZ8GgsMp5B4ff5+jKr
Bkd5q+sLjhYrYfZDmXC9kqhio25zEXVPmn2yZkmv+o997x/CIwJlOxpmDhwiKpyI
DRWuNKuxrror7XvYiLv50PesK4BQW2MtPA8RguGLvV9xRM1QLsSzc1v14CRnvnrx
/P4nWxdTId6xafD2D5RX2QJW9B28gL8NZBqsG/ExoPUYUif7fO2syEcft9EabsnS
JHqZeox4BgBDtz0R3RzgUYwo5SkmFoQRjd1sLClMBhuj+LF0LhMuJ+SPfR4daw59
RAjXutG7k+GkiQg71FZ+l5ct3sYivVwxrevA+FCTXIRY3R6zYZvYsEtKbbI9DgIY
4VQmbo/pGDZItfqfpTeqt0sTqFEbcteDEWro7sOcRVGxBv1qGa6udYUp/0cybOZZ
Uz47TlgVMfFlCHdiRRgfZKC1QMv9V1CxYCP6aJ1q1j4mDZEFz6VmMrmage3OctOS
OPCSxipXrJe3KX2ZhPfIfUsCZRQE4huzoJ0zCeFpOlQ/a0OTmJ2dmlBSTpmUnAO9
0dlUblvRbRQkfOflZhak6EOmWZSzSK2VpzmLJTK3jEvfvOKuJRNex4m1NwxMjCDk
RwxyqsipSSZCm+jeSqTswiKQuBovGHTFVOEM5tNQiSFfh6qIRkJ9d+zcQ+xgeg4R
bAHeI/L3zLEkaJCVRjNkBHzbGZKwP0jw0Lw0TqEG7QLy7b9QLJN8pXp66ahfJcmD
t3gA+Z46FviJGfXRe2nmR26whNgiN6fyQd2ygmEKVNscfds5QvSO86HLV+k2ON3p
MexQmwlDzXZss4Yv1RKlE5B3+bJ/zYj0T94P4vgt5+HpHrA4xoZPQrrH/na5xncR
lLPiGpHaAXoqxa99rGVJmZlbmRzVF4ppEBTKntj1OktL+GYPEqb+NNEF29PDGmIX
ulT4n1hgcC7PhNsWtQKkG9LAmTHIF1/NWwlbBp1G4SjaEdOWRWMgec8musWIaXQV
OHIqKK71NaFO3nrt0b+2eoxoB86KuB2K/QEIrQoTVZZwLlpIK1DOP7QvRjiYS3sO
ZvfmvNQG1Q105mCKt3Bn912RwzlpnsUvTIcEtkvmFcyGZ6P2EUvbXhNYFtk6hUcj
XTpB/RcuX4lJSjxSGS7E63rN5sAy12yj1e+ADUXketz/hDszYGhYv79+GEMgBsGd
bUz1Qm8uOx8CxFTCrchXbAY97ORp36SIcKOJ9Q4u6g52lUyL59Btm8yabeg227E0
DOKZbPk4dqTcDyhtUQ8Oa38SdYilm0xq5pkKA2oojBixqgjLDX5VQW+v89FJOY8g
/RnwY5mZPvJ9DrXDvSViBdPPTKjXAvzsw/r3eZrSf+PEPoiQzzKIFX63tHoBFG1E
BlCFFZ8z4/7t5Q6MktR44mz1ugbDZX0ropM1suID0d/KI51Mc0CbNlc3qEAb2Ws3
HO6fx4JUt7Y/9fwWEo2P2QRYkuoThPSvrxQMR9gDLsdZ07zv2kBmg3kdpN5hO/H2
nYxBz8ZqfISGde4osXmPOQMfqjyJH6YGKYAadqKe0Crk9NscJoet0+MMXL8emRAl
Pb5RNsl7F/kA56yPihY7gKWSkwpgnEo3yHG8mJ/ydFP4L+veYvKLhdjBLbnO2ZL/
ZfMg7cARlaLRaSlWu1C/2Yzv9xM2Km7UZKhsngSB8YcUDV2An70g3ol8rY3bHbpd
AI6MzgY8fBfrgAxsoM+uPFbDmc8zwKZSUJnAdF71VPHwzzUbNDnxmQCJpXP3JMCz
2jMDo3+6iuzojH4HyKN22284f+8DYyXsLB86T0Qzs17u9ij3D0XH3lA09Nc4g4Yg
imjStT74RPntj15vTjkvTqV+1Q1cXwK7NZGL+m9g28nayxovssumFSL328oVHT3o
8wl0yo5g4tkld3scV4gzzmEH0uxUy98E60yPmLcWoJX7PBnXbFaPcNGCVQGql+ad
Dwbl1aIaWzCkzOEqjADwh4ZZbBSnWdYslcm56lboArVjlAz7F8KYf1diu6ZFdPN6
yhtIpw4H+TWqIKdmK/7R9dzspxpBWFbh02wWcJssj+73Q9qW8IXuuGpwOmxcNQ0Z
4BXPJHDjvIWSrQC0klFP1zOFDBq3nHBc5P17W4PxAf5VbZ3+05hjHT0bInlbYXpf
GurVdBdZiGOUBOIF71bhKTYaNlKqOTYMWvShMt8MXfmDSyXx8n/6JNmLQIAx9ReZ
l6qWQftSmguRBckQaxb8LxY/pzBMPNjpaCic6hl4Cl0SNXrbUql/Cfw+t8XeU2Nz
H3M0VjI2ze6MRigfqRkYRDkCAYQRUoyJv91JasknPGOEDrbLQenTr3J/MmEed2dU
FJxoGjmJCPTCBJ7H48v8qXodrpd2j8HdwTA5Rwg+dJg7KVArqJ8k1yNQi+CeV1Un
UAy3csaehbC/ZgUlawK5EQeklWhnJNCcZO2sHwRG4cBWrn6MaxE7yZEt1pVTlkdj
7c6d/WacwIrJ2g1CdDNpZTSmZmQk26/uo0PT7WGLuuwJO2Js6/d2O+D9IJI7ZscM
crTt6mzPopmtkZpUj2v6klzAIbemyyFOIsbyQcOXWnyMpw57e6DMCgzNAB8XGae+
nEkjDWcyHCJAvNFZIEsxL11VNnvFpKHrXzXsN/PyjLvAF4Li7OKevbYtuTNTSb3a
XBJm/RVFiBc8tmMm2TkhNknmzhec2FHEkLgsMMiXFLnoasMDqEBAoOQjZjW16r1X
3oZi6Wf4/NKSkVELgp5n1RVo7S0yX0ZyKcfzB7nUljPNoPh5tvzvq4ycaJyzLUSM
M0WWImirpG2cK+9Ds8Tt19z6MB5z4yNzylXMUDpEYHQ2fptxuvoRfQi5EKrul54J
EqmmG/E4VcJErgtSri8yg5BhhfFk9Qa6EgDWbLLPwdMZA4trdoVW3apfnzN/6DAn
cO0Qkojt/ubgTa/VIzOMpFH6f3F+oBhgMN/pziymTKg2l3Fyohmrag8930r6WtHf
0xdctdUtHBnjX0UcJL0anZV0x1pbGMx8mZ7lNmuUUltnhukH6cbvAcxljD2vsF4F
QT0P7f2VFk/PTGZczTZ/QaSP5ZxtcDSTrDjwYLt8CQ/hY+uTyVxZtfACjO9gaMN5
ZGCDZmC4DDATpyoKz1dG7f1B8aZzROK5nWRjpWUav7KmFeMETKOZPSaK4Hzc0/Yr
Oqb86EsYWN4gDV5EUg3imu0ycrPOJjzGLAZNN4LxRweEzoIA4+eJZey7IbZNLGhS
V5O7w1nBrUvTP0sP/giiGfl/RoCpiq/6wRdlP1J11pdmrkIaBOnx/q6H1mY5xQFK
C+uaLdkzXaMuZYcnlmrXQKJJ/GuTqxWH6rp7jKg3xpKFBiNrfauvwhXuJQ+wBDI9
y6hJwcYLhymz+bsjzvdpEdULsziYpyT7NMoSFmEl2LyWsJ4y179Ckgkya9r8jKRp
GS/gLzX9jMc44bJ+AwlFRyLc7q2yd36PKOffSRdx9o/CCS/U/7Iylg7YFmNHyO+G
FtjdZBGOxkqERvSHPCQ9o9I1glT52ZoMvUtdICw2gvoMfmCRoMdRNVcALJvecvI2
2/B2Pg/71a6VlutF5uTeaEeU3HXwEY5ObGBQY8uJAKz92B7WOvYeqlAk0LuagOgh
ypqtfqtXPghk0w7kp6xznyYVJpLOXiCuL5J5yfFmJ++lyVdtjvx3XJFC/I6pf9SZ
1nePjs9cG8748FAQrl0r6U7Lt8y/CO2xGa9ngz90JyF9hmJfIjtzIWyA/qaJhA2H
KSnfOcWIXk14mBFZEscTZoiloS7wLx6ZF7Q7myv+ipGtSLC2oO1mY6hEn/+US5RP
X/rVVIEtcjf7b9zfMBH/eCEawcqIF9JTewwa1gYge9+bJLSjv6QjodVeT565W9Lu
UR5ZyvhpqJLYHF6wopagEB27oa3rmUVbAS5sin3N9rZXxSd/Xq1RosKZRzdXxJ6T
Alz3iKurqVWLOGR78xH11M6/F6NJ+vsWbNU8Alh0WHJYKQ7F0AbHku/zbAiAr7oN
XbfgNoqQ1RoJQi03YYCzboQ5qRbSgPz7W1z16aF4C9FuTAHfMZfaxHw774DUgljT
3EB1OdG0+QSUnZY0qjuDJWDQ+Vdkbxn1f5gT+aiz2zkTfmASEn54vZ9Aetov9z1N
ePgoBC8BpbnGMT+Tw92N5TJQ7O7P9oqsusqXG4oRTj8ZiQBjXUvswWnQJbZwCCIn
Sp7RwZhk56QESkrVI4JSOGMADLfVAcO0hSngKwkJnJ3CpzKqTNXUl9ZmCxleabfA
fyt3zzsQyVNWEPB0RAu1ZG1tKZxLgiyLsF59Zl3uE3OwwKaP4N0dleuq+5TIe7Gb
C1/aUtPlZNZkLUp8iQyBdliQbTOGypFtXVd+X49PkmkyzkaDnn14sgnKmOeS/vs5
hw53PvgTKqbsvRwBcar/KgM/I5R4GlFAgjX8PLFKALaz18AS/TmkZnb6Zbz7igmm
JO+ZIcm1s5ETznX19BDPYG4+ECmHUeRSiL4iqpjOu+naktYVqYnzaCAqdUr3SUq7
ebgbyYeY6nnMuXFu2NE1u1w2/UKPXUK/8O7i8chWtC8hwDizjoEWQGQ8Aawu2iFY
Fe6mpiYIsmA90vMP8a0cMP+aXwzK7XiF6y1MZJMSNDxY9c/yNBXyRwHqnKUrrr0q
nIbETnbnXiNgUlEvSc50ocbkNH+GCRh/qIk0pIWCTuz5Tl94ohBPZMCR57YepbRT
jF3UlPFfUXY9oSMUPEUpQ1jPIXlfHqD+3sz6tWApQP9yGqbS2BVodzihEVPtkVTU
UCZ8G0sZjv2Lv2qBRdiXljZ6xM5O8LDZx0puYQIOnQQM4zNIBWeo/HRfqdu5t8l/
QY9EOyLn+6rAFl+tgv5UkTCX/71JLTYSYZEVgoOonjgVfpHMWGB+jKmu62nlMiz0
J85lm+zEMM0Wp5IA/CXoZ/252jvurkRFguvuu/QNF3DU/Q0ATl8yAs9F0LQO/gPh
rs+Sed1ykUs8R5GvdBRMHj7XGmtyCqVFdnCIqCSko9bHPz4LCopJO/41McT/cw1w
+tqxdfpcl2XULC+ARZQTx+03Ipgrh7SoCaMb6vWvipIEZRP2PR5d0hsRESZOfMxj
ybFq3fSaXQ1hyvNqf8NRRKcUPIa+qhXdPmrplr+DxNKXxCZryz55rb8n2AsvJP4c
P+W5MS7K7yEWPnWaw/Ei03gi1iG25GD20/QpYhu/HkdyeDD7LDkT5CnZF4uec+x4
BkQbRxYlUCHeJ4qE+IlHRUfBqj0KMXvUooZSU20FS3vuPGrO1EqhYGXA4TVZyKeU
YPZBE7u78QQ48c/xdR8l52qCVDnEJMGl+gT0si/DW3WynPLWDUEMA/oXAmy3/b/T
vAe/+VM7WNo8JG7OAJVMWpKOsDsRsUl1RE21FaAcS70uKR6iaigyIrA2Ca+NcPd0
QZXlSlkgo2wJwB+oaSwGACw8xCN9/qP8lm+I0xDRDn3ul/HvB2Fj97k7Adzwe7o+
8YcT1LpOdWEYVVPZAFTFlx1uBEtOeJzsCiMp+D7qlowF9l3+xQkb6twLOLmgml7/
Y6ZYZ4h/Vx7oTtz4VRNZjtt3/9dxx26fAJMSsDVt/zaIECxti4a2ADWe8Ph+yeWP
7fWJSNBEzqgKYEAfEmxMzqWHxVcK4thyx/LUlMBeQw0zdGpXYN/0K/KQcOYj0hJO
/CFnGzw7qQYa7a9G68Lfut4fHn9/cIU1hOraxisUBLq4yvVladijZ7pQYi/M5lpU
V3+furaBc/gGslXX3T6USmbyXyqpszAQFix5vwg1B/MtbL3fWdtKJKkTMkp1Iuwb
2bvDOOWgar4nNBvgBqKbuhssg5f1HBuSGlt86ZHRvSv9iDrkhHKT/YFYUlDQqB4M
8Wn15XYia7Co2RjJelaXRHPvwQtQfmykkwwpU/0QstZHo8F1Ez8SdNIe9Qi+6n4E
UWSxYl4XY1lXOsGMSVPcmhH5gjJSSEGk6P9SkL5sZUSuvudc8RNXoanGQLWOtQTh
kPwjtGP1S/PEcEuGBwCRjkwKYsSbaD11S18RsdVnmuRJ6Wa4P9jY4GaUyP6wKQrP
vL2nH7/D/bAjTArJ7FXfKcm44UfRN7qA1AiNi/vq8P/ov9YdKkgD9wNwO4Wihcye
8vJPQxMUPX5/sI8duikCgaTyCs3pbMjPy5/sW5nJJBnapYkCX/ISBQUEqfr5RYnb
R8opfUKnVQvYq6kFDnDFXD/BC4FDoaX0d63CIa478U747RrMbMUqhLiLlA0xaFZq
eAhGl7QJAkU3oDwv4PNJdaqJD86wte32d4ZatHBnHoxeaTQb17Gz+ZIy2OyXnIYH
VWp0qcFLgSFTWzkiILWdRuqgQFS2fcxWi6aFWtaa5upQBYswTr7Y5Cquj6gmnLws
dLBxZCzAnPrjy0T7I0+nTNXHaFl6s8J/6r0gG+l0wKGbbM8IyotU6Pudv8om6vfA
Luv2JkBv2QZ3+sMda5mRd1xN0uqjH3WAU/pc0/2ebTA6hC3vO86mhy6i+bWfvHVT
meV8HZwHDV1J2C6w1xnoKCXHZX8DXEAr6UOY3IZf7nbTh4XSzVSfO/xYxb6xhPBS
b3+4N56PyS0KVeQugSNTRkLlONuyT/YbEW1V7nH/dFWfyHDyLzQpzqjPgrPqXrwP
npHgxhpLLWiFz7a6Z2anot85Tt0qieZd+sM/eIAj3rnlEtrvATJ8w7VY5qNcLXjt
x2wezUzHxyt3LuM5t5OEpUCuXGvPI5f1CT/OsUyzChADxTOCk+fCZ97TCnTEZGRT
5efi1AsmlkPlK8Rtr8fSgI9I+sSW70T15wMgl9inX6Uq+yhfoFKcl2PfikCUYwKr
qM0/u8NhJ1WNCkvo4eBJlVgw5MOfwgnkdus2sasoTycbMj8UBZ12W6qxEyJF1Csd
8FaU585mBibW/lAmvas6gheku7PdWAEAD6hPiFAHHG1bxKEZPMkMB9lj/iPsaY20
sCYWvjAkWrPK0wA0yY+Lspm+412Jp16aG7zsCCuUeItOwSw0puN10CCEB6/yxTaX
BK4ZN36iEp+kfRzfhrBQmh2kmUOREHaT6B1zpsZC5nlgwiAIjH3RyEszNYgifdJI
1eTjzzKm6QVfIE5OUfenvMiXHiu8iUsqohVo0LbFPmzgWD7C8gPMk5tP2FFnYpDf
t/2YMNPF/3hWJfCA8y6VZxnTOACVR2gK5msYoyHYFysTzML3bq/kIOm629T9fXrf
gQAKwtGMNW7uN/WRFDJb1z9GMxGdcaUkjNLevrQnglsKiFXj+DVHyCbQUDqMuFD2
YwmPZ08aHmXTe6YpQ6J4FOEPkjJEuiLUhdHWzdCtPxb0n/spcwFl4bH90UuShZwd
zroTkWamB68DM4E0yEedJL1ZsIijsoVIKMGNjTuaSarNBRbss3fBAEJjn7anEbHd
PqvUsQQvhRC87XdLtCw089gHYIe6js6H/BKV2CFz6BcivnS/53t4+1dQYNzikIlM
ixaNU1YLEtXFSiqp629vxrA2/KC1hM/ndE1W4eixoNRbfR1TkqoBB3xuPp2ICSpS
GTuI+FUvUxxMwfPJp0VyM/Fe4RarUW82RxJYQbqNbrfGU00DpurZtiOu4K7EiH5C
wM9Yomi2KNklHmQi1ECrXcO/O+8HhJBZvaPA6bOWLMFX3rkyJhxm02mXz4OfDaTr
6I2yalSdcln1ywoVBmTALp7Gqa1XH6hlbYwkt4TLsFe+KJWK5hVYY2FRWKTA6Tcw
2qZNwmKoIP2tJggxrSjekICbgaDkTc+mo3K+KzyB6UA3wpY6hWevb/ea79pl3QUo
/QuihczuPICPTyjtL2OK3lVXFaOSZhikUmbdMB+a75Vk0oVwDgYN6OHyrL09GzKc
3E+3c+5NO6reCoat6meNJOI5nAb82hYlaUXAiGZrh2WuWOzkO0LPGTkjxqHItQk9
V763CEXk2A65dxjFGonVodVJTJlt0zwKc7a+9k6l92Dkin7voxgHFOXUVYX0NKZV
upbm8mr5AcahGA1T6FslU7zKC3qIDjZ07LhVCuQe6OmPRoLcg2DtSQL7OmeVRZ8P
K7cvj+25GNDSshJJnmbjeJDPkYNI0TjY32rzAUbZQDC+y/V6C8np8lz9sx/unhSQ
NcGav5jIwS7ge+n4dWtchojZ2daNlULeQTGd6ujn3u/CkoANhqxVyuWG7U/pKmr6
yMU8jH5Nl94+DySBWFQEra9PpX0i6+XWP2C/qa1BZ9PAgb60QE56DrKu9jiFflMF
ykX2tIuLAhJsB6DxVpZFi0ZdTY8IbabOKbz0KZgixfrD8rGc1fA3jrg1+bOfPW8A
rnylgVK+VIK5ZDJ/P7drthUMUaipDuHq82KMHJYu5YuL7Y18Q/zfROK3nt2NnweR
IJWaoi9YuwtdccxlIiKcq3DygenUeNL8Ejadxt4+DTBpbZzWUmd1FeFA0/KyqU//
j+se3mQUgW0hZ+MZ9BoT9Rg6oLPaGbhUF451JD+dwEIRq9iMzBNvBoSRTvcGDalV
ulhA4PE2YR5PB4IPVF0NTGWLnggYK5mn8yEqTEmhfG65iciABw2/PyRNIJvaGOEQ
XDVgg01yNB8bRXP9NDt55mNFB3S3TojWW4jYqmXtHDDkUA7EOFiK+ta/dNLuUp1M
xucgCoCy5zaXI43ANKsjz6Cf1wDOUQRjFsR3704WAQj0DAuscisq5i5Ilte4Bw7J
hQnxGy8fc6tggEs4uQWge1cJi9rClWYE6s5QgC15RoOQV8YAEowOchTAaePragbO
EEI22wadVqp/sajXn1uwlsL7I0Tgr+RuNvLGIaV2+bkmXRpCwmduMeAThGV7foHU
17dzqEhagvmzfxwSQkuRERcBfxn41JJ3WzkYbFg4kjaK+p8t5ypeOSWgiZziY0f/
ufAgmyBM9ExCzkn6okWJEr06SnUGL269jwGn50xWz4aKUqHdXjFAc8LcC8KnFAO9
lU3j7muwkx7Dtjg4sJrGMcb+onCdemR/fMsB9U8+4aRCLAzw5wECKN+TZ8oRZEDw
GpMMdZ426ys7ol5JLIpLQN+VUJkWPLaEttBKvHF3Gk+5cyEuQGrJsS/AV7VXKjae
U7FY8yLzlihRm+MTx1nd8dCKHudnYgD3kOAYRdTI2lFuOQkjuNaJ4F53FAvTatgi
e9OaQt1B9kmCEph926mSnR52/L5j105riCCCZa/WNySyPK4uPnMQ4AgW+IDMkPi8
1AdApqGDLmmdeSCSloLrimu0aUY+aF1oGfUYnezz3BGLtqEBSOOnMC4Y3XzTAvqg
omy21XlKDleInvT7/Xu9V8yyTEwnYxEgGL9OGlUJSa5l5NuOJHxBTbGBsSDul/ws
5K4oblzQeJ3PYuOeiBhOGuF87PbtPzoxxhjZ5pSFAZf3V3eq/dPLL20HeCanTeg8
ZZOmiydc6wgEtLke0Z0uOJjJbr032KWFHirZ+lvHMLtX3X45gHxjSlQFc5OtYUqQ
qMdUfDIRxD4p9MOBBuZXOIkgUur/RK86xrFT+Jn++C9Nwf1D/4cJPZikNvt5UC+u
CXsbj65kvmaGXHQCla/KJUEe67gyW74MuOK2NfT+iNDFHjWxW0Kk42/9SS0Z7vMm
4Wq1L/PgYbpMff9IPudjHheVhFo8VEeQOAcfyus7voZSNllqKrc92wF6d380QrO5
pw36ZTcWwAIK2yhh34UNIZ3QSi3VGtfti6nDQ/jpqKAWxjwOSb+UN2WNAC+1sqGh
fV6sLaMJQjU1tDdQDEmpCEbDLhcOeKi+HXNtg9sbabXqpcq71QnouB6ntWoXkZCa
68GP6TeU2MXY7hfwIHe901zxQf5EoUIHuK1tg9CiuuYY67Q+c+5WlJHGRIVMTCJE
6b4vmhn2eIXbWE7t2vbNOFUJtmiI+lXCQjaJaQC6at9YApqn+dsyHt95J5vSzoIH
Rk0RcMktaKQha6/H4MCYlZUMns9jQ3+eTNlM78pqoOezjWEsPw6wmEG2h+jNBCmX
VgPj+ra7ubJEhnWS+sV8bsOhAD1tMdu3Cqs3aRf4/MZxphS7T3Aom/Y1n8cJUYZN
p1ryP8ui54AjRDFeGnSzFX8ldNPbcCrvGTNM17r63fUzBC3toHxIAaDynw2lDaGN
kSaaT+LDg1RPAp5FZ+sY1WWKHRyCTkhxkeR/PHsml766uPrpJuFNb/beK1jHoXNY
38xQcbb1w+mqhDg6W8hRUTftJt/ed7h1GD1+PcpeBuNICM022F6DGpD1eUCm22AJ
3UPJHfceBNUlKDviAYshFLbjnPjFotzJkeHYW3X+kaVD5sIET3faGlDvnlHHdKyE
YQmw4snoBZkcsP/1d9EWriQKkRSXzYRC46LeZFdq5iR/j71ZDCdFocvmEjrD2051
QhDrtGOnwa4efxCsmFWOk8m1c51wYnUHbe5fxViJKhWqSxBr5V05s6bXI0elnfXR
p81acbLDrE0GnArAToAc3v5B6iLKZ99Udr8eHKINx19CwM6e80ocLwQ4LukxKpn/
QybkKj0cviE5x9z5a34NuAdKI9urMCcvEt9+6d9rNYfyCkxoyOuCyTYeWfFs+Y4D
u1k0fY8EggQs3J+tbyBrSN9c1Pw3KEuMeguDyULUZto3LSXWJdZD0GGF6rBWbKsv
F+askW5CBMvx8h0VZZOQW2BDEB6LkJ/XkC0ctCvfARJeH+5RZ/ArwbcsRIbG6iE/
36RSQGAOKxXIyQ7IGitBand2sOC3zaJ3iEp4TOjGAsKC8veuyydRpCHpnCRpEPWF
TTAAAzgsQoY8Gtv3JhcycfFeXnhfRk+3WAloMULQ42ss/GiUqpnI5rJCBpCT9k/u
BHHamJONFzxL13SJDny6BCgRl/Z48LHLVGnikmOfnFQrVbWxLhG35wHc+nzhKmH1
tcBNUWEzby1WBezPmRIIijrEDcoNXxOg4yLEEqi3H/ArQYQ5PUR8jQPiIdHgbOzM
9e8bKinVcUrcz/3juT1ec3o2cxu8Rw15Y2+us/RFNomLo2Nk8A3iZqj9OV3WFOza
wz1uuNLdN9YOe2u575I+JDWguWdDcVAD6Qs1NjJFNUG/Mm9zrHChHJ83hOgevm6v
xOgIijNT2z9KM6KsofpKDdRsM/PxeHEnfKKF5eRrkKHln7ldvD1BH+meX6aH8F4N
Rbe+yQdFmoGC4qOey2v20Ae7muMeMBIOv3Cv9XroOOdAd+0kIOaiWx2UVYp/9j0z
3oSWNasxDAsoiomd4qAg7xla+P5yN+QA/v0tJieHy85GKzJjicKDf5AsAaiE4cor
b0kBpXluS3j1TZGisl37jUB6HDI+eEDRZc0FxX7Snehdjwl2klSPYe58vMogZCN5
n9ibZV372ZPQQFyqUO6jJQuqyi4A52/IxribZFLEP7VvThvTQ9cdbuWn/mlyvIW3
yMm55+xLyODjDhEcJ/o9luqSAIMlUm4m+VuACQ22HphDTZYmHDKucKTwyLz44BIs
Oc95TPrq2Pc2ThhZpURFBQp48roQotGAwSw0UsV5sIQQPDR8NYzegcdQaYL94fnf
CD1utqFNt0HnIgicvSww6J8uQzRi28zh3OTLD1FYoRcpV2fEQQ/EsBxaiT9H14oW
vZODnBwKQ3P73i9qHx/foVNulrrze/sMKE24/lzUeMrAIm2h0tGrxmUlKfuC9fI6
Md4XDk4QS/2nPOJHtCy/39xSvrTiUsthvIOSjhq4bUfWKTa8jdAuY/0vDKyXTx2t
MgDrjuSqgi0yTb+jXH8draDlfflxTXJ85F+tcVfufXToym3P2g1CU6ydmZPqxj0F
pM8bQkYNGVV+bKwXlg03aE4cia0FmxZU2gOP4OBMyH+aSu0UJHyxKBkVXGvj33k2
oz/4dwxmV6w5ZPApu+SBa1skR7JFYxfeXIttc1hyxlcTyd7S15ptgxrsrmjvUWPo
rsfRcgLmTnNymMfZxMTSbT2F7KGcUOu3w+OJj0fJa37khRQSTjCGymUy3qWckizY
dJopCp5cnub+rL2a2KsCT7GF/zgbhMkI62MKUXv0qEX9VQBSLMtCL5yUCY4cstbn
ghWqKCddx5tAXvo1qDGqwAfECFdAD1msuvmpairM7/K2prQR3+eoELTLhHGVMj9F
JUtMCCdvtYChhPVRlow9SUlaMGeQIFgtQYGDvf5bPjRG0xl/uXUdPYcOrShFznh/
ptvOgjfly/Y4ZPB8yPyPAKjQDJ5afgNuwUjBLqXjh82Pz3Dx9tV16JuSL4GX+A78
z0eTWJi62Kq2W+4/8UwdlhxIZp5NGtxhj+Hs1OzvrOGmB1T3V2x7CM1Q0iJppLpe
tTMkb/cBcHti8Oo5R/rgZjNym5O0pfVJh3GPgUdjJ8vN//N9t09Okr1xGG7mouF6
Eb+alC0sQ0s/nIe+S914+FgfgeUzA7DkS3Gz51huV1lgYbc0iUqGFxDDYKUu/po+
B1Bx2g8ZneqJM26J1pn8RN/nJxeLzbsbJzkSXorMESY4UAysuzSJgec951qX/sOf
g10fqVQASDxrKVVyoHfXrsqh6zawjQORI29S78GXSIE=
//pragma protect end_data_block
//pragma protect digest_block
gg+pwz9aoYHh4HiwPhyfk9ZJpus=
//pragma protect end_digest_block
//pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GvESVk6f+qeBksa14XQwOBaGceZX5t4jAs3XvOSa2pnzRUwxcQg/3owienGxjUiy
qs00ubCt+NZiEM0WLYctnREJHg8ddR8iQrWEaofxYzlbMF3WMzdD355BO6YMfcI9
sd4hi4temXduoNMcY9O/cnP+x7gLtqU8b0zDLVTDUVA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6640)
Q2GY/9BfDPt5zlbDH/GmTliNtnhXd1JCnL3F7xp5KmZlm3zrbeYtUkJqmR3YukC/
jXIW9HgIo2m+WllJvV3FXRfMxxnuCV+RnJxOZHSCHpEOhYP7ERUGF/J5F8K+hKXZ
Vnt7/hKQZ3yw3p1RNrBWt0PNKvN4u1dJpB7AdDC0WqXSwpcC1ZVKxUCnwIGPA5me
xETXghzzpp8hrH0srWeDu2efCPRJTmCgQe+rGN3uoo9N8/jBkIostYGXb5G76Y1S
VDBtmN+p7LnJJ4uJaOT5++G0DsIJYo4bDPaDgNCZmVsL0LipBT1xdnRQXuuTiKW0
/9zT4ucETxd72B04/y0OupDskHpyFjfHXrUcgd7j/Gyb6Dx0vxglKfl9DtSxecrI
Nyvc0WI7/80/oa6wDD1jIajcst84VGR+/stFmwVrU5ldd2w6QB2vVtgMjpXM72Xr
AJ/BKBm7fJH7pjvjT+nzuHR328Ly6H0a7l/upC81RzQmrCLkM6MJ6olSrYJpYiW6
SdK3XGq0GkR5kG1HCprQjbfKpI1qeuljsgQF45781u4t2E7ANbVezbsC/GILg9Bz
3gKqX6kp1+PKD6g4NRuqTPNCE9Hnw/Va+P9kh7WS7+sdwn1VxIfxEj1FAuG+GA9x
tgaz0rJllulC6eV++uxj5FltDxDxqw/Pnao9VJsTy7kBoZh99DWHJfx6oAvwX3AG
zSLNrYe46TuqwQT+KJNapvHbdwKkYz3GNFbeBZFB+WA+FhKoqv6fIlRwCe9W9gxp
rauP+doqcChYcKwpPZ5b1nfq1hhnA6Y6bnZ/gfnqO0/XaWqv3lCFREbwCtu12K2p
J0SO4crw2aVJgRC4AKVrCuTprzoABmxYwfkKjGdyIrQaXWuEddDf1p/3SPdG43yW
tkYueYsvi5HO/YQH4ujQ5Vcn+b5Tr7liv3y8y16Q4TxP4Zeq28mB3yS0kWHB32Im
iwNP1aUPUY7yUWVTPu3NGnuKXPOqEyYBXWxYrQq2SqcBTRS2y6IAJOWAV1jRlCkl
9DG+xIKcvnirVfLEFhITYi4MvLtC/dgY+eS2jQ6JIjwETQPQWLGOmS1f+I6gIgfZ
KWsZn4BG/JvpWccAcL/GFsgR3/vfbbOiP6jN1mswybsfszcE9HT74GtvHF+Qswg/
DEwOS4K2VIMk5KjePXdoTQSuhFPSb+j4NBhdzaqzbBpRXSciHGSzRBGd38ZvznzI
1kBmiUzN5CKvpPBd4krPQbZCKyIsMoivmOEzhSSTLQwenaN3SJqBqYVGVtJo9ehL
Lt9tD7g1Cy5QTct2N6pkQnU7l3XrL1/0Uwb36pn3XmDmkSSiAecRRKeX4TOO2HEf
Ds8MlIExQZEVCd3SzSD0/6XurKeeuRbVyw8zZG+nuMnxP/o7a1LwE5tX5rURXZ/R
LptCO/WZ5Mgo0WGloKWPHQUf8skfPN45G2ev9O/XMQXK3rxeRZRV/rT+eEkoKx8x
OXunLVB/i6kDD+Nj6cxxdSaOLrHe5ygZmnMzEqbVFlv7gfZeFcX7Nk8mMtD8xhCN
qtfsFUSeIXt8tMhjjPQnS5wIPVL+ECzuHlfFIFxibQBzO0gfHNY9c75vS0VTTR+x
OdAlxB0Ux3Ps/3mLHGMsbweeBUlNf775QRikrT4bfFfwvxJCqZJ89LRoOyuIxTEn
vfXofxsCKfyq7s7sQ9nJZmf2KZ9wSys6ULQtt4ONQle/mz+C8VE9wSeTS3WeouP4
wS+LQUyFPMfMq6ch5zbXeRlMHPSLvGG3QZxU1EHNYtCdgyVXKWThqDwEqjbbeKLL
70ken/F1kkVeoz5Znn+EeKY8ltG7NB0ytsP/3qSLiZOQUo/QBKbNb8r1DHxQDwgn
alFLd9mhHy1QKv5R56toiB+S+Y/wIvDajBG78qJVAStSoZbgL6Q6ts2FCHWcCMeu
vvf+Jmrccap0myH5OP4Yec8BB5WlZ/CiBobIZ5J5sDf+rrfU7lJtN787RdRUy5P9
gajpt5M7JW0xmKfAORv9aKk7gWUHlE6QYqnzjntSmebDfIOIqd782WJZNEvvcK2S
5dn9jJuRrEdU4zIkyGXiBsYQlrUt/bnbbdGZ8g/MK8H0AYXaSBU0bh8yHuPdEsky
KDlUguBAdvGhEjM6Tmp2kbVVu0kChx4XxR/cthwmr2WFemjzsf8CVnoCF4rjQEUD
1ozHoP74tFW4B9eEpm1mC/TfMqFg6e97+WUnbz5Il1/wDQIbyDd4c9Rf4juo2A1P
USZcJ0S8JZzcTASJV3Virb8+UW7SAJP3LYAZSoSVvKfdkC99AwuPEbzHR5+Da/Q/
m4pV8iWj5OwISbcMy6L6EA6HoQCeSgMGmUnHLGNsO5Nm0lAY2yW52Q4twmTjiq0/
ClKWWw4gMlaAaNgVqNa/UPBL7UyHrDXep5zoyhe12xlFpKaNi9ZnjkcCp+BayVFR
r/+LKbi9UCu6AfkMKKa7Y71uh5o/c0Ra3lQC95tjBcuviwFHaA0yYyZcMprB2SU3
sDwEWO0VoygJ/IFDYspolm478zfMugq+0IhUKTk6VHLS5QWBwqeQkrGFmI3K95kZ
GVwO8cv66dbVFYYXcMsQQ0rVf+gGjzPlWptS8F4RNrSvzXRdYD8YCnDUV2GKcleq
CARid9wKVXAW81ux9gbom5yTdGrSYuV+DmtnUY6T9wkSuMwhmKQR/KiczNV66l4a
uxNPo0t3Elr4lWBgUAVW3a+ll1evsiqM8SVbNa/P8NKSsJ3MQkKubouEFly97/DF
rqvq8pX3U0R48YC5z23Wq/n1xNDwkKjkVF9JBLSlQt+6tj8wbMMTQ6QyxnnRoPVJ
UruP/1paUPKRr22zoxz2+u/QrrfO5kzpjEpgml5kk37hVFGnafHu1xJ2kALGuL7a
Pukpdsh6Q39x4MQMoVOEfCQoX9Xhlue5cahvOymjxq/4LLcyH7dnItUfmLtl67XY
DqF3/K8MsIbK1HNlS5YmI8pCUkmmeihys0MglaX0/mdhOjkHtxJoUHcyx8r+JHTP
oyuCK3yNLdQShdUr+4kDtsNul+7aYVd731RaWhUoX6kMrYR5M40Tkq/+5L/pvGu8
PpsMqXTVzncdlAJyvloD/x7m58sGcYd8J3I0lVPfpLL1zzYyc0IMyvj/mUFagotm
vlpRRufY0qDyaW3zfslUwi4XvVjGuue5oLNE+LDdorKuDqP0uTdolSR8jH3lts2B
LfX8SCEUASd+O1SNYmeednZs9XQubrUWingslCZVlzTP+mfLquYp9S+yKf0vv6V4
JGBuWRHDYlNRLppGrIwU8VwE8Jt+MTU8ZEF5NIu4E5QBd6vuaRzPDvCoHyhZb1mU
NXIvBtkORHo8zzeJe43CLatA5207RnCByAbVpE0U8+ISpYabUiP0xkE4g366oQSB
s43i3zdUoOEDE3Jx2vk4xYmxMJNhIasT0MxZIckFhQI/+rAnSxPTR1kKc4T00isz
+w130FW4BEFSxInP5j7dW6UHkjf4Gt3KcvXykdTPyBBq7utQoCQ36vl+GHzLdoW2
fezZZ8LUQQjXhHAXqSUTNvMBWEjVaBYS4TtCb3mURxi2tE/r0cqkHhVxlSqSwTR+
kkqisQWZqyQtN30gCqt3iGGcjMpNWaVbWCZpgOY3WSt8bOjU1/QqjLImVTJ5Vb0A
V2JdJNz3S3WBJYLK+kavYzbv82Ft4KR9fJ+5GoXariMUxCiJVmNb1XXjm+OphkIZ
wYQ5XWtH1gwti1MMhTkJl4FJBdyEw7ElRO/4jq+S74XDxKAgvMaDClhl1R3xfsSW
iWtwstyGeal1UhZesC8iEBgGvMU5s8/WhQ/Hf1r0NZHc9xJVF3BSciNuwW9Ew1le
Gmzg1QhNm4M6xbDg7T8S/T232+OPA+j6XdPnNo5XA1gOp6Z+EkURp7xp9M/bFRr9
02CJuZpec/kYvHgKpptorDd6PgaO8p3KUkL3Oo0nWiZcVNk1Ez96Di/Bwbn/3aWx
8aubwgAVNjgjmnsSk2YqOtF2UDS/2ODiFqB7eWvkliYu/5xn+fsc60YN88DEDI1N
powe6pB0f79H4oxc6jl+YDDZYLL66Kb0TzGs9iuL9TMZkbyai6MdoIM2z0yNxYSU
16nVhzwyqsQYPtADUq/vJGA/bNfzh0yspGxIhdqgMIosnJUTrxn8qygVenE84ywn
9CorMtrSPEZpabgd4AlQyhgD0T9agnEZrHW/4JIbdpOa22+2aaaM4qrp4L8OHFAw
IpvfRvYNqxTAdhZzJgWOwi3m3XAyR8s15meTgtbhdIq/fS8DV3d7hZZ6ulSbKnaP
LK4IHImWPS/TJ6x4vjRv5bzyb/R+O7JVGU4QCZjVZ4Qo1On1thaKpXDu3PJGnzza
D9JaTPGW5R+LlGxP1YyrsVb9vG6nt/QHvbFldSkYFcQSydwap3qoToRTk5fV8zAH
u8aP4v0ucc4ahQK4k5SYL84rWs7T9w5uYXL9arWg2L6rNdVtuwcQLb29JcO/9/O3
On18VUgB9L9Po3VxHjDzwwxEhBUA7k3MclcccC2pU4TQo8l1YvAx/qUkmMZbbSrK
OxYbno/0HZRHyKAxbqbpPoZvILgjMyvoGlJeP9Ou/yuggFiP+TjMedLicrloDHlO
YGqid+OXGYIPmAaBap7cYEngEeEhbX0EQQO4Sd8trrCPCvk9qw+6Z7lY56PQQHL0
nCfUTyYgJC22WoU1emIeXQDmcFVTUCd3iNIb5tobnOlvLPpspPMOQaVpw5ME51Bm
lWQfRndr7fiZd3EK+yqg+9bvTfx9JY81RqZgfIdTaBKVZp1qi/1jAfhTSDjKmI2w
muAcMZKar3bZE/vsUzClVqlKl8opcLgE8DTum2kbtxfxZGxxlTcueClcD2+1GJqL
IeuzKMz9wujJ/8TftVDWlQXI7N/tYf0I6Gjn4gdbAT0WBqOc7Wau/4FQydeZfA4L
F0Yx652yI6ryIStVqZpAc9KHFCvzBIxeM1mIpED/cZb+fuSOATyjOfomAAPhdWPZ
ncg6M05YynAvr/481UVvY2lVHwvlWQRzoKH4BZjkjtLGJW+zd7z9HlSfANE6x+CC
nh/Zn1FHEn6NNDzXb49cZOXtFzmligIl0gKMjXMCdjbuu1YeHyMymcJ2QTns3Ybf
wrowe8KFnB7P4peOOXPjqwpkbTz8oSAVzIML5f0gM25aBijon1gGdczer1F8+KRi
/8kfIbwWykZNZAH2x2R6yLs1/Hwkj+97SfhvIp4RJ0OTgz3WM7kXL7JkXDkgWZ8Z
afUqbZGt5iRRa+NU9QClB1+MURaYvCAq3zTxBX8XTsQOKCkJl5z/t6PSlOqsCZ5L
XjiKCw0dbl9Pz/G4VI3cy58qv0kOOmSrSrjhbGOuANqvpkb8MWA/FlmfCLHlhluR
3Tib1+1AL0dyaj14ZEBpVc4mJIYi2FJ8pPImdNfymbNKS+uCGEU0IDhdyA7O653e
l5k20oyAojpoI2DlQPcmH6/CTPTprV06e5dwLpxLcXosowV9dJa03Vzzcx/qGeKE
7j3NGvZGevBggLFVIvuC/zCuGEQfFZfuCIMthcSZ/sbCLxzEdksSsLdThogI/osS
LuO8rh1j0y/KGnSGidTWl57+Q3aXiN916JfQ0ErKokTbpBaK/caeHNlerT8hVjTa
wQdzexF4eQY0z6QD7LVA5EfO5HOZ0v0dhoxJIcovtyf+2P0J7H4YAtElsZovppBx
QZbvfWXWwK/Z1wcpD5OXUoCIzn4x/QVym7sSya4MN2iwjrSv1m5r5oz31xMHyIKf
XI6XkyT96Vow2tuRD1pLTmq28MGnyRAv3EuPzw22CiJZMM2oeZf836DUFBFPRbKc
zxWyc4KxnTvV09xKVRVsCu5k2S+ec2jTE9iztCSo2SFe4Nehe3hVe3U2oWjxgqx9
uGeDZRsHVv6XJdaBuSXqJvHVqoSl/3aM4TwZMj2vAN/uATtF5JnRV0vhcMM0VpNo
6yMne+1WgNYcoJR2NpnLKwNEWZ0BAvOVNeQfTZfMAucALQvY74Sdl8i9+xA6oxVT
8NQJJL+QmTajvErZ1Sg8lnHJhFBJcOpK30+hkx+1TkXXSloM3MpJuwXFEziAG2dD
MLpfsqQw7/9Ue5r88dBwm3L6W9ebCpIftxGP6JcXtjqNhXeHRTjUHuWBknAXxgF+
1ij0CG3y3Dom30CANiaHQzo+IfH5wU9nBBeC8YKLR3bkA962i4fNVc9eOB7gtWD+
tdK0sBuANeTie3VzDCB41ISd/LPM5nxeBW4OtJ7lq2f4C47Hv6haO5KrgtX7rK+E
pV1VUB6XKSoO7EJs0P5uPxpnZW7DMTo0fLnWmjnvnKFTRZx8A2bvvY/2Ot87iWxQ
SpAuvO9gnN854umg8DLoERWuEGMWtG/c+qCLX6ZfIcAyfXyTl5e/suwTdwx+2NpT
lU9z+7gKij2dwTJ5MMpfiT56K9yK7YqMW6u82fswfb5CSizFWVM8Qd+AAAN1sY0i
WEsi6n4g2lPhNBT0gpCi+eoPzJpgOfhf6R/uSs2wBQxwU4KftXQL2HT2j4Q/on9l
466oMcmGyyaD5RSQ13gNupb3UWwYPvJ4I+ETvD39/EzcrY6HmJRxJjoFw9pl+9dh
1EA2XHjkTkpdP7p5cKp6Xv22jf0dPXbjQm9W2F/o7DxiRaFUuMO4s4mO4NqnQ5UM
VX1i3zurz1o1VVCnZNmaRjfVJsJaZoZM4+zk0mA+DXIGeNRzc7w7NiQ+nQyQRQfu
WzS3wCOo+Gp+79pLVF9RY7o9UZkSrVNSQtOuiR2CG/U3lQFXFNcUJZFG3rJJXuem
VfmsvbeUn0kb+DvPvXv7dFjjMFw0WpFSYbUUot/pQeS7eMH9nHpP7N8wg02U1AmX
P7nAGr8rIou+WnTdpiCTWuJ2joRcsq6M0M55+DvraHkqhnsGk0ili2SCXnbO2OWC
CAC4C3o4R2gGzl2bCTxa3QeDVHaQINggAdg2guIOTfuy2J7pNAE0NGq87y/4uju/
SNqiMqOII5Q9w9wdUKNNCNl1IjfmsqX1zwUHIb9+fQyq4iJ7J2WZFUugEXX2hs/9
p80LdpvVtFv80/dN4YmXTtRKP+F4ns/k7uuSWkByAjJwN5U2YbpbvTLabDpR03JX
w1zdWfw8u6Gm3g1dfBvwYqXKi6ght0lVu6dh411fDR1d8FCl1jckw8OCSGwYw1xZ
3cwJagy4Q+/voBQ5kEolt15lffkARNf/LQtKhB25EJputmlwGVphKyypa20EXOY7
rRVsJh6GA8z51/311fQvAltdBYojaSaWfuoz7FxhIi5yOlbWd0QbwPXy7PrHHzt/
od9toaZOZyJ22ixaKy+gH9FTtGkT3YA44POfv6Jh9APi//Y++1SDxrxOpfgBEqoV
qcByLjJF7W7huyNWeCYoSH80md4fQOBEkymTzQlZdsBjhAu1rU4IfUo1nELE9e0Q
POn3HrrqTj4tnHKvepXOHPKGucx2Wbong+Fpf39AT3/0/b3Xpi1cl/5xw4qKQzr4
WdGa+F9NmS87+DnZeCJFTTkb73YORLY2nuDJ8mARy/mKomYLAct8RVxYxViogk0o
Dqo7WsUrIYehAJVMHVGNJZd+bgQMfMFV+ZjFF1phFejT/6ghowZ64ztIS6XkXuA1
EDnrkP0IDSUqm4cOHK/G7faQbgbQTOwX5RZ5EZt42M7YNTsVn38tIZlf9EOiZTvl
SK5ehaXeTP/dw+paKC7CQmi4muwLKlJbghkXBIE/MmpLRjBGs//tBBDXCFlClOvM
kXFNwPsNoNMETNUJIayu94FFa4ON1RO0iabMStcI/CBFPbt0Wq1KhUuPrjWgN0DD
9VBKk7QuuWI6yj9TQxuR0U68Syo8dqxt0Mb05Ga1vTY8SQFHZslbH9cR7u9VsMuC
LETj8K+nXH0vtvdfZ95tSgfYI/G5ACegfbJQ17ZOyAYNQDPYM5/rqnMtSI7p1JPV
r7yO2WvF2/p8m+KVXgpd6R3The2Dyf1D8emGYre4pYYa3HkqQtKZbSPp9ATVcsAp
5x3Op6WXmRVmRi4CMsR3Zo5dzGFOYmSBbTpb86zyCifcg773AZ0E2RChUxtW0WtB
02f9WDIi/UEjgYWym1dB1lr8U+TuQHaHl9FIiy9GA0AdMwH6XhvWHK3WSF7/QP79
6EE949ljvAsytSCaKh2DB0ZhWDsJmM/BJ39zyJop/T//G90naI7vwWbFkU05IZQa
1cQEG2EAYvd8hx0WGm6lbm2HUG6cRwVx7XyT9+Z7X1HZJvHWbs3XXztoqZP4uw3f
Ce4+CZ1cUyQkxZfe797/X0+HodxSCjktK5Q5nKLU6zjx75daHw92poau1Kx54OTJ
6YKgDGCk+g0KHMBE7PQRf+pCXn8lqP3hkbgCPXbz7SMpavDQYiVUqZTYf5MsVaTw
SOb95xImrCKY2KftN3JmnpPda0wQL8wMAfIA1owkWSfg+MmuzFqcMKixV7wHNiiI
V5o1UvKPc7Ib/sr9WOMibS9b+CeWSvfbNq2Brjo7tdnLiAbboJEDoZE4F30zhRYf
48ybUaIkDX7HdYuHltt3cOkDdvv23xeY9bvmPkC3QN7BXzaxrl5TpsMUCdoo+aPR
5Hx9K3ObcIcw7bFIziIA3YPc05hEkUw3FEYnWtc5X4tTr6YDBrM3h2hg40YSNKBl
e4kLC/+Tl/WYHehRAOceoGh/89+X1bXsnZ2u8jJiNK3EPZ+0j4i60ir2kVvotcS5
4AIMJQeRLjotWqgJCv2p2R/ygbaDrnqegr/dR6a4vUVsqv3vGH20Lj7nY8pThtiZ
2IkELxU5fQ5E5Ud/uJAVF93ycQ6X2QwTpdFITVih/63ghSGDar8fKKco4C5j3t2U
EzeXF1UFceiizUdxVRZTKQ==
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
koF67esXH0rNf/ellOoX2qyjVdSz8vV5SLZfVEhgwP+KDgY2xRcVhtp8C4hjPPUfzYXcXa5gCjKz
O/rvCHzqbZlswhElHeM1jZX/b2wDJRq4ecdLkdp5QXV4FXRToMI5qct17bmFEH4hHUj67qRpMfLt
w22+TYlvYYp9BaUEJydGiNf/jR1tWmVMlY1LLEhzd69lZWYJCqMiVpPNgtnfV8dm/IpLhIgAwN9B
cme5Ny09j4s1/yNSnhlsxSKXQaiSQLEwtaoWdYKKcChFuu2DGyXqpuVqI8lNdhFO4057W5q2KzFU
JX1OLg2s5aVfvUCErThb7UhpN1DF69bj/AYwkA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 7568)
lnehX3SaTZWPAJZDQqSnd/Y7/db25dD+GbB27t8vVLHDaPDHsoiFJ1gs4CpzyrRfiNhCaG5q+F/h
lGHQCRdeX8NHA50jbd0gLDuxpyCxF36Cfeg7zjFv37wfZQOUO25/r5xOag/nypCa+z0HvxsWKBJo
KQkBJHdGw9dAKfsCsrQYSLhDyOW6BWtOdTn+dA+Xa4G2BcoGxvkXbvdaaHoF9AsXx0mconWOd+sf
NkSZynFwY5W/mERNYO4Qr+MzBpZHVZt/OlbhWerPZ1wU4A3UGqb7h+kdQmPu/2wb6LTn55jvYViQ
LU7kwcvKvI8HTtYo9yOqTdGjjEa2z+ywE6tbnMR1D2ihb2REEq/lSvLczl+weffysej7cCkRJync
dojlVRywMWjN8aF43fkJxqWva4ZC8XRKEpTPo4S1Q3Vpt1+P91AvVlpu8oKRNCFdo7fc5bb77WIW
Tt2wqnKjenq2ygkoBl+upVM7ZFDwpU3tLt3eeis1OVv6ANbNQ4EaJDp2O/fNJ28XUH1bw1JCMYpJ
D6j6yg/nu0uWXVt+PIfYvwLaPri75wbBHxoLlSNJC87i7IGvSL00UsBzbfcObbQtKTIT7Sxg2mpt
56DUUexn4DU55rTNA9ZO7bRBowF7XE1mijw+v3GTAwYLITGpmLPOrF7BTyM20r4m3Ni/IfnJMe5C
rGEzBzi74FY9zzuhh/vBY4GISPsxmXdccTZpM1WVH8kLzhE9FGtIXzX07kiD3i7s+uGan4D2cOx7
Vi21wViPr+FnDVk/navMZE6Zsu3sJxShvAaFfLlC+v0alat/JZUUlxbKoAw7yXWNdtlDcum1A01r
p9iaRRFtOixCrWSBDsijcN+Mlr69JWUWVi/lw9AZ7k82hgVuyFtpYkcZEGMQ58AB0qgy2dG0kOKt
vluX9fQG1Fc2rgyyFBUq7CIoUXARb/k3qL1+bLuP+1nrg6Zq3BU5SbDfnWUp2Sk40c7veoiDubTx
9+otXZXwyj84ipkrk8FQkeWi7yJa1ueDmW0chGfIahIAh59qqBLWpPAauU6IT7f9H7SpQC/TC8QF
KDd5Q29sGX0jVffIvQzPvt/Ad05UrT6bYXf0CfJhDyk9i4sl6lKMzVBtmQqULIowv8+pHzhHGCpO
OJqpnEWo3cYtTOqwkkaKXsyazo+77qe4pXYUEdng8G6XFWuYpifd/Ye5R2SOcGEJbEX8v4K2Lqoj
c8Z/J9UQDmPZdcd8We1ZfILECfpQyqtb9niaQl9+YmazA4g3y56NvgK3le+Dn/yG52vAR1WfNakI
aY8h5PZliQ6WYbdXGOjpS0mggNOHdqhylfzOB2WnYsyvHsYIsC2eZrBmMbzdVyu551+MBLdz/uDi
A87r323iLkwdmKzJdevovyEJTkIpYcM7KS+qyZz7V8f0jnQm4Qi28+B86vFL/cLndZygWtWOTOW0
QCc/odaGQkvydW31Hnxrw8qgH2Ph3LHI1cgnhkFY27OEYhUhSFk+WqXK/T5f1wwNTR4lyDiClyo8
N9zchpGviSobopWRk6+Ah8v4VeabwXs/r9lnTPAEgc2ulzMD6vrDPGJx9EPTxADxwwS9dRn49wAE
z3mzPEUcO+BRFZIvs7UKE5fE7tdSra0c1f15SqfsEwaFWezJI8Rp2MbaNLIbH0VaY3XJy3EH6Zs8
1g1SFX9XrUHRw2MRo+62ul/a1n9VfrPgdW1Ih6rUER/MI/idPPLiBVd7qefWE/9FHgXpb/9v9EkN
Ae3vCHpa8Fy1mAOuf2rI5n/9vywf3u28LlO2xfQC6gzC1Xw2FIT2dVE8iAM2bUe4AD29wsa0QbOe
P7q0Dz53hES70cw8n0/RGQswqfbt5lUeVh6J5K9kuRY5ONWZghjj412Uh2azsmbWGgOGDJG6yWgu
YsVmqTpKv4IPRfv6NiusUTYH1OvNf8/ZPoH9+2eV2rut/8ZbUFwtlNRu03fM9KymsfrsT/B7LH00
gpOSNEGEvGq3/A3wYrb+ChNWf/Zc04EqvLkLRo5rnZbcUyXZ6oPA6xRDVYBHKM+q1HFQOaifw47I
dKOpCseb2bSXgAvCdhrTwgZi0rMfxKbIyEA12YF0BazwQITJTWO0gMXXdJ6sA7ePy3asW6A9gpaN
gfxxYtLid0VReLf0QNfJkantQXa0S/BXkMHGkVDNg13EmS+W2QYd/4GAPUIsfh2/STcs+9oVT/TP
SiI/3YV1icwJbeGnlnFbH/Wq4sXW+9hKf5HOUyYENOGrG444oMS09jy/uNOQYIZslyi2KFMDbclz
MI3JXGM2TPcL9atqan9RO+gwXjL8W2LSccAclBW2eZ7key0zT5sBlSaHv8nqgqZ7gH03Uy6Z+7A4
wv7ZDwosorRRbs/lofJtWuCWEWTXXbZxvHSdahqAv4u8fZZC+YFRsE4dxe3PIT8U5GwRDuch5Yxe
HNGe9jCSxED/qpD5yuqMwBpfcGIKwn+yZhIr3QPVLU/LQnDQyEKY+vufh9vGHHCMSpqFGbu/OCcE
SaI3MuaCayc7f4ESmdWTGhiEwyPQ2Rczn9JwGLP+KBd57p4LJ9Vc0lDo+6TfiJy0U9bOv+1nZFgu
eNHeu5S7S5FdWlE31Wn+4qFRVi3zMf4TNcQj1SC500x51NR4xZxTvGB0hbq8UvCuZ7Hx9jhabee+
1FClAMLrAMtWGl5GsCQHn4DjVnTrNqiPXmAd+VXUyd2GYLvcTYWkwQ9FqMnChHFR3i49zqYNmVAA
DQM0mcN9ywvLYvI7UTK3VY6NBk0OX+fUI4njGodXWFZ4xDnDxDyf5JSG1YmMFWA8oD0M3rGnHL9J
jchhImOLkSVUCurvGIVd/GgayUT0WE+OGywr/6AbKdVKD/nZ0h+jPB3TW8lhXXOAZoRbbaIxisXS
JIHkacy6BZyTwOlXlJdQRWaT0ZrA/9rnYtkSEYdNqISgCWchO9YqT9+0ZIHaZgAyG9UQgUy0r//k
GyeE00rqkpPMPJ6dnQaaSbnuGuXsb0gwRBVyMnvlbW6OFIyLWwa7I//lWQI3Sy2FmMNgq/aEmyLI
oHVyY6VTS2L9otdd1ZV4pRZH+oOBY49Hlzwx+kcmWjfNVUhkScaPBL8DLqUFOmWYapfWc132tGT4
B/Nz1l3i8ql0Zbh+zwfn84k0VdLeoTp/EOEMsBvgQQrKYh7TLxDuZrELlSxGY7bUNmQaJpPqSkwI
OWPN1LGJZChoDCULv2QkxiJJ6Zohdn5SGOerbIUF8iSWJMmqX4+1G0WXPqXielY2Vitz0gHGaWj5
+GUhfORcCUlyg9QZJd2NOeIWfxGTlN7CZbfjJ2yTc/mpjLYvzv4OonDsDshXDuZH2OOvePDGrkMo
9nt5jTJKd5j3tbpOC7es67c/Lc1me3ocoYCUeBwIAz7O4n4+9xUnH+xR5pG1GCEkHxq9fzQP6AWQ
7qL4j11eu/ynWq7zYa6UwIhxXNsG4nw3VjcylmcAt60gUiD74kI49ayhkljKlE5FT4n2xPGpo5qi
6t8KD2ijZjza7O4DE//cO67x5PW0tvT0cgBTQ6nP2qbtveQdhOaBRsy2Im3trQvi4T1XjRN/KEk9
92eCqzlmvUsIAgLXYGQPedZd2aUHeitk4V+V3GVO9/MoVeHGGA2MZVInjOFbIoMr+XnXX7VqsUy6
DyDD1pq7HHAj4GJI7Gu40ctch0VJ0OWsWDVAlc6EGBI+De77U2su+QhuCJGTsw9nAK5oZM1hHLhp
khWpXBw1e9SRUDzG09OVD4QbNuCQ/2upBZBW6ESAo8j+Wejy7Ie5/N+twfMJ0Techl27b0NeV/S7
d2U02YyXK4nRF8KWp+PBWk34tEKf5zQL8hl2IfhymD5n455qhMSdWXvYe8fKrsm7HgVbryg5m2Jm
aERVz0pHYql0IkaTi5s27NyOSf5Re31dBqALdiP6iz7Ltgo2LreeAY3nczCCMUNTkpt1SVNMKOqQ
BYu+fjFoFroI14O0sPvpsfZ69Sh4SKSVWaui0THYjyrPUD3O/9+3ksV/n2r+5TLOViWnrk1xMk2n
8AdgjQuoi2PoJk/jFKfMB17KUvl18q557jzFLGHTAJ1F418nDb5Ph5y6PF/xVIysX8U83vJrN0I2
UGd/3ftiQVcy+rXOhz/Z7GT5nRK/RH81vZCQD0XjMW5YAsGsYbsaHh4XY4uB8Qzc/zPQYBIPcW3L
i/Tl1FRc+4BhbW8CedSmO9ayIF0SN99JEiKY3fhXW+UV1LBLnsDYG26W3JJ64VCknaHenbpqUDIL
He0SKN0ofY9Lh5CgTIr34BudguwN1Y/xP7qd5XFVJ8ntuait3HPg4YlPhA9Nj3ulnbtNvar5O3Aj
Z6FETWMIc2P5EhQHNX8kTiIIhH+AfLYuq/HHuwyLJQF2gVl1RKkr31floR+LmBN2ToFiLJWpp+lM
bN0KPtcYBiH8mKg/TYsIXTZhaxMSiR3zfVSqotZK5iIAYDtZBsbUXbaeT1wydknyx/nU3ew0dKKP
NvtPhAbvET3iNcrTA8C11tnPg6vQTix0W043N0r+oTIU1aH6n3mGOlU9awSMtv62Ypb3Ogs+qgLy
3T28ZHC9BJBTRpcgvdjKLSe298A9+Jje2dnwFmjqEtMGNEbYLBS3IfV4ha7JVm9V0Y07psFA9dR6
OnmF3aRsckEAKshjK6TxA6qKGoytB/rQV03yubmYtl+lKNwJYi+FEsaHftZMYhQmlOij+fFvMhv7
wgJT5Eh1AE7T+l9UMVMI+4lGhQth4Dg6dK9SaP5jtdsRBKE1dRYLRwCYZGfeR/hrSmNVOZw6bDhb
Jx7LujMntYW+1uWFLf8LNB9ujMyZu21Ixcs5jmLfjtjbYRqOHFyrATBcCBjMqmjSNenYmV4a2l3s
E/9Y961BvzfQqn9XKpS9q5yeB8G/iY5XuO4zkMNMc93ZPj4iEZyEjR9L1y7bIREvUZL2QQt0wAQ4
yur7wlrheQzEfzbkskycat/wXSsVB1nHlTmG5MUUO/c3TYzWr7Bhbj2k8mq6siiEw9Ve4EVvqW19
+lm2KjcHwwScRmF8+DdSTprUg2ZzhQG8SxUQwpmD5rXhaFXDxCsGQpZPWy1H45OOewcBU2XGYoar
FAvr1WAg3bzP/a4mpWJ4noMDHf3uekovMyfLePpIIMY9tMbREEUyaUZklS27K+T2pUO4HlKmOpFV
7lakx+7Zzxj43tGbQpxozswUvzfV43yanGrf8tOYa5htx7zCV5xOpo/3ac68NqTfL1xJ97HrAKeP
snfh1viDcfy+vwtNrHtdbLxouS9siaYlA9uPBCmunhr0X/qWvpwRT1pkbpKNmZIg1E0d+iD5ollC
jxkHwCIdmlL83EH4udr/9zPWSqQoddMDV2zBbh/WAzfFTVIQjccdfaYOXVvzOlZyfL+kbo5hcLd+
op3GXKfducq76KprpTBzZp+MpsWGNBOxFGolHOUV1cbYr8vaCS1XPiWavNPhskZ2oYwdmcu2U9Av
sZ4NsNkYyY/GKBnmYgQAiEvR8FUw7mnUspIFBfzWlyK3/H2+co3zBTQc19ml6BhuHoSIif1+FVNL
kgOMpbMREwv0YDbcz2GHtbA6KE6rhM3FKzGFRkNytCiWC6BycbFDetZqglisdeCMSS+ukN33sfFk
n3wbelE6vGewM0T9yKVhCIKtMZDUgsrdEfZyoCa0Bhed22ntSC5gGp/05AAiX+j+kmEBlIhy3tXc
y3k7afTHxmao37ZC71toZpHLB3kdNByPDrEIe8GXWr0ZJXixyHV+QLTtuclv3x7VYs2nksjbjSgd
vYFDIA8HKJgNN4lT0G6zcyZT5uiNAf1xYlXCFz3ULmEz9ffSPF5ws7VrmCE2XZ4yDnWV29/FE1Ud
v0Kb75u26x7NDYL0sTREwHn5+s8JDpDbsPeE0AUIZL+Uzj7ZuKKmSDopAUG64iuxIZekxptZhSBN
CB79P4QKoUqhx6PcUg2fOyDPVmvlKHox2FjdIQOKHBVeupO5uvkmzV5/NEw0XNEhOzWyUtZ32898
I8x5zfOIkzjAZmiTzEaWfIDfwJhGqL2UXabC4shsFPJJPpXEOdh4DAe5JQyc1axycwwIozQjuBXK
s55Ioub+6xadJCOOz7lpQpeIoghgrUuS6SX1H03KCB0ioVwC4XAIDSSDnfL3m9S6AFnr/ItQuHR3
JgajSvAQfwxNaXxQLoMWKuMwF0td50Ll1qJqipvl5x3SJordhHZagRoh6JiiVwQrKeLvQV/lhxn+
PbkVcN9d+X26xsX3vlsZBcSsZQMb6SEBVC1bjo+8m95LUp+O2fPVJGMFFKVYYs+zejLPbqhdWhND
Uj8rV5uJORsapkvMgu6TdK2B+zOsPd7YfZeBFcpxROm/KdaHZS+z1rEKvfUlONxWSb/IutqULPj/
l1FrbBRls1xyHFjpgXSSDXzooNrmGMcv4Ilz8DDHBn8JPM5u1UGRHqwwDGBX0PNs9JTuT5JhevxX
7LNaDs92mkOwAgDSLicY74BUj4375GN+Qv6pXoNpA5sX3qhKFTc/zg4UsEP4sanF7XZILIDiMEa7
9jVGEaW5tSymf/mdwxQJe+odrdYDHM5XnpIF8SPJRiOKW7P/RBIrdQTB5ZN+6cbB5mtwcy4PAMmQ
Zpsxy+jQguYlbKsjgInROUwuJZzAse3PBc3V3Ksj7xoSh72QTy3yEpENIOYGg/bK83Z3jBq4rCsQ
O10kFRe57aUCN/WAYmvx3UXS+C8yhJnixY6dzDwu3Tec/XXAQLf6Rfdl9N2Y+nDawKLd2fhd23F/
/WhBsjAx4aj5kXq1aiOfNEjovhHG/V3V7iP5sYQQL6yP4u2pZyvdbBIjNNXCKbDhceUZ+fUCwcbA
1JMM9ZdwR3JlJdd78DjRCdd3aoTrs/fyfV0xpOjXK+k60TvzPcl2PjKKDy/BLs2uAOeP5zI/8Otc
NhYxBCV7xrUOfIS31T14CiEurYf4FXb3wa+geP1pVPNinnOFBtiXAHcxy4cxSTQ3V0jbZjBqUwKQ
CwIBL1DX/JI3IiGiM3PXxqrNruJKWNNJx6oLskb3SV0/Gfe7hOnlD61QVg52h05KkSyG0Bo/XwGm
ReGng2upw1ukdS5OnaK/Q9Z8I78PjIrUy8Y5o3jYu6WOgAPLJD3C+4F9srT4S6/NXg7brexgASL9
w+lyR6DSiY7RW9T/CKUEc3WU5d5/lIAdgAtvkYhaSJ8opZTwFuGl5bNesTD1WwiPrj9RitQOEuxR
EyI7+t/nd7eiBqH9fGwA2JGBlWaNPHnvsBAO4rScBxjSNTUwQ4kTxQ0RY0cOKL6D9jB5NyR7feN8
RID6VOKeH9eCNtvAESxHCpn5w9J/3c604yL116ffbkV5szFjYbyxT/K2SyKwSAj9fOW/GlNif0It
rqWr59iepkpRBQGXS84Ekr4dWXOgXwcr7k3hdeQZDl3h7AG0DKTsvM4cDhagkadXQ5XbksNUA+PZ
FSpIByeOBjYllFbSkX7wxlSnmCToiLyPPJcumuHK3fhfeQU9pqhBJuyiA5mnQ+mQFim1EiQnaoNL
9enXZKKj0TJPvvDS/1hXIQiQNorxCt1gIRryNKmYzWkNqQQ5XTtAPJPFQyAwXEj6nBnG97J2Bn/c
Yjkgyj7VkxZpioC9sn+8RdRsHftFZJ7YuZlrlTp3LOD9fMpjwi21YDqx63H4ckuADfRNnNTyXq1J
C2iqSYrtQSi7d5zwDTy2kVVasBM47vPm6PgYIcfu8ytoEdb0GQW53PEiLU30cVqJtTSgpyS5FbZ8
8dupnWjAxADI/rO5MC3/ZqHwhaHVWBkiQiG6TstLGfsoRW9qBpFBho1/CgUe9Y2gT2wTB9AIS3ra
4KWTEHbzEqEd1v0H9A1Ky3Krqzl0A0UvN4iQywoxGBIiOgj4zP0BoKsuxu0T9eL0hJVUbho1Wngz
SwLKqAbnd/RYwFzPSe34SQFFq7JekEHC3JY2zTtUOTlXvGy0MLvkRfC3MgMdxfgsunOGg0bCNxhf
9pyA1fFlYZxToXNqFkoUqvt7xVAKcGOfHe8/YJMIrPpGbVeZjEKYPFB1WtkgrLMnKrkEAyMbj8Qm
Maz5klJWBpIxl6iRqm0qv+WfTmoA0QTLU4u6HgRjiX029J1+7JWqZVkhzGQ6jYHctfaQxqRPfK08
1VeZ9ljnUJfkUS/IvD0qyTniVmtXUKqzhLHrDYWPiT3FnGXxXWKxi1NYNRUDyFDMD+ys8mjdZzSL
HSRa6KtXILc3A2/jXcgycRKDYzU8zztos6u18fHdPOFC5TMJv3IdiT02vSeXwg/CaaxO5/N8MgoX
Q3OILkKO/mzSKI4lMEGKwa4PnPUNC83jKl7dx7NpAzMfw/hyTqafaKB6OtKxIYuE7tteHLS+7Gn8
TO5RLeuNT42G3sor97tpfNCmWs1LxLS3eF4XJA6S+1dVsCwHU0NZnLIVBpfnTjEnQEDT/mMvWGJv
D2PZYy98aqyMS2iHs9Zr10uWaTUkNgEBrGhBzXOU9E2KpK63SV+iQPp7SKq7J/ZDwnzXtPkOBde8
7WY30Qo53N13Wk24DBaiNUCdOZ/KhpXcaQEsciTuDLBOn90Wechmv/NShANFNXg5lfdIqY/Dcedi
zVjZDz6z53rSoTbuY+EyU/VAc2dUMWrjFWgyvmCSbud4s/tQbxZLcua3787ECpkzmpcEsNzmoUda
a0mdBv5wyUWyv+cYrFj16GPH+WMVHCbnkjErxSFXbfrGEMKQ0smByJjaLAfxB8bAjU8sK1Ohm1tk
zy5d0UXEWap0+tH1Pxbf2U54Wq9PlBoeJvNw5gFXb/I3f62t6St/nWT74Pnbg1ULs47OmR3q6zw/
DVd/uSG/NqLH+eucOcc01ks++m4hDz6QmPcB9wAQKY5tiCDIowbEAeB6niWF21Xoeke05tuM0G0h
IFcjJcUOQ0fGDV/bkSWZ6CbldHRD/DRLv4etux4jJhTci9jJVzVuArckEOOVUr4qi9NiQMOymFtK
/TGzk6gsZJvNfinIINycm3tASTgvjVi1UBV1Y45kyzNWfOeRpnbmxNiL8Gu3wrRYFLYk0+NZJUp6
nRBeYhMXr//Z9qXf8zqWx71b/uSzUATWSbRv0bhFRmddGBcfQPC/ZIBGIFjxXWejV34cQH86wUm9
8gL3j7VDAgqw4CozaxYbZ9W9i6lae+vSJJCWFFndy+Mrs1sJIQfKLLImXevOYMbi8uGRs7r18fjr
SiRpo7hscrjq8DkcXnBQJGdv6IzDyIOa66mWJBNM0u5FgwQn3x7hof5N5a9Gu9VQugJwysW7eK4V
AJ16UuiTnpx8NHxDrrsxFpxS0MHsY1+A0ZNdhFZH02kocgJhKTX2aVRmtPUXmkrEuaNYkngg6GzC
S/QsKe4bBqp7fHfPv3mmHlI9yfdWhehXv/2mKOUm0N7yer7ragopcrS1aPk4xTsN2psjbQ8fUPi5
UmmN2IN8P5GLv8kOXqH/05pRdmn27WdaH7g2xZaayi4W7d3SqyAEqydMVLU+fErnXTeXoEMT5qQB
vuiG/c4dQ/iCnmRZ8mO1AK+tDkrwJpOEECE4+Fny/vmNbM0r7S1quiivyeiMWWEqkYEpWObsGWxG
FFFERtbPIQzpJNXoCeXdvIdUPzsKsI5zbbOlWAKHSuSHM9PtDI/qP2gryMFH+N2tcEu2y7BFS8g/
8C9w/+Q5d1Qtzq68BKq6GwiE5uJD5X8gboKQQFLbq6nU/rxCye1+sJcYWKOs2leQ/Ls4bFpJZVgf
iKvb8FjdFhWL7JFdu5JwUSUYwSrXgVHoY5lbYTFiUf2ZWTrg76HuJmJdm+hqN61A7YP2iZJbprU1
i+qt9+vGpzZf1Gx4st+CFB8KSGYf70gKvQ/T5TJCFZWW1vjQQrk+YEgeKCWfzIgBOjMRAv+NbjLw
O4jdmUqlbAEPg/uboqoZ2NsQCj8LEJm9p9cXSILixamunt2RScZXMPuozXdNFcbmrRn2iqKM71UO
GnptkHanXGvyNcq+6kvYFz+4LLL4Ne9hLpW+3fl8NcW3cX4KuQEERuyde407FxiFTNGXfQGI8oU9
7+MY+GzDRXxhuPbA2rc2YygTtP1jVbzkJvyNNnw8Ga03+mv4X2cPDHNTIiU=
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
ECP50VMN7tD3OXeLba6oTZ+brq1IOL+0jfnYWoQpgwYOqPBm6D6tLRw57u5HlgKO
Ql2wuD+UdDGdCl9w0OM97qxJDnCViV1VpDu7Z82a4e6Vs4f6OdkIFqun0ZED3rz7
7aLtvtJ0WUgBB1DMqY8IJ2LY4Cj2472sf6P6tVgMhcw6ZRRc8vUaR+ib1CkPm63F
yUzk32HzofIKZpezRJmd6lsSJSQQxqT+0kT4BGalGUUNNSW4GpYbtZF7PSg2Suyy
EZC54IiOqjItFVEchVwtatmtgqyQmUj+9jjtz6Jt9b4MJE1WJrhjXH01OxXdAJtt
QkHsRBQ67fddiQgYiVtrYA==
//pragma protect end_key_block
//pragma protect digest_block
jz6mNKD2hV5qPLO9Gtn6rUWxgQk=
//pragma protect end_digest_block
//pragma protect data_block
ECgDZqJeHGusZvq+mOil6c7KNl7S0jBuwHgj36+zPIdCOwBbOzr/KjWye+NU6BpZ
n3Xzzo1t56ZGgNgDzDjZs4k8JFEaFMa2pYoQLtCul6878fnlVkKNMqmaKmcc4BM5
4EEeWIbnh87vEvXS+ch8IIdTbZInzV2cbBTg4RH+u/14/un/NxRaIFOc/SDrA/ix
0KNeLvt9SWAqRJ5eSIZeoI1Sdnc7LqzNHluID44X6DHkZuUgTfLRrQDFxzw0lIZn
Nd4+UQD0P4Iv64PCLdpZoWapXc9IQNtGLvezVn4tNIqnIlU2mC40Da0tlypZgs2H
5sKQK4OvvJaRgXE/B7btg5vO8epEzeccEkbauUbQKGQtJTrJKExgVZ5CUTgGcQr+
RTTh/ukKu6VkthFapONKqn3uq2DxojT9sPQv+JEagRoDC5Oum2fzV6xAFLDPO3DC
+gpySEgKfNOg1tB/8l2zAI2bzpyJ8tMsM7m6a59Dwih+7Ylvo+Uxo/4qqifwkbiS
e3GWvoafPHZawQZAIRBagERFMrNLSgeWL74ZOFtmBLO3Is0lcMbcQC5I5eIcMnTD
0LgRLgXb+5V5nz4dAahfuIh8hD9ekzdFWLb8/CETZO7kzkad2dTEObQ1BrwRjv/w
CjPljad31fMeiAPB3QI8LZEHdOANMCu6LgiNMHISw9H8OlQIW1g6Jjcr+0U4xBd1
vjlbZDjWxm5T/eD34bU+zim/oklxNkAPIdD3xW5k/wnGs1scSdtvXkdP5i27lOBR
XcVzy167Ng/ckviDv5aj4SitQHIvmFBNGfF5r3iCv3H3SIp5JjLk8E4Qapwk0Zmu
MbBCUMR9ob29IYx1zfHaNOJ6PqnP0/7tircc+qx7TDiUTPY5dRe8FWswC4N8vcuM
34gY59idfKAX3x3cI3uWchuRpRpGmZEqQxmcqXvYBe/j0/BZ93IaUENFyqyPqYEj
w2d+vuRvh+nbh1MgBvayypuhwBGZM3YBd05TFHRLm7rnXLUM+QkJh9GEsLa1zjnX
WkRsKWTg7Jy/hT6yGRmvi5ALIEpvXoBBuAr+P1G5bNJaqtwvxGsMHZG0DX9xA1MA
xy7I+/uJToVGQZhy8xpsRzTjpWSvNEIzr9IY30t/KGWY2OS+PIA+wVOsOWtLInyp
tAZgFZ1AArOw2wCZQCz7dMdsAqTSiMPGnTlZJR6FD8yx3pMfzIwrj/QlujIiUXNh
01A7+Rg1rbe+YSNNV0t9Q1XzN7zr3eUiaDu1KPQR2XnMQaq1at2Xodpa6cTugCYK
I+itMca/sPvDs233Wfu+hC00MPROJtU++Y7qVUACv9KUKlYs1Wn1fCjvALtkKIM9
bbuc50U476w84vCC3X74nfQV2yLsLqcP6tZHXXEqpEwmt9eRUT2yVCN7Qq+M38vP
dVdBN0Wp0Utw+yVehV61WxjgbMgLibbEt2i/divWQbbEV7T/1xU9/zjH6tZyyJjH
ZAMBiykVvF60ctQI7u3X0c5i2gHlhAJ9R44+ov7MQVQLfvF2dIWsqf18DK7KApKp
/Hn0jMn12W2b7EPKhPQxKnhwCHIwGTmOs27LVcmM+YrskRIC9hOejO8i2MQbFVqI
KuA5eYpbnKkKwPOivl0aj1KhsTD4KXBePCMlB9aMGw6BlGMkVygKPtm0Ezf3VR/B
y6v/VqcVZLYLGdu+xJZsVEV8DFawEmm/uxg7lpr4h0JtzYYpIVNPBnBqqZYrNrlL
zTy6nzv0ct5vVLO7c78m+SKONtOXu+0YSLq5G1Mh/yTf6hyRSFjSHPqgUBk8sKY6
MnwMlHfj8ZLoVBKpUok9allVFumuclxxiKjGn9e3c4xzGHMR8Mpy4OVRHYd5Kno1
n9zmANAVR5qcez4DtRZTp1sopk+8b3T5CwWQZmjU/Al6MHW3SyeAm8H2Q1VoGpmc
FX2kdKh96oG3CUhxykWFIJWDIshq/UzbSxAHp+reuNY1t0A5ARrSUVPOS85H0Aej
IFR0plMGp5xV/rrJHj5KSMv8XllpQSJTJEJG+1qu72dMTKcavCAGGhn58tGax2yH
4skLxX4TlM7AaWz7/W3N6upMpSdqPeJCBs7UNURdCqAqelhn1gNVJ+6ThziMHt1b
8z6ejp+JVI9QDontuAhTLkuw3FRDUt8cEwK3roOhO7CeugfmGmKMVlC0Y7rIXAWF
qUbGQ6feAQMaU8oA7+AU74PQuCgSsNIYZvCN/ts0NNeq0d2X14gvheiDRSP7+o4z
FATlQ17JhmPwJFJe213q1VLcn0jEepxaGKs9hZqMaEwky/FtTRY1Zl/RVk625tso
Fpc2vOuF6Fmb2avf+QT7fF1FijnWrufA0Y4eiK0T63CwoXyk5O9WfHE3YdJP5JlX
yVakdoAxDOzD5IdVCA4TcTqMxIomrTLow0kqZPb7kRXflVVO8Sv+zq1P2vkH9024
t5Ak9a6v/ROLwmDsbwJuOLFe7TJnz0yB00zNm5Pod6o4XnjTJvbh9Cr6cH7hUgzH
EKOpJJnhxNqLdBQih67D1WMb9aSfbeKsMCXchbGlH+P4eFHaSlxaSZZQcHqXwiYO
pquJ3zocqjYDNSwVkkZKPRmGF9qD7TmJqBZWx8VVRqooKmZ0jUXa2Tm7kW9ISz2R
Z6IKx7wXt/u6PYKzmFY2fRKk8tyPH5+zh/4xxidWlE6o6DZwGjZuhj4j34ffWl05
PasI7ZgsVpSIc2VvDOy7aCW16qMLz12cxG+THbPRgYZYMLrOHju88dO6jdJrqwZL
OA4JcqOk54K3JFKQubH6YXZexHPD4POKyzp6VIyUPas+qW02VutOXstofwEckCuq
Y26AVCECL6iSGZYp9PDyLRM3itDM+tGI1q+eCJMa5xOp0eK96a6KZEkVWzYiIBlw
WPRjpkcWJ81eEPXMdW6CM0gLUs4xL+pBs525wVoNt0PtPNDpMfZekFSgyDHxGiJq
yvdJ71vcp0nGfgiI/uFagM7JSzVNkcaiCR5halvwX+MZZVL8V49KJv2R+6O66Kfx
zwekaPMPySTWE4Lvym5DlYXXXeq5tCyvQhY2QxwGCLRZfQjh2i0DSsEKBQwU8ZzT
dQGp5Q+VFoHAsz8KdiL+l8kyjBq+RbUrXmT9R2DYGhM7PyF1mRt0C3U6+hqezodx
CfKKhOe8jDQ+nwtY3wVEIQg47Md0uNm5UATNHDEjcIeJVHBjQQSo4Ikw5U1t0hM5
9x97AhdTh1pUeT0mYuWU+BWVRqN9FI3IkwoQDMsLIdQXMpkAgiEmS1aIInIBLQkn
7hV5fdd3mBEOGDe/vmEozq/AXHAPMFq1yaFqgBdkXQ9AwcRzqbFTUecskzrsJlpz
o51Z2Pf/FHQCHy7R8bCUf+Mbu7fwNAkclUyd82bIpxuwRzDkRakf9vHM+QO0w5L6
aDp2ZB9QfLSInieVpXdInfP9Bhhb5bEM+zPDErws5u/Ada8NuquSxm8EMH83aYBF
9/wQ5QJWDn3PDhAmptA/xsWC5bjOBYqeo/PVJ1D5tA4MceitjCTNCv3TesEu5NF1
SGVb/1ComOuWCZQoXs6yNbOImzR5zy3AehbVQpRKlu+HZIqIAgaP6FzegnKQysLb
DqYajdyQgg1QW1huogHuAtF+NTKKiWDurUy/mNqCEYqwd2EHcNu6EVCCvqaK/h9m
uQoQgEOXDOw2tkiMPYEMJxRsJTg2dTCPBFxZNu9cKpGRgxe3stOMwpUKxkHX7iCJ
ccrsX5V7Z0IH3YogQR/BEQOHSYsf6IjioKyfS6XmTxhESQfNKSI6dXzllVaSNQVs
dt1OcGczo8MfynMMqBMdG9QeL8SgzvOjS7MDdN7WVHk/bJtOcBG2723wIjsERMA6
mFJCf/ZUBTuG0Ak3FuDV/VU5cW8LfX5WRy3TFmyRyA5KZmirvSi5vbqr6zqyBcIb
hr7J89tc3LFBBtlQWZdo7VcWb2Smo+sQzNy2jHyUyUO4nZdm6VB0FzUfmVrod4dw
0AOeaeh38+FWLA3M0qs7TqKq5RCj62BoOqCkTOLmpl53lB421Fevl1P1Sv3ZV77M
FMeDWc59moMw6H+7TwipWTkz2JXSKNfXYd4/h8nsRij/oC+jwt6pLUlQHjZ69a27
VXA3rt/o4UR2k6qWvk7jkR8hhO4YasrPPTLqZkT1byabop9uWsHrRWkCgQeJayg3
nrt7kWx5qw87Rx4u4l3xjMypUJjHHZuKr8wVTVw5K/KBsYS9OeYao7g5Cve3+6Dy
7espYfRQu5VCVfl0mbEVxHYFUrWCr0zDhsBa4C2Kp0qkCClrx6CyCBBC5baWHZXT
p8lJbRLOF1mjq2TVV9kc8srGR+vT5g1CYTtLVyrWPUW+gnyIo/f8sJqcgoNB+XQt
AsOtGWUfh2cdzL4H+mlCrirSMgLDYmj9ekjC3Fu9muVDi+2S+90C3zJFMrtfvr5w
frFkSOw+JWGQbBWCvZS+diQqjSip6OYnUEdKDibhq6eFPZukIVP9G/A1f9+UFjIl
1TJe+NaLGEakiKhUMJTffpeMKZlEUydY5b8gDirMZ2UWIhGGVeGu/RdTNGtXI4nY
0xm+vsmgmDi80D1fFjbbSjZkKOcYGrkdZ3sL/YykWuap9XEzXNXAy8btFqoseUth
pv8jeDelv/RBC6cgnJ4bLaiqeP4h+hMNBEBn9dt/W0xZgCF4/J3hiQzGpCbC5+1c
9Cuj+jQR1aTZkNE+IArAntHHLmwNtdKfsbVMTUXAxm0Chu1Wh2W2TjLhKPVMHxdE
1tgQHn3n28SyxbDuMqbLVCiQ6s+Bg8L3q5HkJWp7U5alFsfzWN35krr5wve22IpC
Ck54BRTjFBtmnWlsI2U+aZKwdzPDz+c1UqCXbL7jnw4tqY9vj0ORc3Ce4s8Be1LH
9E7rGGpvhNMyxyYqHpwTFrOAPQwdCVgrUeBZeZ9ZpuiUz6CiXp25buEc9NcdiDXg
qY9Wf/qAYc6adtgv8qh/wlL79/hzf8ee4MN7e6t3JZEb4lZPG0ouTHWsInOTi5c/
dUWPKjSEx1LeYb+Mpqq2z77y8hixhWQgGhP+uvh8Tsm5YKHll2UhmJjQ7AMDJzZo
PU1V1GhYQnO9UT6MBoGz2ROzDQkXy+EUY0QMex03kJwMWQ6LFLQJxCcn+ZHPRdzN
nEeScRCjBF4E2tG/hz0nbE1rzPowSKC+v/DJ41O6mihdb7BjWJi0IK6Vzorba2tx
gGErawLXZea1FrbLKGrjCgLeTfq8eEmrCSZ4PgBomlT8wZdPB79dbC5oPNJgOKo2
l2YdnAxctpQA76+NPQvLLsDU7oR3fk/CLhyXyMWmEvZbO4mbP0NBAN3+TiG+1uBT
Fjv+VXe21bf00EpsUWowh1PehMFu+CunEV668spzZiNuulmX7VrlcJXeuNjBC05/
aSIAJgYw5Z0+REJY0SSzMVrlA0tLG48fLN4VRpsaJeYfsTyrcF6QSEdqEzfX5DKh
W3fkf92l72auXjq7eCckL6/zQhMX77cGrjpeR/SZjoJ7z9Bm7fNYxEEkwXzx/v1T
PmG37eBTFzGc0Q1/44sk51MgnZ/BcBbjovx7JIjAiEP5Xxk7e7hLmAxG1PQDxzYv
yzcZb7TBKFJoPtY3aDoHl394pwEPXfbG6cntE3+P+fyhdEjyI4GVxaO9rQw21ik/
+WVQvLsPBkDvmG+fC1trvyw7y4cvL+tkGIK7V468UfEJx3nzwvd1hS7SUr8ccu41
fuBi/U3YBe82jtEF4RzGWrZrxlfce3WixHwPBhic/cw9h7pl52+oRyMY55eGmq19
y+Ttkt691gDTE/ub1PlmOjeD1eVVHXWsL3PlClJnvOePwthGmmhT0tAAb+w0kpg5
XZ2WJOrDSDH0hmEE1kehAbfDbbIRSk4Y0Y2GbAzJTeNn5zI5sufPO1LaFH4ZX/Up
trH5hp6H4UCgrB/NXCI5/7167Hk96JCCPovCDGL/0SWJXevPBxTA5YkZ6JmCI3+Z
1yLDSc6felrhMG1mhXyw3aDhAdviajX5msfzVzWKt/vabs61ggrStu/qYyPwfdsi
UWwQ++6PsgZ8DBavjWO0kl4JviMCJkDpH95gH15cLyUzALUqntk1AX20xCzJ/6E+
Q89TRIKnEgWVMhTY4pqzrOsn4Hgh2bS6tP2AvmJF6z3Kme8gLU6MvrF8N8/Mtbdg
3gufvfRKQmpkzPfA/pzRWCG1VjpCb2NoPfVY/DvWgzvOBuTAM0QX7QWk9Mx0MvKp
N2dbXiaKPibBRPiKMcBMK5yuBD9KDttXFCPUelilI+pmnW+jI0lmq0k6R4ma0ZbE
nnIvVInRv7H+1B/l1twj93YbD8XGJ81Tbna9ZV6q6O0zkBgU38JPSXDs6SKhWZFS
5wV7MBm/PIreSRGMKCPCXNi2cqtL2m5TbLvgXRUKRtzhrJX4ZekSotD8pXRcxVOJ
AyUH8NmeYn8mGxk4mGsuPZD/IWZcNJYICC/6OYJi/GUnbQxKP+jRZxTFK7ZfY1Wn
EKHCy7dyTopaV7WpQ4l9JZwJABSvqxtB2BfLRIETyxd5T7+mq3Nh8hcqbGulfnQ8
xAo4Osqlj9WsApzXTpAvod7b9uzQtKcRLBKzd1960k6+k+rSWuy52oOeLMlJMLrU
4N2gZigE+4tVkA/h+t5cOLPBsKp6/thXij9VP94og2RkJc66esf4tSPloM8r4n1E
3OgvNVE8jXzKKsZ1iD602I+g07wpj3MFLUvJB58IAohyK38Lo1YRW+xmXuaX+r23
ongyCGx1jzR9vofDUkbfwOJ/j+EKKVNtbTlUrRbLiAyZDR1dZtmjjRug8WjTdo8X
B9lkUFfEU7+qbS6DtddOzO+7bhZ9uy3CoCD1Lmnq6kZZ+nUQ84WlSFyHXL0GdYTv
/ino7JMBqM0aMqy6jB/881/VAhsRKQ02MZmNVX14OpnxbgN28Ar61KlDne0+R/R8
xyYqrDBaGSbmsQLDFqad47hoHry1e2V3H1iWFwEQGPU=
//pragma protect end_data_block
//pragma protect digest_block
kzjby2bEbl+KFtGZLbKSPKIadAI=
//pragma protect end_digest_block
//pragma protect end_protected

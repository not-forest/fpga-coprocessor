// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
o2/InkgXOhhLNeRGkmnyURTgALGogH3LehlLFporyqNbBfZeqdo/rO08tUzsJSmT0VXOmMKJ38Bo
VQUaGRbqRito55hVIPkPu2VEfkYX8GF2XWS6eg5jeZUqVfGVdK78G1Z1lff4IjKL21GImQW+V1d2
AE/eYY6JQzOOvcHyEZ9F9Jvbz7qeznEVl4iwyIykL17WjsmUjmsnP9QL00HhGLt2iUqLHPB+OPvk
yVZ8Cy8fGShWtg0v0OrYczNDaiK0f3fL7Iz4cfnG82RCZNfVYzGw6YDmkEtVggI4dR4uXwUdfZH1
UDkyIBtPo/V8OiicndIjD9ThrbuYh7SCceS1AA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 6192)
WoCa7S6UgSTcKVAUIlGZqlOtYZTPz2xk3YXAe0QjISFEEsLP+fxi2D6UezpTtBq2jOlHw6tuT7af
0ObD7HnTxLJQsf6Y5wA6NTDOB1wfAwPlA1a99i6jqZM/Dse4PGETlJsD8D+RRaTA5GaNA/iPfeCX
ZrsFP7dK/GvOu+qB6x9JuWYD6zEaXuDvGhn4SmQczk8EgfWi8kd/6CbS0lBinhvniwY8JI7AR4E1
EpPkvsshqul0V9QsJQ7W9dO4vsdtO6UBOC30fBtDzgDSB5qRC7RGQa1L96kQLKywq7UmB0KRyyK5
HxTAN30DbIU/NwiGXtKqUZjtbVOHBcn8PBXLS3ntlFmVhqxtH+3ARvz2aSvuX59XlYDasC6r2Q66
1jkGK5QEg9fe32zheDOYD394Maj2GWOeQiYdllRYW9l6d/AhXelDG6/dwXsgPXoC+k7Ndd5XgaNF
BUuuhwn6nms2WMfpy7ycn0iA5BRwT9K1T8F3DFbXbxEDKsXISNuHR+DG76C127ypUxgXa9B/mm4m
2iG+UjXDH8NsFT2uDyXFh5V8nV/HaW3Ag2vDraTxqB2LVwrPHxKk06b0HNWJVPTgkYMZvdtqin4r
u21Z7Fgw6MTPyjZx363S1t+6lIKi0KBWnld93G4I5j4PUbjcEmJBwXbMTLlYtBqloeFLhQQ9vHUi
tliJ1cxYq04LkRxyrJ7gHfy0lmrNEnzMHxWhGki163VbT5+emkBmYNJyidXlk8E/amnlq+53xJSW
8EOCjK+ooF0NNA5qyyHl064izqPPJMRTAtUgOxRMS40gjYYQKtqDtkcZJALuX266C/4p65xSC9XJ
uV8WyPfXKBKUWeREtZeBCxU+SOEqtYCxX40mqZneGF6VLgoj8ZxLKabWzmuJaica5ah3KJr7kz1N
yGcpgK47zm4boOtrOejANCX+V6AA0CDO6zxFGPtiLrQtptVhZAzcQMQ+VyrsTdvPns/JObXYhy6J
qOMyRTCdmbzOixla8T5f2KY7Cl9LoK5Zz5k9vPaxZFOIiEnD8tmxA19HG/LaAkueu4yWr6C9qUDB
EOi+LS1q9j9EiKYdlYPpqtDu+1cC8mUqsSbt8359WoF55HqOBTbodtEuttW0Q+HL4y37ceZF8dpc
+MYVuL9ALB+QFddfiiNbDlHLCEW3H8OcNEGqxt1U8E0XL+JFrGynH0BORaPBTRQK/YiAKMMJpKJW
lrCKBZ0/fxWKF6EXnWH+FW6lFbNEGvfNq8DBjyrjy2koGRyjN3ZqcWUQiI9JWJ4WEP39eSih8MOq
YLYu7IH9IonFz0sIGIn+2XH6CDPcXT7dsOEPS2GV1g1oahQcylz+/jpTK8t5nQbsSUOkFCwiwb0I
NZAOUD89Ar0LkxhlX2Zo0k4KohHtna6JSEcAuSRZAetGey7COH+rc97alOFcnuCN+GQ7dbcQDt4s
fCl0AA4tTw3VeW5aiHfTYCU6+I99Q3LNroOE+60FX9BroLa3TLKlepE+/6kmX2q530DWoj5ZrDxF
h69DF5gpVCI0LWMmEhiwXsHos5eZcV9OqVhSgDXR7CeYGJ4DDWxNyfeYhSUMbwBhKN8Lw26VX5JY
YtbuNKjpgFJ8oPlpFvja9FzTC0E0VFhVD4CNE4puW7eyLSursMNihIGsoKaYTqyFEXzwKpU6UqtH
FiaUVAkGh1bL8DP+Wd8LF+46c6IIFnXd2F2KEs9KB1hDV2Lz9dNxI+zdaaBISWAWCx2HQ3FvhdY7
LpHPRSJWKtsDp3hSYts1FLh/7Hd59CFNE03EolcrH3r8ZkhaKb6G4IbHcop4M+BCbPRmEveDasRH
tbAWZykoRUfvBAj/ZKHp8GOPW9cXrCkyODsCfz8YpnJh58ZfuKb2tQ+HOWKSAuqd1FBgtm7oanv3
sFU2pcyphOKaVrPjxGqDzclvvGRptE0gkGT2gPCSJitxMXPZf112I5nFvFPp5CVyUOE4Unw3IVXm
QIil/Pls3/k/ABgvsjvEsp4Wx2Z008bV5oXwStzWXVugLksamgk2bNLg/SEkjJaMlJh2wYsiVDnB
hwy6qI9VvzImmuCahAEOKNrljW9FojWK/Qmxc6XfRv5vJTpB9jmGWtOhz+3FTsqx9vJZQkxIF5oQ
j+qxj8wS3EEw/MoOoPsqO9GHGep6+9aiK38II+p+6OQN75OvTq2Vx4jibnP/p1+g9uy52Gs4/Fc6
yqCmmkzAUOJKovCl6bC/kVnZgAAFb8VhvxhxW5wfOg+5SRKaTUKkeAcKvctl1007VieYNwpJgXIv
v34b+kWeQvMopXcXlXGhaQx3YKRYxi6w9u0FSkFcFg7rnSSyh6U8jimZsTbyOwfQ1A68Pynym62Z
4zGkQGXZI2sm7H23pYNBZpiOCEt5bRL7vEBlR64izHF2SH1DSvKIVHIS8ymSdDHAanINk4cNIiCf
+SU2qWS4EAYNZFCBnwJMzoc8qPFXedspKAUdsIsqR4BS3ANUuJnJ8rf+Fnaw20AxJQfj/qH12Ews
yfSFWXj9uKWCKgmLCd8x47tg/6/XMGJSlJxB74NwTy+4jN/c5ZAfLqQh1eCXg6UNjY1+ITSqxQBR
McskBTGVhkVP74OdOmydOFu0Z8cA9i9CUvBxpXu5MCXaR6wxeCsbK3kvhR4EkFU/6PIy8EF2WC3E
6CsvRVRPGLGcyErtvyKvYO+/Qt2CCHa2yQtuDt6yrMlLpEwpGJzlp6zlc3HlAyOlUWscHXh3asd5
dIyAuQFAXGYFrWMoQ4fQ4QAVhbmtNPOtDuqk9AlnIbjjfVUE7IgcfvSSZ2HjWJINPRFyb9VOrbma
WePOEkjKMLH24QIFmaxxQSKEH1+CUa1ozcZBQPO8CR9drTxwOYTjh0fniqQs9EVidjU40ppTi5xD
32a9hAIdzSVjiNlGpL6sx8sfFG5p4jczkn2DF5Rmd5zJ8pREvIDfrLa7NfAmjwLVK3Z0kgEN6GVm
aPrRSmUVGO/V20o0l1CJ5EmwvLGMffpFJKqfCCaa38Au/YLt/3W1UTQ+CWy0LdWbjaVfetn+MwDq
YU6nnXF44Xh6XRFI1Mac6OQEm7LLbGGaEzgQ1iEnOuxsILBxQylthpv/dMM7C2CudBdMhGjZQpip
KieUBis64ui+rPHzwh/fw0+zrE5mlaH8qSgnVMl/lEZDH/mg5ewv3sS3DP+5hcwyZcmG25ui6pNV
P5EDzsJhp+7i3CpZQ9m745159zsE8wykVF4mC8paY4j4oPNvu2JvkdA+7MHf4URfIUQgqDcvn9ne
/42nU1rivBJIGNO+IMFA9JVn8hjR4TCt5r3ZhuJ8tsYxM7shTs6LslUQlN8Ykna0hhvTzOLRm9se
CnbZWDgztXUVkZBSu5sAZPGYeJVSWoi9JEqYHalpjozTo7qYXLW1uQLZC0nVPrTh88TbFv0+pBQA
kdr9x/mFR7pFzff3a+z358XRniWgC5XjfbHOy1m4R/L/t2kfa1ood4oeLfH41he8JByYDWoOU1D/
d5bIRbIucZ+XJ3Qlor+asrbxOQzngRW9jIXIeb+cpPdHZd6+FU09tQvIBk1N5G0NMURd+bMw3B3F
bp+2k/ce3K0R1PcHIk0q3XSNFRjv0VlD6NFcQ+W9KGXn+e4OeqxnKo9e2o5G76bP/A8Om873D0io
juydeOL8fMHmqCHWqE3VNko8QtlR5/fmgQGb6yDgMJqRJTB9wmZTyJ+dYwiytF8A1J3tPJcCplBN
u/WEJ77X26aPZnoBgweFpmAGDh3JAF9AgD667Ax5u5KfYz9Yg3PPgk4uSJWfbu+PuGZ9AUJybzmh
XgT76Jm5heg3x8iz/k2VKFiYjnKUZvZ6wbCjjchX/7gZg3JEB7rKzv2EKk6O65+MKe+44j5FaMaZ
fcE3jVNBV/Taw2CeUMHteVBPALXNPfAf0trMULeYd9onYyZdP+MA6dIMs9UMdqM12jUU8DrfxTvC
CRopiHfMrx6i9CxR9JFi7cl7cgWE+21jdw52tmhnQCy0S+shIbXAO1/Q2juuslg50ITStYE0KQ6B
SjGjM1r0EfjZT0PpCg0InOXg29SrR3r457+PTSyG8hm1rDyk5qJTovAgGFrnAhGswW59c5vxyfXW
zvLyd+c0/ZOgI/tVEZ6JH+Rm8oHkoPX7Eg+dOiwNZg/tBmou7iGad4WbkpckByMwQdkJW/q6xtaY
MuOBQzjHeyRiIOrCriRbu58DtXc3kuDNoVDvXmqL6p90BNTr4enshmsSNKSTcAyiwgZRLC/q2gOK
NFKsHKHLrLOt1fgK9VN1Jf7PPhk2a6yTxYe5yp6cWEmuVxtN+851rKodOdz20zlw2aWzG7nOz5v+
XrJmEDupAyzz414DhcziPUPSdiTUAccP5EOgD0R2r4kRYbHq1/qWUkwJCWSoMTshs5cakmT/mEve
BMmUpfk2pKZVmDxg21AONeA89fq8bcan/H4GOf+sBRk6x1wIoY7bUgqJZLbBfUcFJkgv38myo4td
JD7hzl/QT4J0IFq40171DMzYMQZ27sBJPf/G54Owjnoive3qWsseEFnjlqnIR1L9licxChK0t+hE
xt8w6tr6zjllsTkoVdz87QmnxCcbG0eIHDN540vJwndfkgxzP7W8q/zPLQ5rEw7/ewnE0LSqc+3q
Z2S3hNDToqvG/8A8lnuKe/gYmpkIBwBkAe++7HkTfoxpzpamgRtga4YdYzbFjCv+9XrHrMbNPm0N
EAHXz4rXxBLPHVdaHRMvGdv0CQs/ibQsDQ74VRTe8UpVsIzo4NpU2SlJ7frpj0n8Q2LKNn/0/YWM
ZIyzG9rnavhHS5UP35NQpUX0VFIMx2KcaNR0b2r86I/Q05+MarvnLUDCg1U9hVSg2eVPhau29PBV
HP3IT026nbwYzFh/+EhCEQ2W2UmXGcdrRFPvb0H6DtMyf1aVtTufy6aBWB5Soif2fFoDN2x505Ln
OhCq3AM+Y37Qm7NzCaqAaxejLq6PuTW7N1c1vacjdrfqIVsNpQOqhCXlkHl/+eKLAafUQVoFjS1J
kon0AZAgCdJ9cDgOZBqtVXKyFy1I5Dv0EYAImhDtDo6GFzEMHvuT3opzdsnRdwizyWH9GYrCdiYF
iUDfFXgzQsQme1rVxZlbrJfwoVsQI/lW0AOZLUip5AnC9Z/PnEUmKChicH7o9zmlPeffR6VEpFOe
jzf9rhUUg7xuJ/69H+vjqG/G3wWKesZt1QCFM6e1/zn4mAV2ddhiOoc1hhc9vfrUjI9VthMqA9ou
s2lDjA2o7VOIvO6/byUNakR4PS9ESZ42fguZhSCYnXNC8xYYLqynvDlTRzCaNd556UtlkX7sZzXz
szENw2BJ8AKCvVgFVR0Gfp8nDzRpVz2AS+Q0NL6JaMZllr5VMIe52R4DPN2NEp4aAApwNHHHIWFY
n8Rdqh/zRWIHGC2jpRT941DPusJrsdAY1HB4fRv2ny0wRas76ZKDEibcGvvQWV6rj9VIzFbXm8xU
GbMhCswZ/MrjyyWIyiiLYHh0V4rj5Ja9teTjXfxJI00z62Gm3cvxotEoKB5uQp7DXllJxegZmhSW
SlSscGvh5c9V0W5KjeAWMLOa1L7MMfH5Y1sYzMNud6iRgvlcX0y90ld5nN65hZmG7b/hfVrHEUwS
yjCpaTscTRBM2k/32QyY2nK3VdGdu8sCyelm+MP6wuh2fqZurCzUHRjiuFLkgsY9eZsZramG30aa
5EqOScZbPXX6wQqB7lo+FhicNFbLkcxwMUYfT7w9vuKHGUYz0PoKZB2jsP4E0vhdfPWpmtcoqWEa
PAmn99MujPsuR2uAQXBQwALn1T5RJwm+rJbPYCLZdcn3HIzUauLTCTND9a6EIRc7d0C59MlH9djj
Z/vyAC570JZRRf9vajaLqT56nji2F/zn18yy8vnuWChN/1Ok5USrtRqD6m9waDHfz1NCOqddenfM
Bc93dHrN2zJyOVUaeL0WKRdebHgYtc422saYmfOo8nxvQbgvIv6UuLe8BU07BNu7VyR05dSu6Mkl
QkaLnoxEHXFPZU2mPLH4BNrBHn96n7NA0ZioLtCbaurYn2sTYk+kX+qvNKpWHGjCwc1+TFk5kIYY
hqBc4oGYpKGVTfnCULqU1zWsZ1nSECRttk9ZTOM1Kd8mEIUN9784gIzqlw5xsdVIpNoMNbkkzldN
n0oJXN9KeJoX8bIcedNtJ71UN+Os5Enns1dCtGzmqzGa5rDCd1kOpZY3YXqzL5kcz9VDKzsIrOX0
eYSmlyjlwfrOm+eqwUZSmSlx1/lRfSkz8477mLKmKNRFgIIsBe28qApnvh5Tkw7mShKkzQtRvrF2
M+1TrdSxah/OZ+hJjx75OYTOL8NCYawr9XtUe3m/XQDogY4MSpfHYNUJ1Zi3k6aTk44oAGzJ+6LA
naTSQBgkzFtniHWzRSu1KEh9YfAatpv+uYiTMMoF9Y4z/eWWnrGpQm11tyDnVySKSd7klt8c9iYM
LJ17S6Y7h6mxOkF5llNX6BMZcNJ5kWcK9DwkyBme4qdqxJvt3mv+5ufImChRfzXP+8nNqvVp5zn1
iIRsCP67rT8Ped3qpWyW3F8UQAEfMiRWjBCpelqX1Ve/Xd8HDnYRLFhTft3ROU+h1sboTHMUdbUv
G6XtU00w112hI9kwao19h0/mBRzV7IFcNlcUix57Eg8uTDv6qCYhl8hjDJAvHdWOZLfnWb5thEl9
NocrJMN0ezTGQF7PnmLXyCl69c2CKyTVxvvbPC+bMUGWBJdeO0z2i3BZ9kr5HsVQKiR4IRIu5hhx
1pvc1iO9ZsUrUXaXa8btzclB0ZEbibOGYRQgYqiryQ4rY3zY6Nyf7mgECbepDvZDVolH8ay3gOXm
j0EenJNfIcqNxqGHCI8/A8rucSgtHUDDNSEj2RE4NWHWjrjogIUrN1UV+awV67y9mUKYmSrxJS5G
uRdOCGpxt468G1A2JnVtgZVem2154cdGX8ImlNGBd/4tPYQeovFYFrbgVOPu0/CxAKaubzo1s8nn
1+LNEBxbAKjhuSFMQvITFtQNnTxjskuLFqhWGd+e5w//CKnax//ti8tDtc5C9Kj8JcItUWgqCZyZ
eJylkMgGS1ckkLfJHA/RpH9mEl92hlkE0xqdazhDr8R46KGTxfU5hnfCDihZ3NH3BJt7bUBYOuxR
RARgoqtfqpSaaeS6koyIVZ5jm9FYGzVRoeVxmY2f/9VZFir5hTA4RLg5YnH7NiUHJa8BlEVVoCDZ
OPszD96jXHxni75jpnC86BDxYi2xCPzG/UllzbzHHhEluUi+DrVONdIW5xEFG62kuqsrZRoHCg6T
FQgY0p9TnW/wu+4P27asoSR+WN6qHVXsr5leASclnG7o2EfwuxfTW4x33/Bbw2uod/jPQdwNgVBn
nT7QS8Ugg6vUXRzwsczfKQkwAEJb928hSrX3OkytJYsQbx7ByTa9rEI3+zHVZ0QyO6tcQpStW5wr
4jLLWU6ZikSKI6dwqjUykl/daqZYFA1T7OK67NLv5xBsmEXRDBnqqbYz3dDOGx5j20NGbjwsZgiK
RodNS0P19mTXFB4Ctz+MwX78wpyl5piyryOM2cZMCLw58mJxudNranPREyyXsCvy2QG7IDiytIOJ
gc3tqfHnlagwu5LAeVpUMqgDv9+uULAgexr9BIEF0MkgQytDcwEf4bjQNA+pTaajvpon49UdU3MP
UyaO3eVI5mRR4sXHDBRI1yZoe9LKMethXP901GalfVDXAVkFFJZjs/CKsPMO/nHh81OquIMWvLCd
Fu/uy2+Qbn5OdFapLCzmYcZ6iSLjyLtvjKfYmOmjcs/lUv9fI3LbIINjNS1gj0NPRhBx+Q9F6Orm
7/TQ5TKIs4CaWLcLBPeRNIPz/aYaf86t7a+ATD1JmQtR/I5V0fosc5P1g47xmbq54/BxQ9UAtVrL
8xjoqx8ZThEYes/7aiEY6GdCJT/JIc1paLZ7034RvmhvsjHBl6uhdzRQwjEfcHwzECEehnSYSy6p
fnlsYNKStOZ8c53jSSvWNYsY0pjd4ypAzTjdPF2DOfOKoEajNs6/sDIPbmB2MtGsUy+QLJ/Fb+Z3
acISKUEmJdrjjsoEGWhzpZlqUE8agEiPayyj1WKGS8ZCmmZDDgKutD3IR9Iui3VlAM91YWFpMUbm
7mMcvESRqCqGvgWGI+ZrAOuoykFRxr0X+qGzpI5SLlv9TS9b7NSsh3zW4xaVdGiNo73EYytf7lKx
n+DeCG6zETpYW+s66Bq3JMOpqDeRu5d15izK0r1Y0uRYQkRc
`pragma protect end_protected

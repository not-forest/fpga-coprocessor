// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
RtUX9VW6VStgk9HRuVtWiSt2BDpG39zqFmS7dCxUr6Xvol7apfgsD3aD1x9q4k/i
6BFKeIvacqBUA1fuihCCE9OyJq/3HNUQGZl1qjEdFXY3Fs4HsUBYgb6FYfBa1GbM
eXQz5V4wfxnd0Ix3597qwTqhCTIQSp0jikUVlfc6cj0=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 6192 )
`pragma protect data_block
GKcMDVtSyZGVbMHqvH6DsoXyrP7TeXkhaZH/v6tB9ZnUew+MHUWmvsN4QNbpimO9
Rz70paJJyYYiw3WmLYGohHl5aekJ9Isu7TmLawaiJPKUhL0gpReJ7tjwclh8TFGk
qPgqUCjj8wB1KsA9PBBwzmvG3Ekx+ll9QwNYPtYEqA2FFBHY/jocHXTYDS9A+2SC
eaBQk2b+mvmKWq0Q0c19xPD8xo3mwsUWfdVR5avROlujfKj4n2Rks35NlGtWj3Rj
MRywHBJPTY4ehqYs4C1Gvjxl2+9C4c33KpMfK+NO36PIPK0orweWGaGohUSCbLoL
XvNnWBPt5wnCSWKVQ5RaGgL8a1KjBRJ9sNPTdxXp9mmIHsfIeN7lfLBw5pfzxGQB
xDwDDjx7yUcvRCRS97rs+v1XM4ZhgoP2BQl5DfJpmp/0fhlF7Hiy6ilyGg+HYJFS
MAOFbv4jxAc8UsAQxiJKqqNQyEjPG8UKvh7Bb2aTCo24EoMSKoHqJu4tqYLfq3xL
46vMGOGXsOi8ELLUDv7blnNzP4f1Kt2sfyC0HLE5biGAa8NqorLYTLF/ZWn6Mdn0
GC7Oq6spak63v1enQSAG6penE9Zx6lvT+R1IgRYGgIs6Gc35C5MynQ4jeYaVUS3A
Rd82RTV2gWh6OXkJ9Ekw2Vsdk7RwGoUz0EnNepnDdtEUbOu0wPE6Fui2CF9UfRhM
eAVkIcB/I3Q06IhbM75qaOQZHWvYFyoKuz+4KOGJ7YeoOIMEeWAri7/YvkNZq52n
WBbtcIy60fxm1QEA8Vn9tArTanN4R9ItaZGhujhSbdoVVqt6b9qHDXuf8FNVOZmY
PElIrZeJ4y7ysU7crdDNA68hFRW3uYyHZCidd0m3vIrG/mVHFY3QgBH2Qwjduhh9
dqq7+hKgeWUuew7C9iXFPd829mDoyGXWbQf4OHG6olNBTLVGvj4y9gGluInigA4W
5aKlmX5s25p95l5Wnh/0lSm7bHL7pU0/ovBUXAHZRSAbN298rYtIXixSMW1QyepQ
fM12BytCgHG16SB6N0jbmLV68cTvxtm3HWHEZSpTpfs2Y0eT8KchHwPfuZ16VSF1
bhTKLrB+znFe/+PH4tgX7PWzpFUqsqLnPxLXZMaO1KyJIUEjRtTcuZ7LQ17yEbZk
Bbhp3sGy0a2AVFhkUEajr1nGCOb1x8KIf6Y4q8grjrzhKoDF657hIZYeaSA0VKJB
OHLsQdG3stwR3sBqgMM2D+WLRbuz3yPPvCdc5vGQcWlNRtSPTF9OIyG/o2kJ/uzs
FACAV9Mt13JzFj+fKLYrZVFJPhXYbhfkWximHj/ikHg2sO7KBIT89EfchajIH3cD
wavxSV6q29xJm0yiJjaFYTlK+NA0AfJDmzgVyltaGQVkEPZUcDJ6zRkP9ogTglWm
j5v37MURsJtikC62WKDoAt5SISDUf2586ezfr9kEB+4aczStVpNFIJSSlELN73Hv
B3Z5xCxd98cW2WEGKboDiSBTHAz4lBgCOfXBMm28t7FR7XcB+DXFZ0j+L4Ax+vlb
nalXXHlICgT/0Jmw0cK7wmi+ZtwgVBK5I9dwPg/H654REqE4DVnlg0CtdifvJZqb
SYXBXFV3vk672TkaWlHPg21Xueg6NcxRy/IKGQPxmdFq0AHxfCUB0ET2rtBpGj93
Nasez6cRBuwlUmSEko8CY0cxmmrUa0VI2iZHNN4YWnfqNpE9mhVcflvk5I3J4z5T
Deu1e86u83BbJdzLU2C7ObQErqtHA3LC9EiBj9rszqXuxC/PaFsABH3tpsg/erfJ
b5y5u0elNIONZXeG6DU6XeB4Onh8wuSt6eNsloHYRetKWt0wvpVs/tMGdBv74tS5
0HTnOEijxxBiUYn9Y5UhRPJcNpscbnfQUm8gz91MxZqUObTrWLG9Oh/FidrNb+yp
qzvDPfNvr1hcVYf2+N5STfUWm9YDUaKv8Jo7lEWallCTfomK6fLS8PjwCCDXMT7N
CHalx0XwC5y+stozbUfNFtvar7RUOeLjngzP89dsl8qIXh6JkKWNATzlHrDiPLVf
ZsSZ+VJsIYqFuXyaVFadohGdIyu9BTKvb+fo6WOWvsDIOGzj8Q7CNBxc9bckyfL7
5YFcigkQ4Ixnc4HJDzronqrt4cIO7DX49J9SJS1vCvJH9uid/GAuUlH7NmHXqgnU
TN+Uoyhle1C1vhXIj5hy8F42/bHoKAt8Q3dPaPbB2mvDm/Z+NpCkwLXImX5iZSS5
XoH90p9pir+nXuT4fQiD+DdYiSgGd78X2rYL+p3Ew3ngQiTZLdPoUy2C9fLz1lVb
sIBduBBwdm+LIcdFedl5FSIXdbk73+WTJVU+ewl6RGQxLbos0hj3tciuMY4h31Xh
fwq27j10kHw3jhqHpKvD98usFFS+FDwClW7Lap7B+8kqjKXQNezDn4EctZ31a3S5
RxN1EnvACRc2mdCfeM6EnjCY8bhiQHaZA4+707pTXHddmff8hEm9RoLLcYTS+Vr4
+b725OLkwYZAx7jktU4snAA6nJ3Xnyr9dKckPft0jS9BayxG0BDs4W+BHVNm3akt
Wt2j4JArSqvlcjwBo18WoNurKDF9nA5UOpsNqPbyx0k77IvwNaRWMSPNtn4p6KZ5
EEPlGCS3g2qn8e7PRTbl25hQon+AFzXkqi4p3VMmPYjiuYT/txwt8R6rvc55ndA4
FIe4R+kqGMP7it+vYMn3b14AaWor4ukgjV+X5J//cEOdAJ3dN71v8JsGp/3Bq0jz
wsCQ58t1rPxlDdVrVsIBh2YGGFbcVov5r1Hn9VN5xdh/1K6TpgjRzz3WBzetszfV
S6WYRaTd3OQ4b2dK5P66z0UcNjUKMspxUxWZb1fflxg6WE05YqA53tEGJv9eKjeg
7OrfOkCahWQYnBx0Sgc83kJ69NLWNW2VDWgI2OQfpUykoPQb843D/rf8rKtS2gZU
aoGCY/ojRIPErEaV03CWZ16ZQobFLnoLBFDR0lElcgSAadXNvnLm8KJHr/5JMIwZ
58j36IAycBDYdfoDdQ9ffI9P4Y1W6q3bIw8SsitOo6JWeQmcydFn9SIBxShITaZv
ShgcK5YlO4UdmpAF/vnlk1Jel7OJoh4O5Q1UNHhqMQnqjBO0IMQ27ibc+v+Ww93y
FrYN5w0XNlCa5SvUTRSEFCSpTzsKt4d4I6KF9ytvitOofAMff/qM/Aa4yakhVy35
SkYtNpQpeevTz/GS7WTsNLeID0pPp5IbZICm0MRHY+2kUcDAQ8pFWg/0omK2ZO+/
J80jIhDLdSSf54gN3iPabhbNA3yW33T4INg3aiYERm/mFNpMfbXETpyLdUmrnD09
yf2aLVDiI3utgdaaFlI0IuFQoSUEwKOBnzlWZ+uoWxjJDBZOrRhqUovYrFf465xi
92ckH0DGDXL6wPeCFYUmLr5XdGnVrM6kiYe4H7zUiUQHNR4rD+8daf/K7t93+ToX
53Ja9q0SKGYJxyeS2DmqeGWiO4hp9dUUIWfCW6sQjNQonidii03ZP3Sm/LzFtKB8
AxVmp2n9IFIb5YOjGLyipjVtnUb16t9wvrLWG29deNKgAVk2flNHzDYwHj68zNKi
QQKX3ioZnOmnhqT3ksNnA54SCI26DLY/rDun0OMYwwYN20LQlvHI2n6G+2Jps5jc
5zbBgT++oPaIUGnl1ZiMbDU6myvhzll+zE1Emi4c1v2FunjMMfUNItDUjQrLNLbT
Qm3O9HQhROXld2nOwhcU7P5e9hwCMiyyiuGuybbIZvsD+EHuWswqCt6Zd5TRI1Cv
Fss8WOVQjNk8xX5W0yliSlWXd7mq5LuGSYoHtIHEXiMteMaMBOi+U9tbAdPfhVXU
RTJhc2W7sIsFffFXjRQeX8Ru029HRQW98wXbEQPTrSgRCEdP55MjtURTFrc16lK3
lU6hOMosuG8ER7ey9K54R7dZdVdevZXX82cmMGTe4RD+6I94WesTjvi+pq7SKYCH
AG170WDpdkKGZYKvPyC4JS4RbyLkoVkRbH+TPbiRw3JtTnb7zrWaUnHCsA0Slmbc
5nlV1D7iYldcsBdQ2HLc8mZ3AQeJTPrwlj7ASxwR2Oe8iguWKA+usm29yR5vnUhm
x59LYlNIGytFWzUAjHo5MLvrdxXkaxn2hPfCKtUNu5fxHD8jLtyVh2CPpIv/pyAL
EY5IbQSfeWC2zBhE//G4lW9099mgGC8XChxKOE7Em0/L0PX3/OP0VX8SNC9GleZe
WgO3VXT1riHHPgS/99TklTgDLFT4JCkN4ZEB8oGpQq9A2vRMqZPFixLFvAesvItF
FbidDHON52/grf53D2n5HpFFwOwXUEKFY2jzcVtqwq0b5xF94DyZiDCr53jdIWIC
OWor84N5zD+YrQQ0m7zTm9bMdCe0dcwi836/ss/EQs6bdedUQI6y/NxOsUyUgp5P
eqifx3vXPT4hObf8j3us/CCDOX+ySbTy5MsURhPAGlbl2YSl/rmoEZDGixrnMiF+
25J8+mHqkBU9+h5AntQlIcM/SC0v3oVNQDz0Pk976Mr8HCL0/gKqEDeJfu/i94V6
vTptKQW5ytoyo5+8b86hBbCtVleDDGcOfCu4z/Cov0zXHlK+nVCz7lr7y4969ep/
EZYvSCwKhfC5gVglBXuNue9dIyTI8y/mpaQ2ZZrojLYCtYKPfAuColSlfzB7ZqNF
1DxhvA/CtsXrUQyTyQQPCEgHs0BHxkFEVbhll/fthJ9C4jEwyyMkWRv2s8+ItRkz
MTuBd7X1SDA9YIKOXc9MEYScal0J9yZojzgh/q5z4/P18vJDXySm0H+Q1UyIcO4i
bbI8mYx01SjgaXDWzN5aCQD9RwvtwjLLw/XS1n0CL8SgDlapgzUfXKkCYYPXofXC
3PFM3sm+WCHnJVSaBfeLF6SrGzbpFD5j2/OpvI3AACOHo2ooDViMJc6FhVw1KYFn
JcpkYaICNqfVdkJwcL112Q74pUP4awZnO2kFWC4r9omMbL8oj78zKO5r+6dkWRlx
5RHoh2xcgvNHJC7PXmVL076YuFQ0sJbtLFFlg8vlw1sfvkqHdRr8nuDyo5kRXcAU
tH3aJXmOaAweAKrmDgXhBLFXAwqxxRXTSJcKU7U7IagsavLYRjjVBZs4/LQCeUy8
xYTqtqCPH184D020YhTnI/Dq99siaP/1ILSbdWvqztu4/SNexQI0gs2RNZ0ZB3oC
fF+QphllhrdVdi3ciV34tMNh4EhM3n7RbjH2bXG/305yIJ3UBKHDD6VfNG7LZ6Gj
oQKQLI6RzrtiUCsLm3SFBKx759D6sbVfco2AqR8gVIvFZ/x72jAsADCVAO5FTLyg
AozPYUiCsUQ/hRuVo2LlUy620iBvpjqiIlm7YMgnowm3fq7P9J6xvP8Bnvq/Xtm+
njQn4KVavcJKybX6aSxQx1qYAQdjD1MoTDN+B6PA/sECoqI8WP0sENYRn+nd1V0b
NzIVM12FIuGOSuPulnLdRPJfrCOzB0vLOfvC+GgDGhUF1zFgpuX3Qh8oQFuzdlBD
Txjzpypjhh9i1zwflQ6Gi4YM28Tjplmp6D+VAs9TWJsNYvqApMPJk44VvSJcVoNK
JNCOaOoZhfZyDOZnyY0cg8M6Rtrcq4XUNJecVSA47E0l0UBenGDUUD8EMJOJ7pOk
PhYqofVHK3GkK2L/KI66hZfMfmoES+Ih0iQ/TA7K7JkDo/MBBNFY7EvAZXA2Okzh
U05Sthy7cuqXUUp9/ZlQtg1UxuzpvcFQ0ikIc+e8Fhk4s7sZOJM4oymaFl0/VPxK
qdZU1WpXdK+P/+8RRFAQ0UxZ2gd2CXZJBVCS6wA7HQ+YGzTe/mfq0z4xsAZceubW
yoWafa7N8xZTyNWbQKu2wb2CiDZAc5PtBrrnXrLOvPC/ypRQ+vaTDS9AATKLq9Sd
XBbbuM+ZA5xlcHQH6JE26Yb8RzI0/ssTk3ND5h8652c63yd1dmeOne/zamPBefjF
awfWDU1qChrQC+3dmzrtMQE51BM0K5hOeIdEQhCwjfO6P5gi3SevidExk38MSi4w
ieu9T4r6ZemQtrqca6rbVcPzpp3FZgboNiyaunJ9BCVKVSfMjvfGWgmk3q89gDLz
LcHS8FAYLhs37BqpbSGTu+uJjHBqtLZ0nwCHUgzXvPbwyg7RZCX+PbS8Ouaw6Fbg
trYdLuTscPOp/pm9PHnevWdIr2cAiXx6tbc+6ezlQoD4liTNVD7a5//wb0r0GXQ3
7ZkSTERUmV8FgbFUMCUntIf7iHY2Ptn4XaPkslcMOcJ/5xvFxDTE9qKC/vdqQmUm
Liofz3LZ14UltBc1e8ODkORYq1JBBrffwsLq7vPjlGwKwlm07l/4yWklv7yTAj1W
qsPbTcmyVauieFuYrJte4l9gMT4vvmMZywRQHvER8nxFEDgN4Rwmu1/c0gAwx0bV
i/Srq/TztscBx0RoqtiI9Hw5nVGfVYuqswFzKVPMno8wnnXNYK08sGil+bQzZXwD
RRvhzXzSLtLib9gUCKcFPa0DLXrbEzAbncnOz6smSTdK1+xIhqhy9LOZfgSPaaTU
mHhcSovB2D0nxS5QqsYEX5q6iNV1tShCm4AEyPAbKE4XRKusqdZunhiCpupRkqeh
/G4TMwMHcjPq7+PeWzTK0+Nck7LaDtIYmgJAA7Nz2F5POF5EE/pfZiGX8zD1YOmQ
9lftgBPZbxkA6b8n2S9LZXXqD1jphAfks49Z4yLucN7BcojTcoTFYdV3hRn+jw0A
3SheSRm7+JMAz6iiVJjDSG+CIuYdUbd3eRuMYq9d7WLL0cSsHkPQ2/OY4zj5Mw52
BAm5ZKqchRO0x0OC65DbAU65DfF7zOCIhkh/xKRJBzaX/fy4eVX4rrQ5VmOCDb9B
RAtsB8qMSoYC4prqZ2aqpgtYJmbfcLyL/wnor6t4C6XcILZqRbpk5/qnEJoVE8uc
Kt7NzvynD/Pn4fJVlNjAV4wfvmaM4340QJGKW70EVeZ+TIpr1sAbVTo+JoO+m6Fx
c+TADW4zMhQgXzvA1xhA0vdAPlphGdhGIH8cjaEEhedk0XziVO4E1h8u7cxwPhBR
CpqcKStWNj1K6STMNaBq/+S9sFjrlkb38WWuTRO3KKJrdwKEByg9DoFtqqJjRvcU
Qc9s5aoZ4jnoMJICG88t0fdDs0jcAsIm6//lMszRzNIuA08mmu/J0J+fN7EwbIqZ
9D8vPrPyaNqJabcwJKtT+QRfrCXV/OeTP4vzr3RcE+8dhg8iSqUhRSQOlw7vySje
3a/b7dGUxmAQIEwxPk2H/uQSFv8hRwI8Rr8u45Zp/ZES96KoUQ8xhWTAmCKKlsI0
iJfj0LhS7NKxOw4RWRn9jKOjy65bczba3cnX0HvjB54D8f/NRAJ9FXJnqnQOPSzj
e6ypk1AmW+J6tBqFNBO4ACBAlGD+Nma/KjdMOXBliemR966sIvJlkrFiBR2pXWcI
jKVrv4GbdvD350rO0BKfyz94XG1X8LrYWvsmQsE77dVCLNViwznxf6W54o1P5Zo3
So3xVcQOaN2f97tmlvYdMK0r8VWj8WR8GBN1Rb7AzRWYT7v4s43VoBCGqyf46Q6l
WT53geTmpsn+wCSnsk9C3tXjnSjWWxcKeJ5odDdcGntqdU1JNZSO7CoSecUBN+6I
ARfvNB3F/mqo6XdZfY0aHMT2OQ2WLIi2kRVmCueDE62YIzy85TCWWyG6R/5J8UIT
RYYpFGxeMBUR8ylt/NhTXnKvF52ilh+r1Ov13AuNdO8uWz6fgOUG8bfzI4nMibKL
tLiNb+2qJsiwgjlI9DpZ/ljFmRDNfoqTP3/4cIv5kdMwRqgTon9PXmUzDAIzHT4L
f9ZPKk/t2UVcg1jSgsmiOMFejcG4yA2lCpb9rccF3oKq4L8Ss8YOdogUdGC1yz7Y
a17d9aJ3Cupt7naflOCVSgLZEc9gSE/04SLd7c3vS9XEOju/p7XKSKrILp4QAkLW
HWLjbG7f8Soz8hyAr4lYi6bjG+W4rcDcViQOe04eEKZI/C1T++e1swDjE5WKWu+2
tP533X5e4bgsNPQfBH7OQrtRcq7h4svCVHI9ymyxIeuhjcgOd31+jOm8FfnEB3Zz
rObhzQaWGJFJ3HILwHIP+Lv7T/JVXUAY5Ih3dYOkBo2zP4eEzO/I7Uvz3ODVuhaa
irCR+fwM6Ch/ckBl+1sB0m5kIYlMuxZHMi4b5T0/IW54bjNBZ8YOUcSkwmnFeu4E
f9XXfwz4DuRFr4Kvtys2VvGG77Q8HG8tivlw4ZcgZDrAp3gFVuaWzqfE3Reco496

`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
CN1numPCCGjFBlyIbgqT82aN5o0GVc+BbaSFRUjsEew897yXd4gTfPGZq9od4YnE
ghWZWk3UR/+q/89IO2V3oge1cI3W5RwVdLZqWnYXkoio46VtWfyThvLkC72H2lzF
TfuoeL2vGFGYhkPdy9U/HsltlM6c532QsOYPqqeJUb0wXMKraNYK2ZiN9pS2RRzO
kyriVTKLuiN3x8NFtZiIYv9CFAOTVnPdLsQIo398ngJ6gcVLamP7T9Veod4lHUfY
NiJ3KrKpEMoptbS0siAN/DndwN3HKvbMulO8YXg8njeci7ryGdsiUHBwCTccPTOq
ZpgdX4UuR9Ny0IKkSiMDPg==
//pragma protect end_key_block
//pragma protect digest_block
E0/7CHoTttqCGSz2v0jQciGoRAs=
//pragma protect end_digest_block
//pragma protect data_block
u7d2pVRu31Ga4MXvMs4BoflBBpg7gdyN95hla+6vMMqkc68eaQO8P4bKi/a9FUm1
hytPX73go6ZNclduLss3HdtgA7Ee7WAiWxh/aaXtXD80m1nrYtYIdHOeQNbG/kDt
1O3WLGW740PYv/r9+k2u3gfGUwttR5KU48WB80HUrbKv9HRGLbwlE8r9cqeyQ7K7
xYn0N4n1nLjx2IoeBjJmueqIXnprODJsHZRUM5Uj5IyxGOaxEbSh3h9wRfyuwosk
5DGxL7eIipJkg9i3scLxsCvKnhk08+j3lDykrxfD0K+HDkjSOtk1VihQHu3QyAdV
/73N6ZEgpVneNO0k2RdZ+weadLKP2w+fpdHvhE++zdBjQAqXmnmwfS223yUvzLah
aeypHWXIJLqAsmR8SgCt4bRiRF5DN65oz7F5rPIP/IiFSLW5A+EFTdxYIwjgHefB
z1Aus3Iw0N6vRqSwiW4D8OpomqLr4mz0aY3q7COjuna8/Sg7e0HaTNq3eoC4MXM0
Y6kL8ifUsaeTxh+aoxleDrxZKznNqbkXl78+ypM5nNOdp087y/h0hFrzqrPoBXc+
MXi/Fj8MMb1tKCrswkknJNkTqQZ1OtHtPUNyLdOlCbhhKVQR01RNk/p049Z3OYXZ
Y75/Q3u9q9Pnh9SVRQdYV+crITXMgp+JkggDdK62NKFoXXQG8vBQLQ0FuwO6njEA
zWJ12eMtSzGplqs91XhHSkp15nitzBojQKu3oQZlUhxnU21IhlfJn7ZuWbcjJkHW
Rc4KfbX95TyzwalIhigntB+S3AeOxX/p0ic/NYnJNrY70dEd5TqtXaLsFt4fmFQZ
1X/55E2u+2kldp2zSgun8sRU0sxC3qZYsxHdVIgFqg3wVkLres7CyMMc3tkDoR1M
L1DTGdf3SEY8BuBON0sQXfQfReEVsJwdl5Zm/t2GAGxHl+jdcwI0kUJNogAINNxz
V0CqijMv7+ZGOKW/lHhTM2smwWNVbJxFdiRyz3o+IPg5ks7xG4IZIhvmcXX236WB
F84Om6yBXvWod6PkPQ2XzespW776h7uWTXYnRw8WU3WbSAGgfKF2GPgn5NuqWfjY
9vkYKQkjXFDA20WQ0nq9O++unqFeAtNQdvxbWGXZKnSFv27RrjhIoJZ3D+D1ktlC
dttguRbfqIiJm6EnfNNaOaGUKfDcvfQs2vn84wy1seXUCYUdUW1r25tJTlVbdkxs
34U00BMMz8/VnmqxRx19qIYwFHGIFb8wYetXUGxEIG8fEYlxGaKR0HfGLVk3nFzz
LT8pHTsZ2rLB5T9hfW5958p+DJ6M5lq75W8xpBQqG7S5ftuRjAHZkniPQvVGVvc+
pxs4GQyYU3gPzjlalI9FYTUdlt3h7sLRBeSC/xBeEBK9ru3+yB57ljZRDPl8rn3X
NXg4mzD61HuTQToD4tx+yKVIRxHEGtld7l7kRvNeq20USwVxva/VG5PxOLIkYskf
ud8DHJUTIIRnlbCU0NFVPdb989zIYx6WTndxGFi/g8FXFD1VtKRdv4VpnFK8GPtS
O7iiRYa2/0g79IZrM01sG1gZOJzYESOnUSMY8Wxl4UrD/1+Z/GkJg6TOa7VHKmUy
Yq5Nxm9OhUpbyaaHWGGUauhQSAuc2dfDM/pwf60VF0I75qbEaXC8dPPTY75mZ/V1
F5IoRqxcM5INryPcgWFyn49Z8qY35D9PzZ0vqRKfZISfI72GcljFMUbbVMzVQXlG
H798EhLzsIdTZFS0vU4bPj2EAfbTgFP1++zIMTY4UiUBmx/voVqmjNhFkd1OtYIh
PJdZHKR/QtlWx00whm9g+NO4J8z0jjXthDxZWhSxnVypLxOY6AVvymN3z3NcZLHS
qGK9eeDgC9f+v4mABmGHF50jOkvDG6I7/Mnk49DHc4k9OxHVgID1qNdvsXI7IO2x
ogzyD94mD28UFX9R4xjxkBtMPKxduEgnZ2OrVsk9dJvHQSwi+CIIVG97PHy36yo9
PW2hr2dPgnRVW2vZgGlk7aJ575bPiGSSYcLL6L6cnXvOOcVUgC8uK2iSydt5Oa2b
OcqHMX+WfR0MMUJWghvpiy5VTnmiVT6hdhUYfOh6o3tLethQMi/0eZ20ssFg60kg
goAn4/hXksPV46NkVy+uXtG1CapJ1xreKWMy/kQ8gW5cQudLDGvFH21T72krXa8P
VKu5MZFc6sZ1qfUwZgiUVadCo6yT/c5VVZOto4Vgkg2mdclFL7pV0HOyEsqlBqnV
4qTQ64lWgikiC15v1Mi8Z8MBQDV72jKsCT0lBWj1ySce+mgKpN4Vt64gTgoK4FHV
1RTzeipeZchgat06tF70Mu5Nsl6dkprwTVLXQCZ++iklD2p7RTCAua2DuO4BGl0N
sSMN5Sr5l/1v0tztOPqqrCqlBLf/F1cZvXwLXUXs0Z7QbLqZGtC7NcjlSHp1aLZT
t12zXJ3UdZufwcWdDQvVHmhLXUTslLNNJa7WYEGT7arZe+i8LaP499m+htsBRbPW
b70qJKjrGsq5jjkp2eu4fw8ChnEyU0yO5zToWwtMwF5OuxlrVdIOfgFpnxD1Wqb3
YEryg8bvMaS8Cf9TRHBrbdif/2LZC+iOwFycijBiihRcfDtK8+qf+T9F5ddZiFDB
+eieEEv+FdhgH1cVr8BVzVwI5GkyL0yDQe8CKHKKF0PiNsBia5Hfipj8etesP+ni
fSbEADilqNuFGrzhWN7OQZ6r+sOIGjZWG2j+JYFcib97pyoRlOfqMOoix+olDTX0
yDLeY2LVrbtt6Keecv6DhT7zjK09ELYn/gRij0OqSVWFW8JfArzUfLKqQd9RNQZu
59dHKe1LNpXoJmjNld6yAtc41iD5vpwkSky2niaqbAPFle2we+/2vn6wyTX9Ldp4
MZ2Bw/muCKxRsxOKv+S2BytfSzm6qeXrcLi6JajW2FNtVVilsZ1wCQurD4WUvS/t
FMlpCTMXA1CJ0xZzm8qr6B0Fzpv2CVfyv8MpIXUDxbAF02zzp4r12m3Vy1eXPZmW
5IRnpfznOwxWCVFsf+fKCzCush72v1v6VCXGRiVLEBLM+cdnpow+IWXBMlc/akhC
a1T54PFVgrwSCEYm1LuNcU2K/CspUoq0LTixeWY6YtW5yXslEQFeD5IU5KOylzll
RHBg+yqaIPfhkkyb7heAplcTSZ5yt9wXqQuF8AJmajBiytmzffGkVo70eQotHMuL
Bo1RWB0d8xew1CqQ4GnTwQ1H4UhRsQqel7vqiZPk01rK3w8B0I+5QmAfa/kKQwdK
AAhsO4E4mGnh8qr0rgVzDkrEWUbrMvbMnj/cW3vdamroRGmRMVNopMe16EjbNtvX
hBha1YjYlMlz6yCkUkbVc4OS/Bo+K3My1L6wTiK0ZAFuTmIdsYH0uYDW0uSZcYn/
GgZRsQg/wkY2B66S7HdHry/N81Ltpn7z4f6p+0P3ZkdsqcXRkH2KRxTphubYQeXy
iCUkKf5B1xb0Fy01uEKsXXGIVkkCMRAkptrtF7tKl74I8dtawC/y5e/bIh2Wbh7F
fs/mkX8y1Tg6wRLT+5UQzyfjSIq1UBO/JhlQBIoz9D5Vy2joGniev8X1xS3HdhXj
Lto8GIa2/Lu1ghFKZ4zVYe+eCLL5aHN4o1k29GoduI/jucCvwrD1M8Yk+BNlLqLy
zq9+BqIQds1b5SHj3FJlhfw6curj/v0tqEaGmAi7ULHeP1tuu0aaTdCrlU6//0kQ
hGNz09NPp9z985iNWndWByG+qoV3av/UhGyY6K4ORyQ01mndMSZZLJYMEXqwmrQn
ijQxbnkwGJ7bTtbyh0oOeFgsTqbbLrYVg54nmcHDjqads+t4hNk40gXIxexltLEX
V0DIAKCb2NwvkQmLH3UDds8s12Nh1v0trGa4EdKzchsvtSNcjpOATOS6rNhDbTqC
4PZ4oMQaPecLPxTV/FYlnRx2rfl9RxMUEvRB4cHMRGStD35uIDzQatQweeC/xsli
KMqiBz65SfAgEEErZ3gpPFpZVd3Sp6mNOP+T7VqdfUN8RK9f5T5B2tYFC8N8D+w/
7zml8BPRNz82GU1LdbJ17akrh0yGKn69gNmCjAFHTHs9n/IzE9QORCr8CSmMBBYt
vrJGuDu8qohsPWHKbdxkrvq9vqNqLjfkgwhueQJQEYih7njdAxNHLOVnyxZm55ny
nHuYqQiIiHE0LHZWGPxyCkkDjzNu9d3PW+FiQpEwYKrtZ3ps6AAKR8MkYK3VpuHR
mInX+nb3wKBtUIg1e26Srt8pdYKJszNpA22JXvamJ0EidbWBvhvM0hzkq/7HJVDh
BQe0tROC5SDshIiOzr6J9rM4DKbHP5Q1Nyz0WhpIWso8LNyHRb+8nXyW7sLE7VHK
ItHN2A51dfc+5bAU1vL9jiQwm/LcYJcL3emX0sbPZTW2bDTioNFsEfPyVIu1iSUH
RyKB4QcYCPJbyhQwxm7aNeGaHu+66ftzA6F/efocAbc6luHY1onyD0uLEFba0CEg
SCoKZdTNVWAV8J2b+lUPALy/vKa82JdALtQK4E+IspPfaF9vqwVhGtR7l32D8EkV
uMm2TFEt9IcZ9fNfpf1icomZNVk1j9WuimE/waon1HL2Cy4bwVaAOv035yOyF8JB
jwRikBFjDSURQsrMETZa+NBdD89crIaVVSCpivsOA8NILdz2seBqBZqCPndDMsNM
UPC260vs8qHnETJt71aTw7PayonSeB4xpr6bTsYFC5FV3rQ5bd6gIoplWTUbT+yz
TBJDm802/lID2txr1a2LQ800sDHUHINcFtSgR86qnzmfxunyqiWxaUJ+v+UakdgU
B63p0wlqDoNIzXKX8rf0fC87Qekt10WvMTkjrb7i/Rtbp7747QiSCmaOTjAgCkZU
8FgeIb6F6bGPtn5RZvim59ZycDM64nnNPadkRCsBPyXW4Ghn5qvoY/0cA9EmuzhD
rQlEuS/S4qNz+h/ONnWgUeK5CMRngzJNDR/nccHvkUoEX6/qTck9kvSvBRr7Jqyg
sWnbOH0lB4vbbvvjrJqC0Pqwe7FCDO5pz47NlgufaG7tr2Xj8rkYixBOURwmBS31
MRBWjxdnLBbBK00BZ0Kv1Vbp4dkG3bwUIhj/6gsln+tXSdpIjnaBZUUyQSK9eJ/J
arJuDB7pbxjWYL3c8Gmx1FigVdhkcy6KqAY66HTAwjQbgzMcsvwKoDB9SqCDVTWc
mJnNrq9vobjhhNDJZQTTOelMS7laEuUyN31Bj+VOGndjucV2Xu5EzTyl4dO0MB7f
Azpk7rowXGzfThYv6tDTdchrP2qlzOmj4RKsXWwjel1AmdIRvPBHg1ytGmAlcTSJ
jovjbzyjsPwN6N2+9uYCwqRhMSZDJ+2LRCRg8TtaQx+Z65HvSoZtNlf/mQ36QGiW
9GH4fUhjFyGMlqzeZbY8n+u0dqRfWbpcJX/UszvLz5Mux6DoUCbZNk+nUZBAOMTe
3KBp2jPhGJZsbndzANWRGgGGbrYOZZyXgb5t6ROJufoij66VTiziZ+sckAicSBK1
lPcnA1xxSZ2+GtbI5HOou6voTSNkiCB9x/37G9fXDBkug7UobxfdRum+gR4YYHJm
7amDeDAqwJi/981UYItni1Xue7VHAuCcLs64/AcGWZcrYfCQQrSeGICc3BprBra5
YphzpVwJlWUw7bdSkhUnaV3Bsl6q0RucIJJdM9mIjfDarSPo4ESNjqBhYHweNh0G
Gvf6pRPngdmpqBcPCKCFFsebTyQ15z2AzYL5+DGUXOTypjTxFrEcs/0G8HSKO/jo
WIUiKCqwEpNsmEhRpO153sI4LGFdme+zpgrq1a9jpYJPCUp2Bm9vFPd5q1wjEfX4
5N2qjVkih2r0HqTUn+8Sx94zGOZASCiOpCMq193Hm29i25KAuyg7jfRnTn67cS91
nBuBrsg5OK+bhQ+4M1leLSS+TS9QiC+ySw024JT+xOyHPdoXRK6d2ZWEWaGOLUD/
204QGl3P6pdNtsb1OVfijoiGrZj5ZKyUBI/ePaQ31d/mnqzYZHqQj5aLHFBfhXur
LVqQSQRk6PYQMVoXAkfi42BhNIk2WDPdVzafXrm+P4hzOmcJsptTM6nnPfNxns2+
a/qfzfpyVHDUgJlyJhJN7QwFqG5dt6X9j3ZzHwuwlqYvx99h+Out0yQFyRV+om9l
0zMUhlE+zk2ueF1+6dnUm71qb8cOQWWhj87l36WQ3uu+mcJ7BR9vfHhTxVwik2u2
Asi5qG/mAu+Dll5/suf33FmDCgX+fM/9o7XHG84NijAKojAKL3z65h2zG/J2/x7T
S/r9gOhLBQYqcF3B5LWU6J+GAgJiOoSiOjAur+SRIGdpImdKRfT+vPE6lbsN3G3R
aGMoPHCEDG9ae5OyvnmItRwDRslRrNdxr8Ls87q+HpEKE8Iq6YzxppqrGIBLFkq4
IKGGbS84erkG5ijoniYQR2W3eNnEpVgYLhSvcL5RcolVGoiSJidNq3gW3b7V2IOb
IZExmGP31hz9hcGNNhcLDz7eIud1zJNyfjVG9CVlIbvXe8L51+azvLuKf4WFW5mF
JJ6FE6LwOgll/ByEIvZEFB3Lk5548WH5WYTULPF64k2ctUUt0wZhBNbYPVao3PdG
6j6oz1DS/l3gTCzoEkB8DZXWkytYTwUgXqCZ9O91jB0Kx+8LZI/b8M7xXLyCFk61
iX/ASN+uvyP3lU+9CXrY626+M3nEJk/ZK8VkgSB5CqCT0iplwXNauumHhZlMT1NL
awXEMd1X2P1P5hILID12znl/cDJZX8OgFljuTVhkgT/tP/qjPXcqLrmcdcPh5InX
wxkjDSZ6NpxWrf6OzOhz8YJ/CdjOuepUAo7hglZwFATJ9lcH7fHoOLgxvnfxV+HL
D4c4xYPt3IsX0OEO74Myb8PvbgH+AVhMUwC6s9duWfZdiMPKr6ft03USmerPkOsH
vch9+VUliRUmQnr1pOds3wMNRMxkIFwpDkf7jyBS1/zwzIYBhgW4k1q5bmZ2znyg
YCkjNSRozuqDYBmJ2RltNKjIW35Hm4c7lw+Mx0JyCcf4itsuooVIg3NFsEZdVrV4
TfHS8C8dxy5ZjAbnCgHknKXWclyRQ8TyyoIEe+yn3RhLQoUPMyCwiIoQm5t3IfsO
07gavdimHfVxm3Pjq51OCYuGpd8MPgWa7QLgh463rv/zadebhJd17zDRHNyPrLMq
f+B8bt51a5TZ7vEfBuK6eb35a8dN23HakSjMMZ2h5+qRY0R0zJBBVhXebN3Y1/nw
2lZmUn2WdNkkFFV+krTg88wAP1z7kQ4Ohl+sBE6lW+VA2KkkPBTbylQeEY7TWwZS
8wdQEy3LwezOR2YGNndEVky39mMf8U/iP6iFzeJMh5D6SYd7OeAFw0mYC75L3wmq
ILXd7kTwv+CA/HO1y39oD/vqG6qEkqvYt67kw6TFqJ3BVa6sf6u8r/EtCvWQhfdV
dUQv9SvRLAzskp1JEHT3uAQLw7sEG1ESGkD2Gwvz+AddBz4H3HVib1JKJUTU+Hsz
mjy6uG7zGn1h7gJALVW6ThHhxL5RpnSpg6bVTFRCkHlmbXnZ9cmNX2RtrWgDxUpu
5c0pGKUlvtPWFUhj02v1UkJtpduatZqQrKIEa/u97C64wh0Nkwt04E2vMITQuSpn
OMGR6CnCcMyY/QJH49LQb92iOzDNWaV8XepijLEci1d7QoXXWp6oasTpnf2qCBl/
kTGVabk+9/TvlzfCVh+HsdSbcTCTTeU0IW8kcK/9HAEuobH8bEjmKhwekivBitU0
IoMEaMinusgxIdS1HL5ZN/Z8AS/1Ocs7AG9ecpqECf44KRXVlCl6CxJQOPbL1y8+
/Jb7yO7Oohvn3Ucd5q4gCasrU7UzqZ/8d/M+ANQJ4lLBYntnaaMXOAAfg3KrX5LW
4eIkfMvL9UUX0ak3E/gWJYNvYErgkhf7TtssmSZ3GKnCSl6Gbbtw+I30kJZOE4yD
ZrW05Yja/To/BH4xA2oyIEvkvlgzv4A0SESrdVF0VkEb/trj1KCtgO+OO2HdFAon
NUGuf7KyIRA72254mc1fGzjJNlCI2FTlh3AE1MabSrTAwV6o2UgB5DWDyp/Zfg3x
Q55hsRxcYB3R3Tg5UyVLsEihf8KtRuseW2QCRuiYza1KVKuhk4pmEwkupEXmr6Uk
+OIw54NvgSnlBV/ftDfR4NdA/asCB7IKRZV6lcRGNES9qZLmxDzpsA8960/cpsR2
q2ue+1R61FOGwPHzlC93KF81ubmdZ2+/Pbjbk4sEGtQQYMP/bqIUDUyjzOIj0wYD
Pk/7gn/EftfIb48CjEp4WoJgyCss4/ZAEnSB8ze0liZV6Z1FqUK3Ma/BDTLfIO88
qGXUUqu90KrYY6X4yr9YFT2hWDQtYcZ55QH4ctf/6yj07nhTMCYSgFovANyBeRNQ
scxhTCrTOuPp5SLnD0wEfEGTaD4dKeNinV43mOFyGrqpDeH28rFc29eaeDg965s/
BOUYUZNz0euP3kqAKxV9FZjlmZ3316eN7JiHlwXdng3tXSFOEnyHZLSM0b4OVD57
yUL2XRI3hPMgph7PsfkKRN5PPnC9Ujxk/hxk0WYUcgiTglWzsdDIaqhFVsDIhUvR
9vcH7sSpFgj3KWE66K35+0MJnCAsXr+IuX0Cl06104xiMBbCcrGPKTthglssJPni
dYvAagGsfGU9nLewTIJ4Od/bYer0469v1hl3Fu+lVfXg2hMEZvZEBU4r3G4O3Xy7
RryLUjLa8aUr/6LKXsZcksvh/Gp5TFCe00exZEmlcEsv2s0+TehoIlADYNLg+dV6
/Aa9VzM0nNvOKOkYIUtuvRN1CYLifCtnYNP05mfvfO4LGFBJ599xQGuhzwKUd8mo
0RyVBJf/K2pLDLpPHEQiHysKokMSfFxSetPiPJMWoWlD5MKjuvO48tJ4+HwfOLPs
13g+jJItwMQWgGZITOCvxVMHO2mH5I5mkY1ClEtnoKNpYehg1VjCR6QBmIhwvi1x
oWt2c+T/NR1cerLs4y20seVeMOAj3+lgOuWXh8IxH24Y/o3toWgbO+3E1XNmu1ZB
caUkHwc61ZJ6mAp5SuLLv1UDYJSgx0jzK/3QxwZOQw7DFJPBNZZ2UKl35dLsXiHD
qvL+22xUbgkGnG1YZhrJdNUFg6It7Jvnm5QGr63MuDndvmobOulXZdpaoGZcUEEO
QOf0hQRieIHLsNIbFaQnf/Ev+1wid9NLTa2t2gq6DYk7Itodd9epUxzgnoICwmSo
dC3uWmdGC0zHaBDCU4SrUkVyMZHZr/fIQEZDKnzOkrEh5RDhBasypnVdwmB1sfki
n9NEzyneOIfkNgttXK5c4C7kYds8V3xeB9TULM9maRRTjHRdCiZFCQjVXGiSjD2U
SD0AfNMfIxALJGYM6a0URwCSCdF3H3Vb3J/GxpN6WGcTFkSncs2QiZTxQ/k2KX9h
CV5H1ZImxHYsbr4pz5AfFLnP6jbKQypz2q+DOGT8/JbywQ76XxH4xuiUqWo0Iho+
hBbKe1npAKMfKerM+NrRML1pyEFQfZVT4pqSTrA7AR+YUN5S4S+qmuyof8RmvQp+
FPYVbmLgrjFSkhcLwI6Idhsqv7yOIAaUs5gJcJFnTCLLk2U2RbZy03mz54TnaiC0
IwlGg5txBiR2zbeFQkd7GTsz+He5Zpurl594W/4GZSainoMElpSKYrdJWuNPI7iV
/P3X8IhECH2eUQZrIMANUzB90cs4KSmmUShEVww35iMsDF5GIATFOUfNyh21UAPt
eGbH/Bp3iU2tQ54TwifrPqQniYf+p99Fudw9XjoEBrH+hmwX5xMQ5Zm93rIu+16o
HhdnaWie5xh3bekYnpXGHbhGahyAKpDqqVBC4z5zBv04z/JtM8B0XeGpDeTENRfs
laqb0E3BBHdI9PpsCsYGYbtT/wsaCYWQlcU7+i27BRcPQHpgpwdkvctjsiOmxRst
RWk1UXXqsgg98KE0O9rVrWdLZ0Ctybzj12cNMIzNtjm6f30IhsYB/LOoAR4atTsi
yO95zU05S0X78a8hA5//RH4oSAoGreb1kMAvuxmgvPYd3lHXzi2S/eQaJ/lcdRX5
SFDFD0b/eA9tzXlI5Tqb7n/lrQwIXe5aQ2v+5nL02dKm/3jcgC72JLRXYwtsoUBE
ymbmOUzRFJcS1fbqx0YNyrvHcxsU9SZwFmv49xFHX9qj52qlJXDjs4wGqZYc3Q3k
UdyYVo0Pb3TdRB7BSi749TbzBlCxGaKZVYpjS1eDkK2f+4mJc3y1dmVzFgaX8zBS
6mDBfmZtkUkkuEaDiGyUvMmcWyDzO5HZ8rwhd2KmdDLhXfSGQQuK9OYvespdmHl7
93WUOHGi+JGOtoadYEiy6Mu0bAOROKW451oeDFmhXOdcsRKbCDdOujPe+dXBZEdh
bhqSxnRgVzO93fDqz8pbcbyk/9TEHmRTceqf5UhoXDuvFc9lWpHMoYcuIc04INkI
aG4GTccNMHmNc3XDUW8nq1zMFexcpkurbzAYh7xmLKqDUGgh+levLZDUGppq7ify
Qvh8P6uvMJ/Um4Pb5fiwOO/YPnLe4ycxrXR9F5edP4RuE9L5sPmzvQM0quQ8Z1em
hDRotXGwYD5WkixrXwunKSbvV27gBcdaYgJv9Mf+pzEJygAf5NxtNYSFAD/yCw9w
vJx9PjUsp3qavxJpyBDJ+UGtgsrlXyaV3cZk3y/El2nS/YZ6a4Nw1qJ3UNzcp3Cs
JsP4zPujY1c9+vANUC6hLLRermolcuKNxmZoc8vqOlB+YBwy+lUFCbvJpfEruv1r
ReV5NrKPpg1ORufOr49ERIUNcB1lq5QjMIDz1izYLUopcO9PXVpvulFzna/AT47L
zftUT/Crd6xBO47lAjLujTmb5V9i0cTRAPDAnGHVgZDP8ImZ+Uu80cDLh0E4EbXg
qWOtDa21z9TvNgFM5umgYs3QxOooL310cUZWWH4YXWq6CjnqDIGaJUuhmVFLTVjA
2M71AuCQj6vzvfSxqktOi3WGx1T0TqjKiByVSywMFAzFaACCXnKf2JzHRQdHo5fM
tba6Yx4p9TGGTq0XGPSn6lxm2zpSlSj7h6NRs2j/2AEZLsl+6xhnmf8/2n3F0Nvz
aAsx3F0lZFv7PfJllc5lufKsCY+NlX2I6lMZuOlm5L/zkd/D1B7iGdHBeXpJrGmF
mKltNfIJlmh1JBYYCSsCjWhoWcDggZKwzZ4EoKDR7iEjcUvvWpYhH+gBNIdq9eBl
U8YFhY8qGElRyoIqtsyCGTqMJhFiNZeX8/5MFlXdi3v1TVcx4iR6ICfUeCsijIRh
YwWbzn2vSP1r+lQ0PofWla2QeJ/RPLGw6VK95OZY5bDjpkDDFt9zBkctZNXhArZb
K9wdqV0Lz3xw0TmogF29Qm1K7FoKcJKcHMfMBX7on0CnyFQEpEnEZWXjtA/QlQD/
XDa5E+2mYX7OCrh9Yrk0R4kC8cJzQsf8SQ64fOy9oBgamGIcozvkFmKo39YFIwQz
V8S5Joe8SSdD/LAs1e11uiiuo7UhXElRwvkQDb4Cru+PApLbdIzuE1wzMkv6U/8K
BSjTYWd0OC6siMFyB9r8F8bjVyQKMiOktjAFOE0tAi49/SseFS6J8/qYSjwAtkKz
2gAQ0Zmg8ZqeAx+n8uDPgH00OwD9QgdHpuLTRqtIS0VwAorydWfvQ/n1zaTuQ0PC
ZBzZSFGfrBL8ylz8dwA6KksxH9fBFGm7e9aCjNzGI6yHiSfKp/PTzTYlsUqPjiK2
sNjCO+NsRQ3qPE1GJPi4j7pzso0lo2bnN1QF8xl0AvjMkdJeT9mBTvBPHnN3+BAA
0AR5lP+v9IqFfSnezWt1UT+RJOPz+iKCAM0pjpt+azvdre92iOuyPVYiurXy87wl
k+45RNeK/UqcYlWLLIvCeqQMFmMky49MPj/YcVKfFEVaLLodb1BjS6noMGZUYsxV
uwPU49GV3DGk9ACDPpehmm/nXLYIwztutKLKkUb7vimY1clEjrPsRPnF/FUsBBSg
Um0eM+5+V+LwjRR+tEDxGRPtxx1kh1LhY6n21KZz11uUpfPq6EIfTamfLlOTMhvy
QUhr/6UTwgiuTEEzZiKAsq4Mb3iyVecWTJ5Bq+0evB/ecZ+1A7nr/S2zUlV9fJ6r
pFaFMxJQNXdLdd9TO3xoGzJqur8ViT+PIHTSAGoBGrZ2SrkqDSbD9j1Kbej1q6zn
E8Z/qng3N1ZwMUleGa+WFOcPJQBQE03uxUQJwmLmG90tw9XHQKMJlbaEKTnhfw/L
FPH3KEcB4MdWQcC9xmz6Hg4mX941pOvplZ6desmpAHzX8ig1W7z0IUdkUtAqWOqp
4/PyTYLea9fn4eeVm8+zNBWthVps4pKY8cbTDrHXrM8O3FlcTXUOo/UjcSPxhCRU
Q2qhukWNl8Znp2vAUVwj3rkHcZ/T2M8HexrwDhTowEompxqfQwphrw3h1A69eQko
7TcLkTqqINnCxpX6XI2Fuy5WxJO++aRwTNhljaydDFXoz9NJi3DlWUgTxkT1IGUl
N2aAOAMGmAqjuscjWP8bPX7+gqekR1J+6txjNHQ9r+BMDIRDysyyTGpmY+1D3pMN
5g/NB7jvMusxegmtT8uf8Dv8SianEBefBVuureyhfQnAuactxDn/wTajxQmUojfl
c+43wjo7VeIhZw/9ZRzcSDWzN7NPDg2G2786c1ZtOh5CsaCBMigsugGlneXbV0cH
RxqFeP6ueUOLft1WQi/x+Ql/nCXlf2xcqMVDTqjMxCD3u/1wbhlEioOrOJVdEgYY
jQXa7qXUkTutBAkXnZxGEwXBpRE621y3VQ6ePdwd55PPOTsTfzb7x7gKO8rudhTX
6NhBhBUe3O/qIrRXIFvOUoSiaeUalgyCuYQZTyEEtomyb6EMJWPf23z3wuJZWsWV
BynZQv3C+V3jcff5GMQzy2bRBF2uF3lw7BrHC4YHKUdGNFUZUmaAhxsg2OqcHRdT
1vcAhAQtn/5KwQF4XBv3cwpDb0yepPmlC7NwzARwjglzi7ifBq/bH0eycJiFTvi8
p0xxkODq7ju9v28OChm7pBSjEi0fOt6zIITKYdb2rMRDhOf46tZHwGDTJ2xeuaDA
4DTpe00j/TeTJJ71JHYsPvmLICiuJUZsFPfnqxABbZvVtbYV4QnUsshQd18B5bWL
XsSSfd1y+y5J4pKmZirk47JZj2XTtnZjP7KkH93wU69eszb4yBmFBETYMQnUsQEP
Y5KW6XhEQrC71V8kbbiAj9Yjo8GWR23cmmsCaGJEBC69iN/rv1aR/041CrVULqLP
0FGdZSh5/hl37lvXmZQcno3bpA3zjmJAo/i1Wd8zSmLanv6VaeoxszVcFgbyb9tB
9CzCSJkUpra/P8557QAHEjCpypK7CVqIHgS/BvgRqn5/AMSVQKqBp4bfHvPNlE53
kaYJmqu6ZvwgN9NnMu3rXQxNpJt8SlbTZ+pUgWHSxC3+w9XloLXroCeWZzmgWjTR
eh5Y/3Q54AccfUXAma5Ks25JbLxwCR/4f3TMrsJH0UJT6B3vvK6IIvxyk8relDFh
zK8MFwRRVwv9SGUPGoArGQOHqI7mwFriKy6+QBi8Xc779ej5OUMHU1bEbpDgh6gb
X/o5PvOQSvJR44X00fKNTUJGnEOWz49vf7LTqHAhYi/1d841Kt/9YfxRI5Evt5rJ
97OWdgs4cadkMlbfEcPdneF4lUlkrFZzbvvLsZHEwB7hXzoHmFDmGKx+Sv3hgo3P
8rMCOW5pVS727Ut4q/rBLZA95+ErvBuGGY0FjW7rcHUOklDSMtTYFP3PjeH4TogB
mxZk0U2aQA57ctZ3s21wwUvoNqIth0ev+XF0n3V6lA0gQjobIf2g2ifrMzJfYptA
swzqTZZfCxu9lAB+g6xcoqT/iq9fVrvB/3tkXrz8XHHNwBoTlXJHnXSvRt5ghXEE
J0zVwFBJiKFjivYJxtR7jXyWKKhcCJ9pQuGILSGQ3sf3lhJT1V9Lli9NpRx27faz
vsHMayEjc4dk8ircxLF9gG6fZ6B0fbjqYCKp/XCexSAQMy6g30p2zCRjaIZiOLa6
oWdyUKesnuHdGEY2+Ks5MB90tIQCt6Eu4UZA4AEsmGrS/mOFamuovQFSMCcLIVDy
NYmr1cApVU/Ge5BGn6TtDaMXa7OsruTcrD+e6bLiTwJblv3gLqGPmQthQNklSOz9
QfgewyBjrO2VFXBKqH1k3je7ww29alhHfn4xF79p+ZR2TxYbMkUP9mLahHEMS9qD
+bz757guIpvLmES+rPFk5I03KDEzpshzbdkz5CRdRYv4vgZUC2m2ZjNOQFYpic9f
oD0MAhkSikJj+pds+G3nCcwicWghTxUFBvznxg+qbxAiiH7jNCm8wgy4/Doq0VXA
iFu17PQJ6xJhkE6ySOBxp9cYWK8qblN9JRwYKmSa0gX4iH4XxQdQOq0o/0vXvuaP
bP9Ei07n3xYce34FdXX7cMhfZvBLG0xTcr36JzoPpUMg+gUVaErrls8K9KYx2MZT
ZWFMRqnEZjnJW5sd+dqR6Vp7g3tNB3PwIPV7U124Ya8QtLgDxMRTtxGw0BvSdeV3
LdjSusqlNistTdthQYpriovgQWILtLh9h0grRQPQ7cFIS/fYXLQ1fwdXiY/WAmuk
TyvBCSz83NoHidL5eDGzc/ZD45vUV3fXLi73h8c587aTQ63yrhaBeHePNvVyzR5j
km/07z2YmvxMvxXLMI7nlXw2Ylui8l1pzYtWx6j+10j2UyG8zh8TBk8sZxFXRXyZ
85hvdsTmvQfL5IUAudbc8gczSp58Gxvf0+tnBWeTaIADs/A4YdmCtSomnfvJIP8W
CEKkM0BtYZOfBKpybbKEOCqZVKyNBye2MVsnoxJGFPZb4MN1RogHuDqXEOFaFg/e
Ja045JJtiLxgAZeurbehI1YglGugIO4wlVs520SKFWsyRYW1uMFDcmr9hr1WCPP/
yWu1zgEYQBCbDn6tk0jURT6T53nnRRtxdSvhBzCugaKKkQhElv8ElzTyt+W/OFpF
vpR8VBxKYMzuRc3qTrTqEbMTuGJ3nBgPgl2DbGUNyFujNvzz8wevhQ24tps/6gEX
BiVYFpraxgbrAuCKPmAnIYxnv6kkFgDZ3RuSJqe/6GXKK3jxh2AxhSdMWBPmmSyA
An17SfWDhqbuTchLq+3ouGAQhVIjWaULTeCoNtYLobStbML7TzS27qFYwb/sfDMh
nO+VSsboGsncdRFzsXIB4C/0kUthRdNE1QdYoi50DFcEb3cBVVGE55g/w/smTu9G
aJCmuuW/Izh7TeCe7OSBcQiBq+2f8aWGA2Tb/TmzjKgh01ygCYn6/ofYq8Heh569
PFhg4vauetGMVRZBttALYcZIu/47dTmgC2lPYZuqIazhrJ5axrQdwAApAHMdV8Mc
7vtxJDe/DvchklVypyTZxI9ab4J6NLKtrk7qll1pvXzQs78eA/u5g4W+vpeQwdJI
22LNTmeYMIgVwntZX0A6Djx2rdrl4X/PVeqwo1sQ50LO0zlEOQ/KAzoJc5M69U7B
vbrQ7RiZUTDpTJ9hBuDpuvcLzpU+CzYZbV2zH4IWqIiHPD+ziMB/OEF3Vp2g1T/e
n5YLSv3vudHXw5DVL8XJIhmYFszLciQP8a9EGpUCQJtN/zZvz+GjMttvhO96no1q
Z9y2m2XvaZ9XRp4nCnjgOQXorWGPC+S0oUnuboV1XBMGgbEAnQYYhIOct+g4moBB
qF2bbdDVg+hVTibG/Tuj45YeRJ9Zf9eIxOn16R1mSRBieIaybEnpHce6/afg3hHl
Xkn6C7Tn1PuU0JauTFiKb7hpMtRrfQz7iFHdxr+4+iF9WZ6j+llqVPoy6qpFdOAO
2DYv6pVOBS1lEUGXPuMpzKrPkJigLGHI2WvFSlZmsstVQnbO16rySZcB+8JldM6i
Ba/oz5SuyaquCnva5NYbcyH2FdFs0v7KGMQ9S+5Qxbm0c+DTy20VhZtpj5B6vbVr
MBJ7NlgX50BcY49A+s23aY4IGw3O36Xz/O6qGS7zNPkQZyKVjb+MUM+3AshztppV
cEXkV2K51+tAE6y57qpwf9d4MhcPGi9JJ5Vpy6gchQj6nCPtt69VWWf5bJ408idH
JMwlL80Y3VpW8Zo1CFn8fFDmNdqPMMtnUte09R41q18WjU1xRponwtB6Nz5NAUQ2
jWWmXvRqBKtDnn4gVsJ5M54XGRtWLk1onRs28CdmiEcX8BZ3j6X2dqlAZ7AaJnCT
yzbFSumcsS15JmIzCdwE3cT31anCnRvbnws2kOK2ZPtmCH44p+QFqUsFPtUZWfdF
qItn7FFfp5PgUy3v7pbYWY3o9PK35sLxaAhTrzbd4+LjNGNsbIJr72gTjm9cz9eq
mHuMKUL6dEE6qDR9tIJGD/Glm0yx+9j34dd1G63WaOAZ549tZJtOLF89HEs5cdlS
4mxHkfZj4trIVuyBf9FAonjM8PgOM21oywq80xjWb/vtbOAHY8Dq1spN6lXGlRlK
aiHRcFA6NmCpup9T7BYlP9ru0/Q5BXfN82nhXIAnH2WnAhZQmld0d/NAOKtq57Da
Jgy60jTLsmJrp3nCjT5t80W8Ah7nH7tdCGSvUOwlCrUB+jNDmFOYqKKdSmiLuxnW
FWGYJr89fS1eNeHBC6E7DOvScBd9jVCgdY3dLBDexb80TBjRxdZV1HtdVIaszzaq
zfJ4oLumQiY6UHzglVKre5dWy1L+m/6uB+E/p4NuyCA/YemasxOyXrfhelAc6s42
JlEX+R+SF+SxnTHfLc7dpQgIl2HBv8CaSeof17A3JQntzg++EcobI7CgpRQQlrhW
nviw2BCJnVfXvuALmuMi2X+9ZAgKB+Bvr4VsKvH6ehvLgPzJzCd4nSZdw+610Pmu
VeU0Uo9LWpbCephJ3svMhXgm8LZEMEvX4lJccB8kLWYQoWYStpQjYcn06E9btXh6
2SExraP8iLbHUSiwpRAJLKCRJq6x627P007SrisfBZzGJ/wohHNqD+6bzVXRHwTr
f57+9dfa3imCjzb/upudtl3bl2Te0wCfeeVzYZUkQIbc+q16vkXyZ2P7h0yh14PA
GA2b/dKI5VKSQzMjmnF5+2rG6NuozsdUesGYg1OyeOpQ8HoYO/RR1W6o38/IH+kv
1Oql0wCh0TPB3N9jY9alB0sNySA3XnCHH2p3ywcZ7Wg7PjttziSHhZ1DLasMbSJR
Cqz0MBkbMKXvcs/mPiNgFTm7TqYmcGNKLmxBxrrViFeiUQ5ZC2IdPDrGVFgJWAr1
6s5iB/IcE7mkBSsZV6BHn5b4GGnH6dv4eshKYMxwJ3fEblKCIubEhn9Mz54GWmFt
j6HjXNDcYTHaG40pTtVKTro7Sm4TZ9D+bDps9DdpzuBJkK7btBn8ZuDBkUNnYxkU
eMZBUcEP4IdzGzfzQf2PrFn23GPTc/19THFLF/PKL2Qz++2Wbh81u3gbgW6lnuqj
0r0xrvr8cegeq8NyBSWUgOcfuDl9rn4vTBlAztQBz9g5VIX2lrTjSkyAF3hVKJhz
91zWZjO/TAjMVbIbI2P2OHx2HBva16D2DY8v21bPTUmx9iX3cA4+/Cs2o0lKGwJ6
fW1vJOWlHeCs7BAXoIWcLt6mgEz863KicUdFpEEFq4Vi89NLTMQhm6c/VgCD9T2B
DeqMPR6IXXUb5fA/AE2suiZVIzJOioChT+qnLg+6cP/aswTOYTSpqDKEtfCHmLx3
Y5C4UrpQPnXhsUe0Gu+lce5NNUVvwmeQOxk2rOGXfgm9C6Dm2i2ra5oSe2wkDemv
+dhxb6Nvpj1F41dDszdfmTcK6owtmF+9g0Lbu9Gcr74nTTgAm7w+IagOWZtrl06d
ZauhM0LWrfLBNQsZhPmujS9fmXf575iSIaWcT8BNaUQXTlCaYiAGp0EPWUP4fnpR
eSXi6bh2nRdLFrlJAimsKyIuXS9nsHxCypBp10D3LVghNEsMyd9x6lQ0xhKk4rSB
MO4xe988tMCB2zibxAtn3HtoNO+d7AD/feyOkVjsj14067dy1MAHEn/8/67KFRfB
HL9LYRJp3u/zo1bG/IoOF24FPFxfIiCmhFyeh3TZSw6Jqq327UG/w2XS4P3f6G3F
x5Tjc1J03aERLYwabnuk5w5cF+gjsEB2Lf8vOk4oJn+uFDltB51GVked2Xl65tRC
WiV6IeBTw5V9rYU365BOOUdegzvUW2HNe+pmbi5HprSRP28JUCThIaQPvJRbOYe8
SMi7vnR01kjkoux2PRTKmtRXveZINVqFZV4kBvB84JGTDveD1l/9/ZlnHhwEnGdW
9NM8LTir5BJz4cGUt3MDIFPZPWr63keR0CTzut8qEmxrBpzxlpYlWXUv9fdrHy69
DdhH2fAu7vRiFVpK01akzjJekeAmO7BQJS/qAWGk2FSroE0I0uW4eF5kpfjLUtYe
CDI1Xn2QeVAPnWwYWMoQkzy3A8q9kED1j3rgqgCKLB2qt/PEYnRjjs/HBLdRQfNo
pZTJXEy7QK5HFVQHTkdBDVVcxRuU1HK6D8bPuAozwgr8E9uIDOLiCvtzAxLHUpH1
u2fZDG09uvnnmd0kRGV9YoaskL1Xuu3Rr+UvJKsu7ltPhmzhqDQcfFCTFVc0r7wC
9f6VkrYbSYkmBi/uWxajWhEPIMRCXIitLRdcmjedqIPbuJGXQUja1MCXdzGfmGyT
1/Xr51/BVWj7EhG1TkqPF4P9XHwSW2dOljIdfNXYoX8tpVBHfC9QtyKdTqS8Ynf3
zOoJRl4HyvrmeepXXwH8Av4DUe9uWOA2j/DJ3zEigjXV/aoc7armRwfg6G7l/1MA
us6Nzz1PTqS/ntEFlSsODPtLZAHEi/1yc/FHJ/RVkq61hZEk2gH7WucHWDqEKmgV
qRqZIljVg2DgSu0EKakQNnQNj9LDreb9hunndMhKGE81BOSUAq5zQCSwLGTkhRJI
ZWhPaR3POfgVDs5dUp71ZSrUfJCoXF895vyo4atgle6zz3QjsJ5V//Rnqozblqx+
05cC27FtoySYb5WcVUV8nI6XoL8s5f0SJFfdC173wa4x8VHWolE5O237lgI3XZEU
j/AKQ4V7C7md2iwaXa5DRz42k0hP2J/F2IPT0ycE6aaAwLEyfynhklFyQvITUWi/
OcnDC35lThS/NJYtiZQxNQl5Ihryx6VM+P0FZmKAqQw2n4DfGzBkmslJM0uNaYCd
6w1VPJ9091BY0Pijvortc4ldQv8DV4OSS7T1D2r+lCwnGaFWe2YflxSUWSG62LwF
3R6hLUvodWuX0xcjIyaP6gE0ARg6n8nqzf263hcz/MGtWNIjq6XPY2YcGCBCnRlq
o+2L8huqVMLJi1gZttQ1SA3naq+jMjnhKJkGcpFOkehQCD9VvxDmvtCbQcVTs1J2
VNYFGsLPjg5CwjWZ/TPIHA1p1g6vqyCoMbJG8V4muEe/jDpIFdyCclHQyBke9WRo
8egjM8ruBeyM5mT8AkvVvHw03ygySn2P8Yej/dRW9IMxsVd+e2+RkbRslx6NN8Y7
IC7Vu2AyoNtQPNC6QADaIA==
//pragma protect end_data_block
//pragma protect digest_block
52CRxbWKQu1yXPwVBhjMmF7p1iQ=
//pragma protect end_digest_block
//pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
tea/bDFtP2dqPi1s0mkWqAxb4zLH1WA6u9fL+yl7XBsSU/Ot/u4c/e1VdKRIW4L4ZMpmZ37tOr6f
2dcq1P1YegokMLqJQyWacg1CKdCJsDrl38Q4VUSKxFwW1cqookXiOpDHP+SkVFj5wCASVIbv0tNx
kai9Gl5VffeRFKKrxaweZhBpxRMQS5DL4QWXWlzqtpdlV6LrSCtzzBivL4WjCpcl7FE8nap0ePOk
YNmg3DAUUBFHBTLK1NeGKWe0VcxwL+40Osy4R3slb9Jd63t8ggxvB0KO8vGwQ+V2WbVM0k5wnePi
ZWbmm335f7sO7ZKH40aV0U1drXd0WzFZcBJj0g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 7568)
xLqNMwnl4zBQZvKIVALRFb5kWkEABfN4OG8EO2W2kRmQpxkBI67Yla5rHzbQhZ9kkxo5GYYg/MZD
xWa4S4KbN5e0u/JaF0NjaDcTzHUesSO6yS53UsDW8MfI6iUd0xMi6IhYcMUCa2Kr34D+ftrw54NM
bX860T/ZzymCVAKtVC+qJBQBg6FZI87eYILEP4v++VF/uwvtLd+fBYTet6oYbt5mjIVUabcBF6S4
iwj2TFO+aGJWhHxCO9tJ/INqF9JWGPmkDQpupXJVqZ/JCRDoUQR+bJB09BzQPa70otgJLebUOwse
QZCEaxMW4GYh7Gsti1XgUCKcro3zV/CxGFyGO1lBN+PhF0fzSHxYyHjRlIv7lFixQL5j7qwAbAZq
wG4dYF6T0IPqMQ8dpt6VMF7NCB7Ce/fdJmvNqnhNekZtwWdOvQsogueCoJvAiov3mkoPjfxgdp0i
SNuf7GDA+gkU4Ztbe/4rB3NiiRaIZj7nNlMi2jZJITgYm0ArzOmw0S3+nqOPeGytiX6smymbhow2
kGh8VQswWmHi3Xc2Wor9wa6VtPehazzJTRJXAg4EBT69jQGA2iEuK5njE1KjqVw/nzF32nBk8KF/
2kf48XxRbNPKtY8vI/nLi65McErBKxfUcxClq62NcdOgXgJ4sc3cKJRJJtquSiASDHEqDuN2R/wl
C3w1saacqwHLLmDbKpfb6ZaTdvlvZpaHKQNCA7BWynt8sflqz0zUK+YGNMcqQ7rVG3Y7K7tQfsqB
CW5sW8RyMzeEgof8h9ArmJlRJ1JKp4/KL6fNl4NyHZMwc3++1tTYcpcrmM1zqpxgF9vZA8BMu9WX
rPpdb2YE0cUg7aoLtvucEAmut4pvsVRJzBHioy1lC0qCm0z914pF1wopb0x7f5zPUna9jcs42k7o
N+nk8zOI8eb2TvnteKV8OHddGWrDRNky7+d2D8bavGz9Sd0EbO5MVOf30nTDvE+vsiSnbCo/BeG/
711emzCuICK7QxWxVhPNZ89BDqe73Vk9BRaQ6mhfpgm5uRzq/BQTTpFNTysqION+SJOvz4Raxw9r
UZz7zj1nRajCNzG5TJ2OJTL14T/6EWR0bi4KHI1ORRCl04F8j06oJHMWUHfLcwAEWGJSdzuZt3tH
k/0drfafqDmJBgXSKMjmL7Y4iS/maTVYzuWwfSWMzNd+/eUBnWx5RwfuXOQSEsJFH22MS3weay2o
KaqPR1FDebvvRf1PjFfooY2YFJwWugn3uj2zZyjaUt/lq1+M95N9wCngcWErLS9XCFnelexVp9Ky
mx5kfSw8dA+er1tLSOvTNbYUNH6ncrUUxl1X+nOtkY9sXqLr/21KU+jpXYWQi2FZLuPz1rnJNxdu
ifBnF3KGDxWNbEN4ruRhr58dNX4Pd13oVAyAG8MCjOGqwmkcLZejRmZ4d1mOrlkGyjpTL9CiBUjF
RGVxPCiDfQAGidja+/BOZrJ31xs6sZiwNu7G/rd429tB7+nalaaRN5qbhVH2pJytCp+Dg8mZCxNd
uLDsQso4x0ZY7WnBbSBXSvT+Wpa/3yDYhZSiP7iNx/ielaSlMDoKBWVHn7UIxmve35W77yCQRrdF
3fKv63Ow+Ms9cguRYqpIgSs4SGe9Cgij3EkJkhDOshrBs1ScEyPeogvnB/iM6nkufkHVcgAKuFRm
jog5TYOMuQEpTIKncNVXRsNQaON899KvpojiMRp5oLmrF5qUKIQvDG7rGtk+Lwz71DTGILJPSk9k
XrSNtjg0r9S4Bg1P8rOf/e3bfK4ZeW2dDqjPy8orazGLDZx9uyGmsgDTrW+R2RfbszHh8P9AFXbo
Yl2x0/jZCwGUByQeJMDeWrmq/gE5aeEpxwNu4tt+gtTAr8rSA1O/skmVA9OcqMWy00GOX1G1yaDx
izAWn5sgs/tkwk+SaDPvgrRGVHUV+FF+yu9BzT6cXv7bYuhW/BaVtIvT/6QSKlJpGT8Vs1AFQpZe
D/FWANW5zY8MXKdLPjJPwUoA2E7lHMT2VxyFQs+zNC117KIGgeHq/bTOKP07KUv68L3vthMxJj5I
ob5MPLJEPWjz0MDNfxfWPQC7UJ6yC+Nyd3CLy88Wyp9Zle70iXDTkEp2Xa/Wf3fLwep2Y8XMv30i
8VpPG9amynGdR12aXhG2HVbmj2PwAIlgnZgnVwIf6tdyyjlvrx/Rk5xSxeo5He7ou5fuXYp8ePlk
QzjYrReTGNCI54LyRZydHLCFyrv1flJaKx2r6aV1LRUY8eYC92RS5icD3dXHJX6pduQyhm7hE/Xl
sWBbMHwjlnA1Jkfc9oU5n6LoogXq4xFT1xYjM4NCgnyXYEoFJs/Yyf9bSNPmy9vBEGZ3WK3UAKci
sf5EZs9wcYttsPwfUovOVqUzcO4px399blQb3HAnw9C2RNQsD6CtGNHICYcVWfQuIyKqHt6ku6B3
1lE8a9v3okY9iCCZj17gux+rvKmG6NtJNYf0u3op1VxR/FWyYLXHN/O218pjG+UGPF9TgJx9Wnbc
1k4dHMvXgRMnToYaO4KSIyHLMGI7zJgni/eM2BZ8Hfb1iBz/xv+XlElT9lFtXgV7/oBX+WJxpgSh
JyOD6ht6mX5/5myLe57ldt9iyyyI7RTMaQe1/ZvwF8G+a1xKqUZClfhDZALTItksdJviVLKFCWW1
LEl2wRHZwACg8jtREjgI1o9PIdUJJKzGTj/ogpnwGZOC+22n/yMSumFQaefkPxR55B/OD1LQFiRk
Aizy5NZpObUUEz+lTaQN0sQp1Adj87Fjcl2dow8tnkFUTqT1oT/WcLwVPZu0loe+TeNhknO7J6uc
N5XOzuDrdu6VxQH68yl4ooMTvR5+T+C0I23FoejRbVLomrEjDjhTWFQ4riI1+w4do6+MUQYJKIJ1
m7swVmFzc9cKjWpXDIkl/CShdW6p+vt+0iOojLjkRkAzGh/IGNj9gXbT4D4s+2rAm38foksAZy+H
of2HXvncw0zxg8ljsnN5RGUnkiP1hBDx6kw498a0sUDLtL3FuvKhNbOPZ/GTAq76hNXPgLPo5KdP
ExrJDxnFCTLbquMq9Gf2AIJVtLqHWfCNY2qYO6LpgdAN9vGHPP4FLaK0rCH8Kx90IrgwJ+swZCfA
oMsw3uLNenJb/G99iL8Ti2gpZZl5a1TxOzB/2GbAKV5FN9HIetQY2ydmuk/iOX9Vq5+cUtG6kzq9
fpGz68WMi7qbWz6laZNLbJ/KV0RbkKC4QhiTSnPljeLh7xVbb/BS8QiY/8x5YB4Qj4uwZHcMRSzS
Qwr0jgMvCFxw+p9uDgcvawuI8y3nX4Rc8T1/D8lChjf9PnrpIyhjuxNryeEEk2UX2crAn8KLUxng
SB+rw7SDbc0s2g2TTcU0vdM1Rnon83WeZHhMP5nF23xJLi4KePWNQ2tXtEBeU4OBSFrAfZwk7E+B
BVUXIpwtjjU2wdQ6bEaYXMm4bvur6u1QNwrVg3oryOJNa6aSC18kQiPtDcnkbxw/UJs19tA/gwVW
sf9bO28qK1EFIkv1Qlalw39jgxWDpjVPkfW+Ia/b/cWbnhR3kCe4Jop0JKmslboj6vwtFzzbhqVZ
ieKcDQQjp/q7puPCoAnk5S4PcA7l7Apg/sVM04FsVGtRaYw9p8vq49Z7wshqt/ZAxfQoBmpBM6Eg
G8lEPQDToXERQZZb49K2w+1Y4b7iEa+StKEWQQ0CFkMS+IJ77Sk54vtq4/4SzdESVMKzVnrAagzg
YuBhhEDkQ9wUWWA21YFebRCpah183X3KfsCqeleNwcCiBF5yuzexCpKl6BVrl0CpMaDGlWrHqWB1
R4xE+YyXkoJVpxWfssydPb3kzP8K4Y0lRioDXJhrf/dwuySGtSzvXycQ6zQ8qMXD7BW8bQNsACVY
zP3gMCLrgiH9Kbpi2Fy5SbWP3uCNKs1bilfi4gMcmZc0VCsGkalwqdQcqBJjeWtLAC+H3CV90h0r
87/h98UhSsBT7pcTApyHShqus0IbShraXhexD4Owk1Wh2ezLxGRuNUQjpDovreH2ZxelAHPwsR3Q
M2ILp8CoJ3vvqb19XMAAcIuRNiwkT0ahDoWvlf+LAMqMxxhlko4HokYwCctcPcQt1UkP0t+65lgX
GKIS4Geveq8aHjo8yRP1WmAhdULjsT7Xn/M+yTs58ACkvgsd0z5MSBZ/fYUjbyHw9M+XNmz0jjF0
Ky8gXfMz4KSR/Oce/AqqgzEhiE2TUUsmE+/LUwJHztB1CM8pFhvDscyA7QuxgsjtjddGnwKopYr7
4/lmQZU7/J/wBppqcoMGEm8WCsfXTIkAC6BU/9ZFKRJWNtwhG5G+BeaTp/Qq03n569k1rUx+aulZ
C7KFcacwPZiE4vALq6H9Za6U3Efp2TeneHTkpikkvacc8ePLp/Yjxqy4HsSkSB6tYmIp4aZuEc9K
n/+5eTgdNnpDZw07jpgAdVxxT/MmKFoaFVQoJ2b6kIduIkyKu1RKjtWRD4dhV2iMlfkfhnHiAqJa
EGd87Epbp/MB3ak8xVD22cwzkuYlu1PilbnTJaBEgS/wsJvAX/UfDeEcBUHEBw6g6tDSMh9jqLLj
TG26nQUVX5pbMhlNMeOysCRTxOgHxLhXgZvO9xdR1Gb8hGrWnAFWrmQdUbT9Yj/2hka763RKGhwG
TALZgJgwqC8/9y9+ENsiWJ4Xx6d/DOi4wo5yaT/HrMLd+ntKPGcEyd4YeYOIAu13wP/94/WFtQPT
IrvYxgZo5dryE6whcMozyxLd/RFtNhQ5USPeM9eLAlYHlyn1ulBIjLYNF6TlG3o18iv6V+t1G8eO
q0oZcDeBSp0dhJ7oksp/hHzgNQQTjMub3o6FgTUqKSIpavpyygNFP1NhwBWGjTtiK7RxHSG93B0J
Nyq2WmcC+pwH1ngXOBcGkzuzNByNYldoNhV5aA6w8M+n8PgmoNF6s+3aXYF9IsjXM7vZKJO6RY4B
FFYr3KoK18PSZIGwxxg9PAn5Ap8jPbdRS/72oUZ0AlganEQL5jEvgW0sQFzcS3N1mZf3kCe/E6CY
EOiWXVhBMcf2kcyblw40n7Arva9cbv9IQ1pMJHxdX7b1MOrgo3raJaCo1ovM/kKRAk15nQo6at8A
VY74NMmRS9skAuHrFO62yMmb/fudLodvKIOOyfkysMmE87UV10rAkeePilvMXVUB3MbRSoKSBwqL
vez6JIZ/sW9rwr0l7ZpshHOUnWi+gSoN27N7wTK3+6VLBUsTUOiyG1wLxzaHC4DrutVB8hoUvrNT
WxcQq0e+SAwOnziW6vZ3a3CRZ6uj2fPwkxSZM6Zui3mqnG5a+t1Rr0BcM84YcYSHr2vZjSESlPtM
DDS4XKbdaiGdp+/cDWUM4zFZgqwf3vKNybM04WTNDUMOQwqCxi/vgiXZzzIxuyjRhufpGKZHjFpW
W5rclWvqHGrvx/yAwJ0iRVqrmONiJeSL1LnALTdV7QwfJddt21pDojdVGRVFTm6ijXUzZFWO/wCb
27JHHu17BW7Irmc2biPIY0JwDHD6aMKPb/KqZZY8Puic2BrzF7wHuD/IOs3O4JECGi2P5YCK4A+y
yaiuwpnB2KUiN78JyY11081qAVvXFeMTNgbD4LhDbVzNZqiupS+6PXyCpjn0qHwxplrlqSiNXhT0
zsazAkJlAmOFN1IimYEjj3Rp2SfiJH8Q55bbUQ99XJ6G9EZde67gweD8oO7wKtq/yze6x1manGY9
pfPtjg0xZT+/Xi3cH9+ViqP0Wji4f941al8nidPmfAKrYJOASzlGIvzfqiP8+tSC/D6kysIkELEl
NiovnTBQ8/aa1vs2dIcq+N9qQPBGyBWbTzXj0DRV0Y80sJKGJadT7g6644EvASA8G9WkXYkL4I5b
he7J0GCmjoVKiAtVcZRsyRMnP9hr9/AOADoCiKeDcJBmJCQc9eZa3jAhtHNeQ/d7tU7xrLxYN0HX
CrmwRpgZn8VxpaqhKCg0gjR+FK9yi7PscN8hKlMdyVqeTDo7OyPVgjYatF/wNDPFB6dcX0+ni2dD
GBseCABip4VfjKXluWuhfi1Llvy4LX4LNGoS2zkPA8530f1hg50vGj48tela+x8qDLAEqLFWGBY8
HZRuCPwpgrAgs5S0kMWJnI/e9bW1old0qmkt4Is2KftRTDlIfC/eFE13NH1mWAzTGjPXBe0IUJcx
nEjWx42cKrPjqwAxet24tGknPJDP/gnhBNrNk3zHN8x8dekjVK0/wJddP14yEBtOCXhRjNDEnq+n
QRsFGjUAA4YsGclj922Kozh/YXu201tjvGf6/e4HtK3b7m2mn2WOMBu1wBLYppinVwuUMl9s7fHN
nGdAV5NtWPHg5mMJNy52Hw0wiKcj3X4M2FZ36QWoGHLC9XLd+NcxdB12iS66lvtC3T/GnadBEsDo
7Dig/EQPpKhnY2lXq+f+B1Qa2Ay/pRFJU19FlNWvKQbelWl6zUNvbhUCjeiUyrmQ8ZJqNBWeOtOh
xBS9ubY2DVehEF9Ky87yXbwABfU2azDqGVjm1+UKANfltUr24gbswRmYR2z2TLsxs0piaFAQ1HOh
rQ0d36Y+ne0+F2p17b5BVLRBceT22Woldb8jB8vLdodRQO4rbPlrrGABfytxJqtE8QKeWf4JF/UK
Jxzb9pBRYWzBqCP5MFdbIu1MXHrEdPgFfOeeVEWYoTpSd5AgnK3nTGeNVW17x0N9atmAD+25ELO+
Avg0FPipat1PTDDbl9WC//s26Ksu0Y/z1L4tB76Wv2gkgvuIVSgx6huzD43tkyA+9UcY8G8hk/50
rAahPBnC3mtQA3i3eFEMnc3RwBv8meKCTR2glALwLw+Z1eEprLlZIzwHZ2yTO6eaCNBminByo7B4
twLWAma99LcK6uhZ9b1uYv0SJPxfmUFWy7kjLLWuGCynYlUeyzW1AkyxuWGzmtkD+4c/96fLQoRS
ex2ZS1WCcRlTmRWAMCAwQplNfRP8IPDTbCO2pDnebn+Aq5H0JkZVXrp/hpCee04B9Y4d6+qqRo9v
SnzoGhSnsAgahfG0lSsy839x+JXGNMr9uaa96bqG9Du2CW+9PZ5752LX0MBZ6CSVqr0kmJsEoodq
KgQRTdm9Hlw3kEE6Z7ktkUQUCjvp+9OBxHmnYSERru56WwUOoHuG+PfA2scHLkg6bK/AwknN0XSt
Eo2qrt1muGjGlKUr5i47Gp9YiMWBKaWiQSOKIkUfygr4iCsMEnUND8So7mMgCnT46GHIHpnGAFO8
GU6ZnV+g1ePIZlX+F/2oly5DE8twLmXNVEL4AmZeamRP+EE8T4TI7KyoFc1J5KcniV1JDrLKS5CF
60z0uDC8WRUu0HjMvpLx/AEUQm1Jvhq5Rox8Ghl9Q7mUdQyJXeVVJ20jTeclxv/5M+R15vvu95wm
mkPHS1TtTKTw1BvnTxTUbB2t57iCs7qVBW1F/bj4NNQG+UxvuJTLOFSypUjkHvBy6ncp3b0psNID
3PAxzXiNACGWCEr64IN7rKHS7lIeRWFMj4+BKDzA9YGokxXG3Hk3mP6LhCX1IvZ8EFTlx08YjkiD
Jn+mYoOf05A4Q+dkIFznKFq/K4Ctp16HxV5yY5jS+edu2G7zIjRd2+CS8/rFCnR/urM+Mq7+IEjx
xxtghegMcIzgDOOk0YY695Z1IiEvyKYzFxlFCYgjoYOVHFjCgIwqYIeOKpejlb53ld0GGWiElf2t
UH/g00JDo98svyY3jBRXm9MH2i5NkJGgr4TX7KWN/OEvF6gPmzI4sQTQvoq2v0GBDgKnJQLGrFuG
fLiUj5ZgyEHHk+X3fp+UNxH8LlBaxD/IaxFN4J6LFhtW8WCGRKv9BGqmbmtt8Rv8lJOv4FkkiKFy
00Eiga258f5ZUAKAmvWlFJPZmT/xKl54FpSaMcOd/4CJpjsT/Yn1tNmKBZeQtxt280NG/mfFzVz7
jCRZveIv+ykKvRuxrp9XPZwdkTIWsPrM74oO9zAj72g/639HFw7qqyiWdMoP7ARSYk5sCcLltgTt
7fK750EjUfEH0p+sUUP4K48ZZPGTL9eXKV+Yd25qNS0Ozo3UBtN7xHMAfFfZYK9gIEAhxGIKJxSa
gdtL209cSkxGPOBgZVJ8qmWj1WBJ3zOfChKdh9ZUfcTO4W2HOP1eUqt69isu6uhl/hsAL3H8BV/B
kByFWEUs8OiR6+AJfOoXd2JP0Cvv8Ccd5Z5o60lKoAt57GKOMBRc4XYF3+p6k1pUO4PGoQC0idRu
LtgPxqzodPkb9tmpiswEpttr0tUAkNs98MBPmnTMT7HHJTwmKiaZEPyRYl2euwKLvOGHTGGiM5S3
xJyOkQ/ieF9xN0xVVLmPYu/E8I5Y/pWs40LlFDm6UJVuesZqWOcqdVaiTS/9emKHOJXIs5kamshi
GgXzB+CZOPFQZrRSH7TUlrHcnL5SdgYgH32XzCcLlKMxNyejUnLNF7DRpk79K9lxWDxlXU4sgFum
XLv9iYp3jEyHgZYN8EVneZTCGC3SdnMfRwMV76ygl9l5tKEPUEdp6ha5GVe47p+d8qHQZKzAJCJu
g7mK38MBEws32p7MCUY2BUPtFYK9xhtA9H8U20pwCrt6gp8KdZaiXXbJi+qDaHoKKt53DBNDnahM
5BNtxLje6LYdQhzMfGwcMw8I67FDgycMQW1czYL0K1GuOvfp6bcGCP+pvGdqLBMVOi6IF4ibNaH6
VeAQ/9R+Q2KOXfB6ATpSeJKbqv2ekzaFRCaOM+pOHRF+oFnIXz2LQPbIHVN387G7O/gANL5Sg2Jl
JvLXJW+5fODi7/8AnWEIFWAVRuBoNqsRjUxEwf7MPL5x06RamI4CnyAoqot9t6h3Sh35Ncu7D9mT
wwOhCIbJO1+se3TBo9//kIGi0CQmUwh54E1sD0ov+kcnXvzUZeBy9BcfPbD41UlfNtyFWT1E72tP
nPlgQdk2IT1nZXsFekQvEWc02b1H7G/omidSvtE3euGLwKQf8WumnGWaPmBCiLIdVGZzsuv7fl6Y
j+FAXHEIyshVTtt1liujlM4zg0VhKcOO4M04IOGGTNADMeM7Q5CEhycXbZh91t7ajxYYokZnqOgY
4Nn4orQvublejQFNRHqvX2U7fCfs2SscyYy3w6ciuc3ZGRqtxBGV8iiRz7FB9a9HaUWwnXTk8/xY
9+CBZV6SaGiwuL+I3h0jjS2ITu8y+PU2+Wq/NRAT8BwQB0hmtT/nqD3A8hooxgYqWX40/Iq58KU+
bishkIxxm9gxomKBj/frKluh6x4kt5I5syD9YllPli3YKY14CLexGdOPfpmC+Jzes9EQRHKHl2Zu
EUHwYYoQW/gE4ShoVTByf4ZHKICMQcrZp7VsFqCYBprB3w6jSNG8seHwGh00Rx+cdDQHfm0irGpj
GetTBI4o3js50g8C7XteWZbTOAjYvMfnfObhEHJkzyRikVYwEoQYV6DNBoRdMgtqL7n3I9ugjBnb
hw+tZU+gYojMx2PyhUxeOHYEZ/CMw4YBManOJTuWp6Xcr1cLfRYeeIGF/b3Y4aRrpc7B4NoVKXv3
iJAKQZJMi8k2wl8Whw0SBeJ0BvSnUVSrbmvVJWaT9LfJxnWuUqqCcjAVu00OTK/Q8j5QyYdcCjZr
JeC+rnIjwZ3S6jUtWgmoXS1vP6eUqcwWOqkOsQt03HpUbnAmarLfTvzLlNb0RjSVmgr+WMjb0mrf
E/Z+PAzjT1SlUU75FRorp66C9dmPODnloSKkzGY4JBnYNvc3km7QVqKxrsan2qnui86hvUQsokCB
NsCFc4cOsG7/qDkk8XZ95xGzm1JvoFMBEe82DTNvS5zxEeoTxo72qrBuJVEEBxjB969OitKYhaZ5
WjBlCK2/RVGQ9+tffHxHrWSmJnN2wM7tE9uB/gqbxEpT4boNHa/lVf6Y5GfmAX5BKDnM0zYZX0G5
TE7Ju3/pPnUtxZV/1pPyvX1728miWGba/hNPBDxkeWwkKi0+hPPsaCZeKdkiz4USOiqGuUCbM1m3
dTSPtsgVBV4uSOkU9te6NKuqbRUh5O3QCd25UTKMItMCBReDO8eD4iaR5dFcmbZ8jPT4Nx4l9pDi
C5DRzUn0GSmK/0yKMg+Ui7lklsQvND7MbU5iomjxTj93Xs0iJzc3FZ+hgPk=
`pragma protect end_protected

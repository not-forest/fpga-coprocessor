// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
SKe4Lr2CY9wCn3UgGdHk2EJyp6Uaw7iZHX7Jvl+5sGftGd7UQSfQq8e1keu01wIS
9ZqcgO7R0sVEkGf+fXqo8IRXGhYYXJln0jmFSs9xrPvUQy+b4HX+Jo6dC/MOuZMg
iMS7I0e2KGVJOH2dkMzBMY+044Ns9owYTEftQr04NFo=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 7040 )
`pragma protect data_block
+BNE/feOJ/XcMfrf5ufiaZxmIgdBErh+4rUU1856Tm4fn1T1SflHwE+I4s84ZugR
2k5Eh8035geT4T8kEW45vLMlzI38YwblqdwmICoujNo5s+pHcEQ1JD0q9JdZkw8c
SRXOJDUiaTiqjpppMqzC5WXyrlR290CFx6cDon60uZ4wExBdpQo04lmm6g5Gad7f
z68EwB3nK2hsVMgERZ0KWtveA1rhOz7uppQqnN0i3+6uMFYNoJbQqL1pST111fP6
B3ad3mPKJb2Rn3l3j3UIK+1DD+u3Gd+T2KV9TQMtHfuvDYIaYrC5P/uu0gkbPQIV
WolboIvNQyTRScbfExHcCxNzVtc851Wd7NGTURIShsqdLxfTTgRb2ZtR4TaWblnB
7kBQlOfnKq4jAhEPAAOy75k/yyfMJTWbhs9ejBbjOCaevYf0iHJ0pwLKYiyTinFI
3N0sglD5k+UUYw8bHaIJH7hEu3c1TqkgjgxetXfnOPCZ/PIJ/U83PycSfbz1FbPU
htuqdtXLUJpOXekpmwYR4MFdJn63VNmuzjfZ1x1GNPfs2pBDGrJ9u7QcKMKW8KUN
lFlo9S1ucE7v1mdx6Pby4U3IyjkaBo/+wRK/jYc2EdAdMs08/mwKBi9B5oGQDylv
AaJjn8dLJPOw/KArSmX3xjsVClWvRtm5GGNoE3vmw92R1zmimaj52GkQsayLJ6ii
Ly8Cz2tvyw9Y6+3FfI+6o45+c/QdLdHYM19rHXohy/WxVgz+Kbe4ega7SyU07vrw
e0FODZmrHKdrpXj3Cm5Vm6TNexjibyRNJNhIy5e64tG9dNfYX7qPKesKCbPOZi21
eWlL2CoMWcwCBJGBqzsKctNIDqL/gLe/SuRl4GJQTVSFhAgGG2ooa1tK3I/eYJv7
VxHeDelpwtUj+mNIoDJlWhmpudzbpAeEE3kiUmAFTdcywdoIqlrs9YSft+rCVdVK
usPPMotYCJ31ABDQO8voJ1TCANKDJtv7bfGw0KTjPBjpHbVE4OMZf+y90acAhgNu
734/TEWHUAgC0dQbYa8YkaYHuCxjV6D2Vax0Y6j9NeJl+RxI2Tlhi89UWwAekVx7
kfJyyWfYBDgIAsfbzeKrAPPvKiQSMk6YZ6ojSLO34AXJqA5lPRxfvQDCqbZU/+1Z
Hw1p5Oj5Gf5m5OyuXNqtx9frP4EXv2GtH8vrnRtVaPWr5xvJtTzuooBXIZ1Fb0TR
7SzfPe4xsx5xqGujN2NjqAypGC5l4f+EAo7dSNqBr253HVkz8jH1UC+IpL9/F+yo
XySnHlRmrUh6RdkrTcxAlNnn3PwslNRVD4XRYxKzIYep8JGz28v5nm4DgW3mcBck
UX5YPpi/5hITxwfuTCSPr3Ka9SJiurmHUk/E44h6nGflVXGaAUo0/wPoiLeCpSUZ
k0n3jzsv+Y9ytKrlrWwv91Oqbzr9plba1CDWPkWoMXRT23gptflpny1gnlx7FXro
SVTURIxxKqWwRIAM6jzQKOt5By3f+C5bS0URgs2adMpdMHvCeGpOxd6m9rnbXKYO
3cEA3Z+lX4l60cNULb4hoIf3c9VhDSqT2fRFs2qrgwGK2tfEdh7hxvGBA9cOaBe3
lztSWKfyvLk136x1kGE+B/cn9wscRftMBchTFaejG85NK33tsXhB8dVDencsfm4D
txw2lrWSGy+kE8WSY4UBJ0YZRlz+ljefJtEvbBSPfsWM68whyRizlCEEOivyZxZ4
PYECzZpcD8T77h3h2J6+WDJJjP2I2HbnyKcIzAtAqvbWl594RU1tjK2IIWH9EeEw
7I1lbXW/fdbFEA3SdAThPuNmLbhssCKo9Mx5c1i4VBGgHABKMQtU7yF2+iCkmRfJ
Ribvn8HO5E45fGev6H976JzpgcfshzmsmQsvpsnIUDwXrYk2YdsN9tIHFTtTCdnm
av0lRcG8E8ZExciX76upY9SKP1HuRdgpNNjvj7ftKlqyQCpgpQM/mSOvJ5R0ALIp
/Fjdq83fwiFhv4SA+W9kpMAsRagl31Dy2dLMESSGgDSRYOGkmZv571g+qqtKqiV6
dDH901BfQ6toInipHkTmGx9zffjLw0R4e4pBRutVEOLdyPRH83SGNKd70Gc5puBH
nmS146+0pCwRwpmHJOJWCAQRzmSEJwUGOK3dE+ugH7VA3lm5tMbhKfKjY7ZfbQ8f
UfoU5arfhviJa0/hSB6fREhX/HPbALwaKhMGHHTz+GioiLHn5W/ZUTkIWnMJi0j4
9nx7KbY9Q9NcSg4Mr90N3RFkRiWT9gJARD8Q7cWxtAPojiG8XU4aSl0OtDyFFpgK
clERQic3Jo+4+TB53HU2PpDt8u5HUtjQV1lRvXmqbe05zNWthEGKyF3HId3kxx4v
Pzr9lnbxY2mti0RPtnK5nzu24x5Vlx7Xh3FynL4hWIbc7ghcB2T2MjII+0yCAbXf
tIpRi3iS68Bh2Sfst3O8CHC/kV7W80EUQMdwyHKUpxFfz//vl8kt/5WLtvJiCrwF
LVxDMFRZioVMUxW6EPFZ1XK3Ypocp5US/mgo7oaZRU6pxVBUIg9kHkh1R3MwdL4T
Dt6xJQM3ovZBQ0Xo63aiDwjemVzg3qKhEmAG4q1l9P9XVV5/IxEfY6FHCmDJN8Mt
4g1crCFuzXeq4O+/DBwAj2rCkWjIzqj0jYfqIs8g3b0q4DpkZ9tXoglSdFXDCsyu
H2M2LfFJWplpoS+w9ubYFx6frsS1Vk5niaa6D4wLLQsk3Zs9AKNN3DWwEOMDl1rU
JzTl/OxZlYHlpmLDeBoDnuulRANkFxhLo4NRXObetdBoNvplLpyX9JHwwVUvrRwr
2loYmQe4Go2dIddsjBC5YzcZI6kyGvJrL5o1L92Qk8cCiOv9Y6O6rOIlXN/aC4Wz
8owKZPOYiUkJhpyiMzrYcpwxjnzLCx/Cd2VIrQpnc1jKgdunb3LGmYbb7VEY9a39
okKhWNY408Y4D4DED8sPILaPfq7vTKfU6AnxKJ7mgv/3UzLuSitCmrRecQ3Hr8SV
Ku0RE6w5cZIYMtoxb1mJeZzYLLlBzqyhQCUfrJ6eiHDfAwkzDf37qNmTJWvL4Nob
+OucNr5rutJiOxiKFLVZWCoffVgakoIeKh+hQqhyt6/VapleelcQVCeTxSHiN5IL
Gohosh6IB8l5AujBjmhL0IIqP2QoSRzmkeAHnNiu93zWJCheTIGRLZZhOaRHX/qI
157PCZjNFOvwA3kVhDI5KJE+5qGwTiqlVU1LuUKh62uclY9LZnAyh7DA9aUZFonJ
Mt+9YvQktoC378hdljKwxYksXqGRq7hf99INGbRqMD9HbVZfl3jxMOvWXmpsdTPm
m8MKgELUw5ttkrLUNppiljEvov/g3RK09JV+z9nFFIX7FvjYMLucjeDqXdkQzmXu
trBEgbrPeT8SZPbv4Mv5FTDGRn5UC5qVenZgRr93omXTlwSPch2uDCW0N2tTwd13
gLIm35yrsf/K2+lWvXCmRZ5vAsYOIrdQ+3ZwsBGe5EB8y10DgJVN+WnLIuJ1u5gD
Sws/c+Tfhtw9dwNShFXgqXY+RgO/OZb3TMHL0wOOrOF34LJpqIroT0N0QVScLP55
9ijD6XZXoOuE0HAFYL3HWFP6VEnCLHNZxOcrAkXz8ksl9kxeIeskvNh3GF3MBaTo
2ZzRvqKMFt5dcOFj4fdrg2rM5IYVVuvazW0oO0xm8QYTwJP69G6ZlvfctgjgTF0n
c3Fat7ozn6R6XXZqv/oNZf5nBTsbC6qVxVXhYGPTAAIIAwBB0a+SfL2K59UbpQQf
kshYvHRsVOVlwTI7jjCq6StMr13ALaASkCW32ukBvq0hhMxgh8q1+NP9cm0FcxTN
Twpibyjr3+qfnHVZJWAIe6LktZAimQaNlw8AKt0z+gbcuduYlF2otLWNqnQ7PQ9s
p5f5kDQtcubqr9oaA5QNsP2uoIc3h1+o9Tt9e5aFfMVuD3VoAYWE9Mesak2Q+ZIP
mmL4C5CowI+6Y9oZo/lcfzkSpT4C6q4/PwPWawZMiDb0dGtjGPBs6PYq1d35W4VV
YnW6rXp9DCMYcfwnXxSp/ojbH56TC89ohMCSLr6REvWWqoytuTQ+HhcxnQ4LDUKV
SDCIU7dVJG2Ok5O5yd6Kg+MsQheehLv5fbd1l2BptqHw3VBTD18QVBAvKB7AfDDa
u2BzqmQQZ9CDJbTyDUwG4a+OEpfNEfLRPfO3EtW0h5FDO5S3fghC/cYRT43GxCok
6Sm3ATcc0zxJ46GJbkyxpkLJ0aPdg7D4Yjw4CD6N5scgk+LWRnD/wSGyTmQ68nxF
F5/rAM22iKHdUt6NvwSDg/NeIkC+uaZd3sNpGFOkRwdlSsu9FvUQJTk5+ysx0A3q
EFuu4akRmXG9vO4RR5SqTTco9lg3yKOVjX5KvfYQ/5EWxjmzRXE8Dg7N82yu3WSt
ra/E9aV3/oBcELmBmwBaGXIAXC7OWLUyF20OAIRByLHI1MVYxWPFLsF3a/j12bJ3
wlrsBPkzPbkLtgV36m6Z8Yn9F1PWjHzP+l4EW9/PWJXHHQfAqvCHiVhaVONGDAOx
0EIzsb/S17ZZ8sXkYJjujPvVAv4YjivnCWWPFkz/OikuCydXlvmzVIgCpWPUL40F
cq+HXYJojdh77Fg2sMwqTvr3O5F3OUOU08sSr/c0yxQveusc9FVEqPANg+IJzYrh
3e5ZHpKOalrIad9n/9mm/gFgfjiTVUQ0CdFgkYfQUpEAwGNkj4Z/v6gn6JZvTRiX
blrCLUwfLfMjKU2IZtd28BFTCpv6kpwxr5HpA3IYPu2uZX8n4iLTaMkwY6Fpbr1y
bg8Rs0EmOGlLUC0nJhERJh7u2Tzd8lS1XwPOYuNrTFU6lGpGlUpqfP5u/NhhwEmM
Nxwdy/ixkVVQF+yvMW26WFdKovF4gQncDS71CUfC4gCg96BXCZWfolRi4PCJzPBo
7UuFaSYEbDtZEy1y4n7eSvdyY5ytQYIdMciq7DTIGOGR7jn8ZJj9wzs7+BUj76Ig
GPhO/pOqR2+cm+FsMP7b8ReclnT3L8ACbjZIrE5KxxEFp9iaYgkzdrlkptub8L4P
BKCaMg4TQLb8EXXhgzl7Shet+SX03jysG329kXyQKNEo1ApoWFNWdfwjO4R7sgOH
oBpR8zrOtDDQl1JrtIzHLSAsbJMESIalnYkkINdf2qKZA/GVQayvd4+et523bum1
INXo/JBpknUYxbyEGUex1t6qOCDtTOuBYV7kkRa3HHzUlgf/4dYEab2qVE5caguN
Y3SzQlNcWFlKGucOiKnZdDdS5hgM8pqTAyCrT2zpoMFR+JPghQOHHFHAEO6k9uDI
BTMheF4tXsBLGlAFv95AVvB/AK9TbFWddrgk9nfhbwYanEZPXYrvynM+ND5ekjR+
kLjOVZcUat2y+fppj4lSOBQW3GIt5TfYH+xYtfflCe9aiVX3Z7OtE2KqvldAC0KW
kSk2JOYXDUtayx1GtcVmUnOl6RvCTxrrhfC0LcG7Ce4NbGvehT/4vkPlHbWjWJnC
NdPx+/VsDGAPvj5KX3A5IAM/8FCYsL7QmyHlU+oLI+1csxesswwHcPX7NJZsVMQM
IxHKEIUdMv7lVuKOdVGIqoMsUCjoCiFdjPZeRwsDZnkP0RwuVkeuuSmPHYqVZbTD
ahUZ8rqNcGm4PdWZynT6S8MIQtXh3OpY+MxRJI6UpzbxmpcB21xC7XnPdnPNp1WP
LMUciu0aBgcv/zk+qXNtudZIbjPGiQ6qyokutXlv5pGk/BU4V2CXyXULTaiCbZJc
uvc241J34MEzN4pXoEbyb+F7OoS7uMfaXcB59CMtYlNmEYQGemnZe5QhCIjsFJXf
r5m0RE7MWkJ44PJKoM2/LjL0r71cQ9nGgz0awsQQ2PZvGtLM4nOmiZ7eC1LImupK
cTqpkAlPwxj4Nw46Syzi5O3R0Cdxg3/1eITtey9TgrAVKixKdaR2Ai+DHYfhdxQE
PIOv+zptAdRdaqG3TMITPt8ILZJugNh4jMaSujqZhlfG2Wa5pDy04K5ryvMX91B2
yiRshnOoI1EKB0H2CVIIBLVr1fYNnHN1wBgUj8gE8FnN0p1pJi1XJwrHsRVHi7Ax
0pjq9bC603XArEqwAPa3f6PH5cEFaubwhe3W/PmTbXAGE6jx5ZePDIWBOyY6ZQp0
KRFpAhKs/1G1BL7fvMsuILf+8LExH7u/hR3NMQz5SRWJM5mIbW8MNh3OUdE/vybW
RIH1YzhKBNUosFjBgZs+7jS1MhgSu2nSc3FVcorUzm+s23jn9T2EhdMLXqrSB7eJ
s6wtVtlMz9rqrgpOjl599A8PlzkRRfIXL+YO+WlVCP219Bb1mR/V8RRmeAgIY0tw
2+Hs4eM4IPFMYrax1aJJ1tGT0ng8z8fawaXzUmx2I9EcOp5WhY2fz8NPBse4TqzU
Jz3mbIuvy4TCgk1VrUtoUGHBey541cdswz1LDZFkdQzg2aDztBA8T9Eh6ybrkLVt
BZNW8gf/erKWJois3OoIt5INQd/N+9o3oxH8XRpUH41HJvqYqzohztsWXOUhMYku
92NMUZPcqJtKawUWyEHrS5vHK/dAfGjS8MwfpgkW/urcv8j0DPML1Fy48qZJlwvO
D2BCcvuM7sF/aNTkr1RJe+FBVhW+RRyDTzDSGh4SdnZlp/NOUaa9Dvin59OUqqyc
LQo8V5hwY2vIppIr9AM0w0eMRfopQPpReJiv71daTb5rfCgyqcp4q0wiSTuEZ2jV
l4gh9BxbKzGZEsrd5BuDxUYqCW3DTEkar/wlxVMw+CJP+Jdq4lLURDpwURBIBjvH
T53r2cKzGzbtz/jW7ErRh3VEl6509MRMz3zNU+9A1Bb40pkAzNCiaYEK+GlU+Ebo
6uShrCVjA5N0rhfhUolQTsQ+0rngZxUalfZHjGoxKI+rPjnE12ATgAHV9BzbDGd+
vpWXQ9jqYs5OV71JmujVRtWQfOXWaLL13a5S7sgzZc7Bf+m9LpMqiwexTmL1dJs6
DB5Q1i265oVzNADvwblysi9nes9iQsbH+qJipm7aGyPRJ6AuLwqBusWi90dxpEeo
wthyAl/nk50xPSTNFnvF3eDJSi32akcEQ0iVb+fG/fvYt4fabhM599I5H6nfS6AD
9xCAmAW9QQN9ClAINQNfOHMFfIPRXrIOsKT9BB20c72nAaOI3NS+XhDLHafOJA6d
DGL12rGJm6cAjdDHtj9ZDIfIa7ryWnb5nu76IhylFK5gfT3vHy0BihxZl0pmvx4d
FgLaA5h7y4PBiyMaIIqgW3NQ86AJQeA9NF3r00Hc105m/mchaLAW/fOF6wpaDaHD
FZr1Ug+WVQeYhinC2kYSiUCZKEj9qN9sth+6ytlMOmORxnrS1gCsa/3ocGxnOjq4
0rNpy8lVM7HBMHfmtx0iwb57NK3OZSF1OQ7mKE6v1gnOwiaINQmZd515kzCAMqUp
5qYK1YFiwaMIQn0K2jH1q8OO8N/xohXrQ19kI84dTImUYE1m5AHf81nYGFAFsz9M
oOh2UlBx7XPuE/HjzBqjOZyMG/WHjF/WSybDjZeZ2fl6MaFl674zOCOQbO2MFijS
hMZItQ6kk58g95AMYIud29uBGcVhmw/zau9W94Fx2cukKfyXKzSitcbRcnuuAueL
6EAeyFoZYgh9vr48+aHSUeiJ77TxnOw3lqmy2w/ng/WNCUmi/alWzJ4kSAyHr+Xh
YSkXz2n0ZGAFt6vy3L4AFk1+eG/kPTUeT0qTzfhcoS1wtxl8rEgJE4zh2pFl34u9
CoaUhytd4fuCR5E136NeLt291BfxzWypJjFEbKc+7ujb54pi/f43Fy7eU80Hfjch
WAHVAPzA91u+a3OU9+WJPwAiOnqrpKZrqgJeoFKYJJEY3YlQWEL42Rd4qlk/wzVw
lzBoE50aIXO4yvGz1xPl9h3CLzcV2XzYk8yEcqjWUW7Dd3xik4XLYeEpjeUi9gsr
UobJsakYTKgtT45BeS1ayeL/PgJ7RTucc3E++Qs9S6y/PiXN+SnD+yN2OUkUEif4
/3m97tbh31Wk2VogfPzKdoim8bMVwjjHDdA15TFBHBLDXMOR1rSqky8hINcoeYaD
FNxwFIgbGuscSU6P4khBLS7aqw1/GeRZZttQuI9I2MGc7HY0bvCh9u3aSTBgG/dj
x+Ogn8W7UH9Ou2ebmYpjjL6Eqd2HZMiDc3Mb0Z4od/LwIWkjKUjPtw/sSXsgS1OB
bHV7TLmxPD8cKztzSgLnGVaGQHA2wuzSaaCnmbBTr2aUOj57D8hQd5UY9KrlziIg
eecQIhnwSSK9jIRw8StlC/sj9/Zqgg5xoCIZnrpXcTrwui4ZGwBSxTJ4zzwNxU2d
3UxBKMLSjUpL+ynLJ96ldXXNu8mhzRAki/OvJR5WHV8jjiM3ql4sXMh5yYkVwqYB
dAqTx3+R6oRTPwv+tZcZwvJXfVBrxSlxVTxP3RDwhRRKhxWyXfoAirlmuxTksY85
sWA64rctJX5kPFVTg2HXXKc4nUUeG1ybGGERYHVpICShSh50n4B5USuZ3S6MCMSJ
3XWUU11wztB/SImwhLC3vjnW2b56zmae+HTeTTNuDizXcxlhtaU7W2kvdte1ji/c
XkaRKtHlHRhHYZ1Z8fuUSXev/yfF0bbSiljR2SowAOhjJUSIzvI/RW/By7kKxScc
yldcDx0ty+5YPifMxeycn/KwQwrA5xRPs6HIwEbAfnosn/kc6PgbTtWW6AcAfBLE
UTurJoofvF/O+1agjh/ULm+PhuunJV2wWms8pJF+7iiOo/LiFDAIpPoGfC7WLayi
C3W42h2Sp7goQAfdpew9tS5eItddvwnWZZyVmJrWXBOkA9ASc2vYprRSnwQKPn89
1XMS0h1qyczzT7kjF6JyzDovy48Gdla6FdBYyIInAKiQzCvjniTCF3s84zopb3Z2
r9JPzpD4W14TDDLyoEPiW+ecE6wM4CxgrqbmwznSvQdMVs2PFNfx33C84oV4xCft
SG7KDDaGtFc1QiDbOwF/5XAsEyxkh2zAZNdxMOPQqSXVsmsbfh07jizTGSHg1aLA
LGNs4vTLaj/4QgACtG0VyBqO1muoUbY5OCQ889fYOq5f863P9kFbEwp5p2FdUFWn
ahVM2eWvkY4L4xo5yfmnFO45chznqHSyBKas86ScVr00l+a5NlQ9Xu6FUwLbtpxi
vB2lVz+d0y/8R64/JE9v6cfHdHuqp9sNwnlyelePI/OK4jIAA/h0KT5NGz1K/M7u
fJqIFlasebe68eaBzCwY1+ljZkf9utFV/lji+4Tf7V4z562cmtIQCQQ87YD/YM8u
eKWI4lrqwOlfh1JYRhjBlK2AMdR8Vy/p9z1/n3fgjs4eDrIfcZlxjipjTyCfLH4Z
RnL8vs6Kpi4ICGPCR0g/NxwG2kjbtRVDnN48sHUaYF8=

`pragma protect end_protected

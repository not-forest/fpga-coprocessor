// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
TWAbBuewMbgYaLri1UdsF5gNFSSDrj3dzdlwJizytTs4Q+CzXg6LyRf5WX2soJLo
D3e9Sk6MGhd9DTUzqfkS4su9spK5IXh3ZgqgEQDfXEmamJZCNosIFT6nRaxCP+LV
I3nbSrK0IFpb7iFAuMjdcYCwGwAMRKNrR4Up4Ny1MAat5arbOdzQDudL8JxlQFWS
VNz2kvmYRIyENmEYNI9/roYfIJ4cX4Zz/bbgTroucHKuUa79ubLh6uOlF8loss7g
LVKLAUXOs2tcyv0mX5ErnkgPl1446x+oCEpiG1jT6bB5LM9ZlZeYimIDNgkGrG0c
CliE7KCtkCQfkJuUR9rJiQ==
//pragma protect end_key_block
//pragma protect digest_block
8BMdcMnIU+rgcvZMdXypAGgmpYA=
//pragma protect end_digest_block
//pragma protect data_block
e9qPB0WE5d3Ud/XJq1gvhnW26rjQucFaWJWJegWCAQlEYf40hK4XJizBYSyU7qQ6
M2uItFe8HAyk1lYcZR7k789lE1Tgy0pJ3YRbTUpfAzQjsw05EdZa6cShZJkGJGx8
58s2y0W0EUF1BFybwqndTQYcwPL9NP1i+RD+eh043PtwUrtg5WvpxaVB66fOEzv4
Cu6TK2rAiXhNDpfIRSi8eopK7DdmhMArkEGHhoX8AWt5v3MNXh4hOLr5hoWmXsdK
WcNh9qzPE2/BTqa+w9f2NPP0nY/kQ6Jl0d0odJA1TKzGUnsq44DtlMXimfV1fV4O
TCjxZqRsLMeMWlCYNt9K/lftG+UXYAMVnxaI55qlXkY8JQOpzHTws2LeKK6cr9nK
WJSyQTKe3ZihK2bTMg3kSFT0Xou00PogiTIcUhadwSk5npa7XfyR5+U1Y0s2NnRo
MDls/j/qiaH+praouv/t8yJpZ5nxUxxR7SdP5B1KdzV9SZmr9b7v5hjnUIyz/cqB
09GOAmAzIjdiMx+OzngVyYAXanMfJl+dMXt6urBx0Zx1Sxa+HmiUFii7ouwgMVp8
lTu3Y5Lpc7tAm+Pk8gLPKXv2LqfxJpZ2VVWg1adXjKBJsbYdWKhGA7IAW8LA5iem
s/whQg5TXGps1OKJuwb4S92bG4Hsm75tFGKsdVyWx6c2pXya2dCGLkw5jf31wRxf
pOp2zxfPYgfpqgftKg8vdHcHXF6kBdwYD0Onr4xn5/ae4vQOrboippVQKsr0jx9b
hKzhkwKF0A/CeVAykF97KRkroBP2LJgdNHsnTuVq9ydV1rOUGgHWn1eLVDaIyywf
oa84+VUKWUZcUZ6D72rP5hV2T4yXyxK7YrPoZ9Quon6r4ErjMQRDjEjsiQP1YqJb
DHweTSQnjKxSNznFe3VW+jPckR1zF2LfndDiLKqNoB40+l/dn0e9B/Aoe8CYQBMq
ItJAfTs+BLF0E8Pi5bs2j8oef9U+r5+XmvdVZ1wt4BQ+hPhJT0rnR2dqN9lSV8Jw
Vb4o2cI1eG0sJ7lnijKzpkUh2i3zaadKMxeAbCBvCjlMIV7rPDQJwflcCuv0Tusx
XzRJ8/dhV6GRuk9upRHyHoLYLz+C63uvKYxN5m7q2xxmHVy6owqA5YrOG8q7KgcI
fFZtPVzCrMdgMozMuy3Ah9kQ5dMtQndpCvg3U8SLoL8rL23wQ3vjFtRw0Nxy9sSJ
lfBBOpKs1FHjl9hDmoszMC+to99NisorCPNilKRmG0hQ7I+ICBfAd41ze+q3hn6H
OQL7oVpwaq4TJ25ZL+9Oki1XT4IJLxd2ef/uQULEwUqZgJhPjPDR9IXmaW6Go+Au
rP92NENLMeI34wMf4HRZfZuKjrpZaIVg7WUMr4rI1qDbP6+xFhBC9drJNC5TQBzL
edqMAwEpKZvhhleEbGBiw+a5Mcm13ZHlgz1Lmz4CDtu1BCauxuXX+t9OR9XnO564
H9bwS+jI4Pzyr3D2oFwCdypjMCLOG3h7JwHIWnx+ZZtop69ibYfEbm3RyqN6iqDq
+2om+BNOUePIThKCB/fbSMeTOOCAz2gNwKUnnR8xb9jIiVvCi6HN7KG79liQ/hDQ
DTkogSIf8r9QIN1CgKpGFYnMuFaOPsHvmdN5SvZ97EKs4lha5wpjdWHkRBOMPkLL
enlX5FLDsw+5vIJ5TRYyez2lqFCYDot0IYnMvr9fZ2GLANADJQbSVwtbS0ZFuL5b
z3FKTPmWB1yRvX++TQE4QVnP8YnZjbF2maO4nbPh8kH7OxBgh+wEX2jxXRnX59a2
wuIVGrfBoe/mssbgCNgXc5SYCqHnBVZOXptAQs9MbJRc7jBp3+P/2AEkNPGHxjXM
oFhmRHhd0NO2Z2ip3HLj6k2/C0b/ArdRWcGEye0CX7OK+XiGnm2C5h4+5eH+IMno
6mcuh0ypMyek0Ph3yx+o0i3+C1xgHoRXNs+NXbI9TZLYZFQu87WU2Y6rPOuvQu5T
0iCMFARnxCXZo0dedRmd/A4augF/naalUg4FjKMTGhRw9ODfr0htZXP10RQuinUB
DHCMDmbY0/NLhB0bNygrZLx18w6v0T18S+tz8404TYicwZyjGVwmgydumppnStqF
wBFGqnsx2o3hQ6d1eVkrjLMdSBFAGfmmu4EP/eWFc8xvW1yqs6kTCiDxRVfqldDw
MJ1iINONe/YLkgUPlZT8iQQ2vTlb28UWMm1cyC4r46aNSu95ZNGzNRXn9MIeygAA
Mfv+eJnmHLzuIfwrNAQtNxFAMUpvlPr0V/AizQVzOuvRHkCtjHFcNAoUPiM/VfoH
S6J+BBm/ljJUGag9xVDo7Xv6YVP9UB7b+Ep/73FAAesaXLfC/clNlQf8rhLzQyhb
CvdO5+LjN+iDLRf0I/KtW5Twl4Ue6e7RxlzdPDeYH69D51ZKPweWZYvzILTMgnwJ
ZUXabohC/PrDvudYZmRUQH18gxFn5SBjxeX2VNxgk4c4ntml47umSmuMm8oK4X+5
HehZO8vr1xi08oy1dhvO+rhd+bBsm09JEvXaeabNXm51IFMbgZxYOueFD5TwWo6H
gvvuo3QN+OtfDksIakXdm+r6ySiHHS4qM4girHHIA/d0vi8yRrAtRRXAUfw8PmUo
vmigzZXB2YOCfLejrREuRao8fHVg6N+wHbYySmI1tup/CEuJ0wiDJLei5xikARo2
XvwdsqJ2QqZlmRCN8iDbu3R/eUmkHfCXXztr+98lOrBJV4QeXdzwDs8kskJr0i2Y
4nJEajw75FPfztC0/WjXfY7l2LAlztGDYqMffhJxCLzUjbtd4wSm1PHKoBf14H7X
xzPNPIIhc/PM8lPGaLGBp9ME/smWzU+8cLTxWuKOJt/oEMaGhlnmvQhrG6dhxH16
+iUSGfL53OAhDQNyDFCBzoBQO+qUk2fce6MafLaQ+WD9NsUImQJ707xCmUXJG3nb
KzJmWk+FJeeqavy1asn/Qabvct8ulAs2sJqvE31ZjOF/uG+pUtRgr6JvSVYFET3Z
4hlMDcy1bNLUpJxAIkKXyi/waQGhWoch0j6G6+sOk+Sg+IAgxTibWG5xIXv/4C3l
ggSGq+fQjkukHUjM1x7ODn0mLxhqRIF4tzAYDafUgzfxwvlrc+kIf5Oi+XZIsGL5
z1e0bmP0p3SCom/iJLy8NZ5hLmbp+Hae32YCyg7GrsA43adxNp582bYgTB4veaqG
RtLIJAYe6B7IKJM38J3gZ9KSn+UnbsGb31B2wNKWw4KC3Hgv957KRIGEEd2Grpjh
VTadoWW4FFtVId40AZqmRic5fBh3x+WMDX3fSi1l9Wf766tJtYvnz7T00OWv/2Gp
MLQFdI1Jw44zPWp91EqG28tIIiCkBbY/bwgC+UJp9Wy2xVdfKD6uiHGp7EcYR6tH
1qHNa5qGq+KFpJ99m8kiYAPtHRnl3E3N6G1rqTLAOINjnDokPCWbsIpOCuNpJOWI
myJMTfRHtWH22V+TsyK9geJX2wWdQzaKi2YwL+ge27dbp0LwLjO2FYW19/zJHwOG
cyA23w1lc1S/lkLjkaQBapZY+QQcwTEHL7Hjzasxoi04sZRgBdCiVqod8Znup04i
2BDVmG6QNFWEOxeXTvOqN3H/DlKqv99NMLCUKgrK36HknCSxCji5BKmKAFxgLMAg
PCRTJCn7F0Nk+BbXWfZepDShS7eAxuzL09Ohp/pVNhNs8aEAQphJjAg2rASKPr4P
OlPYs6AjWi1p125hE5bd8qc39ohmWlsnsrqamF63kawKuAfqXx6e84fb6lciIjlA
SDs0E/QDArfxniupBfKAUZNCMPOJTKrIOh+uvsnHc3dcCTYybdtvTxrf8sh+6h2M
VPSoaWbJmWBgARgXU9RT0Dc+A8bP81CJzJvRgDzjWg594zBlhkqD1gQjuWVS4lkE
zyrYlK8AVxH5lstLIAD7+XHXZLqHzIgg5auaNMkFXjzbZ9/vrO3WZx4DofEPYFSg
jlG6gxF/G/Csgez7QTrnPdsl7zInrNeNnFItE8gCRSN9atQqFV25H/wC+oMcyv1I
bXjP/Zr27se4SqYHkTkdMgaGYIG2KkIW4yrIunkuC5O8N7twJEijmTN4Nknp93hr
JAgF8KIG68DQd/PVz7586jLEtlfyV4Uo64yscaUtDuYEC8XQUg7KPQNDwJkz7r22
D4dKRMhLjQXpn9r7u/juO5XP0rLW2gfknnFr1JV3Pd7XZHP1YYiirUY+uaa7xSlV
jGxnhhF9LWXPuUfKv5fWamevHs62fJqyYXqcvc5qhD9TUJ8e5uFQoR6xZcAhTp84
V3DbdmkJqTDWXUr+LzHMcJqthKZhPxsncjD1dvj7y/l9c9erllX8HMFIlDtlfd9E
D7vH/26NKLj/HXKwmJCO52KeI4tbJj8mw43mBpIfz4gb4H4J+Z9oq2bvDe0vhUPl
2JjKoxF2AckgcVyjc1g0meun67Iv6PjLeB2j5kmwOXb+V9ddoAuw8lUUNwE0iQfY
uOjW2IgqVpNAi3UZq8fiIwcqUlE1e4RXcYfgAW75bmHOErcfZFrDOM5n3HBF1d/g
zwZK664pY6jaHfvawXdrZT5980cz6WjldKXEuXBFNvLdZrxNUV/3rrxKXD7Q6OGC
LeQf7i2LcA3W1X/wXkvuGeeKsmhcJtNQ3IAnwkBsb93x4I2zCHsF3zts+QMQ4oEp
5TGZ71aGGm8WqccTtoUIsT0cI815TWu9Uzg2ylK6JPGVP0Ap4TS7adMnJ4QLqQtP
2eC1G0vwL03sLkkrD9wgDF9eLGbrhtweVXqyoktlMSvdUMGCJ2NZXjnc03SAqUB/
EfH+3G7GLv3usxaUfeC4in8700jlIe497M19xwxLrp4zPdqOt8sbwKGMXxMp0F+2
XKeOd556XkZg+tt/0iO3oDDrDbrNx4E5zwiqeSlo2GiquyLEJGD7RTFaZY2v9Swo
n0M8BjEd790jfVyTCsy28ML2qduLn7ITW+W6z2NlAdBv6SZNPbmN93sIuFlTd0X/
JGGbF1ISKgbJzql1lvkCL5+vyuQAqzkINm7/IQOV7LnHCq4fpdmw3d/WdFjx/FJA
ZJGWBQcKmDXdRM1ZU+ErJ3g00rZ9ak+GEZ2w1NfvxBsqP92QOF7qA6+17d6Q874m
tOLPuiY7wdLd4wLjaABYYQvEwVivFOpLArmmQagbaOhc/toe0geySprNScxgc+5Q
6uneLMo1GHjBdJq6NRmfm9vv3HTksxlToVaWthfFxlUjyRD7Jx0OddPJ4OnSIqDD
aIFTbuu0SQPFzWKAnK7FebtzwHRqAyD+NfYIthJOWcfUabUtS3sBF76XOMZSYTAb
vTOKNHbL8kBJc+SdEY7yeL0M1LGYn68+q78zCIRwST1F1f8tPUQIDVhKqI5jxk0e
EdTa0jzrQIMgFiBGWY7UDsl8wRr+Cdp8vOGivchUPGzy6gLL8ElC0/OezUAfWrf3
tissqDdy80GeOEU7reQS5H9EYeR9pF+C+Nb2BeXkHm71v3cWqT+5+NwxnzztnMkJ
8hLKbv5Rg/utVN+aDUaQarZ8WQem23tp2Ao9unMWBAB9er2pUDUg6ITnhaWnhlWA
KC9Nw15RHAPf2fa7yPH04JxFdXmlaTbm/ZpgnmDGPGsaSYZY011QBaEFLWOoZvZq
s8G2on3lFXYVUewx0ty4iRhSIfgq2ZRR+P0ecsCQtUMeXr/jKGPbyWNjh/NQMPc3
8MhE1kUXedclN4qk6zm3fXGHApa3fp6wDhAHiDsvPRMA32jyWtYtZLp4NThF5ThO
9EKmJRsACPOpzBWDjcRw3Jqok79shLSGpwIuBGXnjBlae+62pAo5TYi/UiBfFs8U
uHfpnv/IWZIqeCll0QdpXzpZl2OoziGmd13ZBW8WmiOVKZvfM0GTaz/reV3yAS61
4XQ5B7FLSZzE6/zWoHHCbHhHkWoizeVktpeIkCiczXA1krW4ITCNfEoZ8Di4KdJJ
DS1KLYNwRuUPusLs6tvnBJVa4uNKFJ1wSAaQ/2pBf0VZO63lIYYKsIX9YAGjH+6n
7TmVFtipVXJdV1VyMeitm50jL+C5WBUBcyTQx+mVZLy1pKXHNeH+IV9v7zRXdcOX
rYdJs38PGozzgv6/THluzn1iMRaaASgeI+IKv5mJCasgjGJHaOLwl3D+c+7zahFl
FsTpj1+V/Oho9OYj+4stfCbs09r1K1vPmAGIUHemEY2mB55V1QUTvYSMKtw+lJ5Y
8xpSqtpZrjG9n4xOVFxV1OMdD7Eg/LljRQbCamFcWJPl7UTRR2l3h3icTwTscrCS
2Z65MX058p/UVugD5BSk175yCVckiJi4CRxCHYebunf4wDzlXPGbkUIYLC1DoJOH
awdbsgZZUIiPc7p7Yxy6uWoGVztXK3u4cl055gRcyMsZPH3K0n3cXPXgm8Qst8xh
sMQU/7K/LEio86nnGUC0qItyyY/NqVABBValSzHtciYOVG9hRlqmsP7QB7F+yJY9
/eKr0wTBtki4hPdyN5+4zqFS1qCXrw4pp3lnVvygFR6035wLiKN+NE8INeV1NB/O
U6giRSIyYInQWZGOUretmJxVtA+eCPIAEI1HsvGSZWM5ZuHLefPXsZTGGgvIMG7C
jcxLbn/CQkWRnlPxaa1BNUJWfXK21hZclhWcKxDEGw51bgUkE9+l1739c7I2JgSC
TDvsMD7LmRy9xRk3wRM1d53e3lW30FYDQ9bT1ipZ8SYTOqCPSYDWMXcx04LgGZxy
CXXgn0en9MSFBrPMo8C00g8LwOKCsVPjezC5+L644GnKdDFpKQanP6q6qrPG6Vmr
uwKKUkLpwkS76FQPwvYFzwfZnYS6G8KaZ2AOi8ytJsSAmQIOTVXpBks7+4z87wRy
Zz4ZVLO7ZLT093t88gH74VxoGA0jJkUAA0OjLsOIs5fyBu3uJVMUHcLWBm9cWz9a
xUaVdqVtgHM0LR4DpJVjaV71AOHNA0Qlwu4LQEtAWlC/AKwpfSnxbq3BXUUT0Px8
EQmivEd/HdXZRWc4AfEn6OXEIuxsX53x1JYJnJRt1VOwp3XSGNZytUSSybDr1mxt
Zvocg5bncYt0yhp/JRxayVRdAXhH/A9VnkD1o3kszgTAUHUW5OvvouHAh/kOLhXj
eLCi3POlo+Tmw750w9mNEiaaUM7gDvGl1goSmuOD/5LggPRE8sxoveO375kTHBJu
8iUp8hJhPg+Gm+Jl48xWuAwQ3iyycZfH+1PgzAS3jwpGeovv3GfOWxcU+1epaWT0
D/xKcH/80geQSZbn1F3BHMaPy2YU1Lh9shZ2GALFAEd8o5hBrRmhGxlJU0/WPmqv
Yb6b242e6576uaRzMg1sUjWRqxQ1jm8NbR7ONueBSvzSNpfTCvKLd2SwxR4M9AVZ
FFmYuFQZ8rFLc0nAeQ/kZ9XY/nzlMrBXQxQEcnCHEb8OxIJL/qkMLpTg7N6zqcwk
lUGEorTrWPB8aMeMxLR/E55U3h9sb7dGa4UV7xU2MAv9oJnz58qKEF85nutg1KT/
ip2b6EunKwaEdOqxBYD44ERB3000HcviV/Cn2doD6p1mfOSS8byb1PxllEoqTVc4
rqEZt901wdtygCcQ3ZgIQ4KwEk7cDKzhBF+UV9qbypfEcwuNzYuBEkQCVfTYF0FY
l2Jv4CaKPdTNi1t4fHdqIHdyzl7wtkv9tfuWKeOUsPVqkXwm5AeM7IAWW/WkM8RT
iLxtqFeEOWWl4UHhQSk4Ixo+3VGsrXVjLyYCVP2LLexoo9Gx52OOXHO3E1jHOwbD
nYDlwznSH5t0qx2DNPjCCjqgv7Rum2py+cg0mRS3FKjJ9XXSBBfCunMPJ2TuzLdx
MpzE7yE4B1fx5FnKXJQnnv/XLZPdq9SPZuFENgZ3VcvYj2h1s+rkghWHF9EYwakN
jtiEsxPHE8hwyTi6qv48d0NpFFomkqcpC05ApXpHEL02SXRvfpIRqow+n7Xs3PF5
FesNUdD68yAIx/8oZN/ROI3obfijIBtVKWx0bdy5DNtVS7KyTgT/rDAiJPtVHrXb
mswUWQW4UAytilfmTe/R0/HBxtHs5Uv52/vjFHGN+MLq7cAXhEln4h5lZiv29jX5
dwwtRzNroPwcIitgrBO/SmxCLrXCk3QIZcnBYbm4cukGCi1B57H/RRc0rgmno0vc
0H4viVT8jngaDAydKFceg8+xvCyAD8l12DyHQQeWaJ3xbKArasggnv42q71Efhr7
l3TgRygEuq9bH01ayrjj4O1ZqfXsvPl3TPRmvybAGx7i+k+8X9LYTIfkbp2Azg3q
l9wz5Nz2sifA0zcTBN1s7mdmR7x+vVuRvErtaIFd51rGoXLNhPjdKg6dEDQM8pZW
ySmArakuTfDiE79xkbuB5/Ha6QUFXZ+eL2zq8s7WNjBq5OWHF2G+PzktOR1Z2rvL
QwdrkAEtYuwOwv6sBZm3jBxwNGmNKebKOVRHV+V0xsCtQeUKbWS1NnkjObLi0uxH
YuzB4VIcFyvmaOgVJ3yPFhdK+B7nn6oXKxchfwjFI1qRWFTDUw1X76LXdFFLDYwV
yzbJS8nYmOB33Ycs3vOWpPX23HPh2nLPCGrcYMZZNoo=
//pragma protect end_data_block
//pragma protect digest_block
HKyXCT6W6oQAZ6hwn/xn7ma69h8=
//pragma protect end_digest_block
//pragma protect end_protected

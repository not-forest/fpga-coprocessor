��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���X��f;��on�# ���5"0 �T�PL7T�0����Ǿ*�Յ�'x���!�����*��w���0`>���M�I��M���M�At�YY?��w�/��
��D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F��5�(��^��Ěכ_�fK[��Q�AU[�MQ���;�g0t��=#b�ػ���p"�t��M�5�49y��Ѣ�N*�A|.BǑ��mad!	m�@ք�e����4�ww�T䙃@��n���AT�_��ߛ<�4z�)�[\0���h|{��=�%�-xl.C=m�C6�5�'�ڣ�;��4m������7��SEPd��a����~�I���(�~�t��]�N�u�Jeh���W�roj0g'���p�k#�#�����ҏ���GA�+�Ы�m����^iWJ]:]��f��B���Or��m!͏OR�*��(�h���nŐK�����;��)<#PO�G�
%�ʚ˫�su�~��RY���Ӫ���=�5G�d.��\֎,aT�F-o��:;��~�:����Q���t��1�V���ab�:/�4��"a&kޏB�|1���r�5�l� @A��p�g�Y�1j�|B�X%���E�k��<z7)����бie�T�D������HL'IF�QM�!*U^�Mb�;t�)��ŭE�;Qӂ�j+j� �*��V��&�<��n�H�ѭ,6#PwQ��]�9���	�j�R ��f9Pգ�pj��6���@2�0E1��|Yڬ7��
	�6sLt�G5�+u���k��#2AE�
�7)}K�>�B�쿹���d-��2i܋��z=GaL�]��㧁�G%�D�x$�6AT6V����"蹑+N�����`�_i7�:k���	��W��@(K������v-f����BVfD���O�=G���z���F�����~�	��Z�#�+������������tv9�4x�:���LXQ%tW�0%����3�k�V��/�,�ŝܵ'陘0�G�tt�a����5K�� �������O���[�Mm�:3�=��)�9�q6�(�����R��g�\D���H���ޞ��}��h����r=^�\&p<�I��dZ��ݲ�a�S�M��W����wO��r�oi�=�I��*.X��L��ۓ��G�
HO;7�1{g���2w���HXƼ�����晛s���
y36xh��S��x��k.�������0n�DԤ�J�K�q�L�^�֔���@c�&�� 4]?J�|��"���Sd�2I��<;Z�9ɛ<@dn�����@L���ǯ�u�+�׉n�ּ������u��M��?]�j�p.:�\�я���z������Y��~�ca�\YZ	F�U>D��$`y�ጉ���#�0ĮR�0$F�UA~'��3�k�ܡ�EL���k��{��>m*�ǿ"Ô#P�u��A;W��tV���(&���O��Z��k����rG(��Ce���s<�x/<�oe��kQ(��=aʄ�<���2k-�'�"��gx��Lp�{��&��=�5��Ъ�l�f1�Qi��~t������}��ű&��N�ÇLc�eqB���k���u�M��`T>��h��G�Z_�梚����_M���j�J�a��̓Xq�9��b���H�)u�8YK�^H��c�%��('��:k�k�I}�������/e8	��o]
��@Ԟ�ZF��=�O�V9c
�ݖ��S�������G^���M�J�W�%X��������O�-S�l-C�քQ�_�eơ	
�+E	&$��?0qd�|�+�o�{�yJ��C|�� )�lr>����b]���v�ϊ�J���������L2#M��u��EZ���޽'Pҥ2K.���Ќ�\��D�\q5�)���{�z.hm�ÞT��!_�w*{�ؘf�9b]���ʄ�1Z�s�*�?��m�طx�&��7��n���۶�m��ߢ�c
��}���5�.�<-�
��z��ȼ�a{�h�=���N
?4Ƥ�?��ٖ�����~���������}7��(���p�${@IS�mN��H�0�S��K�*3�V��EDE%[񽷗�����@��:R0��:lϥ�gU���P?�0?�&��ʌ�g�v�� �2WǤ2��c�S��r���!��H����)�	���[�Y���ZҁL���
Y�����M�4���E���#��s���(��?1j���ӣ�0-�A���?�V�$vE��Ę�5��
�R��ЎB���f*�0O�0�Z綣z��� Y���������rB�8y��l�j^X�=���O�NA�YbF潅qd�@�9�II�nS���Q�1);�fk.Ԍ�W2�������n��)�ޥ,�p�J��,�UᏑ!m��=��&������K���^/䀊�ų�s,���$7�������
j� 5	�X�:e�CB�-��ue���+���� ���n��L�;'��p͉i�k���ӻ�z�&���mtT�<�2t�,��!^�+V�P�Df����%٧����l]I�P������l��b(�ԃ��DDS��?-�^��ǯ�2} a�h8?3�R�B�5�PA�n�_����f�k+-�\�*W�zn��:�i�[uiVy�����xݱ^.�z��Y;��eY�z�{71�r:��@��M%ԍC/�+`/�:G?���-�a� �t�i|� ������>�c���f9 ��Nf�*X�E6�v)i�H�k=�Up�B��c ���3��˕�=S/
��!��m~� �7Ų�t��M�&5��������Ddk�S�ۜbN�*T#f�) 	���y���!t�nS�?���ca��
2��b9��@W�UX�I��w%{�?��`7�Äl�l�H�j���Jo���
��EAӂ�K� ��4m�v����孧�:a�km�h4��s��6ݯؔ� Ȟr�򒺕����$0���ڝ�&���P�Pj�6��l����Wk4�B� ��R�縇!`��[%l,$.�<�7_u��F lJ�������D���ɝ���cNf��stEM����Kg7��AיW���'ӻ��A��������d��|�s �2J3���z�����Wr5���C���V���!� �.��mUh[�뽏�d(�Ӿ�5E`d[h�;*��f�ϱG�A����~N�q\��	
~4�lp��J��Q�_�X%�����)D��vP'M�e����R�oo-��X�ѽ(q.q�;� 68WB)��dEd��Rt#-�a�a��<}�yh�t�����yD�#���B@3.�'	`�����Ԍ����r�f�����q,_E%�H�T���eĭ�Q
:j
N��� Qv�x�L�uG��;r�Ғ|e��){%��U���p��j��fL�6��㇑�Q����}PT�vJ�^>K7	3U�/��"K͇g�X��aQ,)(w'��\�\j����a����~���Vb>�*Jw.F��>����f��m�	�+O�(���Ĩ�ΕmM�6$&�; ���Ʃ�1V�)׽x��D�Fks��3E�f~��,mTAi	���@Oº}c��=�P���Զ��CZ^c~wd�ͪ�p���]�nx�+��Ry\7�/�m�=�Qh(���e�d�Xh�,�@�W�	{�,�AN�����!#!m���vml�Z�e?��K��N�w�\v�m��	���6U��/�@H�5��mᕧ}[9
��+���@�xL�J^�^�ΰĉ��ߚ}Nq���(��n�Ď�q���㣕��uQn��o��o���	�7Ü�]����ld�������i���rF+�55�|��E`��?��B$.<����p}J��;ۿ0��|���s��4t���K�Y*���Z,ƅG���^g��_kCg�t_��l���Iʕ��6c^���c9yn��.l��;�._?5?v��>=�83}�r�����|ׯ��QÓ{<rƲ���v��E��[Q�����9!i��~����Ɂ�D�J�� ]�6���_�̷g�����l����ZE_-��NFJy��Gd�:!R;:��?��V�aj���Y}��o�Ю���-�==Ð�'\h��T����W$�	=|��J���y�$�� P�Ҵ��u��q՛��㴇Q�{/wU������ё	C<Kx+X��N�`�@�sq_٧���˫'��n�>��d��X��3���)���B��"��N����LV�&i,l�q_���Ur{�ll$Ko���B�I��;�"2�W�B-�PSX��4��?�i^v'����m��Ʌ���E�>	�>r�V��^B�>��'G����9`'q*	a���Ĝ�գw�n��}2U-�)����ƴj���P]�� 2;��E�e�4��WWXS��@�!d�I�nV_��*�g�2�*P���KH?�N��V��)�`�_�GơA���y��2%�͈����~�{?)��$	�������e�E��7Sj�8邾�v�7X�-2[Ձ�kr4qm;5T}�EkB��L�Cw!$��?G�3���	�Y��A��
��f��y�L���<�Fy��,�A
ؿ��Q/�ދP�zj�vT"��jEʰ���R�O7 $���/���|��TF�H���!zqi�J�bRk�
����
�i[�G��$��J�������<1���Vǵ�� )b�0��DQ�� �}:e�����
c����F��O=O��sx��/����j�S�	c�.���ĵ!�;��dB�/����O;��Ϛ�����٠�D�������-NZ#������.ψ؋�yt� fDZ<a{�;�^��Ѡ~��Q�X%�ǥ$�z��YQ��r ��N���2�8*��҃���X'����0�`��>�u�~�Fqo[���1WܵD�H�� ��&%����G������o6�`�z�߲)C;G 6?�s��0�JԵLн���ɣ&|&��4�	���a��f2�5X������`��CzH��"�Y�Ӑ2-��A�Q�zߗ?��?4Qu�M��xQ1��mFy�P5�D:V|n�_�Pdt�E���!?mOԄ��฻~R�j���ֆ���Y� ��n�z3ylkZ�$\�yw_�$6���ܟ���7���m�_cp�g]c��d ���_@�4m�TuG?"�P]����'�-0媏��pT s�b��0�B�2��}p�?9M)e�(_b��fD�e��9Ғ��<j�wO�$��O�r�S�6��
4���\g
��nw﹉;�Ο��Ճ:���T���叕gӜ�*����� ��d-�� �LH���zɪ0�����箿�b�p��n��r[n�\�E�c���-k�'/���66�AN,��~i�7�+�!�
{����#
// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
mWekvgsllPFOQKrpSCMpMGCxLlbEV1sd5bej/UgvEv/5nZbSK1bRrqEzlXSt66XF
P6DjZETlRu80mLN/h1ffhYBoHrh8hdG7gsuwCmRqjxipNYqxbA9dOxgSp3wWBrNB
ItRT4IPAqvBJWdgvDjkB31y1tie039JTsP1n9iDw+TSCy8wb4U4N+5WBKjwZfdvv
S1K3WBuFCW1qdPS3m7+BttsPF70o1PlOnaWHy+10eCjQBQLrLsL6xYbHldQNrPvy
MFoGOJNrWN3r+k0gQBW3vRXUXt/jAVe7CNbgjsXg12tT3M1GMXOUWH1AHJciZZRz
eJVfzhyIlTXA2LI3gCSpFg==
//pragma protect end_key_block
//pragma protect digest_block
qgxe2/713GT0EGIoYo2aarIQljc=
//pragma protect end_digest_block
//pragma protect data_block
ry9Tm25fPRbvX4rVOnz3vKxS8YTvlNZDxG+0hs3WyL1JvXJvfloxm/ePmsfaUr2/
kSqG9mliadHC4DbolTx1YZHDKVrD45z9nN1v/dU44mzky8aXonqvEWI7o2uwKY0T
RHhIRLZvPwOld/sDVKItMCPTm8LfYOi/PMoke/vDOH1XgHlubAByJ8Xdmb1zmKat
aSg7yR0fMQwUvmIhADqCtEZ2WivUbOsa02G2+aVuzYUS0lKTgehDvFCJYq4jnEe/
/3KHetEYCvz3EXH3JlJDBiVDfFkqmgsAERfwRzt8KWN7hekcfNVzE4GJeG58vqhE
Grr4e6+CgQabGEM+oiXI+1BejkDJ16AJMNiDCzJIXySnCu/MFmubx8bEIR2A+U3e
nd9zTsJTXgQzEvm+9TEL3f26memIXcHSNCez4BbxVHPB+/e0/cKkmTQXwWxUi/60
0xledzDhQRvzKytY5dtl9bZ+3AMeNC8cIpg0sqcYuvHK1GCcxBmvPNu81gJI2WRa
3hgR9qiWbETKOqih0NBTxDpX9slUsVhdyc/659xe037tdZRC1zp1qFDPOwCcIylV
1mAHQ6aZGbgaVUCb6AJxz5hNnOu0R/W3Q6/PUIAKKGBMCUErQFwVZByrIteRF3SN
f08zgno/roeumAxPrr0c+lVg9FcUdcxdlWENx8LmoZbN35ztc/8TZCU3nEWlpPtk
AOFkxY8CxX8gZVQSdHKNOFc8S1FkEblsfeKF/gFWEHulHgPK7z1LVBi9vvrKkkQz
ByjH0cXJiudY5OxlLq+Bu7eufoBYfyBX/++suWBBkpFz5jdg3Tnl2B7e5dGMb+QC
UjSiujEeirdoZnKeZiV2gxXacU0DHAGS/sZ12V1Yw/u0SnAJ6koej7NPvi2G07C9
LqHnDyQuCcYkDGcadfvyhMs7I3SMzd2LBc7IRrUilpvz+SltPxKfWLGTjzDaqjF1
6mW0n+29G/5c7Xa0R8dGphH21ix9OgMdXiPzHBQi3xHZAAjCaFxsco7EqRcBVKM/
7vDM7X/lPqg4DW3gEhrIKph368+C2HelZ7Tb+D3Or449Ry401GW4a2X5qvoZS5b7
l21hjSHyADZ5zz6bHXzpJlTL1Ck4V1URBEDEBvy0pOwzFp0JIp9AcJfG9kN4LtzD
Rk+dNMAmK5jPWLFevNy/Ddb5pU44GtJ+GW/+gYN1ABOShNO+djz/sheFWLv3E/To
YfDFNluZHkClZcSrzw/E0ZGbZ3118BIBr+poObpAO4NMrWkGmH6jLn36C5yJZhOs
5lx3Fjo9TxnUeAAEcf6jVe57GrXM7k16sMgG/fflmJXo5xTDeoTMMClbbltL164g
jAl012I5FEqcx12vWC7UgT4QzKxKKFv4A0SeTHkCR/z/hGn5SDK1t2YxlBfMM50v
tj5padSXSDBRGafc6nhLrCks2K8MGcGoDbBuykgkHsjDKPFskmgkjQedyGbAVBLq
ZK0jrgxku1uC2HBKzYbohTd5mlO2dS2eiuXfF+rseQ5IP8WRH9ZN6dgNgnuiaoFM
owTI9EDmr6yv2sR5/tLfndwNt67TM0wZcdoQ0wugPcDa/n5vQHjEEOuIafts9opr
yr9vupIV30tXKOQgJHBvD62s68VDMs7uIt5cB/WXs9a5KvpzLLBMPDO8iGxPdFSd
wn1l1/dA0WV3rw6vuxp8p1begn+G8/KFdLLZCi+WKeZx7R+FEGJotVaVhD22X/5Y
zEEQsU09BIxPM/X5PL989PYwCodlt+XNYaUDphqbJvoU4AAhOf6TBqMNTl8wD6JV
yGlG6nOmwvABQ8cfMhnt/JNl0OAEL3SkqN5/gJlH8Xoq7W49Us2tJ2LcElU8AO1X
yLD8gSC05i/weJISVZnCPziyikyNYwAx+24SBz+GKro+SgiJNqWPGMyyZ9j+jauO
pEe5gtsASZJhQj2KLucFAWVj/CehPqs0FqN28XL4jt+kqEZWt1Qlwqk6NMlXiabk
FmGDxnP5JW31ZrdYsG/ekGZRse44d9I2buNOc9PLolqph6MzI1zo2kkMFlhXgNir
HF93aVOpYdK9tHwvPM8W5DedxbBTbNrav1Maz1BXl967+FeNnudOhmcb4JTPH++k
3SkZHUl9TbihExxU22E952Sq5W6aBAzaN8StepXHrCiDv5ygWSEklVM0v6nPaKhF
pi6YfanBbifcMxAgahB6esaT/TgLFDdkhok5dRWg6PJEAiL1zvgWpf+qp4k1uDc7
zAUt/+plZAR3UbWCPX+4I+HhVKNK54loxkhi/4qHZSEuV/uL6nX0gAm9jYrOn5S6
+xFMwcjo3wuwgqeQShA9yVQZ7IS4a3/v4MVbfoxhmKjeN53YyGtcewAqIZsEjKlB
VdzMbuK3NTesYDBUpQHK1+w/pD7Qzc6m1uB/VePbX+sSeSAKmGT7V0huCxpgu9kp
IwSidBdMfGhS+GoYMnR9jtzZrZcIdn/Uz5kA7ZciaIufKd+Y32tkOyWVtJPaSDf1
+xotnNr/bYZKJKhAOUxW7RmH5gK8/yUMhqVLopx598RlmAfd3mLr4y2RFe5oz3CL
llLb0FVbhHcNqy45g9vpRtBmpDn/HEL6J1qE9PhS8MH71T7rEt7dkvLr0ifatSvy
mjL+uXKIVUhSjyW084TstRvmryIQX9JzUu1pFpSoApcX1g7mPJ7MDoZLleVTYSyn
XL2HCsXQmjbL34lBkHbzG51xR1I7W20L3dLY9LZU5oxh7R4MIPRUP5eHPBWgHhN/
zfG7Hr3t1if0R4KTezfk12RDdHti6UofwWsP6PZeCbWiPGq63wkqWD/bvUCELMtK
UAPgFUHHe/4IPsGQzKT3gX+lq9d5yc/pj88nCvq+F/LOuvuTSyBwQd5sNEjbFAj2
1FQdrl6/9172Sg7vq0wduDLCsRjv70iBElR4Ekz+V6ePNV8//gykn0ivZ4LEsT40
xPZn0jYQZ+yVDtbxV/jxCG9/ljM398fYI9ZTMzfUUsxusGSTae/2mD1pSNk+Ix6b
9I4e4y590vr00XCq7gRfMI4YA/elmj+WX5qxXy++QM+IPXqJKI5emEzYjp6mE0Rv
QZbnpOg3nADVPxTcPY71c9GFrCPuHGgtR30BbUa12YIeHRfOyOkMyCPy/R5t+ZCu
n2Z9zTAcIHTwDyJ64U+ctKbX4VAuuP4sOQLABRyr8icZbg4oXN6ZJWbUmxKq6WZP
aPQWkU/BkGZszP7A4TEsy5OranShNxI0TCwK5ludQJgePhGipojNY7L93z6fPRQD
yuNoiv0Dkppu/YZ1hSWIFZxCrFEfMg9gYYKOTujUkgb6eKMQ+GDy/tWW/ZGFu4pt
l6KYIg8SMJmLYZlkVH9gwCK+e5TSqRmmwly/gipVbHFkCvn5Yv8rCAKB0LGhc7Eb
oaC0g1ymclG2dPUJAvjr0v4j5zcwVtus24TdPQEvb3qjIqBRXZmgysdbKpvTaDXO
6piMP6/TtZ0ymhwCgWUMo/IPDAPMSwNkfVYHtgYNVEZJ58c1tnNkZaYnKyH+raTv
2Dl/qFyXG8UwxiIrNifl1AlZCLdCjYh4ZGMDblHsYcXq6+H8t3wDPSHHUGCyU1ca
SvIBx+jN3hw0fy533/fQuZgFDtcevJw5C9WGBKkU2d+HnpklFQFgVYywPatEBXlx
GaiWs6xFCmLprYF4JdLnPsCbIYOe5FgYMHfwvtFSt77TuQlaEa3M/dRfYnxCvCSy
g5R3wZxopU+56TttlCGuI5KNBpJ3gkgrCVH9xaV8EwN5sj7uP/76zTRq7x1me/sJ
Xxm20n/G2z5D1KziMnmQ2FXBWW0KNsImpnV3VwkZQ8/RIJ/zFh7QL2edgeaovrMB
ABzIa42Jflq7zNkl5F39QV8uKk/3DvwmNHi7p/ECpYICHt7rdgWQ9lv1/ZLnZqT6
85DsC2mJCAO2r8NLaRWpwXuwz/4rzTXR/MEuM5kEo4eb95kLnIQQUUL6g0OpcJzm
QIXmASMyg4DJaWETqHIFu2oOV1+z92uOK9s95QnkEqFMnWPWRN8mgqkeqpkorGux
aOSGoBjdMwX4XOsMli12sG1onBzoV7gLievrs1llWfO6jUw9TrvUOwjqamkQLl5V
u5TzgF47p+rAuQ/HFo3DKAhghubb0iZsQW7/jCTO+u0+XZ4jyJlXIWrz8Yk2fCWC
SorPmwnDFbP08NkF8+TgXuTu+Ii0/SBFvspNN3B7v//uJxGk9mayiFXrKn7ch+vN
T6jbaSfDyXd8N0SxDis/9UBYLh7C6gqDncn1yEe0A8UZXbKJlQJUEOaEHGrtwCIb
lhfmtHuMzeart3zI1PBisQ3F1mNURP06ZxpA6gzR0HwH3QRtatgZrCUyNTdh5Iu/
9hSh5/N75NkOPyA/RtLErAVFnpljpCynvviwN+1rTqbCRIw0f9RUEsKviKhLoaNX
EqpZ3E/lV7fP8t4MX5NKc8VHJf4JogiG/wgYiVyILOtm5hNomGJAyApDS08KlKF0
Gr4aXpB0Xj/c7Le7fizIqPkMPxNQ4rpploJo1erza2RO+0AJy3ILmADsiRZxDclu
kHZaWxQCZKkWXtCrgViHAxvXJKhT7nWBj+K7RrYd2i0GKYV2gc47LJKy/3IsYpxY
bJRwssK4uefJkCxNM2YeB7DPQsr1SlUH9PwOgj7+8fOedTihO82AU/mwR9Dk7bgC
JhRChrGZZM29XxJ+CyL0AG/moT0N435t+s8qTJa0fR5jVmXotfnHm59q76DN075e
qwVrI5PMOouJa9mjhxiro6dLRzwHxqyYEdJOW/clZ60lpG5rI4PznOcTeAy63r04
66Lbh+a9ro1nXyNWVfQj2Y6ETBvuS/w3s8tSHeJCzxhHvayxdkNwuTPEia+SWRCA
pUZlCW6dGQiSe2mhvC1MrC6ZLE9KxPlXaRUFSAoY/WtYEqQ6PHvj9x5a61H9FQhM
8C1v3EN1kPLyUsPVlwFb1m/U0qiIAmyd23zgwDSOHVkZGVdHH5JnzbrMj0nMv3sz
WOiZbf8ot+sAZoNj5JjWLbbd8DfPrcRW6h/eWCh7IZJyqloVtOt6XwMThOAQDNJB
HLHBtDTwT8sU7lAGoOtHjXQz6BtvkXLOC+QHM0mPN/njO4AO4rU5pnn+NodPhoMd
kLbbiA86lAuaWmA3n/08czH6FoJvg1TTJ1TzjBEQwp8QX/PlGfGkC4GQcfolYgzO
mYAMNB5d4HQ5fIpk7AbtPeFaOfdPK/9tR77Wq5iugmOcnGYDSo2RNPBwLL77rPyR
IsB/YO5E57Ld8ivycUnR5qNqYctDUqUCNrgVUEMlwHy33QhEo/+uqC5MBIGpv5lB
RgyCyBrPygCxTamFsZdujvCkw7j9stkHb6tjdsHJdosITbFI1yXKbf/mGyw8R+LO
l5p8D83Ng6awzewrEE4JG5rwSzG7klaUJwVH7imIK0VDfLw1yVujFAaApj0sx/3n
hkCM3OloIOt9W+tfiow3HZimaWVzhEvh/uazl12US5+jH4mjzL63yhE+160qkCZI
5+CmuKHmNZFt3f6Ksprmkh/tLz4XcAUdJAasoriIUXB3Hv+M8uGmuCs2S9tgzsx3
4KUBTZMqh1xV59vXoZNdZgH4LWbaz019ml18Ykp8krrMQfwCyQ2UzwxvB0E44Ers
pzNqfYIu63Cuh0emdcCPtJbGyZs0a1Qj+NSD+2PreRBxsoB2dOYA3ln/uDg52mhJ
2eth2EiN4A/Hl73WETpAZkAAobfZ3BQwfz8d7TeJXQGjU4ufdiA84DROtm/Aio5J
7cL55x3k3veHL/48OZwMsE8kgdg3IJ1sWvH1CwW9pjiBR9AIvL6W2z3lqxwQRiMa
QEo12fhYoIesb6UTaXOU290DXnfk52pcR21v1R2WzIuAZGIaBMk/OFhQ4v3ymGD4
XppwEpmjq/d7wvYRqKgFwdOW5jU9P9r8ekPUG8NUq8RVkAhUD+Qb1rLhXF7RsYSU
gvXx4Sxou78VlYpMV2kpn6zxjq4wG5Co40fF1IlZ2/k/bGWzUL7toyh/v2wqkgYW
CGdCLVYFJiDrbOsupQHlocYMfmphw9RqVHCeXOsRk4sVRgJc1FpgUH73YkOFP5NL
AwWj/dWWZuQUayfT6iL9KEdz+ejFunpMrctaZBs/Xq1Wi3bFBKuJtUKvsCv54U00
45cpsJxHFanfjwbaQa+rNp2jSceApHuVdBiLcWW0uKMz1Nql0kmK3Alm85LECMO0
4Ss3WmwF+Xd2636DKi5GL3ZswMgCX/y8hHNyyCgVLZfYB3RRv0lmtCR/gW98VR7z
YmUTC1t+98urnfT0qLSf6ugWsxtFho8MzrXZ15v6CojVh2ZgdSyjfYWXAnXzoSqP
2pUgzrqNGK0SLcc9ROCYCIlNYLmjRRb0/G+R7fdKk8y0G41Eum/1siK48prFD/QK
WQb8paQHl73VCz5E1WhhFRAjvFO1PQNWvtjRBNDkR0bYxPzgCA4sxBkaD60np84q
cwhsB8OSHOTh9EEypP+yoKYljZekVXH2lx1CW/OgOs6tqRdf+0lw1ENpX6dd8blD
CbohvcSNHbdo+p09wad3W6hJpU7OeFCkVp+fj6Y7hQzZQcUOMPDIfWIEFQ8wjDh1
B4U569Nl7tQvwwkFPFQSxcXnbM+hhr7U3eio80j2zsTI31Dh7f+6z4XhYxEDcTw4
H11OnZkWXof7efVdlIBH8GygtpdMy4wKE1ov6ffZqnlDxph5EHh3DS/At98Lat4e
PW6qkkuxGv4e8B8CrxcheobGX4rtGGQ/c7/MnBjH6jB9A93iqM7gvZEm1ywOR+Pw
710LSGqxcNNAAGEC4xf6n9n9Q1q8ogaN3fJuLPxvzGfy9r+PmQI0J3aMYU9E+cMh
eIRoHGzIzPR2jOApvBmmAlYf3XS+FXrxw7DMCV3+SDciEnrzAR97esOGIofNJGO1
ZNpNNaILAS/gdnHPiiCUfmLFUshwxJ4Hwj7u/vEvR4lJPA2oFWYwytdEtAcuchf3
DqbF9f5WY+x2RHidSGlVQ4RK66WJlkR0Go9s3AJL8o9iwp2vs6ZfqJUu+W9wN5+v
uULjd9KLdDIaAeEjmlYsbiuVl+qBJrOdjGMPYx0X+bLBH31+MSf1NmUL3IgP/t0y
G0sm6aZgBnTjdCAJdhBBtHIKnsaZYa/thcWcm5d6+mO1qAiQ9tldkzI7lNA8c+zY
4p72GIs5QEHjXnMJ2z4aTCbIhRquCMxTRUWdCkfLjXGl0UtaAAlN6aFlrFAPS58L
MMDI2PY/5bPsk8+NV8VGTegCN4iRt+wfbcoP9TFw34wg8/byVi7Q3Ti04k8Ij7pi
MzuDLOshrLlCs9SBqB5jVR5GjKSAS5C+y4pxcMP1iLMGSvvYPhdRqo8bpTr0hERa
nVWUoGodbtTzTQSzTQZCxJsOFYmAuYE4RuoDldiwZ9qh9+PyYBAx9qKitE3/DaCl
OSj9UYCo6M5q4Y/1BjD7HYlSKYbMqvIjMECXvxGdGolJPwiUomW87sHkCBoEgwyH
RfgrFDsXX4mZhyxNraiC8q5H3pc2cSqanlO3kX+PZYlerd7WYZdHKHNFtvclBhHw
cf0hPdH8wX/IF/gB0QjsBekf5KpiKYJj+NyPNN7vs/m0LC0npEwEuS0eS/OPPX5L
yEtp9dG7UbEMvy1C6zBPEU5nrwSiW71ozUvDq5kV+Bda6x6on+1EJ4FFmwyzxnjC
pao782x1zD+VGD3ngLjKtR6eaZycJfqFwU92OPgIpiyNcwNA4du28k0lkVFct/lz
OPGwTKxA7PLofxpcjl2J++pUamOb62QEG6303TDYSpr8v1eMSAP4gciBegVmzzN4
YpVxPnJmX7SONHNwXXDuf3vKmpBSFLT723XGofZLXMub6kdlTorBiG2T2meMynQ1
/pS4DN/NjqKWDcb+y5zxUCnkLePHEWL7tvHzYLKE2UWQQU1A3g9bqLKttInrPjY4
6r6tTOJXw15tNHSypBHmo4D8u5TAwZRSepFrUxXtypMyKrzcDiJ3BEXjrO6M8tFw
o2GUMYfjrr3K7BdV7TlxlB3RxRwdLCgp8SLnP+DeiYNiWMwGx09AYz+b1CqlA44h
bVGAnnapYCgkC0zR7Fdcvlp/dcZGnP7wsEIe6IcpQBSq2wnl7dHTgkR3dq35kpWu
121MIENGyc0MYp97QPiONVFWFgUvh1Dk73SIyKG2oGjTnped01N1wGDJ708cMlZG
yOFY3kka7h7ubhnFy/akpIw7ey2rtkFgsUIxbeMny2oU97GhkjCrHCjU+Laf0RNu
lEAQFWsdon2ti/lpd5u3Al4pQa9TJlYTGuwxFzFR2FeuKAv6VUdJm5a8lAVZ9Cvl
u/Hq0SN31lIJ1eCfXPD/kHaF9zpEz1XxBXg9Zm/uLpBQABLuU8f8RIlCcH5VHlLV
jv2r1jXqqD/DoxL7GCn97kCSKpFPIHXsUFNhuATtgd5/8FqCxHLm0TXk6QIFF6jl
9eaOVkp3gcuB/M7pbzLcUVwNwtn+rZT0TWVy0Qf/YVAluMsTHA0IWafMJO//NBqj
pfu0FPku4wOvV/GFL6LIAnOZMDfOQYBPJZDJevIn1nKARZxOq6wWh6Co71wmFOZa
BF9lxHDsEcgZ8dg1Rf721lRrIPejUC6kmZUmyAfXzruNK8/NLMfGjFAjSKAq98D3
9QemQ3qsUey+G9vL1bfnSvfWNS/LAk8Bp31W6lF8RNfDcN4wXlmMqNtHKKurQeyJ
cxI8FHcHWiOSj67xDu4p6n1f4+XayqUZ7N4Dx+D16VdcWeuyLCxy2qvIt+pi19BZ
qUnbBjqvDIss/9PBXWJxrppDcM6lOWzOn2kW102zyByKGTtB/lSJ0rUvMUdABAuW
q3k/sWIedROwlW4lFcnxhksBszgqExi9azGF3+Fk+aBx7wFSvZgse6iTcZ9vwBr2
npkhwVWpM5ClA0+mnrdA+CejUvKMcCnbHSYrMxc4lj7Ydxh2iuTa96N3oq0HJX5U
PLzJsqvr33apTdBTkkIkuzARITcSJKaxthehceci8xDmDNdjEbU+JONCzRTXAVe0
yfXOvxgjyJEmPSW+nlvyTHAJEDFVVTOWfEW2EU8poydzpKNqP5EtoqWAj/p8edzS
PLJz7WBVJBCTwmXwLh3OO4qzPc2GYcFre2nkeP1L1R9HSku11AqflQRLPgjy4TB/
JNatRwO8KTqHNsdW8UzQmUHl1jveh3Z9iw/lTRTY8t9Zfzbq1btLUactU1+IQWDq
Hn8Yc7DqFr1ENA1xhLkKzrtIhDDLvfGwE15uWLWojRV5AVoYMOJNIu6dwKxkAp/c
j1JJiQU5nL5mKx45Y4ey9DnaDzISDKE0FIOV4EvBcZwTp+Nmw5/zoT3IObMEHzE/
ptkvhi30kMODnHyIr8E81udR8D0+xwpO7ZMRhppNQOYONh3fHgUHnhZFk2Ng4reE
i/EFP3hwrHQH50b181vEDfAD1qfcqohMQ4KF781bK1osGDQB37E8KKbQHFBy9+na
BhrJ5azcvgSNuLi4YDpRchGC0RAF3cdSh4br4HkzSOreoZalsKxv+H3rEUex9RZV
Z5nlXhjFSh4MJnBpTVib48AJmKzg+TW1VMUbR+pM9OFePIvRXqSN6GU/OWaMj9qf
HNAd+ljHAGoVGojc7QEiM2vg9nTZ7bOOj6VTGEqDWPmR93NEJcGtDG0vxhFsKgt7
JoxThitVryDQhtxfePxpHDozwKG/2o9dQiK340KV2uU+7HeM758LAFt9LdCz12YW
dO9szt2AgvTgfT3RsM1hZW4WIbECU/IOw7CwZb35X/4TbrPNkGvj5o7X8cySDg5E
uh6Bww8fdwJUFCgbZB+LeXVQGfl3nqaSWGevWjc4AL+cUCA/WAkQBOcQ36XKjYV0
dQw7mIq2CEQ31fK3t3xKYcxemO/0nJHq9rnWU2xRmj1bnBt7IyKmyiRfNqQdraDH
V8f8q/1tZgFwr3xsayTJ42R3o+ZcxK31OeShPtm42ECsU5AgdR44IauoUEsaiXO3
ENA1Za5AzmAS1Xwol+Mh/cgJ6C0Z41fBHDWmFWxoKzGIOhqyeOwV83fPtzOoUvZf
cAAgSE/glOJQx3rk1RqFW8XxjAqoKyPbGE0ZXe0VkiurJS67qNtP2HjD7hW8FVfn
gXPcBigjacpOmBsLRP8A8lDsGTl+pCMkmckF3kYS9ExbbuKaMvShBm7LOq63029P
KEJdCDIijZV+kui1dErX5C5sr0UMFG5P1OPmF8JB0mz3oKHYwCPRntDqWKjG96J/
3xmQEsihR4dRcUlPoXlI1zqjkt+++z/9OvGgNZyeyloc1LLT8UeoprE3SD/NjYH2
nQKiSA2JG8P9NofYjSlRplqHLLsvAF+ueFKpwbBPnELM7RARmzEJP1oZOiT+wzP9
u6aDOBhP/lcFXvMDKRN/pXsbXpwHbLnbib3vUSrnSfauiSCRd2V6wVMkgAwI/TXQ
xqejX1UzTh0VHbl50Dp21XGhr6S2kbPPc3rTqG9gFq2Fn+Z3cfWzmgoSVu9OpuY3
N/EYRt+DeUR2BKNRr1vn+xtudTTsTFNFpDf+jDdxH92VM3S2Yz3+2n29I7KlH0KS
o8rPejXQVYgdM1wR4Q2Dsb1v912O/lvK/akzQAS6Ssfk21+hiDYwXQvbOMvI7Bkm
Uo20S1KEb4rNoaphoiyISRG4JNac+gcEcvudSPpHg2jV9eF/Rl/aoxy6M8Q3Ddv0
RrUCOLazbYCLP/bFZFFcIxo3RNwwzEyJimf3aKB3rLAh51yTBh9ZZJwjlDDFiBIx
WqMTU6dV6fHZB6go4V+wfrwUZgHnnMwHk8p4q0NoRKhq7csUqGw/Gj/4icbuc9YY
93EDw0PZOgh9Mo1iF91i35Q95WmpbRZ6gzauAXKiMDPkuCoHG+kGgMj9lizGHFyO
0i53DlKld5MOkpZH7cVRAUJrN2T/2RwjIwCinDoC0Yz7ON9h3POuYMuFADbX+qZq
Bh6h3kHuwrp2Rk70bOqRsj+qU4Z5Egofvr0KWfQKLp2kXUSzlGfz0zfwJMiprKih
5hGMLemTQuavGpfhDa3TrpqZd3N4iAxrdHO6pAabB90acpnZ6OPnhNVjkyXOTb5u
MuiS3ddbWb9w4vu2vCJ/Ej4Rj2umCVxF+hpfLDfZIYMV8uWRW4Fwb0IdpMhNE1ab
n9yBFjPB208KhhKXCZrxhs+1bYFdAmoQpb2saFKbaRw/maBgt4njBWenCBH3PlHn
+pd7B/lD1+BxHGlnxtsyuhM1sRwqYXbtWgHNvFsl4BEdZtV3VEAj95Y7+pGNPEac
aZ+146e4Tfsn9T1ADJVZwEspjAz1qtFqlM6FFU16Or4dDbN5nlmJhgnElxaUzNVu
WQWNkZOLxwskI/oI1Fs6luaq7nhj0XGCC4ZAY+ODvVoRj2+OuBEzmN7av5VmVPOr
UAsS3143EwCTU5Y+mRp86XaS/k0UyUkD1d60W/Pkyhc/8/SLiJh3Wh3NfwYFksK5
hIpzmzjjY+iioL19d0DEf+L+4s4gS2mbuei+8ENHkP1od5tZdx1+6W+TjP+lBGmd
TdK9I3lHd/LrTHnpZg+omFxAOISIwgSiwoAP1ONctizuNBUImWrQ+N8e7Mky5Qpu
KTUXNkXqb0wBTjrhrQE5MAdzVmTozw/9LlJGiUT9YXcK5ja/Zt2K9GCvvwmNVLw9
shSk0cNsKOWMD7NxMn4yL5GXA1H4Ab7V4KtndDaEJBDNG+uFDwF0Mz81/NVcmfbJ
E6wqoZ4c4mRxv65jlORhDiUcAqmKt+Yq3AF/T6n2iPh2SPPd0Z8h/WoIlr2EJEGC
CoBaY6jhIXWBLwlP7otk35pqQk3fJ5clqbh97/hDBjAvr78H1qNw5WvRzxnzKgx1
WG7h/5UK97lEKdULEqpmHqi8oDHOvpCv+EKNMTqwaSmua+368cyiWYQ76z4O8ONw
vjtQWidKA96TiW3KD8R+2TND7V4YbB9/D3fxG1ANb6+JfYYdG8HgMi9/x5Ssextg
cB8JMTUDgFUZkbae575fJo2dgtmWPRxhlcllE7T+tTUAVnd1FGWb07Rjx4McEYkU
l2NiZ8RZDLH//FgIbFXqXiTtP39zOgnD2Msjvgm6L6hnEJ1Hv5h8X4G43MUW8+lx
mQZijV30G5mGG9LE8hNRJ6WvcY7wgaE0O5tjXf8XpmOR024bvb4dT19O2I+u/fDf
S/1jWcYFylz9bzQVXmRwLWclwgHtKWVVxpVsMksL840ZopT+CrIWxtBCTsjvLLU2
+Y8FSdCMA89poc/BmpRYanfAHZxlT7oQSp2pol2CBnC3qmLgFPuBmToSKfG9XhwV
AmZllF5asbMXhxEvdFtLvq95dxOlG+bhSl85fCsrcyQViPjfBgea8PjQxeDKi9ls
DteOx3bToKb9ofskhWrj2CYR4Q0dKBg2KYsZgY2oJw5VVKO1kVmtAwQ7k/iYeV5j
P/Uxks0Ve6u/5jzbLI/RZKHP4tWMNnoTnDBo+r/7r8gZh7frLbQn6B27gYxgChjC
ct9uNC5wSpHblzh7jlRQKGMBvV8vbzGciQZ9RC6OLi+0qEG0vuZF5xU686CpFD9V
3KZHtklZXEwfMHtkxpQNC7sM5HzZEcA5UyYQE9LhhddZ78Qtd8ieg3YSiL7Z8ipW
G16VXfp3mZjjlXqcXQcIdy/HoGUlOO+cTtu9QKkull892rHwpIsRLGaMtwqRUenE
IehNIX9GmlBNjFGvUzafM4vyouVjL+vPvDOnBxk1LvbzYkpV41n3r1VCmUFOOXZP
4lOtDt2MpprCfP+Yy8d4jsUqp3leucjuJ+E2QPCP66u6iEaTRZ7q6cQ81tAA/em5
P986sskG/d4cvl/3HWhKoaqYjXZrNgz7TATdec9eGL1J3BWcBYCC9kTJYomsBxf5
kRHXUAhsVa0wML8g6bEKKa+wVfi1ewWxm5o6I3/cTVyEBXOHx6aCGCFah8B4MiR5
Bu+A2ALAzEGYU7ohSUVbP6jlJKEJa5HXfJ7YU29/2hjniPY2Wi1WvMvgyPK1BZ6y
AiA9xnb6A9CTZvHAph1WFOlWi0Gc+vJkrIDkqs77xhsnMPMAuGDoz207fKZQnmgg
2eB3GEgt7SulfnF4wuNTQLcEetmQ0Q1j9RVsH4BJZOJLDD/sRp40iSTDzio/v6FS
vj7FsGl8H6K3tQtiOFSW4ysgGBZLnb2Jeh32ugrjjBZB3yLMJvdz+PbDR0POw4ON
vhlEoJgnBqyOq7l9xGrlB3Ls45VyyGrsx5xY50k4Vt3wCWJJc5WUElMfDeFLFhX2
xlxrRIa/hDFXidR1woT8PNq/wDdG4CijksDJZ8lIoyJZwrTicPdmEm4gJdqNfSub
tt2tf/Acm6+Ac9Bcz8MSCl1tTwsNJ2z3S902zn1jNGD6yTv0MfPejO9A/J20Qszo
rQj9EdFz5t7h5ndc+FuE7+BkfpcvW0YCB0DJ+smwJmsSMwbB3ki3bqjYVshOvSK8
YP1l5gJghd7WuklNibmS1LNmIhvTaURnM2GJRg/8c2msrpMe/dUG6lIJy/dJKMUa
GDyouX5k5cBKQWQZ4XrzLnMrc2hP9gyD2DJLkmJKFXu60eZqMP/rL5gy9jn3E+R0
FokSrIG/gqWrPkkZAzNdPThGdRNT1P8d65F6PO67FvdMjdZdD7sI3SgEn5YIxgSr
69oLGeR1c83YeSyHm4KmNu/FKAr0aR+rLIxQdhKh7BHWJdqURka0+WwqiAoqemC6
Hk4RXPSK+W7lqmJMebxwKMmN75BR0zA4wN7AcKlUj7AEOyk19FNCLSDxEIYBg2Uy
snBSSzgzlttIdgIQi9mqd5NTlosARyJM290Y3i0622pL6Z4yqi79gkLlP0X0gjK8
fQz+rF9K/7lDrwDpDfrSFYbrV5fJchTFkMTsHCcFRfs/KC6lKhbOcSsdD2wNg5A/
3ewbBNnUtJ0Q+FgTlp+1r0QGfCNEt7yUyyLH8lBjulnS319lo1P3jQA0K8snDkKh
pSVu9AujIux0isUXOPAtUlQTKZ5jOxn20sPZNOE6tTROjDEbgcBLQQ21be+aQACj
qxsHZtwiccWrC1eIiQ5wYIqAFhXM5B0/ZpvkRlU5V/r8VDQx/GzqgQIr44wXYbA6
/uZW4YGrdYDrrdhzOQiK3vYNOX7eLkHozIp78+/LB8Wp9z7O9YOSLpok58wpL4r7
SSREVT6hX/s3jydJlftTYznQ09LW742O7beLddqI8qScDn025mbKcSuSw8KnEFgs
USNfxmigd8U3t25NtFxSnwDBSip9xLtGjX4PvMHlWH9JFHj6ODq+8g5+6OJL5UYd
wpGMjrdnNCoUIzkKq6tPSvRvk9xrutBi6TkKJ9XtBhkMcGYpxeBALoxfC3L9spry
n7pbNvlkKmB2RICuzFRTHAKqZIodCTx4EJg+aNuneWYmbWxK2vzeP5MxYodCoIcM
FcGb0j5Ddsv0IZIiYa7Jc3c+kASwfOcIteOadlTfMbIas0ykM86A7jVZ4C9SsDDa
pgi3jWTAt/BY57x1sY7+D3YsUfLz6kPs5qToA9PReiYkgRc66mXu6NTek9fxuxdw
/uUAwc/sSQKSnU4U9kmjFm2QZECyQrqWpjeRhisXl2tohb0zhu7btULwvsuTBX0F
373o3nrvwUKFS1ONUpdMjzi/8aae/PGVSiIIS8DX6mTJNVRGaGA/qr2MRV5qPOtZ
kADJiJRNkidcCsHfI6gHbJ/5DTAM4Sj2EUTH0R0iOzw1vex1E9kE8EucpXqpQsoF
ENgZ9T3PwS1Sr7WnepNjcBzWE4cXS0g0aCBNfj3yBFHE813btCFi+l8eZjjLw01i
t0R5v6YGGFgcdgVbsmGiQ7aYj+lk3+3oBZauRt2UdYg7klwoJ2MZQtb2tmm80LzC
+/zIwIsX16/Vag3fXYIFV0u506so/6Dvc1dqz9En/SiP8lcLp68WWG7CLUkrcCih
TZHDvYKsE9QgmYOQBB451hhGyGGWKBPyy/KF9caIjezc4I2Sl2w+a0IUPUXlTwyN
j0wgsRCHam20zkStm7GX8LiPL58sD5vYRG0YSukrryamh/03UUIGHLwyjTO9/bLX
7O3Z0737tJVoTqx1SmrjASgnCaIG8s1j2mtBMWrHnsiE9dw972w8bs6dBpd9wyFw
TUudcCJ6DSCWz4ZgR3U33YzL0SfagUxc7u2ErnvWx4HlDEFdkKYnu081PXKsjK8n
tRewIBXDzeHWWO0AV3CQI2A3wTrofMqrwyDfjkI0J/udXNgBC0qWYVl4PVyW93Nk
HKNNQPxqKlxTbDd3bl3BI+awSsKH+D8NA+H2e6YXgoUKvZ7uip6JCe2dod3FjWJH
BRmcE2Q+wqUF2fvFryx1wyL7wyhGMNBR2l8IGV5ozzU5n/vcNCD/w2pKUGcHkFa7
2c39mwA0kJZByI8M6+P3w0hR8lojIndf93Gwi+45yniRa5z2o3eItKzGa1k8iJfX
hLySblR1r4l+Aa9ajYML/1bODiMJkx7U7VaFLrOmqwIAHS5GTm+g4zz0N1rAPraG
FxSx9TIjgvgMJKWJsJSUhR36/oIBpsw5iW4DPX2+MrgVeZcivyoSRSO5Oh79M3Mb
NtpoecbjJeXT1lRwvXkWDMEEPiup+UIVVs74VsiOpjMQX28nesjZRiHCJt+yPxNs
g/Capakn57xQP8Aywtx00b5D7o8TgucdONpRheMPOnaYmhC2jXR3eDNNVeOpeesP
uKuVpaUDJFfCdfkBE4KYvYhJTe3pxDgH/hfKLq08vTq5PQ/CNADkp7YYk2ew/IpK
cNvG/RBSNhCUVPoLx0Q1z/nnQ+5R3oDFFkOSmu2vqLr0QgHo0jtRJGytRuuw+G5U
hbSmT+NUHmn3ClC7RHetfNq5rxFMflmJzygw06FQ8DMgai68kSSbDN26TDu2IBGM
Rg1tC0LWut6ghqR+QJEsQkElSKJJQ+XyJdxLE0vYsiXIUFQRHQlIUwHLGmFcZ312
/m2rZjQUreIVYaUbkLrPNOtGisN40iKz1Gg6ml/bMsK+ZU4RJhxYGxXjgbOwGWjS
rqQU1sejwKfuN5guthvrAD/jx3Ibgpdkhg8QopRKd0YJKhJPeaHuxghvMA2JBaZ2
P2Q6kDwQFhurilHp780YhOfALfHu4wBE3fWJcE0YT4xgyElzq8IZq9EaaVHSgmiU
fmwEe9YxlTZe0FtHuRJiWr/wosndVC/+BabO/zkmBMUeHU4teWUh88A/Tiy6sysG
Q8xWKWDCKRTdA1uTM30jRUW6gg1tWhmMvxhg/b/coP9SMOMYRBkDr2VKOWIsyj8R
FLGp0DUNoU7CH6V5p+gtK85ugVPIg/jKKvRIU5LjwzJo8+2X2DnB4nj+pzirWy89
/Lu2KAeetcZsR2MkDKc9gCDDhOGOAJrpV5KV1HDvqDBAApGQAxWBV4jiUv5cZctB
FFDmfG1jQmKXRLMGnw9z58UnZnbLFgHQ3lnYkD3Hcga6t5ayJeF1HN9txyPGOV7U
d6yhVq8nDFSWIdM7tQuUVUV1dG7+VtDuvNOI0sMXYXQG6IMoA1dG0uzhscomDngj
ZtHQPy3AgZfJpQP9dzz3h4Rmzp81WHMprJiCpGodgTsoX9jE3QPEVit55avIxpGx
sBGrdGwZk2/u8vsFonsHz9Az9qygJJ2SIktP/2YVKkamXeBaYVDk8993HTTvDUFF
8SVtdVRrq5PrCPbSL1wpjxV5NSeoptDPz5tgdsQj1TWWiZ6nmfVYgoyQazSnzluz
a8WJ+AjxN7D0i6kIcnqxZR6PATWGpIJkEWnFvzD3hix78uj8dDk/uGm0ZxQzsslu
pnkI35MtAmVxvrs8KJkoaeCPQnze7Di3LbMMPTmQWwgomk1Z2yOIaQrk2J6sHkYA
pLUERAjJqnxF2FbqTosezRjwCpX0k5GuMdL5w1SGSajm6v/BUezoJp28fCZ3+o6J
1JM7BmXEQ1D5k2ce5SvhLKb2FGmGfA+HMinfrstQjnxgitSPIfzvBcnPGr8utzRn
KQZH0iMLqRreloWQrYkgubLlGNWbBbZrZb1Zw7dAILKHHMcNbrTBASsl3tSAE+P+
mmU0AF7ztbU/BMDjc4fkM3bq/pJ9kpcgTDGj2enBOD2sL/uQVb5LE/R36SxXQPyt
6gW/zsVq0Vp4zZ3gtvhQr2rbyuTi0f9ETHODe6lB1qxQGEbsRBsn6B9JyjGhh97A
+Xf/gz+fbm46UCF2qk5Tu3svtW/FEslayhn/TJYbdB1WyI7U7f7lHncL3UUkXvdt
R+cAanVQDKTuxdRjrSoKmT43cuPIZ9yZLwgi+9aubC/l3ZlqLLHAwc4HOw88M52s
f0UuxiF/Z8ieJaBuwGdTv0YRV0gCWPFVZ6fwcwd0wFhRjdXGom/df9APkcu9fK6X
4dZjW5hdBAVCcegSxFq5wzPuRlMY2GvFj8TIROpKHfQrjdu7TFSPjsTlpDTMyT1n
o4gCO/Ox3wFYciKCmoXizmmdgpIvFgxT3mAknjG2wrbNjT8xYenEAKIt37vKy3Qh
9aGrrK8jnxJn6V69LsQHRoP4heRL4x8v1Dn+BdpEas2GzN6MMboGzppmlQfN5B9j
trQD0K2InGstTSfJdhm6lcYhsH9HEEtFl4Sb0JOwSukjAZUrFMIcgzmnJFU3TbSf
0gyHVIw0gJPfO6ZSwktX01tvPekqaexbd7t3XQV8JVsOkVhn6MQtfnpeClIMidvH
IAaGpwCVQHAI2K81blvVyB1BMJ11W1EUdnQMEYytLkAVz6dazyTVqUqoo6sCqZCi
xJNgO6THo1k/Dtwn7wZEPVfDlcrvQRFfeBUy+D9mNx4GrXJDTALcgbGcw/WYD7oP
ZQnrZJivRH5qkC7DyUsOS/Uq0Vt2BNVKyLGbGZSw79JKDjOT+VKS1PwiBxnxQzt8
i+DM2c5IJ+/5ZWsTw2OIBBfEIW+U33uCzoB0Z1JeiryqY1E02khosVA0RG8E/MnL
63Uwo2dPqEBiUQz5PVtSaO2ruIFZdqivU/knUuLXMKKqQPAhstpn6TD/ueppxFYv
xHYu7lE2kKw1Vj6OXwEiNw3wsYJsy7bazlrzRFGya5qJ2D0rtS/drh8VKG7Fj/kD
Bq5kOZHNoCc1o/J4fXDO3ZEa+hHBpGqOBFPNeJlfHi1oDuVmxv4avaSLZyCYtyru
XTRUCbBdPNPwhsDJ3rN2lYd0rn28audKHgi8uXhum9j22o9XE3E2M1nKOzaulzPK
ONZ2WjeObNSeVeVpf8sM5fRkjx1MNDBfub5AkC7J5S/SolZxajQD95qJR/gfOQGK
77z3LKv/J0dauD1PkAtwOhQfsQP1D2z8+erAN2rioGx0nzgrIvJiMd2XX5+zBDO4
69WkZVrG+dtzYb3CHJ5wsnf7dEB7vt3GMCEsrNc8HzEcYIauWeiQSVwUqJ2fIO+E
WrtQlZfyCvg4MPsY2FIWlgbe+mgtzcL5rnwd545A8g9oTEyjcW3lmOoGohm0OUAt
nbHXXqsfwRfgGFK6iZiUl+jrM6s857ONNSNoySL+V2BIPzovaYE3ty9wf1ZJhSci
cPuDnCdY+7mffF28ppRn9AT7huGYho8uLSiERcHlVvAKynuBvuCwqRemFxtpEuS7
Phv9K4SmI54hdoO653YrMYQYHEnnhY3+QPbKEO+lls7nEtvRNYyHFafxc8eE518j
t8vKanN/l6MiBkB16uXHCSk7Xpdi/MXJlluJndxnCzN+30dA/Ylq9HlC/F/EsIWZ
UENVDNqZH89Lfy190I/EhHttVujm6/bM8c1QHqiIhat2ZOPfzGHf/UMpvCq/Tspj
zHV92Go0dMd7uBveGQo5EUNOrjyU4toBPTMpsgdYDQ4aVqsLGBdtn4z1MPx/Dk7j
0CTGmw0qiLbB18o7lpr2XbXL5ioSL/oMdqU0htdH+d3JII04ox/2nON1i/SawAPb
DG6qUg8bfM6zRoNVLugFV1S2mPAEyuYDb18jj5GemJhO5y/KO0dMuaR11OL7SRrd
VHsjkPR4/Riufhoqzrc2JNuPuKtY6SpmkrAkLbZxAatJsGvlG5T/3Vf+3J4psJHQ
vm8ypDbqP9Ny2fSAE+Xa3ChX/I+KcwpEOt4GPMkogq2IaH7S0LlWsB9H8qImOleJ
JSOh1LMeh/8Uvg94jWynEYfd7cd2WkfAXYmsa6EcMTpEUESYMOQBSv3kdJ9KEaV8
rZQgf26LTGkHwdY+PmACA4F2fc2skV7mRh0nqx/ursOkvAw6WmET+ski8v59xuU6
VJcM8R6UaZ2O98RDRJ5IIDnbyt4/v7JpWc/OcsKcqW6qPTYVdRejjXwtjrcsbN8Q
00nOCSJ2oF9D2GZaElikbD6TrIG2rsh1jsXXiJzbpqkZeEY1z5Z/NoWtWpKJ5xwT
EnoPgpSYXL9dRMGMAhvfHFgsU/Bmwd485dKC4Yq8LJSW4uWG1DgjMaiHna8iklKr
wPy/3phLSwKELArbAfupMmUyw5FXS2afNp+/KvMQ0l3D5k+QuFVrmXTZA7Iue3xI
vpPBlb+HKYn06XiX2MzSJA==
//pragma protect end_data_block
//pragma protect digest_block
bCnaM4bBMYuqLQf8iIYhAOlZKIA=
//pragma protect end_digest_block
//pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sWxoPTA1LIFqMCesJuGD5vIsuqIV6FtX305ws6BkKP4k4oVWnt8apKwVhF6Wr7mP
De8Sf/VRuNG+h4PvwHbYd7ToVC9nIGqmezSrhLsSJmfiRxVi3Yh5ehbaN1ftPstD
m8R9ftJn6nIR5hKABnMaQpBKPT3xcANiEIsYFMaIdew=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7664)
uCSHKk4mOjfWT0nByr2ZP/0p7jGVgcZFQHi3+PLXT34DW6qRYvWsfesfxezc6zMe
d3kfKHjxunpMMZ0uz5GzEE635447JFN4vYuHsFRGzoyT7KPvSkybUplgwckwTOOV
6HlzAxHuwkpdVook3k/DSbL9wqagYE6fHuBySasbqzU0K7gyLIkI3Kwcp4vTGASu
QAxk2JUGtPtprSHWXqFSy4b42+fgKr5yv69gORWf2oeBPiPmhqb9UmzOHDtqh4Md
3SNE5TBVwSGtCdRcjpkfrg/igSN/CxNw259IEurhlg3gBJs57kqG+MLydHI1C8Oy
P9O8owedvZCvLtMyOQ9zFW3UZB2LLt6lk3FNbYE+cTgGKVjSK7rNJgDG99ALUO4z
qckycIUTOgO8YPwjrPWuHu0K5nAd8q3iZzexbDyuinGRXapZQfEMtyE9RTUeHYai
j0Apzu1Povz661hi2StwcyHA03aAtUQaQywuJM5cde5VozQxEtY2e6PRflQd1lpP
M/TESD5KTqfVstqTByw+GA5FaAn3+OoC8TjctdaTu+F6PrWhQnLBh/Z6C7tBoc1J
g2I3HBccb8/iXKrsE49BZm3IGLysJwfcA+Zx0SZOql070CZArvOk5KsqKiwn++0B
+3bq7kaXmBEBc7zphqlK29FdJRCbWyQ6Sh2vxlMQnUd46xBlzGRaQQJgjPe8Iwpf
EMaQ0vgb5T6dvd9s+0voQUiaXo5cwovXrE+U7CWVzmaMfG4U5UnZ/te5bIqXWAcM
Uj8fRF2aZMf6E2oum/LeDgos08DEVPj3Z6MtiAFsLrNOYL90CuPELMDqG+F7WdNd
6VbeVe9hX+0PwXPqBrbE6fedZre/Ob4VFgqoLAFwCM7qO0DzevqcF0pr7KTCl6Qq
BgmPpS00Bbp070O2zDqdRjnsEuBVCQTxhw59f/w8huywEcOKarRYFYeL50gAHr3n
wSmn5iLtquz8nm19sR/mKtJOV6PQyHh3KPfAc9f/2VwUhLJYOZkc18X+9lRVXYBk
jBTJjYhU1u0G5ZrZsdtZ/BhY8931lrlGDZZM8o39GYjDEam/AIFfuff0X5O8Jr3P
286OGdsVYB94M6RrwzaRcgjJBSSnD7qvfY8PL+Eh6zvmvhWX1nKfAHELSGq6DEpV
rvyCLYTs/y6uQlsQbOJsuqo3kmCEONSe6Ws02qOkXlRNg9JL9B1ScKk0XjLmFik0
6yIHpALnO4wCBLrfbSa9CQpl0EFzmFaeMW8BKzQSjkGQUXKZq+Hah92NECAfkWO3
HEH0Q3c+xK4Tzk5SQhL6JX+GzEBVShwjZbfE3uuUGqddtCJoXHQ75VAErc/3wg+a
fkDyPsX7V3YlxFtvJZ3Otna94yJtR4AkVZ1D/GcP0mTeGT57Aqa0te3KOLJMw4Vu
fhupu/Qt3yVG8sfO3aTa8mC8eQ+D1YH9+bxHtngCnRA03wh0WqB48DPLlYTOxBS/
NDwQaJswFvpWFc1Tnn2TQuHa+6A1R9LIGVgt1+/H7LjwDG3QNl8dY357ZoG6lzIF
64GuUzxbxqEvmODZSkyX6FGYjbtkkhfs22n2UmbjXfmFsyX9jeRFMfeyJo+pUePA
PDysz9E48UgicdUFeYFkjT5f+vEoFiH+afHBmwMWG4AEL6e6sXwta6/qY+XZCzWW
Es/eKBiNCRg5tBypIILau//ukybKUEyDw+r3nPqYGWCS5NeRvA2Ruix1r8ODGzhM
A5eavPzGOUjwH0ojsXGioYTXpekzG9CjFGLD3xCU4QHIbMa0GUXEYmaKJlXGT3hP
ezQubDeNp/WCc0ob2rUvbQSHpiN+pB2ezTHyC8IZasd1jt5opdvjMrF6888OFzgA
O8AZUqv1ncZkAghXoOp4k1W4G9r90qe3/3oEDvZXks3qCpRMGJU45z9hsq+fqe4o
VP4UsTiy4jTmTckD8B9uCQY98o8Hpi7cHsbxP+9qjsXbm2iLEhis2nqY4DkGxU7o
jIW7zptWVyLmnc4qDswXiEURmEUi5YTmB3N3QVcfQUnzXqkZULtbr7dBies81bPA
GvvlWtM5VjTUIR8MYD1GvPwjioIN4QE2kaUX0v+aO/JhFD/KaYfjRZTLSIAm0227
1G0bvU/esqC99v6ARZwdRzgh8TdGboxzkX3dqTPTeufAp0CWpk3btQX8yCK9Q5+1
eiT2b7Pd0qGUW/YBE6gVd2kC3+HTUrW/yVGBt8lX7dIQZCUTvq+lO/yjFPRlOLiD
T+b1PYLLGRBjbIphornqlf5QaDkorikMMcJeSuPutvn2wPAOGF7ccOGrmWdVtJqN
7mIC/4hjBTqErESiLrLMqA5o2rkYMrxfhY/Gu8NcT6RrGUlXr4lPaZnq6rSEFZF/
m4zlYSr2YPw+rde7omfaL4Szb8+djkC1raOrv3lxzIZ2sGKn/Xpi9ZbCIMuXI7Cm
3n02Gc/T2wCKeseJNQDZc37DAGuo5aT94vhaqfIyneVErSDt0KVZDaNoAVHxOHiQ
uzhCZSsjwwMbox3IWt30FrUXeuGvACsD/7Twl+Nu0X0iW/QN+L1yaIG2WFNCCnF4
aRWCJ/P1lZdaZ43ckYDhTP41UAWRn6yk8g5oi3+6Ei5GM2WhpsrUIs8Qn0DpSOaT
IQN6jTAafVfAK4bMfXp+P3HV0NQn9yhOqqXBYBduSdL+QOqa4umeKjDOEaCqHZ2F
McTLH/sd9cEWMm0XlnlCY8ai0eAwF1L2Ndq3WIMgZ24tEw3yuam2D30EpAi0TOio
rBeqoXEJ26BoDgoJea64IVOta1VUibDU2w4SwedTrG8GFSjimDqgF0+RUctH5oDp
wu4yE+kNZMNlhctsWhYWuzBuMBT0/rTfo+PF1BSjPtJZoV2HuSZpZQoetWrpvNP7
rvWEecJBepbCR34Ym8GBaadcyIgMGWd1zh7nrUQehC42kmY4hHjQVb34ixnnVK7/
i+KztINu+k3FXfZJW12QjUvkAfcgOWvPCRHXJk5C1YWpvg5ouqA0alKFZAqB65Gf
M8opWifNTJwC+6D1K8Vz+L2Q2MPjWQTUZ3kIPjLofnIn1dXeg0xnOxUUYpc9bDnG
VTvW8TkgJLY6v5wZC0nJV6hQq7A3UT5MpqLsIT6p0rM1YdbBsKKBTaGonRuiyl13
oP1FkOLEBXqDrplU5Y47heWBijQWkwIHdOmc6k+EEf0t4voGIxYgGP/vAZbgCNwx
4Mu5el49SbZFJvPVtx1tPkLQr8r2PpmnZeEWSlsooRDyEsTje7DgBK18HjTQTeyH
6iu8ZshmpYSS0yr/wIAl7EUFGHG94S5N4kEAbW9Jm7L1axDq15xSsLQsUtO/naY9
semZtf+YnyuKyai6dVeLoV6rweCGTkQ0x4yV0H1+KCEQUgsVkV9o357/Q6bXR/Vn
iy6GKmscN7w9Zg8B1RCp0PcrBTjTlinjjEYYEbA3abT376DvuGzODYF5193hpumb
eWZiLivijj6649DkMmJ+A+qaSMqenGbsqL7p0fTDtRZKOD+u0g2h60/o2eSZgeh8
LGQWmjjYG0SAeZnayxh/N6KseZDjwZx+C/Vx3ujpw8P6pNzgTppFTwxII+7XT3Qb
JDWe9kEEns3aJIDY2OtftmZ0MyXXtYPwkfvkCj851FzJ2oAXPKiwBW/qkZHtPZYS
IxfDOkTSOeZYx+mKj73koXckBREiF9gT6oRzrufOdzUWqhJNyqXd3ZnMDnzVeHpb
VrCY8e2A2iZBoGZmP08sJ47cn1fKmHD55Iyr31B9DhYjgF4XMFLiAj/1DN7yQyB3
3y/cL6ljc5OweADAFitUJNPBkC6Vmtqcug89lLGDLsWVXL3WI83usS3kogwqTHt1
dXIaWsADyDejjymdpUKg3+8NlUBVG24ckhi6qcZPQ9e9w9RkM+Zn5KNgLqft11co
UGgbJsZfVE+9PAUCWMwaqQMhsi0l6++nxbmjnzdkel2nadP/+tn28rwdCe+PoCQQ
BgLp8VPBCTHUrgxhTohwvgrRcjLmY1ZUdXUe7OEx8SKYJtzfO8WWR1fhReVwvyf6
VGS39odmBNRg849eS/tj5z8xmr31SaXB/AgzuDuX7lYSeFD8/qa1lURiaqFUVuJx
/MyhMqaK+MbEyOBt00QjkX7Gs3XPIzwRbjwO8MS0BoBrLa9zqDhJM+FWZaTU60iu
t/NOkqMcphUoh4ulZilDGroiT7Oz7YTcqUMfvpGbYmOO/KRQHNjx+GFyIhUNNTGI
RMm6i+yaxTB3NzN5QHmfRzshLeq383hqeGY5bUGa+1tmAO1CnlU/2n6NSM5vWOpz
MELLp7u+/cwmb9Y981VZ36vNa4/VBoajMa3d/s5Lp+JwVai/LBVo7kxLJ3KBzpeM
Bqog2IVjw4FLbHn5oJpNltUNv/tvtfGnAygPi28adHxi3gMOfo7ppyoF24VGcrMN
+AgyPkK/pGkTL3QcdGwfPqi9SGLhse994P+WcNhdHZDRZNgvzApiN68vex0r4WkC
Z/Cyc2VYbyGUhoQil+iyoLqISX+X3wFPpo3q+c2x6nK+5V5gm4J1AcZL9k0uyZSg
pbtf5GCWK+YjcBpPxPZ2D8sswGojOdor/5MEnO7oeqT9rjIGk/6tCm1ef6QVPuI9
1Xp5ltXGoyiE9VR+C6oEKU/UABbxlFpYQwyHA7WDHvuE6n854FgMl/7/oiQy/aGN
+jeS4EaD4+kjKYRKphH593N5BXRjXnzcw6tn8B+QNqYiyJTRej5W3itnqx3WiW2K
8ozLYIF0sWo9oi3ZHqNh8vNRuFJ94Qkp7HyvqLEH333nbazD4Hh57xGi1A0YCXRt
pxHjUVu6UV00mGR1Ul4ucyQj5FztkYrfS5TqAbgUH5yquGlP//NyHJ6sMngqUpno
/9Pbo+3Kuqc3dORH5oZ5APg+wZkuRK3LjoCowVxjzVG9CyoNSmDEd3PeCrjRyXPr
mIBv+0Kz1/SPEK2pB/q60CNQ/K64qiMG6NDWc0xOhBa7W56mF30ty+OIm/mVfWSg
7Wn6HNn8yh+0rfdDP77PZ9ihnSPP2B5nn037v3PMCSXnLhIaT5b+HVZq1a0h62CL
8jMn631mfauApXc/NgfA/WTUynn5J6Woor8gUWyVvKx/KNH+qz/llwCYoRICwlv2
5BQeKz41xrfzE3jRXQexiHFpa5TgeKfTZgQ5WM5rlwCGqGv81IztKlXBE9MjQ3WC
6qE0LNVtx+k+Xg4yaeWFmmifNmEkhCfATm+MMRzmbkJeBKO8xLcxLSyvN8689zc4
83LTkkV20dY8/CXlsUrnfFUe5Pixpjr/8gGGrIdc+dGnR6XAjRdp9lD4lEz4lOnZ
P0vRLlzln1O5lPRkeoPflU09FEuZ8iRBy97QAa0XliEyBIdnUvWT2RdGfRO8f4pX
ml8xefW4ciKSYW6c3V5wW89X0bFQELNYCLKVer/mWlkQof3igxtHp0PH3eMLsf2J
SZtMWWZyLgJdDSeTthyLNdJIlXkXsEWR45SkQGYoVJwTAYJLjiVL2CuQfgg1DGw3
wDVfFZNfeMLoNOMQT4a35i31wrxCAotdcJ5jawwu3PN75gyLUeXgE3hQDHl60edN
zP5EdY3eQjNDimf+5cNc8YouXdCQJSNeLEbaUmeNSrNHaxl+VsAHYVYXPsxE3Bkv
stfytkywZo3/KeN+G2kWyeCmHDURsgtYDKklbSWhwo3EFncS39tTGMyQJXFiURpE
iC+aS7Hggvlq8rYyCI3x8sHi3vKXjQ8qVZYFeTcB2TBGejTSGZ6ECiKr4kQtUXF6
upOXpPnSjzvvaGbwLeFQ/mFQrAmd11/5uEAD8fs7amZC92HhvHsyXrxnjLupASZA
9hzcMcgfTDoH/egV/oHhqOYKYYgHw/GuEeSjcGwaV1JLAAJcZSF/zDOgtwhI/tdg
uDsIw0LDeEesVK/QFQYlZUQJ6EPjxDkZ+Q6efH2xmy6ybeNg9kjsWi8i4+cWatui
+ENaQQ/rwse4CCmsd2vYDzRmo7QKqy+ru/THuLchIXH+3fyAAjwJZTtP2i6zAxMi
qkl7ziUnoweGwEkjw1CJ2/zUYrvcMCycUz0VWoFPyWfQVEODgARCFVj7rZiZknz/
/pfj6FoDrd4UyxYAeYSGPOH/oBHO8ff6AIHYeVZ777c+h4kqgKmcXQMQGS9S1/dR
259XfwCihvJvNgvXeS7QDixfCHoppBx6JSnB/VAKHnW1EviTC9T0iIS5KEG0iY50
tTbMnNmhoOXJcP482GOZ9tpL5VQrFVDMg0JLgCIT+89LTyh30o7ip7kQeeLw/3pj
HkRLeMzBYVetfFBhZuJYbNV2O1bPleb5qf+gJjLRvphhXngzEZ1HoviZTuiavaxQ
zICm+i5uGl+PQY7U1beARq83gDQW2Ym8jaPPHfLFZFDFMdygyYNvOq54V6HwZ4AF
ai2kiJHGzAAmJ8XvqYmIkK6iBlSLEfB+lV7iE84toQhA/6g6gWhPXe3uQ9CXGuWy
uCHHIGIISNo2vdWIPgDjg/CQPXKeb2pfCu6nypTMT4HppGD9e8McRx8O6biiQw59
zCg5RxILs6SlIBjPBMJS3PCBGMUGB8rVVGPdF/njvguDlLdBuHVTIYCBHRmMuSS0
SruLrUgZzYkrtwcSxWuFxkxyWBFbC3YJplroDHeK/g30De8hlmp4zrIZ4iXwDiOh
/VEHIyiRejh/WdcTxeQEigeQD96V2XEUbEBxGPobrIxN8w9G4+G//DzJ9eEbDAIT
tBxr2qJ5ViyFBC3Vsyp+xBOqn93M5rs2WDkhDSG7Shp+/sCAqNwG4Swz9IJe9fRo
0Epg9AsaFun8LAe0cUckZdcln773v0eq8+rC8hKM8AT6919D0z1zlimvsug/Gh4U
R+PvYnt4153jSEiGZRHFs03G4fpj0hQ9RlYRHJF5HL4nXz1EYbACdJ+HbXuxViD7
YsFq7ot6ETJTcbdN9vTqJP+bITz8ckqenkdIuBtWvwi6IrbLxY/U8Pa3bvL/ZKd8
tROEtZQgW4azZG7nsvZxwwmEFkeQj2p+V4lkXNol3W2hjbQG4vgATipzZxv5aGvr
qdnUcaJ/R7TA4orG2DwdksXV/1k0yKoKmdQGk34dI/fMAgypsVZYEjInhNs3SLZH
YJBp0ypq6fkc1P/dvbhLc8DqBnLThNkiN8rlwfusgEwa+uSxw+dHU9EM6HMzA63n
qboSTqaIHHJEp0BX90/RdjABKlT+Tv2LLTVEZO+A9IT1YDggVk+wru5e4P8mZ0pj
rk2017v+yFAj2psoMTqTWYaRLOUdb0+pV+dz9yXjCNQghSHDxkHJxLqDyozpWZfk
j3raPER4OmZXWRzNDc9Sgvo8CI+Ig5cpOO0TzsSsPbjlfcwX1xeAGtsIX9YIfXQG
pykecEpzHzBJX7sQNItgF6rYZvSATHpetU/G210skB2rkCGzrQWQGThhgjxo9dXU
Xz/zFSVkoumOzqGDbNlg24MIIESpul5oBzQizE7zp/JBtSNk4Kvxb2TTtJNeD9ph
fDUXrBJ4newzb9ebUHzpmCrIkzE937WfM0b1+2bJoEqzGnuWJiw3lxlthPZgBZdO
qkSoIZXqm2RlgLBdyLw6QuPYGSOcDD9N262hZdFJIbVQhOyyVTw3Y2Cht6qN/O5f
G7TNPkC88aEAmqeYTGIW8vJQNoB0VxcEPvazub2cngXb079eLMDhogUCv5MS1tw7
2tiTtXVwUCbWaxUUNS5FiD+Y1Oo8ewb4LjIIFWV1v3WOBkTi7Bf3iiMhXXTeYetv
hAkDumGesSO4ta5ObBiICjaXk6/I09MDDg/9ldsd4qJQ6081bNA7qAcMXGeqscj7
LG63GWTvenYp7PTd8rjK7xB9IGghu6dn3RvgOqW7TqLH9TfhNeom5+c05alpW15/
g6EIrQZn6XsYV5KyZYUXqfMlzh9QqbDrjpWLMseD8i6/8WJNFoHUmbxFll0ARcDI
LlVeW+7DgnKX3BQdbuz8abGNvxRKKYeJSPAGnY7K+9j8fciFQlAeVMMjkqOXMHsE
eBSCh25bup2oiK/6opWY3UmhoEJPrPEwKQMxf2tqMIAr8pja0TDsm810KfpvvkqA
gQOt+sooPVB52DLQxYBjaO5+enkhXw6G6/WNyvcWw4XQL0d3a4t0mKPqXn9V6Vnw
2yN5FqvI0xfxZEC1ubQNx2zBoOFdckPlsCfmIagf6ZHqVVT/0D5yeCsyr5AQL0DG
0B+oiix84aFz3OpQtqEy/AFjkvSrg09NGiQAgm5ksn8nZUjo9CYuKMMzLMggr4Qb
xHnOjdgYDSMhj2BCYgfnEZCZu4a9f629B7Scm7rbgjWlLBSM7qHWvcHijeJgjofF
Z7Cajt18d9X5IJa0+K4kbSHSEX32nGaxVfngSwlIItRWVixF89atE3Q3QNI+jy1c
6kMPunN6ZkI+pvyoIVZLr2+eptATWheC7KVig7UaGRqgjbGtjdDvNuRIWTTPKGDU
aJuxpoER7MkxJgfPGVaY3dUgZlfoMBABwZtp1e5mKy8bx7ETHdV6wHxyPBXyk4kZ
YHb0FuuHOskDU0AfxWsbSj13kLWUbeFidIDJO80hJ4r8q3cBXVca/2RUpalaDIfF
zom9lncKYyP6qOTu4ejnFQoKjAVm5B5/qfeQ7Uvzm7c3YEVEILlZpQPWEtpdR8WD
nOiqXjLzUXTMZfawjMvYfb9yJQySqTtp+kvkiqoZJWOCZCQhFnRxYJLusDbVnWCD
sg8ekkjcepqTlkDVF9gFCluHNhJvHkbRS2fWd5QE7HVCMDFMKBrHwvGK6y8YwpvG
1lEFtd1lNh7AfBbrwt5xBPeOjbVDcUbvo3BMo9sk5eEXiDmhdnJg8JoF3rBSPzeX
q0Pro8U/Ve+f9Dn9iEFHKM9rPfAZ9Y3GFh5SRvcJ+5ylvJ4dUDiqUUbOa0Fuy6ho
Ux/0NtQmrBD2Fh/eGVMpvKEJtmXqRgeHGReubKP0nwDRglGBYxc496U9dzxTyOAh
NemEpJCQT2NmDEt8afz8/gX6MdG5cjiSZ7QiyHMvhUB4f3t7AccnPGZjAdR+VlLt
vp/xhrgdfW9KIjArbss8NzVT5lffX3H2MWn6Td+33rw08wK7W2OqeEYLVNmLHZnu
BowX50WKe8O9smSIEgBvWMIK/tPHgUvdZ5sX2dRwC12rWtrbXQGKWyHFgUZJx0lh
rWLeQhakx5+tivBhqtznaagiES70HQO3WguvMJZcXVu0aSdh0UD/kJWGi0KtCOzC
wqkOCISi3UMC0KS6y31rT3VAp86KEEOup4lO26NEnuwb5z3YtnwFYskXDgD3h2PD
A1FBuFYJ7dTjmcjWvL9D2D3gdK4gobuQnnZbLTMPrIwg9XGG4aRqiP2Jv/bkgLzM
MWbIyajC7WFnyvlNmpgxOVXonz3p4FiQePw3TgseojI6+g9jAy+FJOMBUS2a/9YE
DcaoTRGvz8P75okx6vHdiKmYO3efZ3P+/m23rlGpfcsT8ZS0cSgskEFyw0nJZbPx
H3+pPjKD0uKU5T95bGkUvTfFpDHBZvfLmCjVP8g6t9J7uIZXjRXwyUKdvVmOE5S5
iR/8ExWFLXV9AYwoDr65T6je+f7OPAagN5v3BPpXaEyP3l+XH9n3awLae4bcjE+4
Oy/HC9pywkIs4jLXel8EFp0z5ou7RVD7ROYcZ7Hj65JpmqGJT/ReavwTOiOLyDWA
2IOqWO6HZZy6Cs4/9yUE4CnjYe4uo1MCSFPDmwRUXUyU2ggZyPM9ZAaw7hLukyLo
XNfgxiiDptlMW3JmsJuYbjM9brpChp1W+KQdxbvGmLehLaB2bmsRDblDaEaXypEy
rRuiIb4ms6bI2mrplP4s2QCGFEcgOhn+hRW/hPZqRy0wS/JRaYAKozucCO4QpGsk
iV7CoVgxo3rR70zpi/oyl0fK4Upx0aHOq6l63Z/+il5NX7VdDd53vZw2rF+Ra89F
Gvfl7A6pcLSS0I9+gpWM3jckWvlN/+9xR2Z0qUWcmdg/HUOn7Tkcs0/WTLctMmI3
rRLqwd8g1j2nF85kCC3ZenbFJnaTf6HYZGHBRJ+IWSajcFsNX0z5SH63hrURqtvs
Ueedy4ewAd1pLITZdgBo+y7EwDFLJEh2Eebz0ijv3jTHZ2DCEuW6OFTfyAg6uuUR
CNk1KBz5IKxDSeggpEoES+vs6t/46tMFObZSkWDCPJBmWcqp5SRNbLjvl9qTNSOe
CK9t0oeKe4B6Qtwtg/M7dc8hJH2uwpjiCVtTkrBoIho=
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
XVzRISZrvDgb2JPlSIYmjB3yZwYLO+cIrNzvnShYpxjUu3/pbobeAMILo2qCxxUW
04zDlbOT0LFusllCc8JqOF+Bmj8wmYxbpXdl9tlWZMe+F14MNpD8/dAFa9w2TDB4
NdkLj+VzzH/4C6VRg8LkTy24FI/9RAOn4mHnWBPjiTePMbeIE2Hds5Ay3LvwUBEl
RihuOYsYaTdk8GIsUpbvNa33DGJvxTTGer3QnqzwFHF1mccgpo4s29HMpYxH1lbr
Ql8dgKoa8qoPMUNhp2VPvCMIWSSF7Cfd+vUurUaNt7wmNY+C+AToXG6OU7Ov887Y
j7TeAmvgdYcptxBzC/N2ow==
//pragma protect end_key_block
//pragma protect digest_block
3qTEhVOmDXV2fMUOoXsOOzMRqTQ=
//pragma protect end_digest_block
//pragma protect data_block
J1k+fF5yXH/HKLzfshFykg52dsiWvB1gaGbnIdeXRQox0Qr/jP4QP7R3WagI/9eC
kQyq5c863tTzCtBDMo133TTpGlUvIOQ9WunbVXYR+vMO54bwVewR1rjU2x4/emsZ
EYIpPNC8OoQBsXP5MtFfRg0lcdvcguIIy/7coXkFlQwDjCEYedavXZzmpInxo3Cu
fhBX5JLBizhYZDN+v3NTQz+9hlWMvORjaIxv5TbouIce3yA6LXSjQKtXagAKW1kV
4srpRNf3uUTQTisT/2Jy8ANfkoG93MO+iX2LImQ+XlMB+eFVCBFw0HPNhes1OlTk
0Q5RJOd5P0HFv50Tu+LAwNUVhOaIIKHaEnKIq0egFygDKvHS988aDALAsmHG4wQD
OV0OwIxzQemRSVdItNXtFA58U14sURTn2iyTEFq8+6VRZsq0hGPZbcqbQxIxNGdL
SfuCsm0TP6TeizYtnqHagvttU8dMfTYLraOjQTSQmsPq3gT4e5yc70376SARX7tV
YS05j2qxrQ8HYScWL7eCRML5NO1cuIdDyqnj3/n83wZ3EdyO/dQWPAZU2yDJ0WhE
1X79VFPTe9bvg1horvntZKZcACwGDQhUjQVIt/s4SEeQGu3Iz1D/K2/gcvv1byuG
EGbdKDDy9fMCd3dWoyNAfTDyZImNU/YDH7khElR9qE7dFsiXxRbYMWyDkp71vJua
+uZ47FOTrS34OzCEqyPufeMaEgpHZz+D7pd0VP51r/CGqbzRbBAVJbYxi1IB6kY2
lqn5UprmNADnwD1rfSD4QDal/jBDCsgmtUJ/Usf4wvQHUJ1U0EwEjUEo5lEqdR2e
LmmNCjGyCgz6KsRNQsaCXN8HQr2xz+82LJWrQedESYS0UWVP7LMZMXKDFZftIVxz
FHtFQlA9oGbfOpscyruSnWFjv9TViJ6OBklZEpV6VIVkPihAwQVvHfu4cF5/iC+X
NX2m4LS4UcdRXmi4cVz15daIyIBnkOkMJcOHDyW82G8FIfP9LFQnbTKNelqleDA/
gU7YCMpARoDwW/N981zo17AGmiLzpAFsURtpxqRMGNrvQx13QEmptm6EBkhMjuyY
yly7zLvS48Tk1NA4sf+f4Ta+jzPgXcCHVKpmi0c+OrWckHFOCFr3j57JGLPLyBpp
xlBYpU22RGFKwj5QSrrkeZsg3N0Ljwe1NB2qPcWeg3D0afZV/blB2fK7eBvQOGPW
7vI2u2QnbGHm5ILDiEWD41I8HnVyshzTs/2wiOy/VB16KSC4Dmw88oLEotPWGdFT
6ywB/x66QQV/VdrCcOXf6Nb0l2zgCIHfwGEjNePE4vL7mw89UfrrI90fRc2qba2g
m4bQK5JLDq81/NLopFHqU/YFY778779ONpiFl6u0Wa/TrcuiqmWYCjeEtuKBvAKz
O4SmGwTJ7RJWst8RlPjFOaghpp/U5UbnUxukErO185E6IlUGrIGWB+86xpnSmoYD
Dt0CxzpDU53GVvHugSGpBQMHNtk3XALw0NdrlrfahPXJnRLqN2jcxpSUjZz3iY8x
eS45wvd0NqnImHrleSwSx95eG5DCOQu0Vk0meyOIZD1xIsyh59w0DjJqoxmx6jdd
0FAfmSxLvaYPhkYpiJ7oH0B9KKtpFMS+1y49LW+auQj8Xo9qxKphG7J4b2qic39q
PDJI8RhSWWH3WJ4YkcZbbr3+PAvhE33r46V0UBvDVgLn3Bn06oJiqzkGL4uU92I3
K0WXCTX44uX9awtyDmMWPZ6NhgQFoCXoDCIG5FQtmNIoRk5um1/UBnLxkryfXwxS
+EcEa3Ud5TqR5+C3cibWLOJ2OOUehzr4+MSgd9rTVXxhE40ZlFP/MSCLxzO58CZT
sGV3s8e1dIwKm/wVmYoajBpqjzzAYXu+klKy/UobueykGXvFaBL6RFjywoGNWxUm
aMcgM8WpPakl9UcxpvXjgOLHqGxWG3+W1VduyeTfRKYyP/b3nzohF0L2YhcwdbNn
GWl6UKTju+xRX/mJ/d6Yx11wufzVcCcfnysQO6XzAtVuT7yqSxQl1WFd87J1p5mw
FNXNhowzfuAigLt8l+Lb+93SZx9s7UKtLwOto/YPX+WuRH0yz1xLstOGUKRsKirh
ne+R1KE+iUKSa26hdBDW2aHKoY8ZutkYajbqQjqQx+QHrrYUlIKyWU/YnDR5bHvX
A9zRiuw/zbwMgcyrBvotxxGgQdJtWwx0+O0o14fySkSppgDgFTk5Y5UGWgbiNJnH
em05AcLRL0OU+t1+E7SqHBb2O8UemRKCLC2ncl4M5FWKZDU1Sq3SnxWwXSxGRNlv
L81qCW8nstT4P5cHDZPJ95xNgueIJYB/B+5itK0IH22GGdvc7GO2RK3vhEM/psq6
MUFzEJ55blCPROllurd+z98GC0IHzauLoRh1cpbw7usUslt0VrZ6MZWNEFF2haCG
Wi9xfzhtYewG4GDi1ZbO97Y2kUIsyi/Q7lfDOjQfs6tYA/ux9ryoC3MQAtDhVXkH
laMdRMvWbKDM18KMjFBW1oEGt0fiUO2Y48T1HmvX5gzEfM8wPT9q/5bxTaSfkmsK
9UcHJ6jlbileh+uJz3XpQY0qHZqad1WXAhOia+p9xOZKKgNrQcnbiWcGMsyrDIdS
DLSjLzXuoD4A3BgXE4ggWlAMOVqdSMDp7Tyw+x8uiTLJGN5ocEXtWsN3+kizoKwb
OckOOMEAHCXFH03Q5Y785I+DJNB09oYTgJ1yjW8svIC6PMwIQMd6gCsQuWviqYxC
mYllxbJ8I/OmgGMID68heJwW5ZLuXrIbrXLKuvk69Lh1W+2VwS6YjOWKXd9LLunz
jEEtOhUc84SphK+65n6sRUV9Bbhzi6nsqRJwA5lOmEIHHTQjgmCTejapOLO0tN9B
szBtMdFICqI0hhqdsBWQlsNYllBOn2ihPjm+XViPi9b6Dl+5T6eFWfiOs3F38+bN
JVYBvqVPE+/d+MtUHhjHZsjL8+qg5cU0sFMl6VkuT8aoJxm0VXgqogQoOs5NdXfV
pWReGZS9bKP5oMm9dfZ8KT7+2oDBcjuuMdS5GaapFzB7ltxBH0omptrDMiBGPqw8
I1b54qyITeuU9V4MaFOaaO9Y568SWcsH7LRM4VfvWfnoW7j8UqITNRgtrcBjUxab
aKpCqrMnxvfE5k355kOWE4K5jA8TP1n3emCBcVin7fKcM6+9e9WDuTPlF7tZZuWp
SPMrb75oxyeuJwzYF/s8HxqQflGLnzHuZ2QeYjHPd1sY/pdf3Bl+J8vuV16l1YKH
RzqMYkpIQp0H4TRiZM9zIsCufTK9bKppkb2QX2gpuBH0iPFgB+eZn/FO+1hIg4ja
KQUzbdYhybxg+ZX6LJ+43i9t75KKG/JGFR9R66gzD01iNvX9PUDh9x+EqV1Xqtgu
SmlxmCNlIA+Ir9z2mMQ8EMW8BQc1qnEpOCucTRHjNKZVtMDA1uewivceU0DLW4wA
YRduVg3K98wMx0ya/+HaEynAPofHepIiZktMSkeLthIHZbqYi70KrROzQl7axs0y
A4+vVzEPrThMfYidBqLIVeFqS++w7FpR4ggn6Xqp0sPjsD0iZ/2xmfxVkJCP/onI
JvQd0FBQNnmaX+khM0rQtKlSWrbZgJeZ4QIozKwi8n8XTFt/G5S6oNLf1SIIOr0p
W2Eb2VQzNtGMerOgRIgHebEZjRFMv7uCaX3RbF6X49EHeeqvAReaguvTEwcWHhc4
jtI9V+ttS898AlzbBoaA71TEvoC3CDJJLuDzWE8XLuJlTkYaGETkVi+qCFqD6tcW
nel7sAWN6ynRKLZNKhYbpp438JnVNz5e2Fu5u1fxIHCS+iGvbPIO/VGZ4WNPdrNk
3l4SPPs1nT/zZYAoy4VHhbwz9xfx0kcVCIwgKdd7M6EX+OZGqJMV+t+0fHunPGw2
QPWdUtWx6b+UB13QjlSxMBmWBVKiMonrSKO7cNv8aPTTeRmsdPmi3EHP5GmZwuEs
fXMaWaKxRqXZQVc1JOCAOAaQpSaJbKhQfewoUfUVWFl7JoIe4EPvalPkP1BAkQ6Q
/yM8wmsKMqbnAZyGROXgDP5n/dPBtxYo/BFBH55fg65sSnwk7i2gB+7aEwdUBuxR
9KyVeAi9xmLjPO75Eg0/0kGaCN9xBuCOSCo6IHofXKcJwmZPhtyAqvNC93xnF3+f
eUmfmYx7zExjhCk8T7Hi918f1dVEukp3gBV4q47aMFZVAKxM6A8GoMxdSy8XHm/Q
mPGVIYfjInjfWNH0GJ//qgea5Vp6Nq5AWyFk3sh8mh91U/OsddMcm2ffCBzYlNEe
ZyB2S3eo/hTuN5tbm9zdIe8sqh4Qku1rXWR7pqWOu4bo5a7dhQqWSuVxGgWqV5Ec
6zeoRCyQI0afU+jBEzfKkcuBb4DfB1KfVEPRUi664WbHzl88QNx16WF+FtUWwfoP
g3XUOJZBqPAFdOqLc7GhyWeuDpUxEZxsa3T9/+uGLZqbUcch5/dX08nsrhRHQtXR
GLPUsrh26Mim/Jatjhl96RG6aPUX76Sfwnr+W4jY9SHciZxcpZZ9pmlO9G3ULY5I
pNjkxHzzEN+fR3EwGCuGezD4aTdR9pVVY+GLy86aoT0irSR5Z5c+QRRPpmxV/KOS
wTirS5tS+FWjSJd+S+B1w/rFR0hORGfeHrJQvuttKu6cniD1LMdHrl+nuxcHmL0s
MtT6JJGOrs0eGROWM5/DIe0kJOKGZRebPULA3NT331qt1vQBou6X3kiWNisbkF/Q
5bm1nX0txcnqdrPn2WH96Jv2s/ZlMX/3F9zMvvcEJD2lQ33G0Ie5Ns4IDqt7Vtnp
H17B7eqhroshGOLv67XgARENN4C8rTX9OVQH73J+ttRFbmfqjQCTDZUrgXqH7X5j
R3O+A2hSqWAbKRMQ654MWvsVUIcU6rWt/wKBqkDRt2DW8VpcXd7UytrGfGwhpCSp
Ke5PeowKrf/owO4g4XHoNFCG2UGnwEhHG1DzUEaIOrg6vD+wWxjROJxPdjcS43OL
z2tWM15UB4+sO5Jm9Uz+f2z7CY4VqiREj0ctsmjnl5js+bH8Ce4rhGOIw66lWF5G
JoI+vgXeyR1UpWEdzWXlmZPrn/WThq3PRBKxg57btUlp1eP6yz4bsWpgsNJfZR0+
hRonySQ+qQpjgc8T+v/isNwuxL32ogavCU3e/EUR4JV5KkXpDSZBtNvWvaNlwk59
xiQ+2HNZ0lxbP+PQoBVUZJiF1tkoDSngeLbgiLlCYNCXBgSluFu52zsNG6wx5ufG
dYlcm6rz7kIth6aXb+7oBxGlt8W+krlgkQSfXf0Dg4jOlNh5u15FHU7lTgrBbqx3
/L5CLaQKWfanAeVHCfcq8Me/JmW/hIMRn6Ixj9oio3u/qvxgU7DkPAavoMNPdvMi
UMUXoHgiXR7vt7FMa4ISMHi02rdbD+HZ7ECSQ3NrDU83mqIZ+CKVyXfttgRTfFu6
WV0kWrImVlzXDAs7YTXvT97FY2+/AKrxVcDMg/fFbgfyfuyrsspPeW/UBkXKO1sA
SvXz40AZZz+jIzRZtWjLrXqJnJZnaPuevyFNYOu2PqMPyOK9pZ1Z90RlGHqYO6sj
tm5JXXXxKMBu3iB1OJm04u8F1/u3N6Nmpf1A93rt9tP7kOOpzJBS2iuQP2dnRXi2
m4ZC9zLpMvj0ytwgQ21u5CC9odFyCYOVCz5cE6soVb3/gFoigq2IP82uQOV80z6z
a4ppP+wSIpJZY264Uj5EBtlshbXSoY3p+wg/sgLTU5V4eWrtiW073yyHNqBs0pXd
AI/CXSOIDvAei6pcshhgLOiB7Jvwt4UKittVrhG30NFGo4fGPprvDPMf4nAZrYg1
1rEGcfQ3No6mCRqleO/+b5wXH7vdqBy2peL7Lj8PvZ++5l3b+XGTPd+Wvzc3iINc
xrucC1iDy24P16B9fsSgp8O1YpgPqu/bGmxwyInKTjo8ini+LUcbCtvbinEza1VX
o3HmRXPKWLlfIaOi/ItHClDQWtQo7KHZIUkvneADNZnyC+11rvBB6feWDKtBzxIl
KAn/Om6NEEd33xrEc5yr5VbAHr8h6fErMfaKFaMUzz0PhJ/J45G6IMVXFnTvuFBT
WBLEJurPt9V3SwIcn4UTwG5lLbRXh1JzjGCb7Vmf7JrY2YzCzsNuLpqm9dvu3zRZ
0uIgiNxgRkMFCANbfaqgJ69vi9T1Fwm9TYG3IUUPDGjjzdpzEJQAiWaLKBKlf3Qe
3fnEgxkXFSzn167uXiFzOomBJSA1Uwsyn8YKVqG+umjzjZ/toa82lLnpIfarZoCZ
0GCyx/KOwibdRuBV0ltv5d3WogcWnBdJdGnUF6rZic5zMkZrL62oJOgHm/OdVffj
N3ERaY9egcT0lGBgj4vSmxjWsLRc8qEq/tHOtsFZI/m7XMZem5Ig2rKSDcPE/kHM
3Xa8ik8AsowaZWhCZLOQg64FHMtRs8MNdmKMBjKWDLvzULvQkd4MyEonRc85+pp6
2TRxAPiXDMXe1IVUBBmxWAErReUywRbfeUXgnvOB6BTlCcTG3eynr82xisUeXJRn
h1TV37/0ndpT9NP5ILOWHDNr4qBiWJHcCWFlCbfszFhWLmfH3NWbnEcUGy7qp8TW
X7R1Jn5MnPXnkcK8Iq+ZOsSIK7R6ewYBxss7SrOtLqMPc1zgAlpJAR5v4xwo4m30
ZxQOCd+qU7+meXCKPcOxedZE5LYcE5UAiWPpWAiB9VNlOHkZUnepYxYWrYaiKbLW
naL6SnyOB1atAqX/4z7oXEwrziqVmAe+dSWov2Aha2E5sjZlSsAxEtCSgFrP/ABk
MI19rvK1Cp1ZENoHp0K/OrVFZ9tilE9vzJZq+iDnwOTOXQc6ZDtGaxrNR8Gv0Y+w
CVctjLdrvo3vSEg0LI9vbAjCIjvuB5Pc9fTw0dfvB7iruvSlWTGz2IufRWoVgyYD
kHxMXR8Tg6oI6O5zpztez5S1LUbFkmBn6rT4W3TG8FGTjy2LAnIYVbnJLXJHOQOp
uTIAj1Nn/nQg0gSTN/GZntneW2rPe7tBvMYvMb+9sIatMMECvZgaXN3iKnxz6Kb4
UJhsq3no4GfkOlhuDNTToMDwor38fX3m98na1Di2I7pyYv2ZYc8K/c3MWFL3mt2C
0rPDiVEgu3yt6hhRTjKdDxT3mdP/ezplie/SiCx7CiXNCGt8TTODY22FqxtdjTos
CwmVY+uvmRlvABe17XNmnF+Z/JYGDjaqSQJIkMWux8UZbFb0FLzZev1eCKAdwwB0
Nyqvl5jrSLCGapWtF21hbAuCp2WRGgvlbHBbDZFnYCdDNoe+W5Q1tOR7EbUvsRTA
tWtv+yJts7gVKwoyGvdOLT/8MKnTQ1c9SrYAULZ0tVug9eZ4TXmS2KFt+CAy7dqL
mk9Lm7FZL72vFVX4pC/tOke3K3Ja5cBUwMtA1p/sD6iHlCvhposW7ni71e57YN6E
anzq8JYXvyNtGZ6IZJD5BcWJUEo1aFLYRjzZtVFeWidBEWFuC++1Y7FCpf7V52zB
s2Rxdt0rzRJ5La3x2AVEt0hGafJaDkh2odCiQH2LnImicbvKypYgW6jophLO6RPv
4TSz/9zfWyM7tO0o3zWrS0Cr552A8HU+6WWDASfry1IF6id8DfmruRVwaDKghJn4
g0Haz2Wa9XK0mJG71hfFTbOhxTC/baAm8A1lPP8so/YpG/UfcXlsl0oa9ZlaHPrU
3dy3C1rYvwlmMzW+Z+rUouVXZl097ezNe+8WtKrt56IC1QZ1GQ6LCkUMnJrH66Ug
j0RJhaTY6LDqywH542DnOR4ZDAwxF1Kdyg1Pqc/yuTYUQMOyPmU0Dv5QWPF6cGc+
rZACmylwTWqAWV6TvTKuvKCUCXPMBdyv5LjBMc1SVyaObcelD5V3101gMnzLuFLe
qHdqOJWrNvdIkDEpoKPxuRlmU6VxHcnoqp9pgWIYEwCY6hyDwfKYYFMwvf2KgaMe
8erJCIz2WXE/aBR3316zE6/bJ2S4GPVFHpywq7uBp3qI2sG7W47WgPStGlQZKAl9
QKmuNzzbCTGpqHcyjbCGxtWb4DjgPpGxfTX3OzE3UcBYX95jBoWl+2yMA2DUihii
jlF18uDkqv8dZWC7xJX8UgiynNTssPPz4P71NOnUuU0OkSIrwaF/WZ9nUC3dHQq2
ekqR4+ifwV+9IIrDsnRmysT9L90mZfVTSCwO5Fg3lazlRzNJ6+8NjUl/YJqYGmjR
ZCef2fFhyNKjn3Yj3Y835Hesru/5YW9kwIWyExHc7Kwq0LGvN5NE6ZXzL9U9S7Qv
BjYJ19F+QHdHjAwojyw1BB4GwnI6sai2x+2Q2Ww7Rm110M9FvPatBICx9DXzEtaE
P2UUhFuYWZJqNKctm17uWOArMXEJt2+CxVzqaGKbmAKzLi0N9hk5tBuEhdYMt+45
dcm5wRlVHtQ2ujo3dw0BfLZf8oxMMEYRmQwHB75IKw2GzihrYo9ix6+qx6iNKHQK
At9GeTCb3vgEx63jqp6yidn5lt5SrQ16HSytF8mtiPQ6g6L0nl/Le/i0n803+2Vl
THoUocROG6AWq9o3DdlZ24WCXDI8LdmTLml2F+G8NJPCY+Yl8SvLWZp6yRyECW0O
lxCgbfQaEdJ+OyXWxlalHVb9oq8JITEjIO4pEhzScoq1j2HQyq3Y/90WNZWZBBY6
7xXND+/2Hmob+8UVbMKTcsKomdJ5h3znckBPTpDWgxH2OfljesAcpi+X1KLH1+97
KoXezULSKIEAQIP4NBVrFwo3UJ1W9WuYQAV0FmbkejqK7sL94CL+sG1svqXEa+H1
1zhupEqPMIiaydV4AX+KhTvVpIQD1M9CUPkWF1qosTUbXjF6DqzFeMd4Ct0uxL14
3L0tgXXqcH7PH1SYSHG5lXUw7lwXdahwX0vc574tp9cntXNfHg4jspHmLk99n+BP
VU3SUj8UXQMHl05JW106BamOWGhSj8G1ZNearFLX3RuWFAqaNp7nQWWfbmK/x7Bd
1eTr2opgIlW/VwfJ800bQonu8hnryC+PkGotWrcDUJtokvO0YK0E8uPHA7WPq3ho
X+7yn8abhzBw+ld9/C0Q7LUM3inbnxxsU2jGd54OVWEEuHNEqQrEqZ4dUIftPYur
0EyDUbG2No+XT78ZTXaWWgkZbcZSAW9fLbx59ddYjaPSMVFs8lzoqZ+ZZOosKC6T
E/Ckn61CAwjkvOyFLQEOYv8B1kl/+9E3Nz1pc3ESge3yb+XIaRBhfY5WHnIAO8nC
sG5qUT8PMxMlo0oYC3g1MrsR6orjf6TXNc+nPkXx7u3Dh/1BmmGHeG7DYW+ONQQ4
s2rArSG0UeCHEricLn45uPaTV6f9Q600Vqfbvj2wURvXsrhb+D8Dyf7QgWRGpNpH
YGxHfRDRhJHk08KJpPtUY132p9v/wYwWiSPLvXJxbpeh4YSjB0gGh6LuFBPnBYGg
UCVSR6taqHYkZ3rjuHxcT/Ej5llYcTcJ7ItLUygAt2or40szOvL2yeQuvXXoHagO
iniSDjHC2cePmVw4eKNo89pQwopLfsNNCY8L+6njr4QatBpxBT27daPO2lVfqosH
eBs5ys0UXTRR6o3MzA7eDgHpIrcyHQsxmsh1uhODWlrfZHcgLE0MABiBHTHMvHLz
xOdaTrv/oRe4fP9BK1fYzQBpwTr0ZbBvnLYqizpg/o6P/iRWrJzJsHu2toBkpEqo
04mAhVmmuIn2EEwduXTjC+QLkCA9tDaRz1O6N0abEh1DpLHYWfNlzEXV1LWsamD/
1dGVLZFvoxeWVYuwTUCq1YtQhp4uruROgX1SHKuuaeYg6GDjb96u3EjMZf+4yrgY
5KDZ0I2qSHUAMO6PLfn+jyQyH7VmW4NyaId5u0+ekBGsc30oto25tiCsjsY2ie4v
4EnPa5iyMJn91qTfj8JgfmnUIOwLgD05Vf8jSMKftPqgtTRC4MLZNUiU2dI29a+H
s0ID6kKOrFmPme26RQXT1ycfokTZPmQI3cv/DNoAIwOcOlzu2rXi+/0JjdWsuyR/
1zophaDq6GPYbgOrtDM0ipOo0kiZ5LeuaZI1DdZxNdAzfZMmHP2ypOYtWcg4szst
3PBCt7fjF4IgwOBEX27rqFYhxlemGcRt6skJL7AOv/35b125D2nvPb5ZjWNpv0tl
9fIm7uKLcbDTMSe+7BhbX79sp1W3ye0QQKeqn9HeKfL8+ZQMGG6MmYzGAPYVnZIp
pPM9AuI64d0FqfW7FtOMX+I30r/Bcj+lSW36BA93k8lEsrFsHFDY4sqrkzl5wZJv
i12ae6jRO6Uc/7KjyQKYIElk5Xc0AZyd7ZxspJ8gUo8f/1e7PnaybQrdvKDhecds
Xkisli6i+/dvoFh+yGC4ZhRJcriocL2Co0idbKgU9NRcOxkrp9JW0pYb6qDhYZZI
8kMhYpNE7l9jHp/Zlvlsi3iLcHcBK577nQp/joJvQMzdEZga6lOK5wv7iePTeIWa
fygOG/FD113RxXSJ49L9uVNKW9EkalmXONReBthg2a511aRuqIOHXDy456Cm312m
2jGNdXwSGWYiGve9gOHCCW3koKdBiMHIy0cywhzGVk4GJYfPj7ZAAwCVsUxeroZS
oh1N/zFkgqBYJB9uRZKuXRo2tbREBVTU5mFtRen0q+TumKFEcXVh5Ba/ZC5zPezP
E0I3b+ON+lNyJ9zxvDjwwM5byjtdL7Mj0qmLsWN9YOQCvUplNDr8JL/jGrmdU11F
UU0EpncyonxjFf5wwlcnKz81ks0Zp3mBl/YWmdFLbuIkpEBCTpxleQvjaXelPAEw
wM3NiM/A2FBssibvWNS60/nMojdojqcrdRg/OSrgrGPpD39/xqQWhzNFSfmutqx3
LmNbcwJUxcgVs/K7YXCLclILwa/0BrNGQ/LSX3r6AazXccKFqy1oTPykBtuNSqxV
ZvuKuYKCGlWk5lE1dYlK8JV0SebLDtmiPFY6jNhGq6TNzhlJG36EGCy7VokUUrtu
p0BrM2huUeJHTgkrr1iiUxVQ3TnZYX5LqdCx42wpGVWevvj9FkOGIbHChZQYloQ7
yBfj5h7pyy+YepXOfPf9xJIjXduucarz/eatkrZ+Dh9boLbrPai6yMWqW6+EcuVP
vNladfgMoqmTg3ldFVNXvkELhfB7Qq2J2Li3TvX/2LoYkT1jhgxIH+dqOil0gysc
vtbBu7OhUMMTsiqtZG3GrxhzE7P6DBDF0OPI9Mg4yXzmSkoLNwLikfhGRsK+0qBa
P8z/DKnyo3VkqbDAZl8pG+HDZtPP4H2j+JFaJaTw+U7CFJ9BWY3xDUvmJ76IYPWn
cAFzIL9Yzs1LSJurzyGkeLkY8vqLbCGvIGc43eYxGd5TuZvXvOgvMpl2VFAE93UN
Z30wOBup7mbPhTu2BObhila4QVq7BEY8mBvLMv5+iNliRs1rQuSyvr4tHgMWLAtZ
15IjO8to5R28RivUaAkIvHFqTwKWoaC8cTygxFaMOy36ccli2vRgZ4dI0bfzkru6
cHjKMEsU6nIE4cjyetSdxdiu6OZXSBcjANXqBXuMELJS/AMQsn6xanUj+sfefqX+
EiMEAhpVIcmdN5Vn2+tCMrBhcwolcWi6C0oeLLQU48uHRRacOsH+RMKa8kbl6Y1g
PetfnAeYgglkt+punSww7r0fbKjO69NZCbqsfeXjXYiPK4ppSlBb70EDnAt4E5Ux
69f9JGkxHhqLhc+Wjl3EJXOzJoHHrI1o/vO4poPQZ4GtnT0Mgk4BW32SpY8wYSeU
Ay0UaPvjqw3UtF8rO1OB/6xjPHq5KvHVuQPbmf3ZzXIwk8NvvNx69sU1rFCggZTS
wpHIoGAOYfCYd4HrZk22qkSOuOKBGpakshmwwItbvXusDT+PoHFp2ywkSh9rcDrW
sajLwmZ9ToDBjr+XRElVGWnEdS3Dc1kSJc82npPEpsByf6cnKbmg32+ligqziAhu
Bd7O3Co1rfiHYO9XMb4lgb26VJ1Q3W4tGhpklgzzGpU=
//pragma protect end_data_block
//pragma protect digest_block
ywwVhS9mrTYiEFak/HNUpEZDorE=
//pragma protect end_digest_block
//pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
zCR0T3Gawq0ML6SAFXo61IRv3KSjwn+3RQfmoPysjMrPElktiXB4+H3tFhprFGGG
Y8n6bFu9OwNqdOlLJkun47zfH3fXI4j/sQvGEzPvWYnmAA4NFEX5uXhstBL4Ll4E
S9TDjK9V1NhdpvnHZhQeZkC7DWsUqWMig2qwAlzOt9g=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 6400 )
`pragma protect data_block
2TuC5ftJJVS3OTM+6qWJtUWyrlyHRgd+S5t01CEGzuETpMmH2SFy90C6iazjejuW
c1BGjdfGRsB0yx8UO4lMFhbqZq4+5+dPILiO9ph4d9ataBRpIT41/eXlCbTbjtJe
wAAfPUZVUsvxaxU3kuwFP9UPXUwyMLUn4l7B96ePtNLKrVzkJi015G1a74ouXiVn
KIkGupzLgWxm13Q3W6sBBuIjVaPJhEyZE27B11pimVTW3VhG8QSKS85dOGkaGPAw
FoSoVM4RwhIcvYcEVEIC1zYeyUWfGhq/R39aHMXNr3dvRiLMF2PYEp6TiRuwI5Ni
Nbfp17j+EKlwUax8ihHv+sDUjnTDgiOgytDMX4BBwQuhC+6eXVEGZCrTcc47Ela7
zBclkYAJehFwDmfQrklgXfkGjvtdWrddH8TW78Yjvot1eYtnWr65GR9+fV8x6BFh
rvicLbP1iPMPHwWJgY7VhmGt1/y8Ckv2wXE3cWfG10yumRgCULzrvfnQufD/QROv
vA4NyS/jQxKXltbK87qIN8C8D4ur1K9DrHu7Jg+e50Yy0Qlg45BeVkMmPwjn1bJe
nPdGUPKznggr9OwCgOGQ9di6JUyK6/medHUS8BHR9270fOEr7gDdPKcnpQVv18EI
8l28KW7sjFM1wNWVqTgqnzn7W8UU97maFnqtZhaWXBncpPU0VLfvRpvveuClyQEa
c3L6KMBBehYH73zCuUZ2/bnnenW8QHPwbfBETZEthzo/zMod7FhbqdzMSyjQzFrk
WduGGnRtJ5SEnRRBfLOLPfh1A1kJYY2b2KkqgJdPX9qYzM35CZCnrapejEuVAwAp
0E+cftD6G6bqjCNUvcSMRpNKr9w3ZunXSQf8neiSRPLuA9SHAhI1PtLho+lMIkcP
QJDCN70SuV5Lg9DCEDYH8uvQlcPbgICbcWJ54WSpK/J5e1CMQWGeFg56k32EFChW
ufipkAZgNUHaRUdDObEKzB9QB1qJuSq5Czk01p9ZhcALi49w9MK8+mKHM7FCA/M/
EBZ/dEZsJapnWqXOa84BQbO/O0j16dnlz0Nl5O0AByrWAMb8/K07qwLpZUiJBLu2
YBqQedJT3a7Wh/irH0nJMSkpKrd8K3pawP/8qcpKnwU/HMGABcsFaMXyoxDtOSvu
s5vj5dZ/3OWqpSj4NzKCUer5lFN/rfpb7QHGzQvuo/xuA3JJJnYfS9vSlPOd9NGp
qEdlpKv4YwlB9sFUjX9vTqyUAMJ6dNQj3D4HgbMHJH4uwpZbZRLODy/7AAais40b
WSGqWtZiLd1KDB4uGMlNgrpxSC1ri9mDsuTga5NgNuTWODn9ef7p3+BGwN+wcwxf
Y/FbpNYOzywO5vHg0IJPxTtUl/vqDhyvdlJYHGBfAAH1WcrYy2SVst1WRF+E6K7T
0t0QXpAOpKJh/pj00fft7GjynKLO4C8Ds+zypJAsUNFyABS3Jsr1cGXkRFupJ8uX
n5lB78mSQauGSy9mrCJamA4cYqqWMuua9+MIa/Kfx6xDANVBh0H+/zyMOzG6WwXN
Cq9CDck5A+gLfQNMuNgCgdswaPxSQ66Gk+tzf800uHaa+0fgovCBYSGNlhHnSqOd
qzov0F2FNTIYl5NuYgyGFNuX4ziVJ+xUFb3KeZYL7T+lVcmrx3e9529nv83pYHxG
gCkEOk/kQfxO82WuTSVQYYjU1oWFRz3NeKxqJ1Zy5exg3DmPMWK5/oII13zBvpYF
QqWdkUwYgg5vgD5UdIASbZUw/0pXqW21guZotWQ6dviR9OILH1aq/7FKLUImd60G
0OayGYOGxcFD+DfPYBSESTlUwoWmLKYZMfcMeUSACV8v6DMnoGaWCXbw3UbegfiK
RSVSzAHXmimtXvuVH9rj+mVmx2RABQ7Em+EHk+/AZulcE9BZ6IpT9QvKBhj6g4Aq
KRQe1DaGpxqanpeCHYomkmg9ISpY45sy8Z+0Fh41EucZiwfbv4e/G9soZxd++iJQ
tFLvJZwuyrtgXx3I8SYlBNnV0y1tpTwbxZmDK82Y1J3OKlF5MKL72BRHPfecxKEx
OC2Uwvtid1VV4oo56kLxjNfBQknM2B/HsARKnh535KEBQyW7emDIpNe3FphaGuK3
4peoS4aO33tYwjNL7gXsExebIsE0jqX7wE1Zsg1BH+D/HAuYGs3HLDHi6GLGkNVX
IU/5igkY2gPmGF7BXwFHpYrn1oK/BuueiqFZqdngkAoFDLFBt9KkgeD2SYYGmuJ5
VfIoFn6dORI3GRW62QVmT9v5bN+VxKB42SqR5fGdFXID65MxUl+ZNar0Thttk3pC
FIikpjWKQC5aICAmv60KmZDl+AqQE6ApZTskVlg3NG/Hq8u6Bi7DKxS36pbNY2FD
Mu9WgzxcVTL2koxDm8KxbeYXvL4bFlB4xXq5TUwGBgd5OLXev0zjEHlzydwhp0e1
WpOwel4Fu2c2yZN2UiqbhanRo18p1xgkximOK5AAqiBwqIEArqQgW00pKgCO7GFJ
kEgHj1vK5tFkdgMgTDA02rArWh32VQUDH/EzL+cXGWc+yx8Qow3kvMYPtVO7flmY
DGE7Pc2frT1Wie7cfhgn2R7k1JghrTTnW2xSCNaJ62oBd+ZtiAGKnRAkb7VpDUyd
u/hyo73UbX5wybWQCFlNZbeNCudCLoO99IJ2uOYlR3SdFbXgttsx8UykdVSgY69l
ksJf4N3ofFoyli+HtbfGHFin3wWak6ipIHoe7x3W/PZDmi+RqYA1iAisFalvOvvO
4pL8l/uoC/SNpDut7FyXSiDFJDA4ZpNS55rcL7dzCJlyyzAODMD1CaLGLE3tt9jt
WwU3Yy6LGnnYeLvMDvmoH119MemSsKOS0+xoWoTbxAR6UWdQMCXL7T6NukWrSwxM
32tg/dRz08SGypVmyEG8aiP4BF8cXsciEZN0Fm+Pq2M0qwydG0+uIsaQdDLjYfCC
2Rbq7ZXGCInjYSxInRLnozluL/Wd5pwX65E7z8YoIZ245uhWRvQPmw0VyC25mBxa
ULebUi0KE+H/YA2v0QIyV0Wl5+KPEyHWvhikjMA/RTuNCuYECa5aaguqd5+/0nOg
gygVFW59crGmPTg91GqL+YTNiLCkth9nLY3oZE8Lz+wv2c2mu3MOt5s0trP6Vgqx
F3VUzB9g8nP4ywU2WQ3dfYUUwp7KXwi1siZx/x8xti3oUfn2FjKWqhxDOTdsse5P
IQ13J3yk1kkln/Pl6do6AKAYtBSyBqh1Ua6t39ULXd/JN2jlVPX5HDogAgMD8JL5
k/iGxGx7O3hwSBVGAxdnjXwoldoeCWX1gWuckvmOWM6QMFysmqsYHR2w8iMIcYth
0jSevJL8z6sVy2eL6VM58wk0qSja11E1OqU7eggexVFodo0z7NdgoHHcas8ROmRp
J+wwzUxEZLWqaHphIOPkl5h+nlqjgjVGQz30Dc08nJWpnedhkyNukiMlnLHAPjvg
yVeqSFnCcxNzMHGicUEVIx8ZLVWimuaFlG8Quu4sXqvCsdE+5s+NfhwV+iat03CU
L8Jneu53Mntimbsuaej1lupRGBK8wsjj08BemF3WUCPvKjjEecpzBwuuc0nCQxMs
a0sWlsaiEx6CJ44/3OLVDlI6P8PLX/PKMSQ6q6rjFJHa5iZy4vYhIqbLfuwpA0ed
zw4OdiWOqsJ6qt/5mhevEOBV6F7VkHXdAA15/cfNQJ1NojsKqP1Mc55HNvgb9erK
5SA8mYEmkFLps+2Ss2ea34bWsQL4uehX3JIZhIU0c4OO+t9H0Iu8ig4N314THaPJ
Ku07Iqad/6+49qqchcn3AVfnvUAhhoiRsgvq1HkAlgPgiI2DjhkE2Zp/94PHY9lt
rHI4xqEUaF9bplK3sw2z66z0kceg64qpFqvRDu9gfM3jHpGpdtc+edau86WAG/ez
/uedC20atksnCX+hO1bJYYdsccD0aObmS0jCz2O2zXooTrPFb9G0ee/+suGwFPyM
nGXaAaDW9CGH+CMYp21rdJBuk+QCLaNu3bte3DLU/82AfqWMGNPDTH/xyrAFyk+b
l63qprr2IY3zX9AvFaNclqcTdK+P+5Ry2QQKLMTSb7cPwYviM3qAu32V245JEwsM
uKQ4/ixRzY3a0K8b/nKZjG55rMwlOadqnBJYJ4iX3ssaYXW9hv74UGsS0fXgPnKQ
OdG5AOQgwrKMfbwos43hI6aZPmzqTUbjS47hc0KJbSGcYFLJZ6QkQovK2Xi5oZ6h
J0Z7dcdTaLznqOX++yXs5vnEnYrIlLs7inUwHg6vnuucsDQm56/qwdDS6qtnAhKI
aw/tp3GiQCaKgCikRYmdFBEAkyfcag7dCu0oY6Ouu270Bs0J/IS1azGJ2jhEtupw
9u64H2ZL22UEc9s9t0xLKZWoGvJhyXpezt/3kBWNrLVAl1L2lNIpvcP6fXOxGaOS
vlx3f0PvMJ6Bkg8vcq/P6ryw1BnPaIPvPWLv6LzfE/GkAF9nN/k5z4WSyWPCjTh3
j0NPM8lKSqpr4nd7J61lTQDYQTW05Yeo9VOyLLfvwa3qwjoxSrD3umzJmPbJYDpY
F6U8ThS0M3eZqd6b4tAYlE9j4+ngHbpAFNswZP30NkQ1t61ZWW3Kgj29O0mudp3R
FDFlID+3pMTx+aergwOf8m/fKs3mZtjYT9Hx7pD0LPZRbbOHisOicvT8IqFPboj4
yLoTVWkdIfZ0GQdG653/qxzxXBlAghcEDvIfLMtGSLApCXGxXDxglvGfxTbmYmBJ
bb/mIj3155iyBgP2vE6vmF6kgr7U8/U5pRUNq3t/rx/4P3gIB4Co49gGywOzWKoH
LKEi/KvgayD+XFFnot+u8wADTfJg8ze0P8VxmDGA3tOYXtP4W4QQ6uip8BhRSXMO
KLfxPnYWUgxhx9SeEt7IvWMhd7pgMzAL2ueb5W8OtOudohWBOGJNvbh5aT1teqlG
Ca/KGoh5lqWouNqNd7ELy4Z1b9FNdOeNaHiReobrb37DaTMK4lrRArOfBzn5nfh9
X73BOfn2mv7DORuf1TCkhSkDzsWDOVTmLnQ61eMk4wCqHIXrng72Dm+gyZTf+H/P
Qrm4wp7E8VFH3yLa7YbY7h3BKlLQGWLW0lBhBPfbdhNKKRnft4UC81dq6vR9qLmj
Rfe0I2lGW4CImrHbR+mfbZJ6rvCgzusMZyNm92eQZne/+EwK8fh0KQPeDPTfyCTl
1DJq1ZMcfXnFZN0LgNYj/yaQyJwvoRPP3P3BPjhMn6ZqkD7pY5L8So1/ntCoL9Yr
E0TOQfpMvhiGfRB9LucKOC1v2cb4gnCuN0U2ZkFIgWODwtxdc1+aMujD7kzX272x
3hY5Blr1PUCx2r/RS0/S1dNGALQe69V0BGyb33bXDXVif5rH/kuO2weHQEZzwH30
e5Nx8kCo+ew6GYdtyJHd9SUchjETF0U4r6qkhwJt8LULxg0VdpbAtk0h7UbDWBUN
jw2pJdTdVaR1Ki8YQRig+/4DOUbe8eg5CTanL11gsgGvwtpOXK3seN7YqjfDegFv
2ZbXE9dUjOaQUeSTbFlL6eKkHs6rx61EJk6uW5Rm89RwLPJNWvA8wP/gvWto68JS
vEB0NSpRArgjFEdr/cphamyWrr+gZ9UkSlRJKlkhivqUBpUZ2rc0XFLA4i/xlOT1
+PyEXKFvaVQqzz0lWGCzvOv4twwDGrguEOIlEXIKIvfIPpCYdowZnsrbq009SEcM
6kIMMvNMumAvmG1tMhUxSDI6tUB99AorgLQClOvb13R++I41ID0A1lPzdNmAvHiq
iuZrDpWgqQcLBlRZ3G6mkfBoaTXTGkeDZf3tu40Sx+Wng4qVzD6rlkMvIHG3Hd9g
JRjwfjQVchnQDmeD9UGG1qhX7Y9lz+2hrLmCjkn6DhoxDpk/VOOIDuE2+Af63jX9
Q5iYS3WdeI1GfBfvX3MePHO+nBTkp2uYHK3oyetrF97gYB6F/H7lXJm9+15KO9CV
hqRAyB9Esv5/cBsVqlIWpNefujm2SjC1I2AFfoQVOE2diy+kbHvEfncGwOhvTIrH
6nqYrbon/x2WfP0rqm2y8YqhmdvTU/x7lBolqkjk0SlyVlk/f+Mb+gBsnoaH4vYU
8dXF6cWIbeusOSjnCIQCFULArpYb4mhkwocEqOdwwiMLYSCHTFEJSKGWMloZZP7i
+sqOrh6lob804FCDmVibdmDVBa5I+P7u5Ie6YeQkcEHpbFsq+9CUgoTlSqnUX+aK
jfiIN+FK2z4kXAhuMBPV4hF2BkM7JfyLM7SxMfTRqvEiYtoOKZ05BDlGaCXm+GzH
lbS0NP1HqPqOuHeSfy8eHJnmUV2HHVCSVZ18V6rysL/+DP7QE4zZOepLXGesQ9QE
fWI7YqSjmGRJ5xFJL3waFdruAQ/JuRKnoGCYgyQTpgvdm2jfdiw23mdnkhuqykGW
OUVwT8udBkpz+kcpmpzFoDYjygX/KFut0hEAF9K6SfHAN1I7UAZfN6ciBq95d2cV
MwUH/Tb97haMxY/xtP3yIgDx+a4Kgmciog0wJDzHCLvdDq3SehheBmRbwN5etNU9
f8B2BnGv4aR0TlulGBYb0pnE+4TQxMN2QcdozV+mrUDVLbfHYJH9Ix+sy1OU9cMP
5EToo+T6/kwT0j2+RBeXrtOaw6A/W0X0mzmB/IdFwXPbxogRhmK7Aot/p4H3SDgd
cNxNK1FyDOiVYtop0twFgvNTlrU/vzmxT8wWgPkHkVPnRa8cD25pKM9wK3Y7LFoH
DG98Jm5+MTXe7AEfVoGDuGYXGRPHG5+hOLaV655n9jNh1SqiHEMsV5KOi/XDEyXq
J9KHqPfS6I5OGnGa+CC1y9SQAGGok9TVsxDzuwt9P0LPneTyBKIlHXZDl9MioVhV
phQREqYIEUiVDGZkOHyOEqXFqlDsfK/an/BFdhIZPKAzOpa9B60++xlqiRS5JAuk
v+lkBtV01K2l/epGoL3hORkHSFYlY9RWC+6Xj+cKv+1RtdoRZDwKnO5WNHu0Y6cN
seTrO6L1DskIYd4pc0fN//HYPF2bXNHrZ0LxgrK6ngLBmVX+hTixfPM7nVUADIPl
VWrTibp0ropDOhAQDKW4EJexhnPFzViQcq//vZMMYTEvBnBlFkqsuBcIR1DEH9yP
9QaaAwJYaY2q126Z6vQsh+NlzQx57a3vy4oKRalJPniqFLUbGpib+PD5mCdzk65b
nCxiZVm/DrRLgENNWpNdyM36/qS1SA2tk91jSPMz6QIUYJPe7/K1/JPUM1H/+3QO
dxxPi9NXNATYrhyjZwybqPdpPZrs41KGm2F+lDGGxDfCKA8SulUVzdtdiptOstkJ
WDl8CugS/UMaRTfUOHBscZMkQsVBZu5mMc114Hy8GzUkZamAP0qP0/89si7vOiAE
LycPRLng8hlBGFiXGkfXzKC0HxkCHIVmwL4hh6ON7xkRBYS3c35D2Zv4urh5lomc
ZHQHOhoaNuidesWrWfTguOCscxu+9N6/pkt2SYq44eXmqCSnyd+HGfhsQFqEIlL2
oYNupJBoZcLralg6q2bb5T20X9rAWzn0Ut061lv3EOMydNIpHd6O4CUm/+Gw4kux
/TO+CtVxO02YaE+AmaeYsgYgLiZODM/4/97EPdLAm/jPPP0yxxEVK3U3ctrFOr+0
lP6kcQ90wMvEfAF6lIvH0iYvglbj8E6okq6DvZ3aLR8CR8ZUpCd3ey5T0GWdZhqB
z5thH7gNTc8GcsVAX1ZGpgcwkRUfFTY9Sr6+EDB3e6eC9DZinqRgCGTVJp1KPdGy
F+L8E3cBSLPCMpO+0nxS+Nhc+SYExX7h/e9oC5+IfDGSjFpCeTwfwyNqZm8IBilP
1TWOk3mIhIhhY2AdgLOtdMppkq7vg4vRMZ0JBgLNFM6zyRmgDqO4mzCUzGG4Brx1
MQ8koGSojrOUZ4iQAse24V47TpwakDaXd/3nhyp645VJ6x4Y1KRa9GbnJ8p0xhSI
PcmlDFRpidSJPo58fYAnsNawb518b04cHQgCyg1Mbnn7uUrEXGpUb3NKPy0anfpT
cXw2vjSk5M+VKjOqP9GJhYyYmEGlloYEhdUt0A0jRtNT5i+xNQVUKXYi93cF8mK6
YelFJa7aIkcTRRoWcfS6ODQElTl/7+vMJleFnhB4jneZOCHNYSo+G8Ne8rbbfcib
SnwJgn6Qt6xKXaoF3iFOesenKDgjyiWYkSI8z9CwVp5IX5VwuJvmGFL3/B4PkE8l
ytF5pYJE7PiN9WoK8HoTrWiqkBW3BE5H4jENiBHxFs00FZwaK4KiWaRxnEhL9Zlc
jLOH/fl7dP8qjOrHzTMxdKNcSd0mGE5Au0yWS9ZoObrY5qbK26n8T9YZbc/7oOuc
GL01qZa0g3I0uAZthJJ2BXVES0yf2zzKs8Vd2wc57yx0SPwwABjEB4JUroNJr11o
GcYMbW9Mt/OPrZnp5bK4l6ssge4a3bsI1ag0ImOs83mEmVRSmyVIhAYkr5Oln64K
qU/EYCko0H4AOE9tpESRDri6IiWdwv6+KnHX8rNnDPMQRZTVt65VS7RbDP8vSxYP
KAhAMwCM4wlJu0DZJu4yfw==

`pragma protect end_protected

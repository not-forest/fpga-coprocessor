// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
ct2nTrrrej44D27oIo3eV4vk0VCsEBQYdRN5G/IVrz9/FuGG9ZVzBJ1JBkAoJ5uG
6tjbt5jA5uqZJ6C9x9/GvO/HX3yEhM9gVkoM2oDITmgMjuhqnA/lVjpkssmda8pE
jAgPdsCCbNl1Aw9pIs66m/ANwBsz1HZrz7bCK4dFbY8=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 6192 )
`pragma protect data_block
aSBz8DJ9vcGUvMShw1fU8whr+biAJ1fMmelT69LOdRUHMUFLX67zANT9kBZguPuw
eM3arZePe+MhBj7oRaQhJgWKtXPAo9Ru9sJpuna4qFBJv0j+JZ6VXwabO880L9dO
TciIU3oknHrL9MmeEA6/p1XtlSIAz7nkMPK5qGN/5qc4UitBSttD1PUYK77ha1QR
EzqlmQNjtRhz7oX5mRcCDY66rDeSyzLw1EryHIwQ1B2cimIcqLpB6H96Gu1gAEae
o/SiGMT82Srk5WY4LLw0mshcQ7gx2yyzQFTiucq+GGhH4iwrjPaLfQaN1fQUedcc
wJQXbLCBK/AM6weDbu8keT7h9e+cFzusSYKMUV7O1wgLxINeCSNbfauIQG19Fviv
0cGi9xMYF1QLWP5KldVoGkQNMTPw1YUP+VyI7ClbkEoC8xHdbX1kdWNzpje1uSrv
aTOTEp83nj+xJfpPE1k0ucLjTiBrbP2hIf8Nd8WSEy8YrqBGey9ChYbJ7pCReZ4g
uZpwiLZGq6n6Wn+a0O1b1VvZA3TioTH3jgezTaFYmzy4BBAPZuq9adVdD2ggMTub
3ml1BJvzNU+t8Z55xatXFRxWiJvdXFxJ0KUqoKPIAs/dolTPQmEuvF32C1ybkQCU
xnko0Wi4WRGkSeV7o+AjIuu66gk8ytmseclyKBPxw8QOdPBlM97GHhqeRT46GagO
w2Bsi+E6pBaOXViNlM/TzdShCd537ixYVO05pHDB/PVDdF0WWJqL7NmbVZwoLLoZ
mWOr976R08PaANo3bRiPcfMqKxRJArjC7phspocP/Wpn2FGkgh0ibyA9AjGhy0j/
5Uch/qD+g2BorLhbyYLf/RhWvQe8MJy+cIzKDgwchvtPC/n74UxXWmpcL1Q77beq
at/G+6ijKVlZUG0j6RKdhw7F4WRLZZDiZHHSljtcdCkyr32rBhaHeGsMLpqnzeE3
wmbeGCTtLDbAJImtY3RR1Hn/pbLPj82egvJ/TMjGg5E06IxLnOhJrfR5tw9mRaHV
HCA/RmNmQK7LmQ6doumxzKos+4vVN8wStLkgApZVPnGK43CnRYSw+0e/VGVa/I4w
8EvsSS4Nwt4Au6B3/Q7ek6ntEgEhskJWmyVyVXhZzg3Ki/aiLy8yQMgLfB12AyZh
bmPSCPJNCiytUX/D3EneIEBapaml4OIv1Mw/SMh/jWyKR6rs0dSLJeUTbVKM0sBV
eQVo0WqGlrJC+t3ZokuvHCQNOa7hPtOT4DJR4a8PAL8fBQwkYkZ8bAuxmturAfl1
PJhYT01146lGPZcakxC+sSOdwpNRfVczLs3qOEW027dKnEgbjygdusf3yFqOjbQW
f1TeEgMrctSPmKyUqkeZm4Gnqa5EOd9XtMySjr0vSl/lI4y6wQkihABUkwCn4fx6
yB7JbmFp5V843Beh2BDx4at2qt4r4in9J1KFsNsDG+QcFYtaHu3Pyh87VZI64m9l
JeuwCO6LLnAaflixH+7Dt26P8JOmPhIfsbo/Ny9oM2XeulWBnVQoM1Wk7s3Ske1h
WvxGC+X+my0rB5ZM8rXXz8PfaXcm0nGXQn2eAAM4XFD3kSdRZ9aXs0thNBTly/+t
s1Hm0kMRuYAsym+AlgpC7G3DvDANctlIE3NoRs/8/FipoRsEPoLBBfo4GB8PND2s
P/P21s3rCDYD6idARLxHB4vDiC15y6dsMiMwldmBSeQjkKmFoIskwmWgnsgPul+t
aNPKNorSJDp9/sS/9hYkqNjMVM16fdMHPlRPD5PRUJjOnpd9HIr4qJ9cDX6zDxMk
mg5EDL8wu5CcfNwMs4dA/aB8BESM4dpPpKj6G4TVLY6F+aodoFg50FAJzGXL1yL2
ggW821wAlWEcyyDQ8kQps1IWqYzOsUO3hrbOcZJUq61I01eS+qoUQJ88xRzHiIaO
bG9vvEy9LymlfPVG00e3/FWCdt8EcpCndY7Vxsj3kght05aoQ2NkyHi0GTQpAfaN
Z8wT/bC7AOe6U521ZrTnqZBotLFHQfwEn2m3y2+iGUeV9Fpv4gaY+EVkRd8ALmN6
Y6Qf/7lbvHnJKFi/MYv+7hAEOHeWecjlJjLoyiqBRGZY2tiELHU/YyVS1t+/s2cE
zxJSLCDXJsQBtkO7Jq96kQT0fp4AjvbVnCqzbnP5wNAxaSSj2dnPB5/+gQDGM6g6
fNmgkwH2U2A8CTXZaXV2h4z7xYrgMHcdR11CJyTEPZudhKi1oraGe46oghrAeo4o
6JEvUaKLDQROWs5T2b/HuW9GOYcFzv7mMCot9y8HSunAfjHx5kJS4LA+9fhb5Huk
w3wqsUoKfv8VwHcXC83K1ne9B2ZRydxOQYHY1Vm+c0mdDpGbjGJu4X1m04/HGro0
UKQ3shToNKiB3dkYN8LyQOUCKYG4wq72sbc5BWOXDf6zMi00PVv+kC0pPytKpzlM
x/6zSAejPF/tOvaMhvMJuEVOWBW1HNKIIJE6OtK/kdtpa1wcBCF23DVqDGalcBFH
OngWEGmQdlIYKojWiXecs/akgUUAqKE/SzS2leV84yzzAI7srIjhLis+Jhil1579
rTPT0jE41I2JpyrO8Edtg55UgUKWI4F3T3ctRq3dArxZpkaUPFUJIfGXwksKnV5+
bsF7ddbHtSvuoWxkFjEDLiG5Wt2lKEU8fO2zGwRSiiF/X0/JAVISsGhQelu5+8TV
kS54BGpm4v6pZHV96lkT3/3zer4e9JavG0glm41MqBZGVVYQDC7JR06VkHkwZCGO
A3j7AkrOelxXivj/0PbtLNpPxUo6aOuknd8DDCo6J+tyDyz1svFP8n0NHRCxkIQ8
swKulhr6aYrzG2f37KqVADEjRCcqtYQwbnbJUNcZg/l24ksHFha4Oe/jJ8xXfJEm
Zl/v9ZLKBmbpT53UpDO5dN1jlq6pskGpafttFY0uY0Fx//1GEZA3S/mC2NKPaGUH
4Cd3L63uA/y1VjxRvWcHPGrfOY5bImaZ5U7e7ULvKeUyRNX3CMn9tbyExrLyCvpP
bJIdXgFv5cJR8jjxtUM1QOF18BTbfmUgbsJaBO+jBWcQLzA4WZVR/KASJMSmapTB
/GCPdX5/QrxKbozRrkdlnzGplgwz7IPFSSdbKZT6OKk5QqU63K5xdvO/GfBtgbz+
AGv4nsFU7iNujRh2BKhRqJ2EosPdPW3ZArK7pws+aFECjLQzKK8QlFkPLlIr+xw7
xFbY13jwCu6sjzjYNyWE/JWsxjHJEMfRgGPdCBZj5j5TmE+MCWZ1jrnNeVci7ji7
fOIEDlH/BNXn68MCT7UeCn1IjRQylGdcFQ23vVcEu+NvgYUryDACgb0I+ju+Mzdg
G50VnjbD50iiAkYBuMNRZicftWT0dAdeREMl2fw6EDxbW33SpZNd/QJxTztbN3YR
3s+BjiMitOAwcvJoX3bLaa76UenPgWqaZZvvGoCuVk/v/GXJyS3oswd4rX8TQ2BI
M0VQ+IVWmDtTGH4d5ElUa87XvtCrWJ5J3GCJacwgy4PJXUNrgvD0/UN1KlSoLJnl
KeMuf/Zty001g++HB9Ch052IIcJoTarCeP07RpgiPxOiuGTwKY7m0R9YS1yjjyss
lXNXDazVbwZTfULAfNvKwDAF4f0b9Q1GzYqTPAm8XfdvjA+KjyUgliieh+0t9Lo/
px8+7hzh5RBIMhgN20oEf16IxXKYFs2ZBld9VBjsGBChULbQG5hdT3+YolXGV7DL
p7NoXizJ5vMiGqFa6NRnq5+G4o/zF4jngGbsdXdFWsRkSew1pRUMoj5g/Ei4roAt
SMDNihOrzFAnD6qh2Myg96gxf6fjalYw9tsIdMj7UC1YhpSgyYfraxnPHTxMJNf6
bWy9wK2YYFjJ9wHO+aGgXrxCL1hy7ezkj7zui8UaE5CwO+bRZ4TargA379Ntggju
R7cOBqG3p72xGtUuMv2PgXG45qjsE2wPveo6FoiNoPWyV5RrL0Gf+87Yf86IkHKL
deOiSE4/2wXRwxotQzvUtbHJfU6vcCc+Z/1BlSoIWprv2iWmx9cKDMVd6g/1gWgN
3zy93AAQNCQ7j8Dm0g/57dGAX0cRE7wTcrqV67Su04f5lz6C1CyhHGxuWvAeAIqN
78HTbF/f5O0Ip2QkINbQHWq3PWg9kEam/lXJNPVkeLBZrgT4tzl6EBa03x9sKfjy
KLesZrm9D08FGkp2HPFIS9/JUTfzPDBQ3uKIIqGFtEGTnrMPQOpKTyEz3kerOiM/
AT15bGk0l/eOE2L6PO8ZEH/nJqUpBiE+7m0mWVksd1tAoprtaAjUgxDiAbmlMhhK
QFJxiJClJ+u8VhWqwkhGCJOl8YInX3vPfE8I4jS53fxg2QPwl3CuiUBruOmfJ7q4
bsROUqCmyXlidmhFIr0QMcGObCZTbASZ0x7xBCuiWZPGaNGaSV3N+RCxWiloyxqF
zURDjp9ts6fPJwZpxME9Ah6DFa1dKnLKmPBZzlqQFbXij2H3JSmW+uj7cN5fSfIG
9yOvQFO5ETrWq/q8vSFnRAYxx54CFDiNI0QSWAgJoCfSJuj4BD3OeJuYvABeQacj
lMQHg3kacINavzvth9iC8sHf/RuHfqn0Ap+tlWu0Qb4iROBE0aXUdPaDcz/zWNZl
R5F/4YB5hXnq67SLMTnYIwJrcZuexC76lxG2eykFG60NbQdCmleXnEAClYcl0nY/
szimeeRS904qpH0qsY4zZM9F/XW/VS09xZj2qOBsjkyjoU45At+257jj6Upxakit
fCmuul+8QGYQ7s1r/vSfpEL4Z29EiKwqWYhbvbdODWyPw2uFjiUSyLZeEv98GXnt
4Hwjb0mNWPY0iEV+RGuN9/mexyEKeDhpCyTNhh/aoocWefQ5o33EaQVPWXLk3+LX
0qBL/to6K0b2IFd3qs0t+fRFVTUIbR760kF8v1jvwFBTuqxZpOsasUARx1cOTWTK
57SWsOWgEuJNYEBIgAKci/yKN9vzfEMNe6pDZaDhjYY0fTaWT/gxhGU/PyRzqOhQ
TKuYJsMo5IsQLmLB4iHCcV+l1oZeJpehsgbvA9pEN1KEAOFFuIiq3wTu+uRD6eHI
z2vb3+iKiqcq5FaUWupUwwD7l19vXB9Iw2Lmf0rf4vLRE8f+EIXdYZbOmtGg1rtv
4hVIjQyHN9LVKIESw4lvnJTqrCI9t+v8B4mFa+w97S70W8vbUHUmnwin41i3fYul
fwybRj+FuI5fpOyX6QkXM2cyaYzn9JbQpntx7LKVPnJTWXSpa3gWtyFXELDtTSHZ
LcnEEDzvIAuFsHVUEsda5K/twhFFIYL19DIEqi49Z0K/W8ARxJt/oH7cbDZqrPqU
V48GheDm7JMJY3/wysnTz8wUjtEe3M5I2wbcScGt/nJ30PF15Ho4kv+DRLHOfZHQ
HlbGNsUP/XPmSP4mz9oVF5wPNFTTKgVne0IdxVRV76bJKn8DAx1/DTGzajFGmRl3
oYoC8zbjnaCPpzTKG2sGqT97T/QA7kiYqFrEXlrgCZT/o6BZ/xfWwXs2opfkL7pU
H71T6uvO9/s0AYrYb9vEN3DOV/oW6XBwRpUNMGTG1p4A9PGGoj3I94dUk9Vbqe6+
vOxi9q8dzkTd1oxtzATDCs5gLqOfEsZsPtkMqrRbERioX5sUJgFYnQU8n78NhON9
PmLJA5bBAFuz49LXvm0r9GBOMc282Lw6Kmi9LBZCV9Xv7p/eGN9FyD0OPFIG0gob
+tVIucwc+NUJV26EVDTrr+IgIWQBmyuxl3sN88MwILLk1HscOj0ECX0mzSV7QpWE
1QmbQzh6/zi379R2IDSoi2yVympkVa7tX7A1TzKShFJg+ueQ0QsuJT9MSuuCVLvr
q43gwE+coe9X8HF4ZRO2bl25OT+3Zs/I2qcWILNVq8r1ZyFlVeamzEqtmsOg6bz/
6YsFAjwOgZVr0M7W/Tv2VF2BjRY/cGXUuiDsAVxzIcw+av5iGg24ACkPvqVr36Zr
wd6v+D+6uCKoAGxceLv8yameyugRAqRwzMTFRkc0qAcVDM8hHlrgJgOwjnj6p/RB
m+ayuqGo8Qq2HO3Dq46aIduIBgdXdbvCXDWmmobd0EhI4pEy4j5YR4bKibolkmmL
f61dhMp45eQnWWRTQ86I6F4x03MTRysfBwGAWg/hg46+EmG7lSE1InL9bGDp5Az9
FATP8wdonvKUJUztU8TTBWsYt33lU4SfBA3UQizmYzWVK3fOk+5CDo1Hpekg+p7L
nAtupcW8RIG+oM5HgkbCoLTOfAyb42GlsrSEz9tKixrk0MDz6iXcpV2EdJ1QPG21
aZ8f7hvj/9+D1jaT0w0OLOgkMV0LDc2B7sstPAUlFRzYlBX8TrUcfrCq6MQ0Bure
CBdbzZu5bGUsjpIB+WWcoA+G5FUI1Gz4sngVmiwmYhf7vo6ZTRPfz7TT35Ow/pa3
mEsMrAfb9IlYiWWIUpt2ZtGcxzAwOBmy7/olRY+nqDtu37w/0oPWGTgW/vB6NA5g
XJPNPcGSN7oc3UX79zz+/ENXgO0P8DZi6UFfmjaivkKMQXc69g5fuq/vxjhs/9t2
Qe+dmMCS9o6CdznJeEJ2/8sFtd8uw8jRl6UdCtsCOOeFMR6gKwTsmmUSszcc8gXy
gSsB59DjTfO1QApmUyZ60IQ0rgGFDZAtVK5oi01igUHiXIItQBnJ0P4jLyJd2qhN
YOdQb1p0iVcUPCWO60cgE56ZLOdrd+5gKxCPPYIRfZmeOtZpq4hL7bcotLefziZw
dyTy3F0IrBakZTVcEui+0yPktlA1YiS0K9StW6Usj1/lJ+RUIB3SaTwQqSdYoF6B
7h9rTuWexL7wu7bML8nh3FLLjXOlasWpX6l+AFrhEEqNqaMQI77PWq0EAmWqR9kE
ExW4oeGLGCDhuJ0av4wPSg0SX1yIoNlVI5jKNgXhVo1rHQ5dD35k4TfMOFNdmCzV
N9QGdwLB0FM2SZCRv4Pvsw2TK8VC2oMfN/GeBMx3L458YO/6mnA5dW8C+yXlCpdA
mL02IWJLvpQndcEonU00nv3qvqWvY9yntmC71AK1l10g6c9bS8NYvQ1ORvrmtQp2
Lw7cE6IOnyWEIVgAHWMu+ngjOIrnF3FYIcwA3FLTslW+Srhl6ie2EHoWZNZtbtn8
FB8ockmvbO858jh1gUCinWw5AXD2AlPtTqruKX77D4CcrUpr3k7lbCw96qyMEsXf
ZjMplXAou/mdWEwp55DbXEj2hramJKHGPUsyjXlo+aVK9m6chYYJ6q7oQf4QWFkE
2ziSYhShRWP7MTxMRHTn/Gx7wCcZs1yTz2LujVosEQpXZOZhjKTthloD8N8t/jWY
c1J+6Wj5RuXFHqRb+c3bc4cjAijjkPia/sVSv+22f31MgKRs3gPlXSEcdSqpe3wb
K8kg7Xxb3PNN2LVkB0xzlMm9kzUMAznuGxqCehoA0BSRl3VNwD6XZsFps1G65fz8
MUP5+qcqeK7j1xcuz/pHGKF/m29jZf6rFo+Hm/T7/PG/j2nbtuZqvef388zC6NxH
Fw6/HJf39JyKB9wqC8Q6TtwmZCvy39+daSDUPaovv0T0c1/5+vsryONg/yN57VSG
8HJqdLkoWCJraCVylVGhpLqey04Mt9VLoRCWUpmH9hHjd9eRPhC/7FvQnNU9j8Xh
bj94Pg7Q6ifSdJvK/3NtvcNPkK0Efzr4JPxBwRP4MXx8KMc0x2cMTw2bb6DgC8Eh
qWqipiMeBrRto7BKKD+bcfpivlhSp9v8HRfBPFyVBg74Ii4dVeDcNlyH9ehy9dEd
WiQhWKaxW9AwK5hE3HUX5wsR5xYoBZ4QKGLz9T8/FTihQuoLYhQKWm1cUB9o57BR
uqvpXEYLmAqGEqaDRnOO59Dt8g+AH82utV9g24Z5FLJF1SccL4iYf5J6PH1PEyFH
ptDRfK6FWLhEVgTSvHJpJVi+IHPMWQwjVcTX3MqARXf7NN10MLF0LKOC2/O2oDMW
Nz0w73YtechMFaKPyPXaPfbclmbtShfCIUlVNThpwWFoyzfzNxOG7N6j7HyIGDji
zAPpmbuo5oipvNP1WJWQAHJS1YD4sUcEVIMCrlkp4Hb4g6XNYrF9zPfwFYrtg/XF
vV15CE0X4NisEdVM2fPz6dmYNTWeAvmqc/FmRLtVrZy3XCSji8Okx1Tx5K0ThPLP
tmXOjUgkmBT6Sj05c3yPBZIEA6slG6r+S/sTwP7Vb1NPtoNqRscgryN2mhcezvnr
Bca3VE9TSVgApN+tCCl1WxBYwmVB/cgPCp9wkGxSlRyzahJEjJy35RQHgKN+61m2

`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
czCxWnvQXUraW3UGEVp7yNWmwK5g2icbaoxXR5bNyaqqQQexIDnearm5MAZG+pTHj4kObYFoOmYa
2ZNrnPWpVw1x39urGAGk1kpGHLubeQ89x41YjwXryootx1tkZEwYK6OQWMkuYp5sXuHM8ptXRU7R
VJUccLpEmS5c/VMdqxbXf/srFVd8zv26uFX8UG6vRQNj4fVtSCJBRdAaPZpxXyAtusHIupb//iuS
sjuKJq1xSFAP4oiNU4uRrTAgodqyi60p1B53X098e9/LY9rPAK6IdDpxd427LwepnJow28cGm/n6
RaRcWxAklBDtlRHwPkyBOv1RMUIWPUpBiD6klA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 14368)
YGda0VHMYNqHg6rxpHArn8TqyQpieRivv7lnr9wLRe9qagnscrerFSCNNqjRnt6DZZ2NQ3cCIIgw
zI74pwnSg3vD4PWv1U3L346Nri+OkJw0gSKdPZbH1xefd4o6BqETwxv33QzbQP3NUQzH2V9US1qq
D82tmObYFWat3vCeK61ws7jjeZOzvBIvZlwzh+gXTHJg9RsG7BB0E1EiiMpFbAK9NYz/ouhrInYb
H//pEwg2ViX5gnwupihYO101VSwzp39L2LQd3i62WxTmcFTp3/4gfhW1wNnAfhf6wogHIe7VSLN0
2QiWAXgWXrdahKn21RBqPi3oa8WrRMQ3KGdqliNFpm7k0T0EBZRdbUAhNTJyjZXRF24hFDtZhfqh
fU1cjC/gSv8ML6pzCD2a6cbjRvmiV/w50IimgoWrWsSq53p1GYPRITKpBioC9ktAfbhuVNCF++6W
OmYdvieRJ87jhcys+uwJIcqttAhRapmQwxGC8I9FO1wVgD3iZe4j6kZ7ROxt1qAJ2Rvw1dxcsv+l
R35i44kP8c07zTWiBErCAGvHsbQz6VqsTb8pKVyGQT5fgCAFOKv6NQ28EmgWzrGfHvLOZk6kY1wT
RQiJezCBR5DMIYWSR4Pzm091dgXipkXvgXlWYD/4cJcKD9pvSpKyHg2iLG8oVCVNeI9sowiprhgi
wSCWOSjkFc0SfY/smWfOgLwzCYI+WbtyCl6dhkSNqeJp3QNmguKj70qOv+cRaZl5OjrS3CBcGjdx
1L2p5J3lr+tzqtPd2vAu2u14BSc+hLj66EqO/rNQEQDTNl2GjVJHuG0uyMZX9fDycrpwp0G1+/gL
Q0OPU5a8cfrOjjuixrX8FvmvOBN87Z1I2I1+KhOXhP3/PR4/X0AG/sRJ5fEqVVUSd0xF4MrEFUt0
IYMrqtbaFqWUenJQZ4FbC8RNihMJmNOvYGOWJC+ZQ35LvwTJrAcuZ4xBPxc3N2j+g7l7ubvFe+Op
3AwE5ZmnzIWqZbMuSoEp2RNaPm0eP6epTiwnziKlvqaRrU78C5v2J+9YjUk89i2RNXISc96nvUyg
uwouLOv2MMEWp+5ai59irh0MWHtrSJYeo4ynksIv4nucUxVblpRNqF73U7hUDFvxoHA6eY3gcaGz
mkgEouJjLjbz8Rg2OI9lL8d8AXUtn3ZRm61tiR7LJVostU8CBvbfzBhO75IH0o8N+L2Jx3DbclSA
+pySIYqGHYr1y1LDpI9TdqKq1PBOjbiptXh/yd6MNWdzZ+Y6YrG7NVswLXOndMRb1vJWBhrvzGXs
djlQ+dy4Covz4GYOkF6uXb2JJ/iwXqkzVZmjBQoM+t1B2dH7QTg0ZPEuDYATXJcwfdh0r3sNZVHg
QcwLmy4Ncqiop641EK90tc+S0tcH5QMzl8czYQcO2tUzgZuzQv7IfX/pzWbcnfc0VZJSHH0PCkiU
rgHJSuE58fIAVcZGW4DZNK3uf0OptmvBdPuQgOOjeLOf7x0MohLIjNOLhIm4t8wriccvslsEYrL0
J11mZ3pR2GPF/qGaxKuR+B3BvjZLijnBlyGyYaE9fE3QhyhzcLoP42t/me7FV2KEPESGqPxAzxEP
2oFq2eWQMlofA6yGzs2oH0Gt/VSChkFKdBLKKPpqd6w3FR1Zu1HX326/uvGFznD06y88oyUFmTeC
+wffCWB30F21l/wCMuJszlqI75ADbAmz+//EVaNsjh5RhvPuY4KSS977UHKJO2pKk8DakLXDGbb8
MC+Yz2UJObL/OL8qUTyDRgLGhxI/6PSzwIyqiyrvsPBxZoS4jjARGpToAsBS5VhHJ55Qf5klCmlc
F8gKDY9RSpeEzwfdnrw+/w5irPf0N8IM++gpD1fcQrJ3T3TJUvYxNjXRkAk2TcmSSxfdRyUWeNL1
yLTEfWOl3D/9WW8+6k6FA+ge+Z2iRseQBFTty+EJoY8ElaxxR8x8oz9tK9mHIomRtidFt33jzxlz
8f6xiqJfGMd3VcTlxnqDQmkiHQiyBd2KiIRFz/4IsVmMrceYat0RCg/xfoUJYnANIiuNaXyuQE0/
jlaub+eC0BmzytGhzEL41XgB2VgHaSt5KtzsIaq4VXgOsYkbThTuURiCAlWNf9Pzbb4mg7T6/bQz
d8mgr0/8l/ykWnuyzak019umcCpYnVQe9Tp3F0zfMTsJW5gHvXbjHMEkm663JZBR7mRfjqnKYtI0
XPKX2N0+rNzZ1hSlZYUXhm+INwpAkamMlQ0cp7/jdWNT5vfbUUacBdBj3/RdX3K/JdeCvhDFD60L
XvDnIL5/69Rw0GXxFyMVzYEAgjPIlpUYQUhowxf1vApCJYY+wSX70fjc1fizSuShrpg7WGw18qBe
uM4L+RIL2WxYaakc0yelvykcIQ7OE+pDFmxl7KHox8K+BYHrY9VXHkVQPEHbg5KlUWzAJRlWPnAF
G8LnKtJc23PvSxzh2yqbMnC9KOBrKj4qIBmA1UYgAp3ZZjIvBdn00V+cPqWqdsXs5QO1KefuoskV
sqhnCp59m9QJur19jDLXmhXT4dNY2hs088ADfcbfkbV3qQ+H/vjYql7fM2to5ZDxQll62wB+a9QW
q1x0I5WWkg0LrZhSJDHsmJxFl0zSvyjd20sHkEDBORy24hxvLLzj+fHYTf/MpcyBz/dMAEGPyNkS
1FhHk5MpJZ1iIsiViTvHE54Fc8Inxv++p9qHxYenYCvK2FIGTycdqQU5NyJJ+57n+m6z3oT8xJ2z
UqskoQRk0+6mjYQAY0GOtv4zmU8Iweb1XPUOfuUh8EXwHv2+cKH1sDYO7UEbhYwzL7TCbOEVs9Ke
4D5SXlbM+Hbn/09tSCL/U6WMJXkNFOLJUHhMHM88QLWCd8aqAjtDzwmjR0+hLv0Z6fUwMWyRYZ5Q
nLqxMN9m3HC/ry2LZ2dC06Mgjb6xCtLwYEYzqpetmcBNqatSGwvArKNklQOBtsFAfGcUMcpzfpi7
P/bTRL8DRYO4BROUOyJHUM+SX52olutkbvmiK1PUu7UrqO4uOdqT6xTsw1bbgV8imXktB0Oq2ZJa
rY1Lk9Wj+3F8q9Bsvz8qPrqEaZG5iAvKEkKipUw/R6f1u5rJZlcPhlN2Fdn1m8uU+3gNucowmBA5
BAdPyGRNRmBuLzksJKwM8yFwumj/zeAqcsVMith6faEhuVlmn0PSs47uOQfB8ryMueJKFBlMrvql
hBvzhiQPqmSkI7O8gbPi1Zt3Pc865v1b2tHq857e9th3ftS2KW1EAnqrQ3GBDqW9hjV32m8adgkl
g+6o2asio04swb+jjDXg9Okc2NeL3DozJSg6wPbReBerF1NxNsXJQlMr806DuhTT9K+nT6ljQOYR
ZteSwYdGMc1FqHD8+tXOYEsTPvP2NGzmjpE8l0FSBj65jdC0XJ+NkpxqNh67np2mKDgB+qz0xAxd
Kq9nDPbeo1MkZYW/DYM7rbJEYnfjyALriLKL8WlVszZmeMD+WlL3T2NNmO12aU9uixEeWcC54zeY
xK12IWlXd5UPU5Yqpye0e6x32b/N4xvU3zCot+e9Q9BEIOam/krPMfc8wT84Yg37nSytLSKwz6LV
VUANIlEejvp0+qRLbzxoHsZcevtJJz/8Hm12MfdIrGqSYLeQQIRJFogmd9U9ShGNuIIe9GH4zsuC
PVCpoNI+HUC2/v6jIDZledMp0tmcRuqMSKKPWct/Fho2x+E2dpHWk5PUnAPT7vP2IFvhbIjpbGYM
DOsUUlapFuPaqjk/4XQseMDvJLFItgheR+uLsiZ9nVQeBB6zgT+G1TyJCq0pNFC/w0Sa+p/YZO5o
hXsoWXR5q8aiLy45QZJajgQSm68AFfqyEQG5U3u7Or0Y1YUWJh0DOjPwb6Spby94bRx0JSfB9eEp
FX/M4RC31MoYIKBzRiuUu1rcpHW/slZxwO21FiZ+MAD0fxykCCxot049W2ayWC4kvbbmLp6PHgUd
OYcZ3phXxa7hJMM7EXlU1LDvie4y8majgsHnLRFzPMFSIhT4KE+uUiK+cDU94hfJlaHfnYdXaph5
gqukbZzCi1Ji8btalcMv21hnNDf3lpu1cNG82CZG2NjxuOWWTjQsEw9G099DUAj3hsCHY59rdfN2
TXVN6/QGfo+oy/p6Om2PV9mPJFKIS7QDiGK+afTgi4JkirX7UyFYESUxsxP6/zl7evye9ya4vljn
6mA8Pb+BYaiYu7creMe5qYO0YS8GsDApII+X1rTP07WcKpp743emKb3hDB7+MUjzhoO1LxePZr8P
kkBm/wd2p+95zw8FYd4B+jtLeIRHISK3Rkm0lXDUcwVW/fu5WyCEGOLWR1zOWvez9X4UGbKVTGCA
6GoMd6W7GZZIthP23+el1Jmu3jLVCE2aGXV1crecUMkElSrIsHVG6CHAiEGn8+a9wWZWq8zwXwcy
NDHAdN0cTwHDDP3+dHc/fYNCPAD8runIWEQXg/4vLztbl2TrHPqj0KdMMAWEUGbHeHShwVPFlbP2
JfzeKq81XplqisvOTR1zF6eHWsSbuHpyRV/oh67+VPZBOfsq3Pg4Vwkrmx9ABF8aJZDJzSFFmrkx
8ehojpJoj1StkOkvjkPiVA4YSw6YBK1YbdnRuesDa3PLUUPoLhvm7+USBJJfisHxz7xW8CXwXysU
l/3fCuKZlDged7qJj8dWb15TMh++j7ECwH2DS9SUw2Csp65LsPG+eUb60sFKhHuy6jh9CLnnfMLH
HICAeOu3G9MCA3aCynksFdt21pxneo0MB9S+cVVuamsDdvrKGcWaUOZG7vhwSnAlPPcrD/LfeDcB
ny6hjLZLOb15e1bHak/aWVqlTQVAd9kALzcyvxC0bexhKDJ7ALMJ1l6JO3pN0bY1A4UbMBf7o21e
pGbyX5I0bWvGYN8BBJJLxLIRSeob/m1Sfu9MKhK7JevmxOyuMjX7c7VJU/3mCLJbn0SJdWeYQ/nV
ejTh0Jua0pv90Rag7mJoQ1Gxkcv7+QcZqpPN4vFxNA3bziJn3MRRpqvCI5SEXDHAhobkFbA0U8yr
OP9xkqqHnVTpLAdqbm8Mo4aaTlfqTMZb9Ou0Dq+NrpjCI1JMzUC8vc58zKQjdNnjOJncaIZ6kbGf
msb4tMeacDF5C0EPihrpeIN1/wbo+Xf5qSM9Dd3Dep8oi7LvJK+759uM/zDV2zin8Yi5ZJJrLhxd
g8bk8geSW3IEokjEGRsQKHSRaJe0sdXIb8TkbT8A+c1aDWIxgNuNvbKV28fefGhSSMVWXx1d/cWN
PnjHUbQ26ArCzlZvmftQPYmf5pC6i09lO88BOOW1idKbu48dw5A7gZ6GMcOTWdDMkfV9urYmZCIE
LIYJeiDZkNDgL3X5UP9Px+RTKT+8X68bd/zvhBgJbxJp1SduqrUh5E7hhvC5Xavg7FjI3XeNwEgb
CTcqE6Esbkihh/sJw4P5jcNqGzu9teMjZryaXh5xVQU0n6d6PGv7z/Vq2LhRpErK8bSRL+xerKxl
gtygC4LsxiWR3E8WnNyIsLD9xANViDrwnLotYqYq/ZSZHS6roxrIPeQ+DxI5gun0Lg6EGPz1+zLS
lf9jkkWahvbgsL5v4XP0ujqZVfUkqwR+5A6b0g7gUumLHhY7QzghMceHV1OzJoO+XDcC0QeCV8kz
sc2HYUJpsDG/9NgigLskQSu2xl+VT8ZLejhtGn6K3Aa5kgp1DsKJDJY1u8a0ur0FIhGeLgVh2up/
wORZ2PYdX2qHKAsPWhP7w3GnZGFzf7rS1G+LZX9NLuF+DZwf1GcCiwztBFJcEiiw96dz5F3UwDqp
B+WyjhSU7LZLJbC2kSfWNGn4nFCpwHkkHEZKNCg9eajHMdyqhc7/gsX0lFoZpHAipNfYK51UB0GT
LceiQejH0OsMR7sQdOgZX9srgD24dV8q9j4ET4dl3rjt/nLGBFWVLz4HLhSJ16K0NDIdrJ8LJ/DZ
58Kev8pMk4U41UB/hHJXsp3+yHMkd9Ph0DR+OTQiF8f9UPmdvt9DpwHY9+Xl9EO2vSRqiIMFNYFF
nmXGGQfF1cO+lHqErI4niryqTHXiSAvFxQro/LTl3ZMmhLf7H/DFjylKGtrdfts7fVrkB0h2CQm+
iZ1g1pRipSO02QasZLhH83H7wXXhf5cEIfaI/j85b9xZaSobz+rVN5BktUcNY6gZmXsMvsekFBZ0
Vjbb3KJQ+RtTRc1qSfzdGcvPcCHnGuxqARSH21OJrOwSa+9nV3sBBVCcXE95mIjFhLs6UKCRjiNc
AGf9DeT+LE6N7ZGHwnJj7brjhClExYfxfguk/Fm3mOJIX3Wg0Zs389LSr5lWxS40bQ/yWtdunvvF
76P8EKfJyjCv+iNn8Rcui8YgV9Zxf+2LX8Kria7O3E2PsGO8k3NSSu6O6Ez2SZenGWtpfaGNUQPe
5psIXmTDqXu45tbCXaQ/7O2Hboahm9dmrSdLwoHdKj/IkmkUdAbJT2Qe2kKZDe0TyF69JGazmEVp
qePU5tDwtDSf7n7pJ56XXWIhHIfWIzmWjWO7LASvCHaaXQLRJuJhlj1DB1FnJCtLiFc9tyhoRZJO
SaMZWZrObGB1ImFzYKss4didUPgjuzo1rxQ+ryHPFUsc8QIjXxtMJq5Gr+za3oq+0m3FYcMu6OU5
Lh3xfSRXpzLKf1unzZXBzRAQ2sfV3XlL6zsfR6+q4n1AdgQecJXhrPPUnRP6z+pridSC+dl2HIMU
Y+M1lJaNkPa80yjK1ISviogdEZi3PbPfUCk023HCuqUOEVpuAQwEX/1sZ3QgxmZ9Hs6RqPtLh+xN
26tq7C5HdNFiklE4RTo/KBL+TxCPE7kzzxNNlaBNlJ7wUcqppi0ZYwkNY0jx6WJxDHiim46ShLCB
7+lOm7Bolw3jRfMRXSZ6o7UwQhxKEVeoMep5EXmt87gzBgBdVHo741KVyn80Tf8750zCY3xeZ7dT
msEKCLZTDDXge/Sb3t8PQ8xQkkg1C3kU27SA7UlYAjY6k6Z1Fwfu3ULtUIgxBwish2MDAesx3kH6
+eWggNKcnIRcmiDpIMg3wBvj7zCbem8OB+lQWG1Xi8qsS51vjnPg7xnIsUF/HJjGsELwZL61DCN9
AwzfwGGN2WAdVpoj5LcKhNq9yDpDL6B1RH1ZlTUibUGK/Hh7IOTrk7d3zxgnj7vPu4q8skZ7aPZY
9CQ/h6roWutEt/ikun4liDO5aiT7QELWeV0a/MOo640OPww+6c1cgAJfazK4FwAyAuuJ9UzQZgv6
sTItg22TdVLrVr8slwHX4w3Ll9eNjtQbk204OjBrgyFh57EnCi+1CZ902DgMhPz1KPkE51H8Nd6A
n7+RqPq2aQ8+bp2pYCryHrSH3BWdNN7GKHoODnNOGp0mvjRTccIHKlPNLItPuCaHdDwzp9w2hSEQ
iSW7pXuii+9rX+/vmNP6r203ECWKE32v0MhwlHVat0/XMTK/bUIrVoTxmjcdl7vEkUIp9GgZRVVO
S9ocorma+JpxQ38VwIsilp6hL3bYUxJFyppClTf0ipRNFTxlJM9HftDrASKIVw43MW2Dz2Q3kMjA
ajCebUatuh+bmr0SPoMvLEjEIeVUTkAxcjobunnM2c4dxETXnPLAvSUjoIFE+7JOTgVwYExShGAc
TgXXnt502PpTjhdXFdOGE9swRm/Tb238E4og9BH0XDIZ5XvApuXSH7LyCV3jL/+dW/yAPSkMpA3M
N/x4p7AEw4xJjNFRWsMlTOfbYgfru9ZNxj/9TGuPWlZyEDDAUE7MVY9Cg/DgtMid1TbthCxKU7Ku
S0aQIxsC69LAGfRmBerttkV9bUIFYVm3MPoFTRmLXI+wmG0UGBk1gWCA8cUb9EoppQoC/CG0h+fl
D+1Cz4CgBs0zsyuz301KIxqkXon9h+5gfYSrvdwTdY8rRy4xlVckzTpOacBliTlikm7uUJlJ0chI
v0rdWbCb5YkW2NE6Y8Stjecm+99yK1il3qnQ75p/ie2omjvtJbM+vVfsWQ8a98l9b1bGNKYrCtIH
pZazQ31n1+lj04cQPbtc5UJORRq8OP+CWr3PWxEiJwJ02+RNHUeOnxR1wxEC5eY01fbcua9pzxqH
GXhKUP/HRlP4iP+TbRHiKGFcQxuGgBFGI7fJ84HMsyT3GgZcR3McZHokvEqjgoISJY9l4d0UIVea
J4UCnhTpYQVabvIJwKmR8pUI2xka2ocAvA0cm5Zd/xgWEaf/Ry3032pM0f6mCIHUefkwBGQevHNK
CCvRWQios9lLppZrrBEKarSO3yX6ZdiCQB+ipaPo/WY99iUrzHSJTKtiqfW6oaB08FRoD/DqKWN6
tFs0C4/EZjXqcrpd9lbK+7WEPGtv0jLYxpP5a3Ngo71QcpZQ00nTt3iwhzFS0OCI9akQpqua4qZs
9zah0uJtNyxR+gQh4GgFnK9S/4WkEoCJFPkGs0X830HhVm7v4miL//zxbGJxooe0b4aUXe3pm3A5
2y3GauKP/sYoUHdFF0vm1sMTlQvRu8AgBTiqeLcsIFg9sZzcZ5uj0+eQq3w8ZRm93ESEzICbq9Rf
IQnzIZYho/2RSaBiCX6CoCCTXRiAXC1JtyjM7Tms3ZViCpM/auFF2RDsCOCLZTg92kiFIb4h8xH0
fprjHqzpm/6FcNGhbrYtXQFxQYOOYhsKYjDQ0Q7eoqBuPCMn3Yw+YoEmbsInT9K0XxgKFRCVFKJs
Bqo7Yz04YNHlgX1SZQkpni6PjDbQaMtaVGiokZO/wcON25qtDo3/8/ScrbZiN/4IA6ylTKa5d5o+
53Jz8MAcd+L6pfc0C2w0juSKw/T3pIJGyTA+kO3iwVgP+lGJqZPcAw/DpH6DDI4sp9sSrxuREkKz
quhx9HMdjcsZEGKH3nCjE7G8pp7LBw3TD8ntgOUKreKW64L/P/cSDSLVvFhwJXf9zMIBEDz6ojw4
XkhsjRjOhKHo809klJl0pUFpPsqi8WqQIVcG1xBymABfoZVz0Qr0Ax0T4tuCI9XR1LsqY++u02XO
wMJ9+u0ZK9tKLvthwkPaHPqufSeDN38nw+jgg57rN1ZS41/Kq8QUHgWejBgH+zD6p055bEYOz06h
lHz9doG56ID46BeosoZDOiyydUM1bxhboQXuTHYlYiCZT7ikCM/Cus+49d2gUpqOiFXh/ZQqfsW2
bKSTb3JC20C65tKLxFxPXJskdbQ4x3a8yl62liyXc6h2X10uEpKSgZ2Y4VCa7c1IOIAUYHPcPUgn
7zqUlDDkTuXrn+1NmALHRkCeXA9ss6bRcnhow0QAXWkvqnoMJ1UULSIfQ7KpXq8s92K7nx0iISh1
RyPVTImEypTgeVCfABPF7f4tdTJrmadV+Y5KYpc5yT0HfX8uzlcgisjkBr1NvrwBaRuuL+o/OlmY
LcvSSuvEhfjgnxp+JSmp8jqiVCayZr40Gj70Kcy4RviIkWjajF+6X0olkyn3jl+9o6HgH2ZwWdgj
ANF+/UUi6SoGrm3JAV/7oUGK6hm6ZpWxXIzYK8cwSZslUS/yOYXoN6fzW4ZO8QibuNyvT3jJT9Fv
lOcm5/R7L+Z1KBXeZyOyK24zo/5F21RF5RDEyqjOjHkvRQty5nHsXubz+zaCUOrRnOahiOuqYlrX
NZ8Y4VNMPfld/If5NEaWqiSiLcsQPBLYS1ieluSq2123P2nKT2/sdByGpZvehxnwmzpCzHGMRprS
Kgpmp8cT2IbGTd151UHJ30pdNrE8gMn2IG0gtpzYJFPBYvda44lp0jh7d3HakD/fhpXxlwUqgsj5
J5P/e82/9pw5eJMDeyyCYgvSTmpmB3J5ZMM6K9rZ7PmZF694DgDHyfEXPOFH6O6/00FpwRM6YeO/
cJDnjkU9mh95SkeTaR5LegWfBhbFokf7l/INWhrwk/LKrwFTDYs3f0VEYN8x7yd54i8KGHM1YnyP
FvF5FSkEHVHPXQNjKb9weKIujPMcJDiOdpLlg8/lcVqypErwGvZUPHMNA/nbKoIaWQ3tRe9Cqw4Z
gwERkJFvpzBnXfksgcDdPka6YBqEVZg8RDDZSMECW1oi2Y6i/4M/kkEh+JTKMSWYIb9xpW6eOoQR
mEqydikFAo1bkS0qD46XzIiPi1sTJ/Ua2A3edN38b9mNIMoz4MYH9RlUdvjd5MRCVW9UPi+0Dcw2
3ptnzgb1C5Pe4CSL6K5msnJ5WwWn7RSpuMH0fKawxcOxbUB3+cdIiITxW66WIDJNsIHxHGiJom72
O72uHm3n6alVJlzsK0yzoyEXTRNLPwg7DtGpBuGS1QFYZPNHHUeC+xzShJHCcb/073PC9b7flFsC
iUJhIOR+bfZM5mcGlekcMUduxqeOUJ7zejENYW5TCyLCmI0P6JDggJX/au+uRxwLZmMCI1bvd2ol
GjjQw7hNVF5Ah+f3r97KUM4ssBEL06yXpPDxsqqfOkXxupqdeUmdcy7D4TNRB5xF0x4c2DbRedN8
4GFWZvxVuXzv8St8uCe8e/Z9UPTeiVcR+Dim+k4iW+6lS2XECn2ryQwxTo1jiBHfFO0k3NhrS4og
eK4hqUe9e5XgT4ppfk+QDGUAGJR+SckZQS8Q1qP5q8W/wRfnyh/5TZLfJoGGSfLbhsa4b2tcNYB2
u2Mo7NVZRPTRdZsfJ2Y42RfnMNsQQc8HOyeCtcvNnFl8O0oE3fYuP0gZNlAcrYEcistAQruDHshh
fF/TEN1K+J0UbUargCMsR0vF6hnFsG0/+1adg8XeL1ocf+4WQM3Haja6dOfAujKy12mpIlA+bBed
d9ypcRdq06XJJbG+J4v86UMufd6fBRYs1Nf053TjSJdqVExM5WKZiAfGZGf1/xcupRiqLYy6IttI
dXfWXpvpaLSp0b72lx4uxMfqg3BYbcv8HsD32iIkEukZuUgCJPKu3v8smQCN+TVhuW1b4WAyaSFL
D+31SgRylpGIP4kztKlYcILZjdsnlYQodC+4eM668q0I0aA2YDRxT8Rpod6IOdaQ0jJ7mfpkWGwT
G1HFwqT47WMykjHUUA0bLO+1ZVzj7I2tTxaUSImvtggGCCtGQQOxukQhhYj4t/3G/Sd4Ynj3ov0O
cZKjNpRjOXH45EaF8zcNwrAC+qFnCql0/OUEahxeHQxrlz9GCvOsbG6sRCSyZ83wovJuBJlb12jw
8Ngx28SdvWusCHVo3drAHSuJgLmD5P5/zIAPDLKo9Woc4vb3FJcaXjBHJhkYcEEIPTsMHvtdvJMC
gjGdGyIq8u2ZsjnIU/Pyi9zUwgULDWPzLtulHCv7Fy89OpMnnqlFeyLpHHtBP9wnqAUacly1CkgZ
BqnGO366ibJi5TodJjEJjmsNIiAVUVZJOtnCG/+JY5XnBz7ro+JwAVIB0y2N+M0lnUi4c4HXadGl
GtWBWTRNkMEUOKpV0Z9WyKgdBIuZWpEpBSSNoVEAqhYpZD3p5gQHWHhojT8fIjWaMSy3FkgZ+R/A
1E5AYY15fUvahnSsirC6R6tCvRIiye4I5WM7fHnuNgZBZ/wED7kjb9phwtb8CxfSnoFTVR/oTPCV
PGytdQsYH+QbVDejCPb5PwQ0JTFaA06gN/XbSfqWfly4cKLIda2+OPwHBZ+zGrYnObPAazKyUKj+
I7Pd0IT+NFO2Vw1xMrmX4I0bjdbJz3wcCmw7oMC8VGe6fqZpDtWV2lFm499Tjzkr7j1TJpdI9vuu
F/TgOAnHxmivV4EPw57vGN8OvaNnvsJ5LrdANJFIp+5fEHozOhpKvhTl1N86rdh8VGq6ZxblXmRv
ze3OSewMZ9ACkeimOGzj3jNXEw39F0dl4A1gtuC8gspdw1PV7e74SS1VRUmgG1DTRvZzyfmw1O5N
jcGPTA7bilKAilYOxlKoB5LzB9foGzutjK4JCC6A38rVZs6WwL2uDOsbuNHpGjgZ/vxjCcoK11C7
zuYOWTGyOdcD/97h9Eyl9C9bUgfZMCUtADhlr9H6uU3ZSvGBC3dr0UblQzSIcIWYNfy5AJdYaQjg
xA33SBFh0y50kiptVx48NhqS7i4UlHtOFCffPgUHEydbV3uDvwaTDfmSNZF6eNNrvBb7C5flAa8U
tSIjyr5v3d/pLK7F3dXF5wTUefXuIp65BMMbHzDlDW/yMBC8P/Z1N15bEkBjkKTNoF3dvtUNAwft
ZOMbg9CaaCXQrWzHw/rjL6dhgHfM3zW3Z9B/9LZF9v3BDiBNnD92tw4Q2E6s4W4r2I+jO83Polm4
HV7fYIWSBctgvBVejjd/JzIHCmrOm7aljoO3HGyzsBpfHzQiC+Tw4vI5+T6/JuhPNydwIdm5frpe
28k3XobtuUdenNPLGuw0c56REhMQBqlvcIHJSpa/RghVbbyRXGLXQwmCY3RlnXPMMqKmqFYvcGLz
GaQc5C1dmukxE5ppZBSaFGV8DkQGOg8lF1pXW7rXL+Pz/luMk7V2y7Uoa792D0zG5r6pL83VqmLv
imueGZx7vocykip8l8bZee/hB0qUA2KoNdSuG8357CNlM4fu50HP6dZkIIWHDWdy9qV4E0W4/9cK
m8Oy5RVySs8NNsCFSPEIfmRfO1w0g6S05jogdcCdUF5f3Uicg6SdeTFxefoqgsjNG5H0yNHsiwmo
W2Db5ZZt+xeTx2fegx7v8c7OwxCxkE+2ECfj/d/C4jWVskjM+N4rVAZtB6odAJgR8pRXdnGhTOP1
ONg5O56qft2hOxvgwaFEKpCuKcf0pj3lXQqt0LeiWHhhn+Dq3ns8K7/FNCA4wBhmFrt1FvT1ZqtF
4wYcTfDs30cK8A4vG2BzMEOclvAViSj7SVXjZgiMmwkhUIgMLCj2tFx42LNSOd955D29Am8tlHoW
mosLkce8g3+Frj8S+35EIjzK5HpdzaxQxmXHJuOmEfnPuwzIr2TkL8COKXAiMDqzWRZ7LXT2M2WP
yTclRXV3a3Htv3/IrtZj1HZs3EEazzp6OB8r1g0F8tBd2cZIQwpiTqFj+wXiiTLoahn/pSnz76gH
zTGvZQPwYGEVp02gWIE6IV7zBr+4ZwtSqCOpefr4odravPry+sry/dUOJuXLpbxZ2+4X7zvQOt+Q
R194JT4s35RVSAUOsozP/xVFl8EbXWg3eb7Vi14/S5seywUbbBQTdW82Z7Kt4Ysj8n9lKWvARqlD
fhioLx8t5KFP6xX2e9WhLGdPlTncXLH492yFW4AioP9dGOAtt0rS4UggOpot5k3TyiiQWWdM9tIk
JRySVSkb63O87YFlCuDgU4NhLq5o+V9sE+mS9btT1kQF9craZaQCAJL8qhioKIGjzMmTlFq0hstH
J+8e8KqKlISDvgVRMLDDzfnopJySYc5OfZ2tYfARlLVPXh87qBDq/XW63fwsyJjv7ZxeJWKlQqDR
iv0RwoWR7UmFqnnBY3fTUe0NdLFn0cMhaGXYlGcAi85IJ4zAL43TBtJZkmOljOmQZoOxw96CEpmS
OF4T5sMsa0hlpdB33dwDmSZhUqOwWlRb8G92QqJ/KihUZYyOK2hlVZ94U07oVz9X3qgVa7RSe4ka
Rzq9lVqZNQOnLSoLgPgG4seOxrY6XYrMvgopuXsodWTvkqPdD20ektl4EFsshwf6pa3sMIRcMSUX
b/d/l9f7MTVz9rteJRBVRqT2tZ1C2luCnJLQdkQ1G2i5X2HvgkiTB+QrSoViulxxlnBGHAUa9xKA
SIBewCtG77Ht+kDILBIatgtKunF9sykEdLqqfa09wchB1KZ78ojjlHI2fwNBdLYFwQrM4twUCDpt
CwrVKUV006QwOmclBh1amUkQaZU8z0PB2WNqwEERQT3QLLwx1Cy1+eCsXf+F78qtvL4ac7x9GlXe
ZnsqZVTlzcM+uCBrTX1OsEeM4hvPFxqNETADfTFJ4cHYbFIT3/8P84EuRw8vTS9PZooWzkHomb1Y
NBM54DQLm6kxkaam6JWLTI4+ge4J73WYPubJkhA62EW5Td2+E8W6LFOKFSHm1eKXk7ijRv1Z2ykg
mxj4UpX+OE5toz828J1oLODOa7jx5/JmIkQsDIVMauWcjyA4eWhJOUHFqQgMYuWGTVhOj/6wMK3B
l01oWfP861UcMFF8h/Fm+O/JgG6j3/1MUw0LvB9R9snOJpvd5lX3mDsuahSmzBKkXhj1v/GPpxYZ
Q0yzLxgeXuBah/iS7AgeJeetnPYqV3TtVr4eDw9a10mRTHJA1YrzaSqrqZaKEzOxqxI0gwGwDgcK
MOvIX1idAdwKwpf/KQPwSzhwnqCyrCjDw8lmOuuIAEImraJyfFmWHxMXcSK+cktyxs4ESsGf2c7F
psLjdv6CnX/OtpVFcCAwjf5Wfi/5fCNX16WwsDWY8YgKHss35q1QtqHGp/ppyILXSvNH6Ew7y/YQ
dRXm5Vql+BNrRAqwweLhT1W1eoxf6ubeD9n1ZsRew0YcDBLV8HgJnaf7qSmETuQjhn76gwmCeLgM
GrXyhN3mYkSXe6SNIDB9V7GKd1ewYQapGN/znM6ASBsvc8Btfgq3RamMpR4+l2YF9TCicfxPkbPy
gBTB05e9LVOIGVhLG7jSzlH9m7Xmd2YYNAKw1I9x5ElJUUv/cSSK/C/bibJaAHZx2h6oydgS0ewN
LKZsjuy2M+96IPM0BzolOBm/7Sm5C+m6W1kYuzlIjXaWFz1j/uwOnjGpRGvbxDVHuszUoOkUJlF6
tQU2LRs4Bbhkiag2P/M74kdnscMi52pZ8yx30MdL9q/orLQeFURF5Pgc2t7jKRkDWI1PRN5YE9Ck
EcNF0/RIq32Zh62sLE6y1APdC+CGpEwpNlqNXL/dIRK80V3Ki+4eqaxQRh+T+G8w5Rb+tNcSKplL
ApX+IunSZn+s9+Q0j9UN8aI8XEJrbiFBCh2bou+iW4So0RUj87CIx7ScRBRzpNCcDDADg0XE+JpT
AubdyO0lL0TaLZ+Wl3ZA7b35JiB9m78FKnUZtUMT0M2GWvRjnXV6mPD9s8zZAUho1Kg9Dx3yttaj
x2rznHFG04bwjV8I19RMTOLtsR99VKSkp9Jring5q8FGu/XUj5b1pi8ycXwCG5+DjemiyxqLWEDI
6w/qbr3ijZDErbZ8IGR2DgxQpdtNvsQBDMkcLYreC9xQ50OwpJvORboE+6wxZKtyKfT5rQcZBF07
JcMQjN4TXquNHPCxKVi5Un+q3S1ETAHfWFx9GzpBi49qr3w/T31JL+x51hx8QGTrgbghIDFcHW/m
Vu/r5ChOHtFhYq3Z6PL1Ijk9qVNPeuKE3Gh8qGuIH77geMWuwO1JtXC3si9FZWGF+x59J7fjlN4E
GIHpCiL/xeZxfOEubXgYDvEWNQbn5Qw+P++WJonuo1C9gVna00q4QTt5FmMDATnVSsnzeraiMVBa
gvbxXqo07OIGwlT/kehDKPKb6iAuOad5PgjMTLccE47EdbQBXDHC/12YJ1b221zR4Y9CVsWRBPx5
ct0HR/D8eCw1jOdcO6hajzkZD7tych2lJ2W3PSw1mMicNsdhS7Vz3lp39527hxfQilJi3I2uepz1
A2IdI9LoJsst7bFwdibpoJuclcbl2QvGxpnMN0YMdnhT3Kxj2gzhfwHuTNiQI0WICrkSQqsczgOx
9eldnQ1U14ThbYEAL4/fQlKyYnhaqp5F2Xet3W7so7rfBLCguLFgDuSNDkx5xP94Zk9Vfw7j+irb
/x5Dpxyw9M2JBWi2GKtXufs1+mVO1e9laevzMbaF99rw/kTvwuM4WkLPKxn81uTiInKUNW2fhLVi
XM36y16GTON567rmPlPkJz87RHkn3HVm8G9vIlF0ll1TJ8Sfk2Y78o/UHrmnqXMp+59qUGjCK8Zj
WpL5W8rVUdpfKOm/IDmMeTr6BilR4usK1NSZ59x26qOL5lgpU28ghF1+pny6nJY5lk3i0x2/Ynml
beUfWp+Wzmwa4xQBMXYUmWTdQVAVX6a2HtoAmASOgHEpHRtP2PhxuHCRhpKgHrIUJZi3crO6MtnA
sJzxVkSsQq9WtsiIJcwa88767E23jadpEncN743QaEskNHL31rPtSSwQml2QUyhvGnubiYiXAbif
jVsHAcBahujSrVF8oSsHClU2va1SQm+2jMp9SqqvW9z0y8FFiSFLueZrYy75w9Q0oRpmvbiplXYP
yR9XeSsv+kSWAe4Re8480uAOt+Ikxys+b3v5wVrNdovoY5xitLgeFrdyeliSDWjGYDNspvmldv+h
8EZiH0wFelgQ0RB5qbre+dX8fd5raKV2YSypNdalg1maDXD9SnDv3jm1LY6KjTJeqbr4gwjbseSH
EbZhjljvUoPykHoDgi9dKI5PTY08XSLPOBNgNegiaUKH7PkeeWcquMe0d6uIO7/3wR3gtRK8wRAx
4tZRdG24Rb6jXQQ8DWunbwK92dFHHKtkmJBnu6gAmlWJViIFYGvZ6YoG1KBGcnM3NfeLYy+sqLRp
820PQ5W9hrnFE0mccdePynukVoZ1+XzclALqFxebZ2Xv+V2NKCE5dfJdk/Sop+9FMOelZLjmK1SH
NQ1KsCUPl9EFMdnTC0+LwwJi9W3vNatbOwzi1DrgjiHIlBp6wk8606+WvZ4FxnOKXOuMKvuEUqNe
gRqekdYZk2omp5Md+9ilNot7x2I81cSRanKq8pGH/B3HNZwlguwXoPMGv1K8zVDrLIPPSBCd30p4
95R0Y5+JeWqWkdoBMjp+HQM2wbRSheLRe46Km+v++NCuecBAAgHALrsHZVPZOvDj9FPVGhKk2TUt
06TmRqZpFKercikYBvicCj9jCtoZGk71ZYz0dMLjIdP9fO0kipcGo2LixV72fVGLFJ08r8cb3ELJ
PaHmidByTZ8+YHsjStxAp4HXPCBXpt1lVYioWsk2YJX7MDwEClcgenr9LacwaQsEDaU8CPoz59lv
AN02KEMI8s+ENw96c/Qmqnqbsbry/8SPAHJGsBIh+jIY4R5KuBQQqhL41ktODJc+hvnnb/3n6QNE
YEGGjsPL3KxNH0sxtuDwWtOmvzUIP4XFd050gxFXS1nc0XHVjS+7+18SX5aDAsRv0L+PRHZX9ABr
yAZ/selPjm1REhoPl8JaOAh8K2JD20E7jGhdx0vH3yy/awsUfSjV04tpgGZFElE09BfmQbiea4Kr
bn3XHmi+rqWMEyAzt+gSErgCAqhen7W2NoyCZz+0LFd8UmUGf0b8VYBZCZtFQO5CcuMDS3SShbsZ
tBj5APFa1cMXIShNWFBrGxJMyYQRqIXgvwT42KZZYoC7G51ygcJ2BRNDmeszd3pY6C41MjxRNWLU
ndoD3YVmFyV4eJ1QnDhuEZ2f55sSKYetMWM8S25uJQbMwLNDALSWz0zu4EgKnmw4FDoZJ4hKVoar
MPTiPG4q/bUt5YnCsVn3RCwMcQussFJp3fmGDbOK3DG3+f5vB1vjbbqEp/aDoYL4tw1GmydH/YDM
PxXnHb3wJOqur3JP2wgTs/v3yQA9YPh+pWGc11espX3Dtzf36I+JlB5DpC5Ms1nhTcTbzL38Dgpo
B+RWjzMk5UJ61G22UTbS5PrEw9+MfH3zAtdw2xuedkeBg0v1CN/NImet2+pTNNXXxbZEI4JEfC3W
hLQxuLGUF/H8xWJQD08c56WSirfY+jO0Kq21SzzzcVSJfBFqvGJeFCqob8/lVBwHhZlTAaz78kiJ
mGO/F48TadQbPpRYOghtWECtUbsK1VQrU1c08EpIEuYvl/1WG40g+QQQbsP5IV78JQFacpCfIoGl
v/9mlevvFLAvzZBGtls6jOcBul1H0ybOccEAyxOiuvy/adoDuiWO1m+X7+Ok24NPDjoVulGcu2Ax
+GmEoWNDOLOLgQu46DrlLYyX/BDwttvUF/RwJ1kbVKUJl4JX84t/zq57ZPTCj0nitkr8WPe6wvwT
02ftGufgwlleTZIPmfy4vw7NJCI8+H10Ibc3x4Qu7m3crRrJwSh2MP/G9l972i2/px7HMcQm4ECr
yse8kLZaMxiTpLCaOj8BE4bGC1BsTn1OIqNe4ikFznGcKO3qsXI+zPkThXRP/mx7G5yFEUlRdBBI
7G3DtyxZyfDJyydvYmQOJIhd5XcsW0+AqJot0/IzJUk0qXx0vHeQ1PxZmIEwF8iW1wK4OzS6/Gdn
RX7yG0f7Rm7mlczW8zF36dXZ8zRTBflpqE23AV86G9rzwH+pEtS09OjtPSP5nLu4yRAIz2XfrrSF
uzcPwYPneeJU5f+PH0aq4zo+dkrFRGtharRR+etFOUc03LGkupviNxcmxxwViGM08eAqrGh5bcpX
rSps+BiKMmU4de5a3XyDH7W2K0uhW+JtMWpIPgElvNqe80WC9IDS046SdgqlDkqyR6yuI+6M74MA
/t6Fv0gNYTtjxp3kESLSSsRCanKj6QpCuYgb0dl1gBQIkhXU6pZ/O96l6daPWtT49thU9udc8x9s
WbsXTS1sHl+d06NJhtJcpj2KhJy46pn9CETSICHGML+g/L5dmFu/Wv8uHVsX+Pu/ih/vCrwW21Tj
ru+OdDwmasms6SzZ4jzJpsHNZtHqNg037BLg5jk3Mgdc7uGlqk1rV1BPfKjIDyWM/nKthkoyYq7+
hgXWon0yc+FTdZEMuy1noFB5uI7bJh+1YOcfNWcp6+FuhuNpqvgr1hGDr7BdFgM0h0N393G4ofFH
kvrUzD5UHmgnh+17zZdlCkNqyE2h04j6ztIfDSQxDZfTPGMkXrL37FNIWIkfSGrI/kgh7xxdF8JM
XQay/bXGcGugRHt4jhF+KrgLJj8KJQf+7IZJLhLMXThfWLTd4nIZB4XScxMf5AkrIYSkduCMnLlK
Gi2SG2AruzhV7DeITv0Ec6iwaMLvlQQC6vW//+LtYZSyejaoLdxyl/Fyb/Psh3BSQFAaGuxEvJA4
K4SRMzxWTjwrs0RnRff4RTxV3j0PI1lFa9yQ69LUNZpttTKb7UDg53MNsKVwLwvWg/czi004btpg
LNe4wiRo9vEEyzfrtCMFGJKxaEqF5WSsW0P91O7Lrkj+KG/MPqzpzUH8Jq3mL5Fc2G2/UPq3uiQu
dk4ho01V8udGSrjGeCRRv0XhIwbXZz7igyM3VVJRGtqhuV81emXIBsh5sgkJDuyqwKCu/JQA+8m1
sjyb9mzkJyR5VOfp06tn+XuU9sPpVN74kJs/Pff5AK9mAQp4Aeag2uHzQGwPHODwsnT71TwUvSfv
uVMc93GsCa1bBv2zBn+AN+qBtaPHpuPlZNYICL/B75nsVkIcBjWflU/tgAfe8iPYw8tkcwoz9FSL
3Zdgtw==
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
kJ6mkUqji7dHfLRMsHQ/c1/hzz2Qpnr2kfwGyMt4GY7iVbhqxMEqlqLhQ7Y7urob
0Tcl5jXN/b/BejP39dJF+qqHvOi1DrfaKd5kMbGVS9uf0+ur35No319qbbrKL2pI
vQTxDly/E4dS0kur65XJFTBeyEtGWIgofCmWmNJ8ZYE=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 15456 )
`pragma protect data_block
kFjfDObD+GW7cxJSLXh84sVHJOAknSPUzqJTrfCmIQSdqhvt7OMT8oR0LBYDkTMi
bHt6ndsDQlqY9uCfEMYKAd+5p0mV0uQkF6a3wmPp0ggRDYwjPxAjIyu3tOyD7H45
5FxZuw2NGTw24XHdAQe19TMkyYo09D0AjX5EMkpuaea7J58z8CUTwj5SkAFFZzmL
5KX1l84j3jckvJaFAwFHvnKKZbiVwegsWkOO0DwcwQmpL9viu8/56rRqJcbYZEIe
YW+U5MkOMvxA7dGMXBySS4gef6ggMG7tegmIjz5nAZnMKQ+RsMCj2x3Vd1aSkGUU
QKv4G5lHf6C4Iik+AMuR/ebuip6kXCvejGmgb2tOq5oKyyTKoT8xAJoN/D6V6TF2
+VtdBVJ8GvVK7/DNGilqJCp+xA36cAjjrwWg4p99lmvpSG+x4M15mFbygiRiB2ez
cuFuGPjye91/BPNaRoR0dDjUVPdpm+nCluInoxl3btz32GC12DR2bEvNUNXRJH/6
YqcZjtjxwgcnUFbXmtCxeDbQQPINxxYdOn35SoA4Kaapp2FtiFuM4PNweDSB7Ng3
oD2UgOjHhlbJMDUnjaLMv7Im6MDi9P/d8cXk8eguy009T8OIuQwNYFvKtQuzM9Zk
LoKdu/pyrHaHWBEsrSY/OUVzlnbNAAv0m2JD7UfxL6KxORfBOgIkykLXzoJbCGJe
vSjmlf6xehtGz7jtLmrG3V+aY5SeojR2THwbHr6Ow6arQgvTXHSudVHScQLg4a+D
ISHEfdEhaUfrenQuCZEHEqbTl2QQW+BXpUAxxiLEMc+7dlAjmDAzziqqJwPd6ISk
CqNiamhfzcGEbO6/psmnsS40Icl5tyf/cXID0AmF4vqt09dWjt9f3uDce37XZTa3
sjz4E968CKaOh2PfzKMY2E5MyKSc8v+tyHCWoxp7LwX1U71llwSW1y5KofIya1Hr
0C8Dr2Icwcuuamq8x9bHeebTSoWART1b1EzqMJ8COElcS0fj2JKynlK3cyw5zOBw
5GGfzwkCIdDjGEJ0EDNVygXCdl842s2KcL4zXIynZWiTTctviZQaFj/731Z/Y57x
jtTYOtR0SkJseAd2esEhggTuT1a92vWbjSbMHKBOZ14+HFK89irbY3jr6ivO8Cos
AuS4JWYRLiZy86lbVlForQEEJa6yrEAPid+FiJEQjD70JHzCqbWY1Aj63OFGpcB/
hiYeuNP8v6SMPMr4Tyv8zMLGRg8/lfkQ9Ro9dPlFlIGvdHxSXjZjioxMuDzmG+Lq
K2TQJJUXan23utbgJuhP0ouxbT7RGWHNyK1jtiZgnBvn0Z4A9nHnMpZ9cVHXLnrx
qqZVSn5J03HlaH9Tzkgr0Pc9yd3gPKm0BiQ4YWGag8JG1mEQ4VaGvV71OiSFcm5h
e+Vn5cJuNANKg1oUrP/JL2r+a91XEz9oyk2HaS7M5mVXIncetIuroKJVYPKWkeIi
5CBfd2vYXg5sid+Sqn7VFam0uYs6LwgbsK1OO5JCupglbxEd0SMg+iVzm6LNrxyo
GYCrGUCpQ8hzSiqdyj25NcDEwmQmVfyyXQtd2LzbZywVExJBr7oLtWscjJDqiQk+
mPRcevzoRs4/MMUxqvtMit61wTI26/Lj3VDs824pCeq4WcAaJCx7SdJo2OGXSGVM
yPFirRAjcmeL2+ip8j+AJ2St/0sdaQMCgAo0GAvbpMDn4Q6Uh2WvwXbqZWzvEP4+
Ug2RIFcatROEAO6MKk4KIfqnbJ42TIa7Z0nwv6c2HKf15G3yq4Wi7jYdWhkMmtws
P9UaNYvf2KDZWe+gl1axi6A8XViorGOnGc/0MSBn34cgwS/9wOP5hLEREteeAQdP
Cxo2KsreqwDW5K5OaN9R3NFeIzICPVbrFB3Pt5ub8R9cPPTB/5Zm9HieX5p1Ssgw
0ob5fvPPCQ+NYBQInrf5Kio/p8kgDFUkiHWWNTMdFKdeY3tGFfXBdis/hKFF9ipa
7Y6+mDO/387eqCN3ghw1ruiC3q/6vzZmAMYQOTpFaz1Xx5KMGInUdu4SeWK5LWD1
BbjZSsF9Sxbd90JTVI0pWK5JmytEnimtclaTaNIugUhmpkK646ZUWOpo1tqswFsJ
CWeM8XXgRVvpOgpqKz1TYzCmTKZwZJpDh76OFCC0J0S3T+9oAoTo0jR06IQhuSKm
g+jw/TSHllojaETMxF31kXh1OjUnttXhaNUXrqhqEiA7q27gTYiCu8rmf4Av7SEZ
xYXWK2YmQGCc5BdMAo6SN5RL5eb5oFKRU2V0xnWZf9SqFUjJpUrJQz1VqaRKfhQa
RZ0VG8nM8sp/B2z/EpRb+9aiWiOX0hAn2/AT+cbjuo3mT0i4IErONiWF8X7l4o8Q
6U+m4PocTDOhUNxDHs1y4mhhbZCrMQ54QAViIxVPQ6QxMCBgMTGXTbJ0uHGDRnPF
HYBlpTF+kKXPQ5cyZbNFBf4AuwyGcFSI7C9Rath8oTnKpw5U5NhmTBYnYldi7Qm6
OVDPw2Je0BDjmpavzPouLZhG3ziSa+dl9JuFKmP3kkGf2N8LEiFWgjhoLgUHyUn8
VrAll0XyMM2vth+oBAT7SB7uLGiWUH0mJ0Ssl0Xlr/Sk3/RfcEJi1VAksHB7vkiX
0Skw7MemNtwNtPaObjYzkckAbuZTpo5ost7/zimI6HZkCHD/i8bkuRzNo8wXsqZ0
8Lg5OB3cPJG8Wqv2G/X7pvO1RXFl4+2Qm35lLHM3Oq1f0b0cGQLN/9OuLwxFIHB/
YZHW1UR8OzDhdQcdUmYBxgC/P3QHbR2/3AUvwe/QLF1pcqyJ0YNkZjLOXJnHC65X
p1IdJ+C+J7hAw6KJdI0DyuUxKzY/Ay2a9xhbFxas9HLlad0mulu+NHUb3T89BknT
5czFZTZz+7ZHbbc5J+uND2CSsL9ADeLWFvzpKG6anZB/GCI3QEHrzuQmOYo38AFa
h50IroRJFR6EyeUobChDwkFvveRmyZygJDTNrnnDG+R+t7PEqYbhNmvPXMfjR+EF
xNIZ8B0s3x0wZAZJ2SJiA2UmCH6atgjHP0N4OLIvZu69VZYn0cD7eyRI2juPwDtv
hHOGUQKJk0Z348P+XvGj28OwV4eyHTeBJnTI7tBy4eeSqxijVosM4NwjBvJiHLHy
60QAFadkrT+bsooa1AUWf80QEn+2ExP7M8LgmCYu+mr6kF+UfKoeNXD+MGs8hJT3
jUUZAOKbvAn7oyDRylz3FBZZFE1K4OyBI9lJEH7KLu0k1rrlXP+otmhSU4s3LjMj
7hgdDSAEGiewkOWoGx0uYezEX69cQvsUGWlyOSOCSJ8m2P4hCUthwUcYs0yFuwBN
nzAMu2uns+r/xAF9lcJDzzUG1q0BP3svHvvg57ECv+kbIQfZTWEnIgOXLw1lzua7
fI7yANCYbsGoLeusdFJf5QodrGqKSF4uU9+0jqUFB03vWOlFfVGKZ5unV+MLj05P
ym67rhW9Bxe4/xVSXlbT63V4jV4epQdNMjw87H6OnkSDYk8wyk9QQ3m4MQOS38KE
KbVFngDN+irBHKHosedqsj6qIWlehFvKlDpq2arc2++U3W2DdeQofDI7lbo0n5/8
Lp4KR+UZhBqogFe76h4fAt49XktDQDM7wATBhzXd5WfyNqbd9Tqq2RJg2TgAI+g3
N1vE3IH3hSgtJFJD0x28r8Bn/6npL+RxxPvnl28UtgUMXAa288Y8BUAIEwIiLZZc
mQqKMtfc4qh3Apq7avES7N4uwFz7m6laUHqc+wAjDdJstI5SmACcMo8/sC8+6HfW
qvDENKPtVk7DdbUO5eUIv1068DaoMVBsl4kX0NkSKjRhQCaPBuJEEEQUU/7WMxLS
GsRQeZCyGIzYIfz9x1N/6nD+C02oOsXHxdC2jw9XRqrz4+yzrxQU9K6MvVppDfGE
fVVw9OMWAqKG/TTo2hX2U0iceGpFOWWLk+Tw1YKKdV8raJe3u/vwWAKinNzo/IDv
Ek1zYibGz6FoWIYyYIk5/BazGjBaKgY/3Bf7c8BxD7VuTy461oADpf7yTjry+itC
wfzAg3R1DBmvwMeSNbynS8JiH6XTe5xAYUBTJBWsIqn3WzkKP31EuC28zmXJ44Wj
Z7JQsgRzADw6qyHBZOLfVl9lX0+DefBfjbJkWdXdQSf3dvgJb+WYBiHeB6ucrH5w
m37vk+n5g1kfeO1YHuszcsq9pcWz75HMEtN5y+D1LeoJtraToUrvTKqMBxkkPoIw
3ihRZjl2Z8oDVx0bPiaIV9jtJzrHSoSmcCjSRiMMp4YBdS5vYXZrtXqu9jET5EJd
EPF0r3Z4rzLZ6WC3l5nl4qGD+OHFcrmd6QsCJM/qaVUkjdRI5Pma1KmloLtSsxb0
Hr/SNGTkUvz+/euG14zu2gOeJuysv/d0ci/RIGkPSKp+rTFljwvcQjPJXrfHhlHH
gYqjiDUxb1iJWtGJ9eE2cTx7M1mUwubMajGxcX4/6XCem36Wmirc3GY8pNWoD39t
RjFUsaWQ8ieBRDeptanZufqagq9NFgNn7UsjdBZg9jrFfJ2DhBWfODveOd+/G1bV
itDDd0lCTEYkoexuXwX6buun8H8NhUL8RXz8GBS8Au2nAlhomhvRpVefra35Sdfm
bFZwPsG8w5hgfH0kGuK/OxICXcJ2Le6+pTQDTm5b1Fghw8FxmcN0xbeL59H2Wmx+
18dfLelj9s33teuyZiLok1uiC6yK85gu5FjA0WrzC/EM/+Bhw8orULayMpZpMPJi
jIkYRCd57kAXaEfewKsh4uFI1FHge6MEPZ2b1qnCCotPsqfqoihntXOmpMU//Ow6
IfoXH2z9SsUqFy4CC6RmhbYPFY9rlYuFifv6gOoA4Hm2lOpLxhXKJi7e/4IUTAIc
1GTriNhXcsxA6vE9zCQpR5ttzVqPouz16jBeqhTkQtNVoRIunFvUtl6VOwPlEIQY
0GSbYukZuqxv6T2y1dtbSAexroRXIWPksh2RTxYgAf9oWdEZMz9EcZRdOoWUB0Uq
9uiHpMaxEq6UMV6avtB0GFvaIrcqiX5jLKEaaXUrC+yCGggx8CAsC49GiYSy80mQ
aFv9+eYLAgY3aQOQvmPlogGP6oMpJcDLkKZm9fNv9m/4pgV2T8GgvGUCyJEUF8gM
KevEbAVJz6K3kBNqW14SOep6YaUXFRb0KjmLIM9+rH9LFvcbtH/Gw4fRCsK/ktPi
t70cx7TJhytxs76dgahmo20e32y7HsbJuweQPu6Q+gowo6lV0kCDqf7KkvAXqKFT
ZibbW3pE6lnt+Yjb9Be0Ac3lAhHnvCmOiBmOEvCPXSVANmRcd6gRHrUmyMckwkL/
Qd1hwi73YygXZWj0xlp9NA9gHffLTDCtuTxuDQiIhnPLTUSs5E6aeLSKoek/qfX9
Cq80/S/BQ24cNeulHviO191NRrEw4lJx7GtKdy8zWEjUXlMURCVZ+rjIDi8AkogI
IutNmCpgk/5WM5Vf6aKCwTQzLfYA4XZ7JQRPpXUuER2CGVqNUqEkNOT758W78IO1
umVV0tGgDha52vCPm9ZqsSyucXr6AhParKE6UyXtiMbWnZUIKHmgTOEgb+fxOCUb
/iPiyfNkPehIIl4g/3ZtW/fM/oVwtLGa1DhZZZr+MReO+UnPmEZh/ga7LVrEQYk4
yBj3xeyKLF5hudtRYOIVT6sXHfAJjvfUWLKPbfHPe8TuODMeEBsi61FKYBAYHogs
/o/lkQRMeCG7OlFPr3+jq2yrJ0kND/FCJa43BH8fwjBMul0F8xPRRs9gujig/7rC
Vle3MGjtfb+Cg3HIJ3JrFC7QY1rVERZFoRyqatP4B7qjXy0XlnFEoXqIEUQZZlwc
W8eiVMRAof91aebqzORqqAps3I/R/v+jzKx6a9eyUNRf/ErJ19qJeKKP0vOPwc3D
0UcJpcCrfMaETu5ZsW47WnL7MPp/M7lR6udltqnJT15b9Q1EI5ijw6IaibTk/LE5
p+Mbs5l14hOD3VugXGSu3IvGWlMh0K9Bhm+IyYipC+EV1oi7BGOFgW9XBcdndK5N
peAMavHe+tU1hEW3+d4FhJ24KAb1tZLRhboiZnmshy55/skdhvMk2QWPqp+lgUbJ
+8JlYzlNYxo8LTCgUtWpId6rehL279mahrRmpCOJGmx0xE5+NdDYwafCAyIgGZVV
8sE7diVQx90Ts2StRTjprvvA/36qKdSLBRWFLs60GZwMrRAqZcLDUE/fz3IftEZc
U3ZbYJx6s5jMVe+imkBng7pl8DLgaC3KAvglpeB+aWvBDpyJdjyyf5vL/nKLsg+S
KTwhBMeY1KxJ2YrEMRhPJijC6oFCF5azwNHo0wtHmomTFQrLYlviJFZNG7FOiE0f
Oi8I1ZQtyGPUXyoyEOrernBjQNgUWYzSmKxQZza9bndTDpGazi97aPpfZTGFnXmL
eVv7MQACfL9iq/ZWPRwGXMI4JQG1rjr5Xs1aIn0FqUKnhh7J57+w4Wze8OL8+DHW
QRkKDaKvN6Qg74txiLIJ7kFQVLTk3VBeISlP4romEoCwEqc9UtNU2bvzUeKqKHR/
dhxsZKQa63pmW4H/R3Yk5dKr+uoTvLmdkY65Wkq1eprHxkjz6qzyjL2KuAniW06L
Icv8j81CQ32qybLf/mselmnu/3uMeR/KN/iCnkTC+taClI0aANXjEncgb3dkLYnQ
VcTDDzVvXB+kIxcyVtVEm5DDH9rwMiFvAdM7HiivQg6O9CbTq4DQ5jDiL09bsAIT
efU0XVz9LAYgQ2FK59+/Co0Nwi8cjRceE4ZoWAFBer/JkqKl/trrnZjy+SaFVMSt
YZBNs/22gAub/m2zqBnXtqsACjzDBNGFjm9gZ79xDMA+hycByON9yZC3l+jIu4Rk
ho6EHNfiklibD8LnIR6wHSFOA/1U/dJ+4W0k3fUnvzTpv6ZN6g1POvP9Pau+K9Qj
W3fR60vU8eZk82pLyqCMJz4F6LFy+FtB1WrPuDKwX/9/nGevNDnrPyCdKnYd1rCn
e33nlrdGespRXcg9AvJkWx/bXxXiNYsTvMwTq9pSjX6yzofWYmm+b8L7q0IdKzY5
pE3nxuI0/gieQSVz/PUNJNIH8bomcfjPu3L/eCzaEEGmdekfHF5Tk4MUsBiF5pqX
+XV6d9kOe6u4uklaN3pbO1XPwIUrILsspspSZIFoUNOuRiqeV518KahxVss4lLFr
XLZXEkUcD3hBdc7NwM+FPvGR3pfXEAxqrF9WRgt03BxKioYWo3KcqXMqFGmQ7OeX
saZWS45eZ+uOkWLAOXRx/zkqNf26K5XQqVWXAyAmClZLf4UYksXaL2h0LUW6oiF7
wUHRFXFLwjK9wYVu3Fq+qbdTTf2LPA4BOBX6KO4n98Y/Wbks8xck9dY9TZVzdzUF
MAHIcX/2N7H4uZe7OQ2Pd0tSP34hvQjr9wgG+VF1KaAMLc+7EFqdn40L0TnZh1D5
FkdSfT+eb2R+0jI2ApJm+pOAVM4ixwEhplsO1vMGNPkahRq2GSyy7PDaaMywo/xt
1RGawul51z4eEh4XUBLjqEhpJfTPFt6mroNFrfZ5ggSwiq7j1q1yFRrvkBoORPav
9aihFJ+tk+4aLkk+rGOGpIvSRM0y36pHw14fhM9tcr10A8BcWwHEAMQxvbEy9Dun
ZMCFDBTssZXNzFVGoh9REUpG8Q2XcMnmt502WOPFFM1sPPKUW/cVOu9QWEOMGkDo
PG2CkX1HnuPWwZEm0HKdEfHOU7Cn/I8B3QPGzYUTAhSgsr6CKZE6UoBuZxu48e3v
WtDA79BFskgJ2AfzXKt2jqzy+l3rLjPoEqVNX1bQMnj8OEIF/6NVNlR3Kv5weCuS
q6CMQbVR+cf1f0VdeGpX8/7TnkalpI1zg6BpU+va+C2nxgyqGz+LmvrqQ5XhlXCG
pdcw1+DM3QAufc2DmvrRUCUm8xENCGxbS4c/sS7TnaeCzdsnURBPipSfhzVVib/G
w17YqvKBtgSTgnujUOx84H10qkc9VNq1VodCcHmkSjrXaLQ/mZtZK8+U0tn3002z
uUIEr8CFVudPsMvRdMYR1b0xGEKmuIkMuDuqP/aeKAkRNc7o6ULTaSM5Fwt8XnxH
f8y+oyIV7Mr3evw0rUrtuZM04xdzn+1FHFdMkJ3Pb0m+qDMNWetBVobAl4SZQoY4
4H+1cFKWfONV+gNNlfwGsTF4gkGbjc0SKzICAhn0i6ZECZChNki+XaaICGS70L2J
slZWToxJ8JisssGgtIoiAIyBjYnmAXwmCWiyUYYSoe49/m1MdjaZAObyufILJygf
S3hsb36aJ5+dBgyudzwUAdWtVM7adpV59mEIEL8COZMAjuW5mfM+1LK5BraUqb08
G0EwH6nv0pUhSrCEadO+Lg7KJxMgFxT0ArCOnSk0EydYHimkzcsvhcIS10/Mt83k
hamPp+RcU7dtT/bK1wlL7gLGTHpQLoE6lf3RvfH2IR3NHzVfBdMDxjlTDFcoQvPU
pYgLT81MAIQWc+wDNNIWUBEgpcSwDvq1p3VskqMBqywZmyE764RdICkP/OKu6hqT
HdFhfC/xv1RLCmrGanyQ4eJDp8kAaliE7TDspDeOqm+qVAt2NwmL2m4dKxder7S5
8kBtwzaNwrQYqiSQHcfPm45pW/wuBoOMs8qfcUTjYazw2fS88JfRLOzGIymiKLJR
Bh082fH1SeLtOGb5zZjY0p29j2cws8NVjEQpHN7HeaYhAgMoK2cwCoFiIeQuuYmL
ArFrSVAeu24ACKdq7gf7RMjgeWJsm2U5z6YbNNhQE9MsGKUbNIexeZl8ruQB1QoM
fYuyq9B4SRCbpsKUwUr3Xwuy2cMH+Rz5PZQANQuBRE27oH1ze+JAuJSMRQT8G3mg
PYmhr1Y4vWzrflyeyH8AF4tNZIv2XIikbtN5vS3TfUZ3WnQk05Ommw7u574Go36x
f4gRFdyDkq0HUtdCZFpSZ6ZI7OWFcb5SDSZnhKQfYcGnLxaHEwuxsc3F2ePiLxrP
ZJ2/NA/PD+oab/egEuWxvhc8JhvALHlpB/Y2Ky+AUoaUnmGcPCscrikrpD+hi6Pz
cRFSQeIi+prVjda/VMxt3tMbpQ60TAiRiUf1pwlMtmFaiBLkQt57qxv/EsbCUbIl
wWawgJ185POFjQ8yjzlVYQUuZKzY+ISoO1O0upbhrpcJbAZjrHFDafoGt5TuQNI9
EVEs/xphRZCL4gk2XTwz+v8dCwjNfW1tH1Hp0nywxWl8MH1tXW5J7Kl0dPwdhsDG
guaxHFcQBB2QaTotPlEMDkZOb5XFM3a8++tqyKIy+4kW/i8UiVXu7yo9r7YfTPQx
nkFfv3QsWlVooW+b58qNn+7wV526a8rZ7xRw8IRB+X1pInMTW1Hanh8xUHqb0QDH
rbIikSJwQLySCixc6rC8EDR5zcaiKgewpzULJAMRGyqXrzvwu1sHd3X5olNcE2PW
7qHVBSKCyaEWK2FxUPc87wCfyUPLtyDQ9XhE+6EFTrFM9ROAj10ZAKUcDGiFpJS0
rCFWUDO7r1IimZV3oetXfKalG4WN6o/3RvR7kSkHaf11taWeY73YVtMGMsYXPVTN
IEONXUbfF7dhIFBhieK43IsuhnYj2s30rtazXecVm+oQMZAUUIWDwu8d87W3Zjg2
/SFR5q7uCtrmoiKkockqK6/ipPm3SaLTVmat52vre103XnL/m5G5J1Fz38qGQkML
ssHKyIykj9jJR17X7lq7OyetEHYR00V8SaYEwGeoqniePIq35jZfBTHuMnxM0WXJ
ddwdzHdqXaDojUj520c23Gxh+lAeZWIiw3XOH5vKNruI0CCtWLTD4wVCFuDO2tL7
HipK/GKdPh0VxzhmdNbx6ir6MjRzH9X6mCntEFq2TWB8k6xPv4SGS50hB230TWCr
9020r2errWAPCuUjoWFNxnNcRcdj5YEANfYcL6LIi2A5BLQVnLMGnpSuiPItWJkm
huFJ4HF5UsM7pl462ayEdRRJxedLJHvFkbtaQZi3bFdjO2nQ/+TAlG1EG+8sd0rP
/3UWjBhtZB9AJ5hcwHsViMReyZFSXZGPT09APxKw//9unAjTnXr9beCjS8Q15ddk
qUHHd29O947YuOH8+dX3X8TDiQmbAS78V2QgIp7gO/lY095NKo7QFu2Xr0VatPj/
XSh9I2xl+TELpYkVf3Hze/N1gMC+h+wkiNiw3dTFz2+0NC8JWBzSvY0H7hBh47Xu
CfVtHh+2tIRZ9AAI0bDjOqpRCI6ZD8FfmivLZ00gxZ8Ut8P/AfYtTbkkfDImsMBn
8jO9HBeI+iTdwKntacrjG9uOgb21vccYsCS7hCGhvWsPv6Ju+V4eOJZwMhZ+7YRT
BWZUHkI3GRf8nRUTqFpRXV1v0TYSDlsrUCQvxCWe4HDQUGxIWGM6XAK3BJUTuQAf
YQ1tAZihipkLuBsaFgqvK8kx96nayYCGFwYzobOomIxII3UMeJ5JFiXsLE0hXYD2
rI2at+f8M3Z0M/vDJc2z374wLjLXpSNye35sN8VKIYtP8nU1PpJ2eM7BjPudtrog
Fvcbb7yO2/DRXKdEy6zhGWHlGcjCt0R9pW6+UXqY96YbsH25rvnc/nTMv77J3seS
OUH0s4Ki2/tZIPOegP/D/rnjuUR+u3YW5eM7ZoCTZ0hb4gytacCktLFyN85N+MpJ
zM5qHEU5zWWHIAvFsUDs2MHvYrRFAlMp5YL/lpOvRLb1E+aUm4TeScElMcPdSFDm
vRthcNCveuwZQeXkRlJoA7qPosLHjdQqT1TAUJnLuojSOJkoP+6gzgz7bVa3mCt2
j1MQNCRiD7TzOa1RXItzvV37tvDdAJpQC2lsr0gxoaaEYR7TT4OK0j6SYxi4j4tL
4lyYV+YbDlkgTZWkgz6WJrYsUq0FRnUG/+RJQlUeIXsIO9Su1jzW2rp1BvcEm6ea
O9h86sFBUjDj2riXT9tkGy4fxMDIVg5mEl7j6Z9R9/TmwTZnRGKQk+ZVbu5c5PBS
7ZxwQlzHERY6xXH+kT7fiGdmy8AncEzKk2oln8Anmonw37M1eFbQuhLzPx7CA3tz
/2uMvzk3+uTgU+qdgtf/wJcomp5N5Mp7ftO+40Inx3qpCbkgGvrJbkDQpzaL9doT
kyM8Q6LoXK5eAS4T6hV923gdJ1x1Gi0jaLiZb0L2r5VjzodHo0fM16OF2ONsM4cN
nW8soIwRmQTfYAspQUIFijJ5fVEIFTCz0jWY4vMpj2hqg/rAMOZGyVaERaz9l5Vc
agnJstESL6QLv4tOWAXMtuPUoifQ1GXmQgqja4t9YcuzZfN7NSWgZMfdWS7kXU2v
19pbVY+TmMz374/2gyMpVpvS8ZLcOxv07npn6fv5y+a4aTNFGjekphOTQgYKhWdb
9af4yUFToE4ZLvU4EDab8cD/vgJvAaDJlCI03AG7J+35NvMLOR6FKAz1NW8B7Bin
4uQxxlVmm+VuPhAElhff7fJInkUaYbHO32YpYV3tPeDIY13Z5BGBBdgP6ZUyVGMT
eTmNdPMRvgOSA6f53QdCNN+ttgBhxzsNexY4Mj0DWaNv8CSwwPt/gtGivdkR+Een
ddLJMBkmsj35GTB1Pcagb1XxpibAgIdgZcd2eXrx2sCleq1qQMMh/ZNX9qN0jEeu
TBjuLPYuWwKHnVPQ0Eze8nU2NUa7Z8rbAXopn5rC3uUB4z2FDQP+bnjg3VKay2+I
yZnoRFBy3tCOEqEKkesZbMLrjtSYgvaUY74RSQZmzHbz+Azm4O+twOYfyKO+YwXl
uwbFXL6egbMrURZU+Piv6coV1rG6SCRae1raHfaTuW14S11WMVciUwT1f2SqzPtv
VqTVtKr8g0Rb6q34LkCl6B+4IS2ctjxqO6xNwoCFVNItPaqNkTGaYdUttjkTrYzk
pyXWBQUy0tZuC/bm+uX3sKcVdJQIy9r1EkSv3wK/iZVyYk4ZmXGKu790jhFEcnt2
pXvUiwPYf3E/b7gMm7OrzhfbJqk/JQLQfXJaRJrGwK31d9cwyCvp6/jaFVCpYJgX
hanAsHQArlZV2dIK+pK+30CZX+lfgpU5lQpU0/TpQb2kv+mcBMWAtCO8qkwxSH+t
fwBPO5JhZ7w/ygonVdj7PTfy4Ir84HQ0M9USrjnk1c4I2UcGkT4KazF9QpoixKL/
/rUES0fLu4SzBcSZaziqJ2vccxFuUQNgofSwS0AandrNB9HVVemIAHWiqiUVXnQW
pFD2BGd9+KwHPq0/zg9L+C5ADdfXQfATTeub9pTcxbPwNu6Il+s0Zdcc1/rBFg7I
NcueZCS2aRHkkZ0qaZQyPhInPwFMAoD5lJF1i3GzLTt8ippvtSu1FHu5z7wykjlZ
tetnUKXr7aaW7UrCpwDehJrPIFCiZdWbhiM6RSfZmZqIwUBAmQIuVsRGOtRkVBO6
pNo5jqgcCjiYNt0w9OQn+xgCI7qZr1me+5UKoBLQ4Mg+fYe2p3Ob3/Zps0swNaaq
fZmQ5otLlcZK1mPmIKORzPDjSKRhRMZanV7R076z9JvcNRwZkGfhxrhnpXJzabew
uOK0kD6fGe4tu4uTLWIgkMCLLV5lwfjDPX5MVV5qb49JMYSmO0TGrPgMQSCeYMwL
ro2rL1k7IkZMfoXwiymCUG0WxxSQRv/02LuHwDaDn3kFw0+jkEB1ryJSyc2B21wG
Mpx7da+3bp8rSNPQdY32tGqLUCyMfhEaDk+XhVC8aUZrLCiYA5vPaOlHiaNo+mot
3PUv0fJ2YJFjeczPy5+XUXqcOroA2dIbLJBtFZ1S3rJHQLRCoKSd+p8aJwGRg+Zk
o7IRZVbhArZLkSPrMXZvHjc3NrkxN5m2TP0Gxd2VgiLbSxhUOZT3fryix17feg5g
5P2uQToGBd34KDODXJ6FkbC9WzUbN1O/I4PiViQtNV+3frs5Hqauv0XKHkldlRAq
fvXnJkQndGtW+BRGvWfcegXtrqvRbWbwtWaEsesanUCIJVPnTYMYi8PaHIRO89Ki
4KmLNfFWiqu4IqzJM5C9HdhqB8d3v3KQmXmohGQjQkPT6Dmw31I3ra4aPx4xwrsM
+TMrielS22Wu9YnGjlD9UgQEmhF/eDWQgtWmoYzFlQoHup4dj529Uw1IJvt+FPh1
f/fwtiIPGnKnnU6ntAbiNxBrZWcLUbeEzkNHLOuDAdhs5u7rs9EKmFDjRlNy2DLv
mC3/naiioinBAC9Ulfn8R2OaCcc6LELWe9Xg8NkvFk/HrrXoH58xL2/KF+9GqhGm
EVBuhOuLjHcW349DSFYCNSPdsMqukO2utJAEmzvvnkuPuzLjJYFWGBeqrDHkVpeh
gbC9d5PxIqAS6m7u7XIQ0bA8JPc/Vqg+gAP5Ybwg172wp9sY1PWAgYYRhEbOlL3B
68GRMjFLvPPnCfaiZb3RvxoGctR+y5uFfvjpdByORmJrV3grys4txSlDJPlbcAPi
Dedu9Wlyu/nLPEF9N6ERc2tn2yCsOGt0/l7Wz4Z1fwW4v5NbxVLtnbRlrWMKP6Kg
dwT+8ASzl2LVZWBrOAzhWqr6UXGW3nndiRdcE40WCy/ouwdlnd8spaHzdhkBgZny
wc+idS87dqiX/Rf3YWNSK+JL8jrBnygg/481uf0A+BkOfXlrNOiiyBU0XonkJwIA
kBWsledmubLmj3qKkW1psO9TL/oWp60tTZA2ZA/AKFhuj7CBa7ZYmvhpTFK3XBtg
sh9TP081vzDEggWn1ls2+eD00yL7F2/N3HUBtLOoFP2qJ9EzjPcLJC/TX/2bKfKm
1V08UjBhhizO29UBSLIF0AuxVIdZ+ra0XZ4Tjku+1NLLzfOxq3kU9nzX7QGcom3g
1Br7ZFXjXSZWf54bChDf1JqA30yOYeryOlTXsuW9xZ9Csuk4oM/nmOflt+jaJbMc
yceiaVeB4kaEObAOTD8Y6595IrAzgVwkeCwoN9Krf4ZaFGinM9IzdsCYFaPwFd4I
haEiNiDIQOQPfvAL1VYnZRvBRC5Pac//iYzgfLfWvRgNtSYaBDBD0dQUEwf3dQIs
JeYvjt0oW7z+Ds3lbzrk2YP8ZSVH9CR0225OPSjpU2+luhN3HGmPdDNE3Cphh+yr
pPVxuOoxmGRgrdSN6VBgtbbjnk+b8wvcFYOqAFbsfM3g3Zc+IK/GHnW/SZVAG6MC
izV+FNSAvO94y+OhK+68yfnF1w3EONjfK7EI6A69GTw5hS/9xksPp3H49/VTqj2i
1/EyLsApH+yYIfR9iIEKB/JTbbzh+e3Axt50VXRiALBn4cLuI2QWRrxljXdQ1OUY
f4zH66JQBzU630nfUjk+cGCdZGJ8wTqL91VzO3LChkfLFAjpeaWvxLuIwleYwZV1
VnOpldxdJP13Yr+xgYyHzzxvx+T92575rQ/qLfI+Jb4A/UtxVPeuFxD676WPGOQD
xQtQn0uAiRFEEyxFdmZLDmPNGWiyJvl481M3DGDpD8FcHnG2j1HWT5uR64Alf4d5
qLYEzod4iOMds/Kni8NpEKdWgQzPeM0YGHW3jwMzWt+16ut3XNkKCnUpApINrkQU
gYXiWMTjSDgM8ujBl1fWn903epd5aVVX4MssASFvVBvKEMK+4t4G0YgUEla3oX30
lhaiQR2ftm68r1lmrgQigeADARKCIbTzznaXut1s75lhjoFPretWXpik8TocndFl
xLKc3NJXqx4Rdu67xOSC9lMf8qsq2pXOARijn8vKi20ontEcc/yxIEhEO/IwLre0
qnYp63JDBXRqgBfsPdHY6rRfSuIVsJCXw+p70F7wizqXDbsIPBROJxvwXdL/1bEa
BFrKatJjsZp3N930CsqcWJ67rB51i1/sGdQlnaJ8iPKkaj7da06pnNY3uT//3t+l
Jlgjpz1eLGCh0B1jV/MU80XQBlsQ4STkVBtsQ7xUo+nShmOPmyJe4jZW4ir9Wf4L
k4Be1muoO0gmCIO4VOf00fr+rxXfh4y6YnwM4DfSgcCAkGmGR7eNb59kl2RTVaof
cnK/50QRCEp+Ej64iW2oIxmD9xVBibCNoOZxznS9JXqTE9USGM22aGkwKsbXsa6S
a+WUay9TM5qvqX7VupRg2Cm/8KMqTmUFiTXZ3v6cshVBWCL1LxY3EiQbfzCciFvR
B74iRu507YRpDX+fzJzn8xaZb59DHSWdFqn32RiSkVAKInux4b7bgtIlVx6zg+gy
F5KNF4X7Q2nXgGXws/kWm1Y7wOk9c6EMAckaxf6K7ytqa+ciONi++EIvyVuFwXaq
ag2+iSlInhddQP7gotx2QSUmjra/leM60tQibQS5cY1bQK7CRqJ09jH0OXixFpGL
Gfw+mIuJOjtm6PTlvjgjsTCqX13SehowDaiFCNPF+adG66ostx8ZgY6OpiZ5kSXD
lc1WLi6Ct8feH39XAtbFRKc5hplGAq4mbncYVj1a6o91IcQjVZMXFx/TWULsRAea
3gi1R0G8BhXFSCzwVSZH/Z+yH7ZhzTtC+gCSfPLyaQ7zHtbClHYg2q/BPGMBThTK
ODtclkg2qxZ6K1feR4YIZCgLhZqNVq1+DtfZXO/vWIirdszqve/Z/cBNdgQhgAiC
GV7VvKZHuMzkpL7nG584OWhwiw23hzMuom5DU2NK/FCtvaiyy4R09OOdZwagGYwx
pPe4kWJMeybq5QL1TGoGGdjQf2/1oGCHODN0vIWqGl0hgaRYcUvhX7ICkPMZSpUL
R8ORpQ2B9Ky+MOA8358HHTmG+vjJ8e5xQ9qArfvfugFdCYFDZI3p8m2VMsEaiQ/2
qZVje5TUhOoCjrOwq1MzTvnB2GLlV7wRPruSA4kzob5pfCgW48/x8Dlx3SUGUKP3
B3EsNtyagdgayjH8clP2lW/mKtIcTVnsqdUaBj/V9318ChJDyVZnJl/andhbaNY3
7XtuErGlfXqMnLmFnjaJ2erSQR4gQvaTiDlqD7gST8ta5EE9a8F4X+O684zZM2NB
fAw9qfY8BXYmh8gxwCb4g3msg2kZABDIznF6EhJkeUYeK3eTVsLBXRg2zQZp8VM7
dLLpBesN+xqx1DOap82Vr5g8KsAFRBUTHMBt4FqGn7RZ6+aY44osJhA5k2QFHYsz
q8Q/Atdl4EMbFXL3RmSuKYj+Ve2+Hvkruu4+uwkufdVxjFqHIxGXo20ayYf+9WIl
HqSJfCIsxmnEDj4B8K1M0XrOOh2k1qehbV83MTMTadIsV7XtPLWzhAx1/dtFcOfp
N/4mfUIBZYEBlOk+N/NNfoBbFSRQ1yDYtgH8iqa7i04QmrhNXSJF8cfEYRRSf7a0
iyzerujoCWXJDtNRm1hQjbQlIWvfRVHCHj0e8AbA66eSuDW2jzCTt1MHqFrWnMqw
62xgweWW9jxsSn6sruhQ8TXR1hyqKUrPlUEjuShLNYyg45bMnb4mWi4muyZiG+fW
5JkG3ZUmelk5xgX04F4vbxAlTh+WGGgRTnJLo1Fib87SbX7eOoQvA5l2Yv0CLH69
0FePzhzG3+Gn9Ahyj8BM6HWQvqcB5ylniB4gmft6xB3JpELhv5xSoHXNpLxX9fOJ
x27Qa/uxfCm3OmCkXtaaMg508qqLujAp89lNAFt3VQ8mmfYDU05OmD8Lt/eNZK3m
bzPgPXnkKpZvdDA+DByE6NNpc0FTL86dcpuo1ruhKFeEbEbm9kQtVjgjDAQzTqz+
MAqVJ/gOT+yAjwuIOZn6861UApTtNr8hf6PTOR7ee7aPaTlnhETuNlgXfFEF2To9
iztMEKj8lnaRubDV22zNuku2lfJtrUmpDKm4Fl9LDGpJRjnxKfOCnHvRidZWKBRK
MoohdbRAqHA3ho2OmyMg+KLsgjuwqWOij4P9NLa4r0jP2Ji3QNYWQIN6/jEzwjAv
Tc59n2+lOOVTicjt2DKWHBHpYo6J59fTcZ54SDis2l83tqorcwWVLgSffl/nvcIQ
NHLIWb0hFG0W1WTHSEnAmU5Yb8eRK6NJejE4WneSRMIS6er/L14f7fVQ17PzbV/v
CHIlXvVD3clZHRWLN3FJqbC8HCPOdeAGXjePu9eDQrtH3Q88zuX+OGprM883UI17
Jq4OiKQi16XvwBd5kihyCfuwGkAAoKAxtz/6V2yi0dGvU7/tfcv4ADCiw6139wEk
yoVek5FzLN9gzQTNzRcn7RzsUB1ts4tK1PQ277+csbRGqp1vpd+Vc3foHflqCfI1
GXhoz7e26EunAo3fmUdx+PcYJLG6pCsNW87fJeIJDCa/8Wh9wnNk0GCf7XQY5qQr
1CJE/6bRT91EV1HmGcvM3bkflhu4PHmPgtjUO3Zvfs5tJu6XK3QabmVT2X97wbPU
t9kYu9VqDntpcbcUzLc7PS2SgzjngZR2GAdq3xcpHBZq8Yd2pY8OzGcwvLgfLpgB
Ziz1qNe1X9ZFwt85Jv3ZFqqP89kseL8Dv5cAsb/AIfHxOBPQTeEhFHqVVi6JJemk
gJHSfAcs/sQq5ZG768MaDnpEvEp7HpFoKpgQIe0wdWCJqHT214/GvZxX1zvyw9cy
sujr47Kzm1Xhqvk7VvMugSAckQi+uKAiut7b+ktwFBXaHsGMcNmeG/HUBSb9piDc
eV8a46igEu/L1n8uDwF/gbj/vQp6wBLceacTeK6FWXd2zkadKrAs1pQAewOARXo3
lolKG3YKcyRqu65A+gItwhduFX9/I7rhOCEmQu6LKWTUqO+NQJHVgTr5GJdgGi/R
MeAG65UqY35gUgDsDIe9eJ7l6jPWXSrdz9wLQyLsG0KzJSHyAtXa1RrMLu28C9lv
4lJsBmmdg+Hhb45lD3TYrDqitdBI1UhS8ol1lK5TG3vimbcZiSvHCS8/9KhnR9nK
ZouDXLLQRI6NSjZROm2BsItamd00IDEatDxtO067cSWgK8QaQX9+9d1Wewwa4Phu
Qpi2QfUWeGcKBlOImXq7NaFAxdciHNhAITKygh6WATQO73wDt1OJpjaFllV3ICuY
kmz61RiWUqz66/JyA986+FhiJUDVilIGEp5ZpDx9xPPxcFPov7ek+yk65XcQ/hDB
sANVwTyfCjl/dO+GJDK6TQLI8UpAelQCnWIevcEKtidKKVWEnT5wjcw+c+Xi1Wkh
LwBFKUKYfbGxpj1X0RzgLk6kzrJ2t6Y6jF0tAz6sK0AbzDMrsT5O9eIKfgEUSw7O
vxeO2hmpRhc1poSmizZNUUZ+cB51tcdqztP5v1x/6UjQ4hxZSUWa9z3d6dk1U1uc
7BTY08MX6gotesWvAPEyNh+3tN5TfFyevDrP48qvuQuijf5LLn62tGJUjGYTBcF4
VifYAN8XAxsqVgGmkP2cwwtMhCD/SJ2YJ9NbjIWkeYPCo3LwVRSV3cxT5Ct5DUzl
rQkBHlojivrDSHAeoK1amDK21mU+1FML/qr2PUlpS2Dq/MuyUPKN/mBYTxXqHlxo
nxjyNjA5+pr5h68B/8lz3LgBdEwcVYF67AaIzCQcczw6us6MoK/VvivNB/yuDmG+
B73l/Yf9OXYyRL6sWeSzW9wby24PYs8hs0hMl7j0KBogo8R5uYQD/8ao9FNQ1jd0
xKBz2sMFjyX5AoD9JDNV1z3tzKvOUTwcKPw3wo9ASHBqtFO36VqKmhyiBjcmVMtL
1+L1wBeGk6TZNw+YmnUSF9GswV50/o0aeS+s+lgVHVz5d7K3tcgUIpyWtIvecco5
czlwiuE7jLIzWuwCYItYlkufVmSiK7y2YpCDtkBIICBu8awSeiz9UGTjwXTMlrzh
IxI1KcI2mByLrnkMyHbyZ8tDS6rljc5NfKbaUIcNogUG9XR1/sXFD7BTNPm3SoJT
LLDCDS4y9bZSFWJgo36EdwkvN3FN/+GXzTePcnwCmylbUSz/53gl4FaV7XrwH4nv
YYLpseHbFv9iayAIXTypQitLHXhDO4lwwEmZ6MzblhKdbQrY9p3I1GBtjoRXYQqQ
c1pOc4VJk0wvyqmK2JjDkGzOeHmnjv99zGzEYq+GMmDVay0Xhp9XimmJqsg6gmh8
qGiwQ62zhm3swFVKy5FIGuzXn+E8Z5puJBOl++dc10q1MGYkoryGnFqypeyP7CNa
bqPBd8AD7caEsnimIK++YywNvfI3KUgb4ZTU+Pyls3hST0Y/wu/qWr8Y6dBwkuCP
Qj8AEX7pcEgDaZeo5smb0QTI4/JxdESUWJfVIjWlT7Avg4g7KITYUHu7NpjuoJOf
Mn5GCAaTfsr9s+vu0ud1A5YkIqaTZcr2jLNcPkemOCjeC8uc78qWbjHAtMmvadPK
HJQYvRHAd2pCPu7Evb0ZhVIQGdJThcgo39jPDbooj9I4eXikRSzTYnqX6aHWDE/I
0Odc5k/OHcrv5Vzu0u43kntiUbO02S1L858TDylcSc8CDG04ZVGqlU9p8ocejwgy
SrNrIvSeEOujNcJtAZQmmSq/vIFPaPg9BQv6HAptdiIqDk0vQ2wO1Hni/34MDwqB
Pr++KYh14KrVoznv14gMrJ0CtCof1DDMZ9KLO/OZAhPeXzrcKT/mh4NRVbS1v9SA
kQV6kF0kB/HWsK+FDw67l0XkrQYNvvIY+dQEnst5MbfAqlVyKzmk6SWU5f/c+Hy2
6m0619hqf8mgGPpkJQy+znHzNWX255xIOkOFbinkRhjwnZocF3M+DueVLzEe9X3j
3RGwYV06ft96UDf+9KLL7iIzsZuQRL08ohKFH+q7TZSbSLi9KxX1dcKPPqOKLW3W
l/qpc8vHMYF1GKBogW8P8VR1fmvw68bMQ0Y3JsYPjsxBRPElb1LvL8mhHq6oiyg8
3eWBV9czlaZArW7jFnOK0b29rfudhXnn89DguURGAuz4zS1E1bRO7NZP1hkXPmMt
LIJpsuFOA+JxgiUjV1mWQpd7YAlzZgQFJRAkAU/XKKhnWmsjPXdT4YNTjXcPOum8
Xa58OWPeswD7IgwwnhzboFtn7qPSKj5s5Dp5MsmrjkRE9kI++6jLK6DNuwb/RTs6
3imdV37PcosUPWeMhZCF617UUYyHXslfbDz62mape3yr1HbA8CMZZgzTvu4qLhhk
n+bLDLPN11bwEaAxnorraXvLBG6Zql8nUjLxRhXJh4nH4eiPhP5mSsg1BMtL9gPW
4RA+OgjeeVw7MyzGggAPo+28/zml/QdoHPyiLBBK05rTheXQiyqBiIurEklHf0rm
6J4sDUdrDuQrvb8LDdkIZmKs+1KcuONcqz4Mq4fvak36JtTwlzl7q5yzpB60y9iP
YX+yaNCd9aVIN9vzj5ix2tgDQq2Xqvj461YceL+7JfKUQ1UVSrkkb0AjhP42EM3n
UwE3EY/ZdYmSMQ3DHgG0irCYvpLdG6nMLkHelU3hSzi7/a1jXhACXt0ON4AUPTcv
xn/fyebXaLLgLNqJ/ceBHUkoEOZzd34sSBeeZaaK8df8dwR7RbS22BLhIMnY3ptu
lVpBFrnyK9445+hOEvsG/L3tspbTPlpB1OWqrEhx0s+vP6UNcG1bwpCb1QVYSjJW
vLc5azG/XORpNmlfhrgUqh5n/r6VKA1gX1s/k73SPsRBQMDuyWa+ywXFcLKjJpL9
kMkQpqyBV43b4z0RIWLviU46ReGx32+MsSNUj01v8NTvStZJRWeUGJp5t+YL0CaC
vmhpondn8mc23tuBnlfwnREefHoURdpDavUVvUYNEgUQWIeTTuNuHBx9RTO2mm8S
69kcNXUSXIzwzDsBICx8XVRKDc73fDbKz8ize72TAXho/fG3oY5pdt082F1aMwNC

`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
ncmIlFq1PDPtgUHRsUajibVQ/fLmPJzBqhfp9wIpoGFf7nGQVH7F4d+SHQQjRjQo
VYzNPOB3M8bUgKd+5sMhJTCLX23S1UclPt5E3BwKvP05hw7L9CLTTZbp6yhFFgwH
i/CntK4QKoKMn+rrRADUBJlrehjFxAhVtRJ61JyoAG8=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 2080 )
`pragma protect data_block
/sbdpEe0rSoCCs1pjHYSolmxLELb4zdouqW0wfSR7hEQeUZ2lWTHsX75knjyXoUd
BgaIoQ2/5cSaFwKrisVsb/ZHTyUr2dMlOTkXXXy1v0JpwNuz2+Gl1Id1qq0Krw2p
mCT3vOn1x+lD6HgzeytfC89wLS9kb/SJ6DpsFKLQhHLlfeyPifjbihvTO1t/Bdfo
ywqNNVUTcnVMaJLnVyTtURmzHt1hkqrFBnNisJt9HOt8xgaDrtNEsw+DbyoIklB3
XRAigfAsowNoLs4v2Tv+pn/8sGna/Pihev6seTsbnRTqGmyS3UlOqk+v6cMxOKZ4
CWYBTOLVAwSDylMaLl9LypKCxe4et72aOaSN5r3P19gmmNvQkkVrTImfho1/bohB
s7MQQwaKblI6QuBFu8PvvxpJV+ICkSBM2DrjfpCCudIxs36WVKKou78o7lSWhY5U
nFe9ZmSXgRGumUxR78Nk2qvVV8lCY0WsOnIW0Yh+uIEOoiQC3RzDIb4daf2d+j7T
FCwsZ7ssdpCSbIojIFnDYv8Mg2VkptK5BwJlix+7TEk8uA1oBlG7XRENhYN9P7Jk
FTPO66IYZbbptyBrtWMnGjYtEtNcaZaVbZ88zlO1R+uaZgZml7X1q+VvcnnVOYTb
Cu9c5qJdTaUfTpIxXMPjKX4muCwS+LK7BV051kKaz3EFkBcc+Z9PMXn4uild82mi
FeHya+s4YyIebw2pdoWyqJs8zIs7VDewefDZr98eeAPTt03ocikCPlFGv7zbxVms
MBFqTYja67ct0wm6NxQKUcCtrb1Z9kULAshw/MAsyF6A7N9AmoLN4E1y8z2mlTQE
u3quQ0C4iCfX8JYdQi8ndKuGGJKwm7C4KCvvWSrB6APlX8gyqZ2gPnVGNuxPAxtP
Kx1t10onAZAY7nC3PYWtWDPU7NWWWdVVWmGxrbwVK3qmbGSLPQcSIoSvVuU8NZ1e
qcQUhN5n+/0eVtRbcNGkTHo7fPG2uTS7pnQtF7U/NwRsxXO3ycyyoiuyuLMwsHuw
4h5PpvnPvCSKrJ4ZAd6owxE1VkrLye3LnzwZ01ybZZHFpLNnqbKrJa5i3uS0Ybm0
yaCGXVKaU9jBuRlv5AFQ7MzR8816zGLgOK3IsK4yITHI3ws2DRJr4hXKkJuwCy7/
oXcSj9w04BTGQ8CYw6r3RSWDykwsXzLl2qZkTZRhX7JnplKjnyJg44dfLAC0SCfJ
2w9cPtK9msoed7H8NR/8bpwMo9PwHaC0ArHVwUycfA/ZeKxPlWZ6aE3XRM+lDXTN
4CnW+NJKtasDu+39bbzzfJIMWOyQ2bUGFHvH9SlQ9EhoX3AronkGiGAUziQ1pF2Z
MeDAe2KltXVpuNEWneECbcnTdJ5MlBv65maKWQ2ayNF3hnLcvozsiL+sRPTZicaF
qAbqZ617hHBG7gsqUonWhpCCVpV5/miiaecDSq1ejomx7nrQ29avsnohtOHzgEs5
kQdWv0VB3zTD9vS8yZ1fxHXkFDVEWcZOAAbz1Jms+X7NoWc6h7x02b9vvn39NE6y
pBP2Ds3R/fGsL7FmgEn0lLCesrGbbp15dLSuealaYd22SvJThVyJfjih/PcDC/6E
6S67EB0REt5bjG6OxrFXTMIhodqhPOz8GOd+ffdbJ1QVPi1MZXa5I+QfhHh1Wo0Y
xi1NgN9Traf13dSmlkR3lRyk5aBa5EYeApR/Y4X1nH5wtU/ZpQtlsqzkAlxLhIdh
9LR0fl5+j66FWZoIO++ZslE5mOEDhBaemTvucsIpkrnLnqc3YpZh/coViNNUokzQ
dZ2p+6Yb83oNqBxswmOS5ZHAk8MTNGweiKoXYUwmw26N8/sYbW6NYh6aBRFWTTTZ
Y73AqQeigOXiF7rt0GY34dmwEacEeeG9ZnTjhR0QIiKWQ2Wz2ihEkw1of6RZ20Dd
GZzIF9xiOsEUyawGkVgohVyc4xsiVE57faNFHDa9A1FR1NANk8w6BI2NzJt+RRdL
Ytm+gJMsdg9ArOYuCnnRDE2XqeBofbIxBoOybtBRjEwGgzQ03MQTy6krkwmTjQ+6
aSJme4d8jNmAI+0SLRxYvDDd9RgKxHsHc+4tuisVAGcPWq+wnf741oJsshcpzNrO
KqsPaHmj4avQzvmgD6SQbeL2JZBlmOSFwbXad2dQgqrVD0MU5Tc+PLUoFpclfmev
RG9y6gEiXfGUhgpJyOHZagLMWek/Ms/8AIGN1Z5nHjl3JLHGePtI9sEv3lk7n9RW
jtrMxS2pnemDcnRwR+BaTFbkVr7gu3CDUm0KNrFS6z78q2Y93PN2+QghVTbsEiHc
406dCkZ3OIvBrmmhLBcbVILahth/Kg948Lo/T/friqBpb6jn4rSgnRHx+kX+d3wb
ZBqoseOTh17iuZ6lMvTmFod8w9Cu4+G4//Ups0x6PvAAoL4RpKCw5K4VaOnhPy9l
HKKlNou5qasSXgHi9F+k434SPoAaHzdh1QDPBw8Yep9P7LPQjLkK3p1bsGwKs52B
8OmMryOsOz6Efgnm4HIHUt78landaQj1o45FTGTVpdgfoSbsv4jKHxDnUg8qXKdt
OWwRzOifuXGUP/Dg/K8m1btW+54Lzk/wXuw23OfgDaQjVZBD/hjwNHDwE6klaViU
+D8iivUxwhQpaeZ0LYwp2VcQb8aw+bzJJtySCMTvx+t9WgDShTRUyjfQZl0hSBT2
EBbYx7avRXkc7RleLjXw0PRrquGIWAe/RO3M+BVJ+pmSmrVtNPOBRlIALHaM8jCB
Jq6Hx0eM4mXv2u08ox69hw==

`pragma protect end_protected

��/  di���s�,�!g�X�������l'��ھ���r����pVFfj4��S(�5�4Hrp$���X��f;��on�# ���5"0 �T�PL7T�0����Ǿ*�Յ�'x���!�����*��w���0`>���M�I��M���M�At�YY?��w�/��
��D���x�٫Tс�z�ά�̻8��tfģ�%�|�?���|��
e+\f�(��:K܎U{�dj������F��f�3vUP���aQ���ܰ&���岟�f��.<i���x��^���ܦ�&�$��;�~Ri�/�ؔԮ���*��r^j}�kva������%�����h���؝����0`����[Λ
	��H�~�\W��4�^d�ز�mZ���[>��?�+T�߾�E�6J�]��|�r��a�@C��B%��C.k�l֕�=��DJ����'�0����s<��=���ϩ��n���b�jc��$q�q��A��Z���r7i@�w�s���D��'��Z�)�
�Lm.C8�{0�z�)zn)�5����D���w:���
���J}i���y�)�u�Q�$�,���B�}��c�@0q9��g"��m_��g��v0"�����D��j���s��et��z� o�ʹ���j�5��x-���aI�P���b�͘�1Zˊ��:7=�~y�,_���W %iؒ�Y��i#R��?�*>�mƕT3e�g�?|/�<?�Ϲ�g�����.��t��q�K#���^�f��4m[ E�Y2��J���:��+.���w���Kr@����zϏ�	DՍ&�w����,���ˮ���GK��<U?Oأ�+,�0�g��ǆ�hk�4
�w�l#{��\�e���PJz��)�]��+�^��2��n\�(G�:��)]�T"�і"<U�c�1RUj��F����� ����m��Q�D{S���;��ie�9ߧ)������o�A������5�XY�_{H�'�'�	m}u�QV���W�C�H�M���儙�.?T\���ۢm�������|湌�#���Y/.�W$e{�Y�	���O��K��l�b l��~�9��b�� %惦v��TtJ֝q�'-���cX���`�d��ƫ{���~�D\��0��P����o����O����B`)R���)��]XFjh�ݸ���"��������� bZ��3]�C>2�-p����Ԯy#ʖxU��4���!��U�]Lz�7<�`E���X�|�����;��:��/|����U4:�W�2�u��B�z$n�x�7-*T������S�"�N"T������2^:ofJJ�%��0��}�s��'�sرR"q�3��~�I�%�Y��R��m�"])e����q��=�s�w�w�TG�E?%J�!ju�@�NuJ�;��&�$Wo�^_��N���:���6��yU�i�vS���L�p�?+��F|��Ա�)U�����|"戍���r�vZ���f��E�O~\���|Xn19�C@�x%���La��
��*�(
���o���$_jȥ>J\t�^���[W��0A�|�0����*m%��L� ��}�1��@�ę�7�}����4�@d߲�	�w(���=c=$(B#��'̍�Q�S�9�-�x�N�W!�]��I9��5PmQ$�:�V��Gq�����N8���Z�@� 쬑�ZAB���t��8I�Bj�Ka�KB�/s��dp��	OG�g~����c�M)uz�8�^��ZL��6s�v��c�� ;�bD��^��ua�*J�"	���R��K�S��kG���9b]~c�5�&LO��~e�ىڈ���e�P�6f�uL?���Րk]Fi��7ll+o�m�!�+�muW�����y�@2`*��F����ӌ�:U�����u\ى��d��rXQ'��x �h<=����~%�`��I�{ŰȜ���r+lv %EK;l�[\s�7۷���4�*�p��(|,x�X��7�T M��<�:���9���{r�m�]0��#Z�#-��i�Ҧ�Q�0����L�߰�l^c�ha�o���k��>/%�|.{��`x� �G�&Ad�D��\}��:Fc|6!����fZ�}CZǩ�Sz����+ۙd�Yyg�W���4Y�r�{m?���	��
F�����hC#���ke`5�,ʚ��#�j[���*�n�Q!�j�歳�K���X���*"������6�/U-�[�,.�e�K�<��vM�\�A}Ǉ1Qψ���o�I�>�чz[|K�q��|�+j��[W��3Č4&�� T&�����g�K���jQ)H�#Ajb_����KE���#�b��h"��hމD�9�P���i����z"����y	b����~�ጟ���Қx������m�'o(�P6njJ�R�AU��޾.�2�i�=���W.U���w�I%�֓�[�y���(BW���������gF���rf�4[��m�����9yi;���f�#��T	ͥ��Q�][������p)�CH-���b����޻ƚH�����x�'@&�ͫ2��'KT\)�L��\�/��QZ�3a�&�@a����=P��Y�3\]$���a�Wݛ�V)M/����g�!
֍�I6�\�K�Lw��/z;�����;b~�O�PO"¸���׸��2��$$���M��z�<"��&N���]�S#mR����Y���amLK9�^��vU��ά��,f�r�z�>~�a��������ْV��~)���6)�'-[��A	�R�'�Ivr��d�~�pL����Y�_9�Tѣ���orG�$h��|{��'����u;(�\M� 34�eJ��]�*������֝��\]�s><��C\�LN��V5
��~��a�a]7
W|�m��k^p����)9��3��ӎ�d�_���4�N:0	.�QŖH��w&�`:�l�B� J|e� �l�զ_������	¥|�Fक़lп����z�g��{�>�̏/Kʏ�p
O��S�i����b��255/�?�m���>/cB�90�hx���?1���xn6S���?�*�dL%vW?�<���� �7A",�.T�a�����p�� v�Z� 	����g�wP�+7n`0[sn�&�?�>#�|��1P=��\ ���������$v�WZՖ��� ��f�C�tB���}�6��(�v-��v,u��1�P���kfW��Jp�V5�L{O������A����r�T�a�$}NƱ��E�v��Fa2�&颷��_��g�0&�Wm�i�������%y��w���^
`���7���5nj��pʮ�"m�z �j��R,_8��2^�rV�:��]�Br�p��B����|��8�f$F�{ອ��hK��,�R�����e�/:e[��jU�$+4���J����J�M�SI ��7F�F,?��0H�<���3<4Vg�_ͨE��J#�ļ_�W�ӂ9�5$�iT��,:�YJ-2����1q,9��߿�^��!�>8�W�K��}�8yH*��������'��a���_Ig��7Ë�����>��&�6cݝ������?u��p�ǚ8�'=�����ҿ�E��"�V�h�zʄ=^:��{-rX�N���O�f��~�`
\��� ��4��2~�}�_�"Ճ��h�-_+�����lDs�u�0�fI�h�ŏ��\|�b`�uf��5���(����7��V�u A=ʩ�(�{KA����~8�l�ȥݍ:ܳ�~�����4�Ã���@P@�Vw�����l�jBDĥZ�{ٰ�+ ,d����,�ϕ���TE���Z��8���T%�V���0�WK���d���c�)��(���=�}��j�?�I���>��+�=���75�6�����2j���̣gP"� ��F�'�%��E	+�?�\�q;U�R�v��˄ڊvV,���gQ�G��df�q�/�ڌ�Ų��mn�<-9���ybQ��������>}�����:�(��P�%wsd����-� ?+�;0�3�K��xN����/�	���.Ȼo"8���_sP�Ճ�
��3A���HӴE�IoK��I*8�X_#��ն���Z�,��E��Η%ss�i�DP��&�z|vm�~�̾CA� �9�'8U��jr�>�N����9S���<+b�~S	��xN�,�5ʹn?Ph��� � �������^Q<zғ�s����T|nVS�g�Ã����9$��Z�Zu��Pn�����B�4��!zK�������H˔�/�?�� �3~?�d���Vy��Gs���t��z$ PD]������Q�^T�C�Ch	��Z�ĳb��B�NH��rKJ���K��s[}�b����D����N��_�[$*����M�o��f#�n��L�;��t`t��п�xU��Ut�>�K�h�Qn:�-�a"X*��T���VS���t�5S0Rp8�$J���%g���(A/p$���"��� 7���Y��W����g�ݗ�9!l�/I4�-����0�8�/n��
E@-��y*2Ɂ�<M�а�&(��+^�Z�M�E�p5x�6��_~˦���&��;�������K��@ny��<r��"TE����Z9\�;�g҉&԰8i����4��/9��*zx��\=뤨GR��!	����j�@��N�}�%;�ḧ�Ϗye���%��J�F�	s�w�\�Ęnk�tN��~k�|��␊����W�\��k��p��@��6���c�1�v�)+�u��{��ȡ����ֲ�;�����M�����&�:4�no9�\��P:'y{��J�l�܏�����<ư�qJ@���|h�zU@�A�b3��L(�GLP��O�4Y�c%�X�P�R2.�m�z��ż'<V�l�?�����������/�<H58�N�Z�B���٘�h�4�D%��i7�p�0�_]i.Lղ~�Rg�<��A9ֽV(j/o���\������d�G�[��"6�j>�,���n"
P��!��%�p $�%�#�=|1޷��f�ގ�&M��~�5FZ9�n��}
�u��K������Z��D��7V�޼0�_����8�ݯhzde���o�+)��f�I$�cm�p����j�F�00�����Tcq�	��.�͜&��Q��7a[�M���M���+�{nw�:;�u�_aGv���߳�"���F:�x�t�l�,ݔ]r}9]��������Z%��hC�����Ӷ�v@h>��5�!�Mja�q`�t���*K��'Q�׏D�+܁�o&��С �J	�4�c�z;�Y�Y�;�|d�Cjcd��F�4�u�1+�]{�:=%���1Dc>�7�'��~锇�bk���Cǁ�ei�B �f����ʰ�r@����]\X��h�L~��ƣ7���ζ(�
��sp?�9��A��C��.��,���3c��CCSgQR�M@�H �8�?�H7�kO�� 4{v"ȍ�:`a>�r�y�J5q\��Kg��z ��R¦�x����ޱ�he�rT4��L6�+>�1c[sJp�������Fv=S�P���^-y+���<��Xe|j�$Z���
�S�p �.�H��Mlt�uaT�$Q��#��st�ǘ��ո��f�����Ēe� 4a��9��cR�8��@Ԓ�Q��t��/E��� �o�:4*ܹ0���Oe�M
�/F�ϩ�h�ş7�uq��7=Y�TM��G�>_�Ah�rc����@�!�ȸ&�F�Zoq���(�m����f��4��ܸ������5�f�Bq[�������Qp8J-˿��0�1��ޖ��>����u��������W��)�y�EtcZ5`R�\ú]�.H �b�f��+S�Cx�H�N�%}�8�_�O�l�mnD�� +-�i��O6��'��C=Lcf{��"�� ���>�	����F��"�z2k�fH��L_�e3N`�5�|Ll�sV�o��)_Ag'W)�9.H��~(�x�4<j���ʉ��?���v�
$�@|��ˊ�"#�
Ҁ_� 5,,�TO�z�Ecɼ��7�|s�۠���2WeL���q�,���]Qd���uq�*��6vSӗb��tS,B���,+������$o���^(�i�+��r+��ꧤ�q4^�����2��M��$�5��g��iY��)�/z��~G��$�Y�����F��dm&l�Tql��v6?����}��
���F~x萉���~�7<�r�P�w��5��#��D���s����xP`f���$���\kL��x�i�����\�M����0�}F�W�7:��0�tN1�s7m���k�L7�e�5�	�I�ӧBt=U�~�g��X>Pno 1�� �m����_�%�S�O�5����}�XX�y�`�1?�\��@�G��%���e:ɘ��Ya�{F�����dl�Qa�J�ɑ�P�i�-����bT�,q���x���$4VJ�V{,�����&���r���
�h T�HED�L�q\�e:<^��a'E�n4��_Rhfa���F�x�W�ޟr��Kc�\&��XSX��vC%
R,�s~Ē�ƛc��W�ܹ5�~���"�D��3�q�Sw��"	I���޷�O �3P'rPz�uv���.���Hc�]��=�]C����iK�t( ����]˽�0^V�*Y��nV@�������}�y�6М�!�'�e��j�����T�lw����d� �s�C����Q"�)V�N��N�QC��(u�ߡ%��l�[�'�,ϞO
mCO�S7�lA���!�g�s�2��T��O�����ɳ]zv�XK6!�>8�aPx�i����mA����	 ����� #�Jn�P��/�߰΃�D��͔<Q��y���3���7F>�}	����S=��h�_!{ � �4�ݜ�i�]HB�2�)�A�)��qRp�X�P��&��>7�!��AI�x��*� <p��!5�CK-����s� "H7X�S�<W�R#�1��[?�'9n�'�C�����M�H���K�,�P ��X]*�]e)�����A�?�bC8��'���3�"�gSo�������
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Uanpe1UXAlQbVLyHHexiGzgf5S9y3O7VP+IONcInmY/KHslFJpPFewSk3sDA72E7
L0Fa98CvqZBREMjufXFqZiGAw3S7IQxluWtB1wL+3urm34mH0xBUjuOjvwJiWP/P
+WfsryAVEOAvw1iLa5a0/8Ixy/dBLYFcvxHOBbzXLeM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 6208)
G9pGzEoB+uTuIp9K1jVduQ13Pj1Eq0QvFkPVaE/Lyt1J3FYmDLB92z6qU64Aagjs
pp73S6F/LQADwoZhcBHk8c6HvRUu4yh6RKKJrCoD8xjqlLCxAeMFrfzM82FbAHqs
JpfOAxvgjyYJZ77giCqDSUOQFCI3By25vagKuA7QIW0dtS16TfINI3dAfMLl4q6Q
cU0UCOYrHyAKVo8iB/j+KQfGKg7D54gMGr0WLPusk7B8IuWA2gd5qASZATaFGV1S
j7rk3oyJWtxZPNSLbYW1a8eRTqwhMn2/jzqvq15L42oK7uqqIOW2RW9yzAgHrgDL
ax4ze6tIJYOjhwi9McWYao+BpxkGSbTHURjHc35cC39I2n++jgH26myGIYzZ3dJn
A9bGl2cbJZqOSQIMyt9GYS/h7PbCWq6leI0As0rRTDGXBUMv6YC760U78ckLsExp
8iy4VYMpsJpJVrqfqvVWdGw3K9d0yn01CHmotJ+nuq/fmy18bbky6RN+EDLVlelv
5sFyBtWKA0ASrMrE8ttgZiAaUUtE898lS0OGTHWxsprHv3EYWXbzKIEhpHyNm5IF
b8NdG7T90MKiUH8F27Eae5/vDJ63cuyF0hae+DxyzvrT9W6GsCcsBKBy9fRcLS0h
xPnms/mnGH5FDpCmSljXve8qcubC6+2iU1j5MX/z0bhYMry0e7KMm/2Sibyb6KPJ
HGFesc6eaVNq6jb4NsJ0aoZPjsxY+7W9KjDkulEBlo9e01KcB1OTqa7IRRufmiAC
TevxcE8vErEtbVvDyQ5JZYyuyWe9xn3RhaoqSy6kQ3ECT1c4Ro5mDW1hFMdtyS+g
xMGEJLNTI5aDF6mZa9u8BocKcnc6VMF+iy0DNnwJeQdVIrAnmtqvvJZ2EaklOXAu
cXZ/5sLYsxS50yVB63tDfhRXzjdmFAftAPnG/MPGsZBVL7qSS+rPwUGQipDqsT2+
xtJI+rB/GEy/iN8J65aSmAcUH1uIk7uLl4XnDvqtf5ZS9BPYnW4xy6QVJNJhTG7u
tQUzN/aauVPTDyWIibzabrxCd4aEO6Aekk/JluLnNeas11rMd2bEvWy3i5GyWjVD
GudaPZe3lJ/9TgtJ3wY7j3kP+i5ClgioneSAt1792jDrvQ1IWynzi69MLoTcB5+A
ob5IoQOrZpKwDVRnuE52C9DAVbDxIer+bot79flirFGfykBVDqs2dJM4VKySWIRW
M8WXqn3Od9pHzTX4W1w4TY9qMp/jWSaJ1kfla3UhxzCzvLiqEtW5SRkiZ8m+qEvp
8SISWBU86BDytjbOYMMprd2Nvnk8zGb4V+v5/DEunWxv1s1t7BjMCJ85uYvSClhj
2br+yhRXyOK8z4JB0n9S4jrWS+c2D12+gSmW+Jtv3dF1FjxxV84CKra7Tqy425aT
suKMoVpf3jPRDYv7QDEoRAEmi4twbSxdGbSGwNj/McXfXKeGrvOAExU8deehsal0
+yrp438N1h6w2hWLBC8UhdgH4C3gXKxR8tulDKGZamlD8XPEgk4qSm8W1kQGqRJF
X+N0bpXhm2rYqfBI0aJoC/MLBWjNixTYYrVMI+Mxj1ffFv+akTaG+XPNRIt1qVix
5l1EEnseoJkGV/pG5qyg59z9Xv0sawN/18TfRIhviZrLW37fdIKkUJVst+UuDzPB
z66f/cSafBBiVPXT7B7smmI4AJQkoq0oaEhq8z2ksfqvv2otj+tXexpSFQwHZ5HW
he1hIdKM2uBKZbPBZiyT8jjjfN+Rz/jIZ2vYF385mg1SFZFMkzfKszrzjJMHcqDO
iK3cfPio/4SPWZlnT3Bt53ycsTaDW0tk6sCRsKN98T0y4Fs9lO04XiOhhCRWwXg2
fX+lsY20xxGecoO1F8Z/6yIcnl+bQvijBz3IW5tmiqj1LFZAt6HRyQkBOcMWJdGC
ZyrIGs5JUujkBe5e8e1fzTmogkZrZOgTro7vOQejCRrOLs8VkqJlcJHP5PEPndJ5
uIncenOdBf1MTChDjk1NjiUk2Cd3obZ5LE5VUicB+krrDfDmGkiyA4uwJGDsdZGV
L2GawPE1PvZLxTBmMdmp95t8Z0FSkBiapkhjKqSX0dmAy3tOelRHsnb/c6+y8Gdz
1/M+sjIZ/nLZdYMP8C8aD+IwbL78eHOLsqveXCw3Sw81myExK1TZjDAG9t9mSzjX
00ZUEZ7cbu/lQQWFNHdje70WoPIUGP+H+UIi0l6Y03UIzDE4lDvpLnXboGmgWxrk
etzWrrRDNbHZsj7JLzbmCjQVcorZQLb38PDP4L6DQfMhLzmYFrvqB+Ky2QPicSJZ
NWLvuxAzNd5oxntytnMcSREcJ0MDu1uldVphC9sTJN9EKxYK0/U80cPZ7FMblu8Y
H9Wc1BsrqAndMO18Mp3p9r+d6mqVIF3NQaoVFRfRcEsTLPorPLmT+1jKg3KqrB3W
oFTh+DtSuLQdGjgLUbR/oOGYjz24ulLgf0UGApG11iEqoVXz//UbyxsMwSje3isN
Mh9NWVYofS5M8CSqJt/NMwwhifSg/6Wnbox/SuaSUfenqetCNBGLOcPd3fBg03xi
9XE/OSicOixRU8lc6Ie7JItEtka/2l4hfH6LwUdRWVbpVsX20Tl0HFOs3LvPco77
UsQ8p+HETYONNaAn3rMPB7gaIPwNPdCseNo4AGrcMYcU4BlYa5TM67cgppCn1f2q
LbHJ/o5hG+nTIT05N6AwRrDih5PDFmxjDu+aPebKQI4HWFn8QIkIpb5R2rWsTQ9R
aGNvqUbpZ4iJxXegEG5rIdBeA+Vi9IGmpe0erRPEXIvC7bYNukztCMC2yD9rnPRp
mXeP3IZeDbP01L0hgcoO3PkxRlPojp6+ryn5F+vFE1rVIgKIzl7ZOBNflKv5sOkU
wErrja3WRxWPH31mZP3t/oHQ25H3wmwSiy7X+Sva5WSUzfUZoZd3y2j4Ho97coSS
7Q1Mq0KW8X4okPaOFSVXdILwsSmc8GhXQeIhTjwC/wbol7Zc+vDsOBM/si86m+fm
RjAtbomGDEzwzpPoPRVp0kjLx19zjzYdAm+htipEA5sz7hSlNojsUxq8KW9sxymP
TFZcuJ/5FhKXhmb9oRvxAvmj1ZQxbBAdEBej5P0aV7RfacmasN0LBMsJzJAosx1f
KpFQAPCzFVXAARw9rHd4ffWvdvNfy8Qb5hd5N3pWfG3RVM+DU+eIvTPaTItmrFua
bpclPgKtN+wMxsB0+ao9HkUkZ/Fhs3TzVRTNCGZIebxarMLfsuV5WckxRENFscDO
UnyOkMOXh3T0rO14JtjmoLIgXBOo0I26nVfzYT+z1j7CfQv2NccVrCozqeV/ulcA
HeyjuzxOgDmInhhD3QGy3XW0z4+xz1MZLJX0fz/6Eg30JaPtsJDj3LShFB/+ut5m
cwU4S+4KcoGEqsaWYMd0nvRDnMMB9V/P2BO41YVyltFl8ifL4L18KxI0fc51shkZ
7sqSOfGRLneckB43cz+INbIN92aoCLshqKHc+SViBk8haWaCLkW6cajGX21CDHiW
O2dUKwtzUNtDctA+jAuyzTmq74J1XqiOJu7KPfYh/Krra6ZE59pjFfI9FNVy3tek
o6gi2tUej0NxD/f4I1i5v3NyCEJnyhK4lPzakjc70JRE2kTj+R74gbLcVZZZUZyA
SXZVNKju0WdatQvfY/PLynmOcxMJGW/DFz7AO6cMPKqdJiZabCNETiGiZFtVXXac
v9D9hRBsaQYzSxU9InVKgf2alJHpgNnI4UiZF2386JDZwdtPuN53YxwOPYmdpC74
4vpoE3T7jxiWMDwDz9Bu8kp6QNra50mmDOKpmgqURjAyjetirXbbNcZ9R9Q2ZoMp
GPzxB71h+x+BVk88ISWCKNdeHes7SmtBsalwmQpG6wo0S+OHTqplKnpN1K9BIdqS
Q3XH2a/x0cVS5uhpITXLnGMsohTkq8HxfGwohoDJpBX0fdC9Ny0WPX7M31uMvkW9
hjuTOCdpbJSmoT/y2wyibtdKQW7L06/yGV3g+Jr1hAMHsc+4RfKu6pQDsA9sdbw/
LiLMZz3U2U6lOCzjdkuwrbwox7gI67w+hoyjuaSogGTByHNjoGchISBWLD+Q43Pv
bPxG/W3FTDf1qlN4i6uD3q89MhGM7lUo9pzBHZikdRVUg1u4CNRq4GLdiDLdBmvR
WW1+lIiA18ZNbCnxenuB/dLjW1j/zHsNlCxFdrUZVk2K5Rzb/3gOff1wQaFb19rk
/xbGFNB/eGBh/lb58lnkh5cT4OSD9MiLyWKUGUqP+ma5rqO3NHXbyzoEM5NMcdis
dgCS1ArENNpurMeAWB3RuOfWMJy6TcXf3/hiRDMEP8abSvAeuhN3LRYLCFgrbNdt
nFaP8g3lT3/mMvWmNkJvk2rgwPcK0XIApYohJrQfGM4DSvnlLj636QUui/vi+Tzs
RSL0qbo+FewfQzpAmKxYfOwg6664/GYiSZdMQ3alslN7UJisQYJW+Jltv0tPzrkl
zdlkvPSzsWBcJ2AX9ZbFvneodlMrEF6KrGhYWRNlyV+XaefCyJjXyFlXQNWxC3dn
NzRH/Es0PDGMg0zzzNDnFvTniCzdFeYGGW9Bb3SsYNw0pi/qs6NlSlMK5cDxVnIv
mm51A8Jj1z6fLlbVN2QIZrVu94yIrgH5MzGoS9N6ucZkUckkEQjkRBK35tXnbMPG
FDuIGgAGGWtZn5gPDULTn/wqBpC6OzMWuwTbo3S9/Wd2A20M7O7u6695H9eZO0J5
MspN5dcMI0Tm/kvTxW0RlbbJW2J5/DOsjFER5h3sHSXa5JAdgI2hro+n2ylh/N47
9U612dSefPLIpR3eKHdjYAqdpTHdrzLWBDDLOoDwf3Tq2TJcwsUucOWQ9ucmi/Sf
OxAr6+ln2GvNU3C5WDoQqmaF9+Wm56Sv/ejINHarcGBu5kNiOhmLf3LoLNKxaqCi
3/VUO/ek+GyAAAbaToRGriVL6lftkYfaXsquMHthU9kOydzyzAQ45zYSOKaRHomm
KH757AhjKiyvkG/r5WVpm6/yOj3ZFLYcnQ9PZ805QydKTl9exiAe7tLg3Bri4rCJ
zXa0EujPyq9+EAjqvu+wvYxj44rN4a8BMscgTSxd8cMyNUJdCUrIqoKzYOGjsmE0
my3jyHzC9A4zqPGoEQKGX/JDBXMw5Hc5caDQGjDqC6zxx+AkpZ3sGPCe5kq1QR+c
LHM2Cn/0yCfZCXO6w1XKDaeEHN+xBb/wTSN6o+5iv/bWNgJKbcHZxtzipSFGzHj2
PlFWJ+BZt7CXpcfZ76mKlNx0E2dGSBj3VtIBZcUE5sW6+d6KmvdcOIHYpLoQy9fC
+WY/i3AqayVhaCvt7B07CKP42R5YmG4UCLVwPRZNnFyzRtpmsnYUBTcyBj6e8t5x
Oq+j5gbbTlfO6GoWKquTck/8dWA4UyJlb7hEh6qwnJagfQuLftnm431gkt4O+2BY
cvZX+TcotpcLUFHec5CgsdNlPA+srEzn3PTkKMa5/dMPPPRmwK7fRnkfUcOZjt1P
yiKIaEEjh3AMZJChr0cKhPgMGRda3VOlsttPDb2BnPqHyKvwVPJwy2UZj28Gpdvv
du99Pi7TxqJBkHRmEFLf1LXF59SkYjuvzDHmpKtamlTN7n4kbPi9dgQDibe03KNJ
1Oc8wJgPblBag/mEG792RlpZVwEtJUnDTVJxAfkSqPLpjWDcAMEYXQSLSSBfEPjJ
XSfBRizNaEgubVL5I2IAYWJF88PvayDsQ8AMnJ5ntqrkWHiyIoEFCKCSjGggwf/q
Je5oOl6RdrkE9ysQFgpIM9Wr1T1/FK2YSq0ip7cH0mF/hheCa1ynhwWkHTSXwe8g
PYoA2X5kDoLOicsZMkypO1UY8iy0h4t6L5TSzDb9Aeg6aFBdFyhtNcdl9QxsR06A
gg5RzJvwEJoOii5fOaQRBBx7/EmrRRy7IiKukYfW9bv+f7QzEswxGQFpqxggZp17
cYcXCiKgS7xAyZ7QOpgCzH5IDlVjgF4QEcEr812M+inFVbEtMe5Y+RYIHAIUAymU
//bHH66WSCjVKfAbnq+lQkwaynZaGubfxbg2a/JDGMGeC6Fj9OIGfXPf4DlZIQgm
8TyjB0dXdChepjOOafaqglGQl1t+YIwNvyyGq3E52osoctYyfY0ZSt1D/+lefgbV
uKFczSWdbfYnuGEYy7ivg1T6B6xX9m2B1BaO/7ozDNWKUOoL3b9E7h4EBsoPWtxr
UjGXoArIQDGSil+3BSg6nf0WFWIDvJjFi1Ew1qDkbwRJQlj+BbIlyJTYd0VCPTlB
qbx/4zIya5Kj4hgXD3cOl9TWwu0n3hn6acSOKoYFOQwc5yGi/qiSNfo/9Y1TlETI
IU1d2VreKW5vqEQIo3PPLMg22VzBpta6tU582z5sPbFmcKhyKren/wnkYwuVSshO
npqbvcO5RjHx6250o5ib7MFlNgtUFxdcwoOHzWOGQqora7TCJfMBhmQJMHfMbN23
+imPx/vnIc6b+rTdJLfIrZhxgtfbpqcOc8F1Uz509pFlMRXGu8zhNC7t3051WaCS
finpjpfju7tBLae82Br2ytAiFq//dSgcvXHMwhN2thAeSy2E9ekGlxvd+OUyTq0S
vtcFMFNtwyZBYG2AL1YG2wDaEh1Xaz+oU8R7XFfamnrnCxv8AOVaQQZAX7vm/mOB
4w4pFVMhZXsLdfhTgP+trl3WSqT/aZdo9/mX/Jn2Wj3x/Wz+y+KbtvLiQP3CDhuV
jysSSMrcgiarAPf3UzPlzxHh58x17PP6QZGvvwia5ztNL2cT4f/trQl+Wq7qzbwZ
O6yEVPUeFMcq+xuCwsfDTobhAUymE0YnqlvA4I1cuWRVqwonctC6qTY0C0PWed4p
mdGbZhXn7kHyJQ8ATRJ7zRuLiDiow/FNi6hrsig96cCGpOg06TOUHmbxZbB6fdNa
SBTV1485vOdVfzRhOqF6K5Wk0kZHGlwATJaY2Kn3X4Lr9BzDckGLNhpWJnRfoXuM
eGR1/Qa9y6lXHNRp7s/1TpcVSYa3bn2tRAMv3zox0xAHXH/RojXKffjkmFhi3D8D
5KSXkwMH0e7B0fuz0TwdWY/zdCxAQsZ3JTVuO7Th74PbM6Vv6RNZzhpUUY2aFmcC
uuixJ/3/CGR8psouGzLvtDFMnMd6bfzB9f53NkdpdEdwIQY2pyYe3TZDz07wLifk
Qi4mRFO72FXpc5AhIbJJnzAMh7VBePETDDYJW4hDoViGcKGIsZyr8UJHaEARJmo5
dLAYkq+R5R0eMRSXFGLQa0atrSovbvA25aTHLYIOCfVOF1Bqo9kP1/0Uhamqlu4f
nzdZR/t5e4KelcBmvI3sAUi3tSFjOnRfRgnO/M4BJ45P0cK3k+CvEPNFsbvrhUw5
/uw4cp2ysMvgcI2xMfIi+tYaal6Ihi+Rm1bwrfqd/80/wyXbP9ivWPQeGY4lrt9o
dq5L352HiE7PlPv8XfD8cBDzmlc0Egw+RouE2ta0n7mM63LP6Uc/91Vxry+sDd0J
N4+dhfUolayz2I1cRthoUPYwfNWrXb044CyuTN0OQwoCCksVECGf/xlsYxr0xOzi
PUFtSxDGDObQ1bGn/feUFzaNytrXfjCvp673i2i+5gUDbWolphNL3e3krUFM+pYK
BFeRckIFVOrVmCdO7apdwGcUpfGD/nUh4vGNUUY1lEueCzqy2KkiMTEirvnYzFj4
AFDW8wPzPwYSEhkwsSWg3U5hdTcyeDSxR9Ai5cwfW81i2BZmR8uxl5j9leSYJRbT
pIV4N3cjAFzOGpdZwNbvTIx+noSof9IChUL0z50K/8/4iVdhFU6/063FpW680YAY
LfQw++8Jibr91LuDGDznVbvpe0isbHICFqaWmNOX1STf53Knz6eB0DHzGfi75pkJ
bjl/PFW53cAySC8vcUCjHfNb/aA0MbrG+s1z+UooI+qq4lPxwFXmabsrknp4bVcH
qrascEd/5Zd49PfB6uRh4EgdilbqxpiDQZaLw13VDnIAzQN1kCcJ+omgdOsWbjrA
KRF/LsNMa9773DTvLPSiIBT4ozBOXw9ifrx33L6gHSxstQWUy/TP2P2TFGHLM1b9
iS2lfJ/kj1Q653xVy3yiR3/Dpt3LfRhjBBsF7EXzWS0N59CCTEVqoHiT5NI2SmDL
r9sA8jXIjpUvV+/Xs9I72TJpqvM+alzG4dl6N+wYLlCsqI9tJzq2RPy+AdHEOZl9
XYLw2ql8htztjIDvubgGkDhFSmVjp2NGHiF/k/mvVAoZ/dM2qBG3C0tO3UsfbQ/8
5agvfQgYClUQwR1WGczmew==
`pragma protect end_protected

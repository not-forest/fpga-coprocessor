// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Kgv0s5KYGrnj3DFxbFCWhLrV5bwTR4wLhn5iDNhK9XuTVf7R3VG7ubO3XN3ezcA0CzZSkubEmuHA
UOk+5VegjRIXiGXEvdHpAkiPY9IrSfpTVxzC2OB68bY2QBzOOWB9RE/O0lTlXFh4pmHd2LqUJnzj
E95/PZVaFaqoX6/X4hamqOlEEyroyos5WkVg/Gp0uaPvx37V9L+Kq4UMrAEuwraTU3IowiuAu+jD
Qw2A34pP/vjzFbj/EKAXxNli7q1qqZZzc/NiTQF6n6W1u9TxBhQuFx+cmfEfKrTY/MaYKLuA0Y0O
3LiD5bgG7y0zayd5EdLl68U9FTC1j8FkLFU8Rw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 52352)
4dU4NdXu0R9mpiPm/1REbfgLEiqADFKXhkZJkYHsAUsQeYYAWh1H4PMdUvsPXnneR3CEaKYzuQBi
fVkgf+2u6PWvzUsozqCiK5qDrCVH4n0mamqgFBybckb4fvHPk0OeM3NJZg4qRTxNPovpRjQaLlpG
8I21LY3M0ck0RFVdo/CCd2oNbssDM02oIZ3HpNhaur8D1RftbVliEZp92ImKc0icxasXiQtqHXtW
dffYdEC8oF+stbPweDLDmiRbZMg5oWoqU2ImwsbObIPFKf3neqPC5ll1xEV6WLPVPRBUMpnDuq4S
ZhlLHAw9zp5Ytf81cnSmL7s8iRV6mPqyPV0fBuX8gihkD87bFn8YcptJhC0iWxhRYY2LwQ1bePHn
nssl9uaLtOrAFtCu3uqe7xirvHF34v43A8NjnvGHwhS+eeY2RcvwQHcgXc/9vNVvQIdEtB5tEk15
lcLAV7DklJFtufM8ZSv4xbJCMxZ/QFC1nMfZdQLauAqmWZO73M181iKaKe60EVkDUo/Z+Zp02fzP
OTHSlJ3eH8Col2fAiwZlxy8crfZ9VDYIfAvr0aLY7vAZXa3n9VeuGIueQmWBPt3zc3zp5JTOMUWf
/9GPNZdZyWy9sD4zhiGlrZQ8CEpZPqWYlwYkvQH6OwICvcwL8gpC1h9ISn2XMwkYnJlut0LCGNBn
nIfFJjTUTl0LcixA7s8w3pBSOTqK+zRcJBWBeWhTecuLRO9ljcO+uiZq1TsgNsp96FE/exVqark1
WPbyQUpU96yO1+9ULFRMNtB6f9Iwcr88dcRv30MkJQU/IC4uX51yXMP5KKmDuvkQJUWDfSLIigyx
xDa6vwekRcVsBphwpKKYkLQV8fsP+Jt7m0z6Eakxqfmt+bJ1MgkfwjlyVjVMuNLhEmqTSFVU5lWM
F2cLkWDoNG/XzkuCmSFmWLhVabBO/yzQ/jcnmV4D626Gk7NQiUXHSXH4qlLYi5o5iMrSWFY8K2fr
nWWyZn1DWB4XIUHm8CbRCgMQ1gVEPraNKtznJvYPjRum1tbarD1HUMZ0dOkwj/HYS5qhQtILYujr
Scqs/kHcJnb3rL6OwT6CfJj9gF4ZY3TLzD0M5CszKkMH16RmJ2cBvFzsjpTJRCgn9vqSkKLyI54j
cROww8ZIxY1ltfsPxdZaH1jUGR5VS+5/GtcWmgFR+/SS8uPeiQ4WQ67zJ4BxscxyO8Iqa3rPMVcU
DanPXNiogtFx/QwZ7AbL4zSWQMqDRFkp1WKVnJlECBmgQtxVIJviu+ddeyR1H5OrnTvuDYmqrL4P
D6Ucb7lisFBZOfU+Wv+A0g11dIcMB4SypCzIlxtiA4ZMzwUIAN0g5G7Qlv5bjqlbfdKuesdJlA7t
Jo1cxjzEkSzoi8CnSRAk0qmDOtS3/I55dmdzAFyFmZ7H6mCf+t2qf0d5nD0oY6IyUybIxRSXBP+Q
wajOONlr5jqLnmrrcN2sSj6VUeQ+/Jd4neotF+oH72Rs6/9ObeyBLroB11Drli/+rXmgj9DI2XFU
+i/7t6X6Lpe5M9mkj+2E5M6vAFem8MoWJlaO4ybZstGZYHt0k10HnayEbU0EzVuZJmndO06BtNIE
QjZKh8cWFnnVtwGVHkRv5Q+P4MX3zfvoDQex+p2rbXweiA8z5R+L9hRDZ5pwtY2LoxsqwPcyI3pb
V3xxmQ7se/E+nnHwOX9xSd93EIgC6mjnEqVFdYVlcRYegY6xU0lFPMA0JWeam4nJt8i02JFkum3L
qk4bCObARxd0jpzwlQPfYIQ/EARIn9sr/tEQ/WC/AvUIJlszfVhPkDQzEHRx8X5hOdQNrGxpFhyC
0FsLU+s4ppn6mmHODd8Ssbz04BX+Lmco7uRNwLIlZYy2Euf/4wmw5XceBOwb26g5EbMLkjbx2Jmm
DMb/ck5iSEZh2E07WsPbIT+nkVRAxgJEWsbMVPUA03z1Kg3TlEwcR3iiq6dVQxPduvnRYSIpGmrh
pidkB1Go3P3KeO4DhGENpG08rsYsLxqljsnTii9N791g7gBT6oU7OBGT1RG26jNXKiLtUHPlaPuK
M7GMgYZgNU0X/TEwxWclP/02pgvWx+zRjlrU9HqZ6K3vp5O7NKLKgYNtVQRTQ3yfng/icD++6ydk
7GD5Cmcy1LP5zFf327Py4hz+QnCTTg0AmvZiBoJWS9yzMqpqp+0yDTYRIPXvUv2nRGZFSd+BrsZZ
dHl5j+rfySRdLekxHtoff/b1CqotEWNrmDhN2nIDqcwrxWMD8pG5Z3A/5r1JHl3rpPONtCdWw9Ga
wuLxMjQcs6xDvQRafDb+0K8D8CM92NSLeYs2kfuMM8Mx6PW86C3rloW+Z/kKaYubMoPrazfJT6jU
/FTNi1uPTSIupS08q1dilaaNzx4fWB5Jwi7odybR9xvYRCBMiPTHiUn4V4Ivs+7l0J26vNYLXUHa
pofn30cfctHnBPt2ZfId6HXv1/w0v//6ipyPoX3vBk9dNCoUCGQlJ3cw1Tumwr6Sfa3TriSiAk+l
AwsPUfTNAaXo+UAO27VB05UCbM0M2k+HDVYnFRkEomUHKC5UxBY6dfHHIjClYZ5B8M2C21t61QxH
KsDWaIkwGsGPK+Ziwe/aaXGC0zXdqd73YbEi2ZGUzDYa69dIyj1y4ja3spLOmP1ZJ/3M/ocXuXx/
ypaBcAdxHoXSPe3RRtduzTiX3bGj/T0CDqqSHe1s6CSpjhBjX/kf7S+jElrylWJN0kjFvip3Kqbo
QjzCJWg0DXVzQ/1NpzAHwlYKt4jbvkzJsbrUBXXGRg3Wm6iuaeMoWUEqj7ea9zqpszsIGSfL+Gcz
qqziuxUAtqW5rtPZ965eJIqze8FBlgYDwat6lPmBZM0HCnbVxPXLjaP9cY3uiJjkEmwOe3NmXeyw
Q7CMXrnvzcMTiy85BewmmVjnx5bHxlGj812gJln9wogLgQaIpOzT4ZqX75BJL94TthP5CJC7c4BH
i/bh8KWLIvEszQNSyzTOINUAL6Zi6wTAk1YXzAg4OhxMRJCuoqjjTnq+bY6BSbjmwJI5hiduO5XM
o9xpJ19+KT4mRopacgHUj/bSFOThLHzGeb/HFUPMAfg3XehhAEN6LrNMuXRF/40iAWO17dlS/L5R
7YXdJleqhT8CPO3rEPTdt/7s8fXMrXaXvLSwA3/MtqoCKWhvJGaeDegPOhqIuh2BPIwwwqoNZFaX
y+RZDOQTaF1iKvoAFxT3hGp2nR6oJE29ZKxXVYIi/oiH/rF1EkSB3QUCI/R0TvkomMLsvNIc1Z/1
gURm9BMTuApp0OVH06QCq/8/uV0XqEpPDtAdxgXAPOXyRGlZ++ksv5O9Ee+Zgn5v+WkSbRMvzdDW
39cbuOfWuqeeDap7XyDNcaW+EYlrmjacmz7duZvbPTfcl64Hqu1Kt2fHo7UzCvrjz65CCwZ5SMxD
BYhgBdBNurnwo+F5cjTrf8YEmWA3d9b70M+ofi8EHpvJQNLCjR9VbApGMsCO54XRy7nsjmFDZ0W5
gDdO3tYXlMb5JcW1pb8Ea7bO9KHApwxz6V92bLP0kaBzG3POf3+K3aGyjnsLYFYmYbCqGnd37dTd
Fo1BM//sJZTBNf8i/9d71NNlDht/rMrwP5uneR/0Ib2ll33VvWddl+cX9+Fs0w11+u0qaAcVPJZ0
QpJJlTtU5qCENVHnnnTuorq1U9wanHt4LH2BGxc5L9xwyR0xZ6DE7stRVvZ3DKvoIv2G8gto+Syd
jZ8iib69EuAoDHhdSodWCg6HTdJ3fQqwIq7avlBeapqGDHQl2NKof2jhnXioA6QY1wvd3JJGDKsT
NiUUUV6wVFKvs/vYDtDJX9nfSeur1oc00oJDGg39CPASX/lh5xbVEP9HDB9sEIOzMCt+NxEL08kL
hiZJS4oJnNnP/ynV196ZtDoacMY90tniLQHI0oG5iGZxmRtpEdaX458Is2tkZsTRhkfBwR+Q83bg
LRNGXrCRsZxL5vwKNKbMys6p10wQqieD3zApJKVHOwa1iu1svoO14Gw2X4LhQrDHVKmZOPxyZXLX
nkf3+3Li5SYSC4vJLRx+orOGIy2zQD39AoBMUjuQOcNXPtyQB8RfdFEEcUL6C59vXNa3pgni1orm
Gpszwt/OxqvL+ZiV3/kSmnOkEirFUe/3JONwsshXEuykR2rN+yhgbTqt8TCpmtkVYsWGyXo08aru
1K5VzjfM7lGKUZxtrTZ0cV+mbqZGQgqoGBK/LnNsPH7VejO3ntq7OLaBZqqih4f3vpNQWbA3cT4m
DnyUvztsK8BmzKX+/m2bRLXtK9rI6Lr9Z9OCCqLfksR6II2yCuVcXFQi2BU0iYccQeE+Xv3SAeyQ
2jyh5Elp0sA/aV76vRN71BBOW4+bzxz649ZYWSmMUGT7NNQXyodY/6asjxBmA1G+g0hQTvNE38bA
lDjw8QY2N478a8fIX8AJuhBQ+fOEnZMpyUZu+5PMC9LtzpO8SKRsazfUv70zS4Zmnt2jRjz1q2Ar
s+yiiI6d/hzKXpbN+bG0wdMq7/kUFRJz9cDzVScVOX1iG5PbQhVLKveCwbr5Kl0N0wH0OPGANfqw
PkgUxZuRd4JomD+dvf+L8Mc8si4aB9te7RSAat1s3oGjhvgPqiFLuYjb/3OXe+xF8CRpAp9sQz3P
Rqo9DgAdpsgXbW9H/orTGqW5XSR8QFWv/6qC0V7FF9FQr5YtCuI+1l4hJOd5fm6oVjWEJXNtSRIX
UTOE9oBqLul7aJC61Fa2IfWWRD+c+Dsp3vBVljdRQluP3YfvKCVMVz7NfmKT1tt4UZDy8lauezaw
p+zKDpBfAi+lr6CC9Gd0EIcCg0LdLRIvSdJk61+p5U1d6AQD2A8jxmvhmIY8f1W4vqLQCZqqtpjp
V6JCqVGmGbGOfrYeaBfRvdxLS94FgIwpWUFO78f2Wf8nwwfOxMXVaEXXTkes0jE0dWPnTc+21EgI
bokDw7ScWwZm/0veQtI2dMKR5dxJJOc+PPtiLyVJ38hV9IdTjqUyVV/Tvibw55owYu1CNrswZxU8
ro2w9AZFKaNcmv7q70tBNUOvv8/QQVkLfyvEaZ2RdxgWlJNBUGZlxHisbBE4+PsK7oZgnlq6ELgI
/XTAlOS2+FPRS17+1CafC18L7pjfQZdksPmXyCTR7A0iyGxO/c6QECO+KmGVDkcZ8/WgknTyNtSp
EeA3vO30vsf3rWj4vAl6+3KQ+6Y5PxEhw733TLaf4qHXDvBLaqQri1HqiPFrPniCx2tcMJhUtazI
MUf3Nmf5lCJmew2oHwy/1tKq+KYeDSuA2VuDzOAvuKmHPJ5iRYZmg5rfSnM3gUGCYwdJHeDLDfiC
mx2Bi8lVN453fblvuU876aK7WnWRyf8oHmRc09AymLlJ8RxEmSlcnsKvY+xMsuAe6HA1hjZaYlUf
AWzneAoLaDhUVxnL+zW+Po6apVrrx+pHosZeaqKoCUg5Yeg/ZBXVhw0noaYKlysmwRh3otwcSVfO
fZO951eDygR+3Bsbml0Bsz0mUQELJbgNsBrRpLY6P4uuP2cjFHnm5hjqG3c+iaFGz4z4u0m3PH6n
n7h+pPdYMwCfaBIMT4gtki5spSMkB8ExR//sL6qq+/XEuQD+wplOmbPgP3fzzgx53Gzg7k2hvyzN
fpC0SZTkkyFXGb7cFeor4wM/Ig86xgpn2mhVgMGhFUNLmw6z0ZkcRwlKXVWmRKv9oW4uay2CjcF2
N9+BWQiPykdQqqg53x8Dv/HgwV9fG3f3pmRFUMGK4UuPbEzVnlCyUYluMdeZthR5Oh29eFEnoaGB
08JYjmXZy7px628HIwnC+j+DeS5T4lF97svFtBk7QXM1LjBgrOy+SS7bRk5FbYtTVzVYvf5lpQFy
fBRSDHt0NeEMjvLOrr/P8ACvb9Bdu16fS/mRg7+KTH943syzkbbna1uKWOolOjLAYAA7VgjBXXRQ
S11zuln2+VoD8AYHwhplbOMs+FapIvEDft2uZ4fCdEzxBlsppQ2bMBJWhzdgfP3ZrJSl5lOCiNPe
vwupz/q3eOKJV7MTl4GF4UHsDgFBcy+bJYWrmHiXNVVJ7N/pHMmYRcevX99HdLCN8Iirx36G9gFj
BNQosTEUa3dTyLFKDRewlcHrPfTKkmmliw6FdlpPC854J7VYcB5xl9JJK/n9R/cJwlErVEgK4ea9
2kGmpgTkWrARTIYi0AFZ4Qzhg3bPI5+UVGkgJ+yyvYrTX5EtqJBnJGe7yyun5rjMKcQSdD+7Npm5
BFvRI3uYz+IgRfaGuTGMloKEyzI+TuHOaPaOz6qVLUZw8LjmEc6YuZcDZqYpwU8IAaKWywZNjezH
7i8SOhJGS9v2QAWhMEB3Oh+4lEyCsBEt7TYETvczEjRgs5XA2KBDB5cjuYHiPkqxQpoyqy760Si6
YHCji4xzQOQnDR6YqJ+L174A26vktcIKH94jY99pIiqAHrce6HYIqDacQ0yE1x6/nRGuNfxQB6kd
Lg9SEOKsn+9yZB/XUY4L9NUUl5S11cEwC7dQAREPEOzIPJ6xpLwGrygPi7X0VThAPkuiJkJtuFoh
/Wt5pki0noAmuknDyiRxD0HmnOrZgtppvAiBShR1PG1mORRAOGwDEx/BRGgUU8mWrR4nq4n/+sWs
csKDMeF5ExW5wxdkysPRK4OKdH3+eAy1tFwob4AjhO5PADl4t6BfQOnuZEvII0qX2fxcVRpqeTC0
c/hiWqZX5OTgoONzy0k3+YtFlDmwm1S82CtbQSKBBTDKzXpGQfTYyeYf+d6WpQUxlx+OV4IKxYOn
P71A7aTU0goL8zf0oO9MfjZhCjTTml92xEsq4H3eMe2qS8RPzmx/twHaGtecBaIDLlu+t3F49vrY
knVfRcgg76JdZTnZgzZ7l4Khzz7Ctdyi2xDxXzRYRO+FQX2oxiBYIaCnivinYDJDqyr0zd3raLAH
QHqYe/l3SyD0v5L1lFrfj1HTwq95GZgTPOeQgy50fdIhR1U6re2YfFKS6V5/66fKeG/woCRFRwZ6
o6m4L4RL+1+UJ4UNF0hRseLC/GNoQwHNNQ2KDG9LnhSK3o+VVy3ZDVr1UOoiCjYvIqPhJXd7iNUA
1byT7T57sKRwyeHTOeJNMqhAv8I1G1VTkqpMtL+M0yMH2cCl+5hWlHgRX1A6mVlvLh1iro26Ztl2
Kdbejqysy+RRi/OrF0VLdpCsqd5JvPn7PGZ7IpQbWr2+h5HVdk0FUL4w6S1+2/DxpwTloCGcebV/
hB4hPnrUownAfBMzn3wmWEq5o9IrmOOUrY/J1UPTJzt4n8U+nc1rZs3Njr+KKRrbCjKAt0P+BSXQ
uISsjqGU9cV6novK0Wc2QWutqTiyFO/01k6qdSKSU8VcQmy710sn0cHIj+8g4hHrsPm99aIzoJGz
gwLjwfxqHgU62bFIqhzVByjTZ3aS1JVIYFAcwUGmdC0ACKACf8wNXKXJdPQ6dxJrzU01TA2usO/u
9s5rTLLz1H+H4hQhSYslc0/lXfTbCGQErn86MS5kCki1VdThm7LkcMHTw96yuQaBsO6pt8jDBT0+
1EbRU2OBXMfeY3sjSsASQbkz+JCB6y7x5YNWPFMgFfFKXahS+Vm1VXfpVfm9p22RM0TtNZOmZbyn
6JGZFPJoZ1e6/cCkhhLaeC2q8RHRfoaYQbuFDd4xV4afNPWZbZTmOZ6cYHJYCKzg5liuUlg09iBh
rjvLbg7kAmr2nVT9wUyM/P25O6vL7T2eOBKYg4TP44RmhCUi3hB94rI1O45KPgvdQ+onpxX2tTuJ
hV+LQq8Gk/ZxybhdYtZe1B+7CwzxGEaWOzBdm/OL+ei9de+DV6uFWAwl3yhP10WZCvLGIZJmKMux
dOxjHXu/d5GJyI0zTGHuv4nRodJRgER9bIR9+8cO1efJe9LqvZyv6BRXZGjutkmP5qZbpLZ1cmnn
eGd+jwPqLZzMNdNwki9XDfCiv5c0yX9kIJdy2cTjpER9OpHPDHMrThtt3+Foz91ZMZJaVIL7FcFG
6iNtw7w+n2mGPFiFE6jNvgJlbkSOA/KemauxkZgdvV62CiAk8zy7SjNfvA0iZllTJOLQ7RB2X1jZ
bqRT9EOO5spyVQS7lC7TJyNydjAHQi+ARX3QAdZT1rXpBnWyUoSJ/GmuCz3nMvRwuDkbPtzfm/J9
TKWIWlGrIhfUkHXGwP8ySJjVOnKWbMj2CNzJm3u1Nq3q7owcyYwItV0BDy0O7KuoMYDzoE94Gyv7
vEbvh7fa1/YrUOGixX2AyJ90MjQA3gdxBkMsdCa4aV2r4aRJSoNh/8JnSFn0Dgev7lZv/J1zRtYr
wFQa7V7EwtGwJA92oKXMiC4kmdqbFkUTpDyL2f+cLd7h28ghzbLnyOAqaVnGq0gaxVYSciAap0pv
62T89Tz4oIwbLZXfp3mo+oQBnZMpgf0U7jU9IdiMN6UQv1lNv4KV0AwmI+UoxMijPCqMYIWPuaJW
uqX1hXU9wSXQEkw8nE2a6teM3U2yJpJnrb/NswVG9bSnpgdKTi/xXF4bLFxaGWJunZ2W/lrwP4Vm
HETXC1jIE10itHGUp3TnUXqGfucytTMoEjWDi6lXYfTQmlrYaLGfXEvvwUNCjPl5WbrycPWtf5SO
iiboCS6E3+9InJ8oMlxH/CDuFrrc6c+xfZh4dq0hKxsrtxsMc8386oFHSMPWPJj4/3Gqx+ncWWIl
GqPw5Rlac5Z+BaeaHMXYADQMf68fiSqRZDn79e5p+Tu6trhMaGyRAWYqWPmBd3tVdooTCa+IPRWA
q3NuFkTZGJ2BgxfrNt7JA4taag0K3tsuRmW5n32MWyU83d9Z8v2CBX0YoQr6OcCvK9UuxvRRKtoA
d9edl8qTtHSxZLRcno5vT/YxnfRXiYpWc+5oFQSHJGlhukTLDEbcxujr14TQ/ovbl25gWJGRoBM7
1IvGf1TxUqESUeES7YQ7eueHE7LjHJjh6FvztnFkG5rWmtPhceW5iB7oVwJa55c6Vm3SISIHKRja
+ALPQgj5dsge6AaUdyDnwLtTASSyRiYHrps5RckdjWPtVA6Qholsopyo6CQy2q89lHlTarfAAdyd
pvyatZr7NDGyrUV7mjzzicjvhxVtKvOJLxXOxI2tLjL13f9xrHXErcNtmje+f/YpwL2hd4ojUbwL
28lT7+ijjVERTogSfHB79BCP6aPFXIyKb93693F7Q4tYTT429qGkhKLOfyagKw8WpmAAaScuhfh2
ROvTY9PBcBUtODUF1SpZ+O1WJjCrbd4UdlYZH6VsFOdcLNLHnEsA/XE4Ocm3xWW3xQBleQ9Y5uwH
1awA26FuggLZKmtEM3tPU8Kzf2D9T0qAjUtnxZBpAZPmwz/Q8I57SBepLup/keF9B+qVjdp63tpy
V0OHHTcGwpowaL04Ld1NyMSMTI2hC4rPKzz/UFiu7qP96wJAbjvUdrQb7qyMRa1px/J6+ZUnCA0i
kwqCQqv7slXYPO9dtA2FtQO290hygy1ixL/rZA7gB46Fz+oYOXULa2x6DoegZ7zwXaa5r3f7dSCV
OAaOBijyQtMcD8hzjRMMI3yqlzhffzHZX3/yzsWwmT/o8OXqh5UNkWicml2OGxm21/dWfcgIzilf
AGB125o73UrBZQ1VIk0ehSzDrdgp/dB5yarECDUrmt4F8Ez6mP7Cd63NDaIWIXmlj/NGONQiK8d8
vAJhkb86ryNXvG5pyGjRPAlNuDxbLEkb9Q88SoHZiJgNqX4d7PlUB3usiYfJ/t6ygMH6X+oWDG7C
wwyiDoBxvMFDmLVPsvK+uA4C3p0ctaN5+awZmpFYzXEmx0YR+TVFVqcBaf+Nd7W3C/DHKXnqkdCt
MLBbyhclE8RExfz1HwO79mQ9VipHCaKMmilBqTpEasbDBQMkdyyl9ILN/O1yx6EBmX4AApzUDbEW
u3Wk6e+tMKTzHhgjJ9WWM+LrYhROfQ3cJkKUNQ2Q9uDv4V5ksg86fOyBKqBCG55VIR3b0xiATZHM
yarTuDsBk5LcJpUruA0ChSnCLOB/ye0SGFTzJQA8nVP4GgFciIVRk7JfUrVc2sM+K5yGxEIF0bpK
jqKNnN2VfnJokx/+DOv/1cg7K0h7bD9cWeSsFdcaf6Yb66gjXsHOkFf0T0QqTDJv7v16Iz2gErqY
lQYFFQE1TCz8rrFwSwXXo7s+9XZLzZxxf9rtzSNVIHqTZbiRlTWyN0xcLFxljpyZzGYkdRnGPibS
sNgl1J6yVqmgAIz21ZuVWPZbzyA+sJQB44hS+MFmuSV2tOD4SJPpZmT2nDi86Ynhk6S4sh6rViVl
RWh3uG6BNHBKmxT1BeWS/IbTuoUaipPdmq0wpS2oaHK4kufTHhd86UZLtB12ebj1rt4+OBvLN1Yh
4RjzK8gpg54L5umT3KH1ORiDKrgitYPEJ+Ltb4MQ1HEfjFsdtbM1njv6SiEPjzQJFb5PmkIVq6se
+SS22i12kwTdcOyYZMAKx9h1gFsHT3UAb87iTAQzZdcpkbSU9R2gccxpmjCH3QBw/ZI5uLLXtiTU
dB5MbNQ5k0EMArv/8jmkth/DffU7NKnkLMY8mxJxShqy+2lyoj7EjW3TaTo7ROSXVNpmSNpk7Dc9
Z46tRsCoUeEjYz5cw+Oy8NqQMHLXb4BMM8xJZGfUmAzr0O+//+EO/jWfSpPtkk+dtV89Ui1+xNga
kug/pC+qpyHY0N8Pe8ZomIcLXS3vMKiO9qvOCEC9iwE/RYxfdAipT1Td9EGfC2QfMDcW3ddDQ3yA
J44B4tdm4b5xDdjSh6LVRhRWknVcnCmTIzIicHRm4wkjYCg2yciw3GZoTc6jTYIQgyBfHJOW8DcN
9Dez5xlA6JGx/fc22uoMUfLkWhyAtg5obVlVVwE6A30Ar18mEj/gdoi+5Er5HFv0hNpQ8U1lgMQ3
SMXxp22rKpPmfgJETxZ4VERnnk6lRDBjsbY7XI8cCGsXCR6sS2N3pzY6LIJIAk1KLHtBs5lIzXP1
fJETP4RjfeU0kBWOfx4EV8I/TvSzv4uZF9MXT9nu8WvPKv/Sa509Ys5ELWVT2jU2LeJxTpZu6t+o
Tzk+CHcq6EomBBXnVvbKxjg371qS9UxoTOVum5Sm+sT1g6JNZjYgNyg+apuiRRs6Ms5lHMdVBwN0
crUgBooNasi1U3V1gPDn8JSqrn9+qnLjzVSvn8lwAjHR3YGPJZo2Md+QG/L9Gx2hefnA6UanmfAa
/Y6ab6aOY2DVJF5dir5NYXywcITo8uqhd3RseLqd/tHRGxpHNGDVOEneAsGTbQ21uuFNfHVCsR71
11qTV6oULNqu5AQkBflGNYDCX5R8MeC2k41LwUNAexuZTG84nP9cqcUMmhoVurWZs4J6zuQg0iCI
4Xml9Ujxf3cg6Fk6zo6XOePEjuMs96cDlird/108dF9j89sjAehKtPvxBDXc5u8ps5CvQt+sn6AP
sfIStn78pq7dJGQmMYBr75yAqL5vTnS16NO6tul3ETg1gYHCoGq8ry/Qz/oM+uoqwcS461A1qglS
v8obHb4mmBO1pGW1k7fj5OLwDPCeVGkBVZXCSMxvoZlx78ih5bBmsH2WWFSsqUgB6BN6Rmjfh6Tf
cgZsvNSXzwVtFheETCzf2gt6iNsgyvLw4/0vXViLO90KL4qd4ZQ/F2HxxH/3einuAIGuLFi5wWUO
CRHfRPkgS5f1fbsrcovvYKDxUUYKLA6LmPZUeCn6NQ8SXBMglU/AtPQPObS4YD4V/uYzcBHlSiMd
bWnUIlrLXFznuwncccNBCHkKoGZBc8FMmIKc8cDB7mCJflQgrXzHt8FuSN+8JovopACnKJmdcZho
Hv734Ir154va2AJh9s/nNl4jiJg1tqg0Es0ITvvxbVi34sYlvUf0eZcw0HsLhpml4YXyKJT/uZVg
YVAdEFTuN5KC560ILiC+pvmnEQMBKpKvBLm1RyEpjDyLEjnKDqyEOcjfiYUqUoTFECLsdw0YkInQ
5lXi/kfLR02YOTgBbmIxTFPdnMYlAo5hdGcXxuuczFMLWhiJgic1VnlVdNqNCTw44KsS9jSUeYPN
kBejdC3nIMa8oS6Qu2mAT9j2GOzdU6lD7+AGIl/ZwH/UR1bR6Hv7gloaThW0OEQcWnK8pp4te0tT
n2/CzkcaBfPF6H8kkbEG/bo9TXEM7v8vnUdlMtTf+vu0/9FY5tAms+OrsPbldvhEZmQ67GEgioOT
IHMAKS+Pbhh69LgBFKctiEJNO2Ik+Qz9MOGk7ecQQ2BUZZ/HoRfWWRtT5ZnQ3OUY/pqtGdSUmuAY
px4XTCMiFml+MDmpkwQtRLy9+FKGhuflDIgXSyrHjfqH6vj7UDWuQI9QtemTer6JG944mtyNysf1
/PnV2/yDhTdCpO/Uu3pVAFikInCmN7GUHBS6nwUhj7iCXNTztB78HQKbAQqu212vcthZXlLRMMfA
l6W/vgIIsUfNoS/TgHmD8BlGrDrp33J4PYKV0GuhiRr7EkxifRMzlf0yhkiS7RNNzJ8cyd0RjStY
YdMHAsSVp7DXSA6mVRPfpycScSiSL9KSxSSdzKhOVbuXsbGY+Srsun9nUt/eTDMYHg3+vAtljUt1
fRmuCfAE+NYH4f1ns1Ln5wDg2n5dEfugHsl9frr9wlCVaPAx7FwB/RSH8XMBLBu7DOf/cgH32vMZ
XN8AmJRziqMuZxhZ9YXSpZp7Jn3csRsvOEyqP9fum0oQPrywhIYzRP0kN2orjnWi/iWbTDAhK2aG
NE0/BiI/Ijeh/iKH9fFvZUQx/Yfjuq9FY5/u4cbwMspoibrr8heZ0UDY5AyfIVyU0nKCBc6Kep2I
YcjrDzuhmJgebDFUViJ3LeYy07+gyFjosWRf2S9BQCdt7kX+NsiVy5FibWwmJzK7iiMua+LGsjsh
q0piBInVKxOBqaee1TrTLouTZrTCw/IP5odUUDbWxC+euowfEtb0C8wiUKeMxmkurRKS4jW49lLV
JNzlI3zjPBq/94I3KiFRxxKnJs8M50TVCuv85PlUx9VuSEX6tL5SZs9WdxuEzP6bcoUGpKBbBepg
SA4+dhIaBkSG9CwpO1MHhpvsPg8jNaUAIHCX8dNxICBF7tzYxnPpSNsAwlvDwiGdaM3Vhg2MBUl1
/2zbX4NA93GTTBi3YPfHy4Db5FyTc46auyxkAWHO5I2WbjEOtXYPIRV8971AueypI3qqlzC4JjSc
quo2lthiO51TUbYx5+mxYUs7m4p8mv03oEO44mVRPTXGxBVlk2FuM6guYpQYYmnmsPMMMNw8pB0c
tiPoXfjeG23MGzWx9uAOJ/21sJYP3CxeKjYlE3AywqW2OsA8bP87fWbfCEI7He2vB3psUwHUKr3A
9OYUefMRS37x/qBjHghRDVcmdlVZuhjCEl86TsJM0ehNLUVdETeAwCphpFa4UUGAhS8Jc2+9IayW
YY4D9rEoxbijBYscZ8F6t/axHONzkWRO6CtXQ9WtgPo84IOdzzdJaiKodypdlAg/U1TMLozGNxaQ
lfvQo69WJgK7d+C06JxZoyUhmQlB3AlJqfwLeLn0FL7mcODXvqd02/OPw9Rhx3xaq+iDyfF4IKYO
ER3vhfS53nLI/S5Nm9AO5a8Sgb2/WshvFmE3nRKumqIRh1FZeFtFmpyYcV5Izj8lxOn2z1DEznsM
088F+TldmIi1QmZBKQfYqtpNIXCqs+r8nWT/qUKdPSjDrTHyGDpCHIgmDgCNx3M47EMmu5yX6F5O
PzZbjLCc2phD2GSWHY6fNjo0+purzusQK0bq26XeEmuCShHJIol+roMt2mT0Rj/raOhTzwzo8QIQ
EaUlWJpEYg295nKSanin4N1SG29Pwr4OpmZOKAefOqybmoZeeBnq+JgooDr9boiVIKSVRPmKap9q
XLP7gcNAOKk2/XIcsoqbaShep0iErMM2XJLZ416pqAb2GJYyo1QDpyWOKyhRo4LujoalnQTgwq0c
YGxtCBKiyupwgQb31AKtCjIdI7p4SnadOi469NQ3h3KjVK7xfHHumBxBJXy0sEexGbusYSp/Vdx1
hnrcLjomPoCqDi67ioqp3PE9cRTy7YM6vEX0uralqw6xDl/m8gWqleErc+1DAIGqVorpYTnEAb5A
J7qB7nL7kkfNTUgAbvRAJnHKt/xQ7IDwi9P9VVKn4lvQXuBeGMOERloMxUNhvSE/qc+UO4zG/S3Q
ts0q3EPlBOgQ9RzTdGNjxOXFf7er218h/yPDkzWdnKzEuF6B8I98LAtjJ3r3xQPLOD0XoO4P1vJ0
aHDmwchzlK5z0J8fadOMARIjWXDYZFkBJ3BV193e7Qnbbsbk5ldFwNNghu5h/izH2ImR9UQLxtV8
kdtD39Oex5kwmI3JUXCMDpiTgw79n4+JQs/1ThpDSyhgfqhyvlPsItagiUnTp7m+N7YPrusntBhA
JDrb333VV+igOaqYX6c+hPGre+yuEICt2RuRvBkJbojZf3qqMiaRDOJn4fqfuW1smrxi/NpDJTb+
aL627RJT88b49yXEwBlyrj2I9MoxaVhqq8gRvIhE7ZA+RUcm/f69QlN9+rKCgcguL4sOD2Marw++
4cY8efYKPos15gfdYKKJe0CNRwskMrreuswfueeYVB2bs9xLlOg75aZ7nfwDJJCGvPnncVZbSUnd
YIfewfGsoE7DtNyWXfd4yItdaiN4agiGFpd7TYEnhrYNAhP0WnjwosWPWJkneOqbtSW7aGTjH/sX
v+2b6foWzcYfM197/pseisRAZV5aKL0w99Bu5aFNXt/qyK9rL2aSBlTfi0TyJG5rYIbUdG3RxU0l
EQa08mlG7Iap5w05Y0rK5C2XU6qFJVNFDZuomxNxd/2+WsLt45nvTvFSo/vn0kr3ts+yI3TgKItm
9OduD08EeBvZyndRS/TkHjplHNPFbk4x7TguFp2I79Kvjp6AOwnOxbUz5O5ABH/c5F2WiZAi2bmX
j2Xl7u1TLfSrEvb1SlMo+ssG5A1nMAqvaa4Hssar0GKrj+Tj/NXjbe8NLWU9T37ljyBZS9e/RCKL
fl2Xnej/KrLt7WcAckoHRQPQ2gHhs5qJ7klgFoDbHoyqXHOU1iANmM8c616JSzB8+WKm0lLoAyob
J+/Z0QuncXSqYNkFgkArWR90tQS4QMH6Z2UNe9+JJpoLdJsVWBpZaZd7s3wpm3nhnZYjRXyD3StY
7so50w0rTm3/VZDN/Y4y76HBOXJX5zZQIveXklwYoACXy1vBbA8rIZUfgWESVhQ7u9GUVsy+HY+T
i3/cVo/8khV3HKG0fcirlhQ1+a/qgIFPPW3mSdouAC0U6QetYCXGwGFNbBGI+4xZGqELhHCmSj+P
lx+lpxxXbA6w/XIRQM/IkHhH1cnq+StxcK/XnYW4AMnm5Tnjqa601472ZuJnfEgRKHCRYl6110w/
/S0il456c1UpTDPqchXd9mySmdY59czfq+Bt5ninVC35Qx1AMHYiDaIZNUk9TS60Gv92/DeDlISd
GHck8TVZkiEPGlUzKktT2jsZANPCmQE2BZgp6It7/1CYUp3yqDC/dM+5hxvhEoox8WbgB8zr4O5H
RtxMZGke8mLscyGbezJUKgFqsV+IIsLYK5jNe7D0bTpCCJAjC4Hgj8C8iBKH3BT/YpExRSbWk/Sv
hYwMuHfgyd/Kz2Uuez57hHacDn0TbayK/ir/ln/zjTZl1RKJoZjC8+t5Go8Ag2TRWPv09tai7GyG
QYoGZnF7D647uH+k91DOoeF67o3eWUz3JgQYH57Z6FZ67oAlfcR8mSoA4dUTYlwqMCOOW22fa/s2
wtxG5/MhQMK5HWnMQr60K6HRLLT9uwoI2NDl24UOutRPzvI2f5ghVuk8EzlH5/k5eUcVjoMeHBbg
FpLluPWV4uhpD68I0PNU6c/2q9N4+CYtJ+AQDQfP1c28GVn3yDikWbNwTKNJvuSlGAsadFAAxbhN
g5tmLeZTLbdddCnG/z5H68ClXWYRKcHw55Cd0hLPzFsjiD7aY++9DY8Izrn3MCdwh2yUYn0VgQnk
R3PAp1OLCCXxj9ck2Qc38tpz9PH1YH5w970m34C35HsClDJpzhDn6aC/WjnVTJZxVVrC4+p/R2tS
UKH/4cJJziwUHryaIwMoZGeXOoFi7Jv0anYOahhfJJTcb420Gt008sVFDPiqWBG27XsSwi7RHQN6
SZZNLcRR8Ma/B8lYLJN2etDvMmBaWIy16Kmr023FeYL/SNM53SaDJkzldqJHrEXXE7/+sIKu5E5Q
/vuqsg6MAnWJmM5rvMMW1XND1x09myErfFy+ulnJmjiKqeVLyNkPNT4Wrut9hKN+uNt1pWTy5rrF
4HJVTcOZSYxvJoxkreJzwOIr43tzJGYCpOaXLIw0G9C0Ll2RH5ds9ecG3JQKWgUrI/B/Q4VdpGgi
A5r33BbshrDDGHNzJWFrxdg4FPdDbyBXNjEZNLSSU4PtLKNR+pjnMfnqTrh4pE58Dud0sW94g72W
tbEMEo3Yk8pX3LM0UpotiWPGFLGwE+Z/AwkI5UQtMgzxwBxchMjFkrAq4osZHLkBVQarI6vlVj9W
To5z74trHQNtbDTpU6EBI6UAwsb/YAxnu8JHfuMFWKBKFdbE7qYZ6VCFjh4M4GXqZuHIBY0EiK12
+5LiPVrCkvvcmPwBSUTeyYYUEh6lQvLOYAFjYHNEbMSOhcnGaKq2O9cdLAcdXUdKBpnEuk8NNS65
uCDNdv8KJ5rjGpaf2T32z0J2b+oUbxkG5yRB69fs+Jw9xxCGvi3m6jynrmzY7Te0TcQqS7+ZkpGI
PSiDKXGwp3bNAT7rg8xgSok2gLKvZ049z+0/5mOHsF8e/G/rsW8M9qgI6vcFLNCSvAzJkBs41Nkh
qgrA/SAFpot0PpjygXcdnwvvM041AaxehDm1we7P7u5JAQ+jAMZflBjeiZu0VNYst4QJI4oHPn/Z
J91OwAkpdiiHnGz+AmZ9cNnCxW/Pw4mWSAYfhtiIKPUZ2xIn3cCMSwceLnvTCDxdYHS5G8G6OlEj
a/axMhWw6Dj77SIrPhN6/X9ezuIXrfe1Z6JzJ+hlkjq+IJLktDBukubF0u3sYNnoymGmgBsxcIZl
5NCwNqSdC4QDWCsAGWmRDmsJw3+s5QM1G7hr2tcnx2CNoGT7/7+RO6/waBDKUqeqo/gWVPWGS9jP
DKLj0YsLP81yESc3O2RSzgqz1a7Gwhs4SQFkhLe7Zt9t/JM2mxDx+WN2GzlWRPZ4SopesqdYIlsE
z5cAI0s4/MjGdtqdgDeFR61yMy4DRL9BG7yt69Fv3i0LppJ9DMCiDDVBBAyLHtqgg5HBtkvthNTV
C2lL5okDMIm49VVbP/Nj3C383hOCQ8XJtXYZMJuB0ktSbIq4Qn3tzPGZTERWw4lkzrmbAoyzr3Tr
1y72Wezt/UAwJHBB/eHJRQHWTkVIoy+nSa5o7t6Tq4r0fL4fOufwV5DTa5yHbHw5iv0n+fHiXjou
nc11ixywISxYCtGxzqcUIl09SUw5zn/z6wflli9svxCcOOozQgBjvcbCC0x5SFwWXOi5pA7msLyT
EaLEaoW0UTyW7PiZbQNr60ZR8TfJrUM4n2uZfWxYh6j/Gw9FYzGwrRAm7S8+pA44AqL4dygGCG5A
MHi+L8LF/qdJAonrttIdsuJvd4eKynDsBYO5MHSi8oJ9F/Kq2eGHOhLUs2ymbqhWhbGpjmpOXge7
lPXBzKjkktPfWB6BMye18OQVzo2OlCBncFwG0MGoz0RmtaUfU8/OPbWispR8JxxcHElxf1Vc043/
9hfIInk+9coRtZ+uHQA6ShsuZxiHAbNOkW8cS3Hqk/H5v3vqUBLKV0BZdUJNXGfXN3rNISGktZEM
fBj/Ob1uw2vVa/nMR9HbsSQS7PhETnNkLv5zyMxrhZf1deFWRCpvU/x1BxVSW5TKZFnU5/4ynetA
XmefEnvKSZ+V9tJUSYPPVcIHesdNSGVrvZEXUgxpKznCqoJz+wbzay2/gYym4Upi73n85s9awYeh
d86Sw/8S6BcwAx9hWPKtq+6F1PgesX+j0qG8AVznHDckveBYn8Me6ObwrcrsIsDYjJ6R+UXMaLV2
21ObM/5jZjJPdGGrZ/HresWv554I3NmdfCTtIGTCihen+aS5j/ZByLjPPnOaZwGlsO9yn5wkZ/9K
0OwEcEuW9VQ5smL51pDaZ52V5jiEXDuO7IPEly5YrjBEMTBifafXqaiRbf0YZwsDER7cG9pSqkxH
IwXWMt/tRB6pILla95HmCtzmvh8T7wtngul3SeiGq9iL/q94/M9NkyJZpxPs7gbH9fyvyzfNO7PY
Q7BEwVmeZn1jnrlX9c3Cizb2klfBroVKc2lYjVvMmy2PtfO3U9PEoJD17ofpK5tfyEaAhZJAnzhN
xht6dQGsiCSfsb4sWIwLv4fpdaYzSm9FDbMP6gARLOlDArnsOs7lY3PnHWFuLztE/Ard0GebyDJR
+CzhCNnVC1WOT5rDER9AfbNrWvLo906jKGBHSdA9pNIuRHEShPKr4VAtXCcX1MC2GOniyNjULr0B
ujA33ovu6+Twa21QCVNEKRJz1BDVouVRJhLnmcJjCa75TnVQZ6srSf8kk/50G4pkNe93KX2HsbHp
ZORtO9xd0e6U6BPh37TuvKiyJ5wxXZN8XWmG28+eaOcYWHXw0JKI+Oz8sOUH7hJo7tFw6c2Ju13x
pdGcHxRtNmSRt2qKiD9xfUnm5qp/50j+eZ7GL2lbAQIBv66/0MpgdKCGyDvm8SwpEuD25xYIeAmM
aeU6PaCQKZ5JUGKXPHzvvsz+8KX31gGIX9DrzwrWO7jddz+F4EqVn6aXGx/OAyhY5jZXZnqGnCN4
IQb27i76+oJ8Y/KjHMABvIMFt3NVs7Vo4a1M/bz015XF1kM9ii0cba7gDJrHzLllsJ+f3ErNn8f/
zRfKH39vGLWDfsJG6zWfFX8h3yI/3zdvFLbRSfz9B6eFdEKHB9RpnqlC91MH5BhPeWLZX+TIKQ4b
9rapCoNhE0vdbzzBtK9iFb/BT+Q/BaneuiWzYC0w/gkUVS9gPf6U7Ro5Bc8U+qvt4diDxQQRHV4L
hMYrwey53GrQyel8nUBAitSrEsvk87aydu7p0pKAGhB78hp319jB7zhPjYP7DuVBhk+2Zx55xvjz
qq17hVO+Ccp81mLFStvQydUaWchJkTH6RF8nSjlXZ+85w+PsNbeeRovbqCUIEqUX/lbAJzdZSe+t
xdMyvs0+K+mlurgIN/xlqTtqj3ymRPuKzjUFjkLriNLlmLgcY6DWARCk5qKnui4m63AmGzPO4J0q
hecbd97KrPUXTUxtKBbrBfDUWYP4+Vhls7j+/J7F8mzSF6EwcVi6ddBeOYrzlG6LKn0BPejq1F2V
bFxJkg+kYDykWGcSgITshh09MCpHN3COmL6Vn8ldeCfgd+iNXt8LWnyUwWI7TMsCXQO7+zF/Yb0J
bIk4/zVFPnAwo96B+bAIrmswapqT09LjQiaXv1DLZ0MEMqISgOw7R9TwVP5S7hRc8EcCwVVdDa9H
YtAPQDCSEyD0eD0pSC/iuvPUd93d7w/gnUgsnT6EXxfnUDrO4jivIpk7dZBBy6U9vKNL6TwGCMcE
WYrtZEh7e1/E40InJBPCZiBZWNgfqNw/ghwsAZpQ//MjygeqnKB31l1tqAfzPMq5UrpcBuvgneyt
Ws48lY91EdQtQNylPpFBzJN1Zb8B289B1rBYJKjpa2AKvdr3kl4HamleW478pN6IZsBm6EXJbZ1R
jwA4JFYYypVQOxBmRli0/rE0xJIf4ZOxcp+TErisPWUF6KGE40w5Ztknq8K3G3zJykzzZavhZQ8o
ETRdmmeMGUblYSIqFNWN3r6Rs2qi8d+nMgomtAR3VKb/xtJO5cSqqW3MueeGg2GRRWhgjAtbmr1j
+ca51vV9n8Iibatgq6c/JXBPywj5SirmsmD/phXh9jtNFGVg43L8atg+DNLXqJOr7CWtSqy4tcb2
prEjR92XQ8TZv9Oh0G6Itz04cH4n3JCs0WwFNJJBvMu/qAXvloojy6V23sKYKJkbmgPDYUKM+Jrd
4JOvZosPlkFZ4lmmKwtESGkMajYsYrscTRQJQNkkWyxkj44iJ1oIufUZKlmraSF1Z5Jk5mfE90F9
xATTREXzWqcifWqpm+TL+QgMwfJ+3ZBA+wIpICH1k/JrLuBkQ7iv2DEuq3jKh8PE0Vg/Lpy0LGyS
HIzEF4/Q26yzzEMO5Te9Ng0zzk8mBgG5Eatbe8XascVoG9yDnEqk7lo7U05/Ty2+UfjQSsbUnb2w
h8ZRGfIhk5q72U8aFjbqkvLzNpiSdYOlX4SJ8O5C7VUEgTSMxSvcQPDHlolGRFNpvYvGRpbRKU22
D29/g7iGCLwtDddDf2wlW+luy8nAuUCbphJx8IPUVZNSTmQbiyEBTUDf5rY74E7atWAgT7ZZkwgI
JH2rAgsu+XAoFfF46SZzOfN5ahaxkjK+OE5yQEmFkbf/tm+X5Ge2IZhtHjZVKLBtKC7SGnfWuPZK
hxadFSqCP71xbPJDA7RGNkurC62zMM2+BkKXRrFYliHqvuWNuygPnYIjfh2xzGn8YwYugUOANFDQ
90GnDFqgyO0+BoVcOEkCeEx/ImLX4an0TPjAtAKc0DfWQX7sMefGlDa1YPlNHdobVhDZOZy0qVIR
OY3bFy8foDctQ76qidleDaiVjH0O3F+AWlW5mAe6RN+1GVz0CS9uEBVCjEz/JQ3LQg5ZrwB6vyZq
jSmb7nODTK50OsmcJnbKUaOh7NHismTBvCr+vdDUcinZKEz9MemN/JbLlAHLjpDckKR9/WTJudyH
iE7ozIZADTDQ5lkM7ZR160r/5Kc52hyK/lfmFX19sjNc23MXhrB6/PfdRWzapr/KK5rAZvQkC8iX
KiNU+2x/dli0xVoC8cBSWNB4RmWkFjorFnXRv35BwbOArYTGAeUlIXvbG4lQ8EweTl+P9yM3m9L7
+dFk7U6rJkcK4nHTpI2/p5EGXaWANynpibR6ixuBfAprVtPu19P9/yyG7anIRB5wDPUkKMtCuFYZ
F7V3ku4MRIMp9/sHrqDsYtNPkoCpsv70PoxPsQXKKYoUnL4rp7E3Rz0UrTsj4C9KD3drAH5t1Rge
Ed3yVblYORLOXtwSwcXlE5+H2DxabUZg89D8zErwJXMX7/FQlZsaMCNerGIpkWqMs9+phb3aw7iK
mBNKAJM8aImn3gnN5kg7B9bSqm2qUBW1iEIwmXBxX7KENlLpGEnTsNGfIMcldnedggb52a5mfbwf
8+X16JCgEZ+4FmmcTB3i21PdqbWfGe4+YTLZtRvrr/rfLTUYbadAT2N2ARItShBIxvA/C6wRtlzH
a4N+vU3u6p/OsU2R2sb2UYJ8Vkxj85Z+ybu+q7aHbC1ztw1uvVSmgkcjT3rfUHCW/ue/ZdwfGY+t
ErLu/pxpC+BvGt2Wa+e/VLT9ryDRJCrO2lmjbcdrPbhloR2t5O7YME5918Cdqh2Ad8Wl96Gn2/TN
+hD39d7Hnd6X6rPnXw7OijZS0GgWxIYQGFSotQ5CxHZMm5mqPThzyi3/CGV/35cYDEN5pbCLCJeZ
Too9dGsEN28ZlKYEY/I1ktctLcVGmqJqY5eYdXUfdUQFHaN7G1lWgCvOtqzSFTvbQ0otfw3nwGxb
yOVNRD3sqOMdQXQc+O9NjZzB1aQqBK7rc5QQ+iuu2pR/8yPYNXUfsz33bScuwSBDwn5vcv0C189F
UQVD1UUDBJXp+pBxroIrzQxqM1/DwLY2LuZEMhSXSdROWftQS6bMxHh9s+Nhe0j+dTCMlyvnvEx0
sr08R+K/1+ybPiSXiuJEG/BFCvbZhxJFVgJxviRuKMOxIOPx8zTBDInbBscHaRIQ2qUe/DgCCeVs
2Nx8khYU1uUNYvDAK7hzPjelkrF2QTOQTkFEQnAwG0vD6jIjL77kcnD+mrjUQ7rsXR5CG3jeyL51
QGBxEdCKgLvB1zOeGzfOLJoCUClqVJ8WsG8kzJ0gJUTC5NoRwTSb2v8FiUhGhK84llZTpy4Fct55
jUdTA1EtpZIw15hqtTZ8MfSb1zz1TMdI00UBbNvPmn4cLYhf7jGPKcZFtj3ZQG0CvEYHdE7+6WLE
3O9Iey6DzRJZgisvAJ31uAeVzSsPQYbbyvYI46HsY8xlqih+Gn9/O0QjCOSwcLqQ9mdTa8qrNCTA
2d/lnp3S4BiBR46npV2XuuXPuatjrk2O7u8whah+K2FNS+VTAiFYDMas7N6EwLUx8Ae80EL2iojd
yyGiIS4+Rmo42jXEPqD/t0rln5Ol2zvbxveUj+JRSilYJkWeXZU8G+qAE4ToVYqQlAHbUklFddC2
0T2ZGEJhWdfSUKpvOdB0WnmXA1EkkR+e/tL8rGL2EIE4xKAZqGjxL1BD3/1/UY7gvRWLbHfX46q6
p1Fzdhbe9symSMtkh+r/YzAqPO/HuvKLcUY323z8KVVveR7T51+8gDa/0fGyLSyw7YHX5PhVm0Jp
PumgeGrZPf8/DdNC+esERHSMZdrL/jTs2aPQGA9b3QQW6+iFE48ro73i3L3DCBTbectqE1OqSrIV
RynifCTWOoADj/60qNCJMrZV9kE4ffVaLvoA6S/oNhGCABrzix8F3sbjQ/WbVO4U3yMnlnx7qKfe
taCgTNcYXH0Jr8eWk0he8Yzmi6Hc9cEBjI/wd7eISEw9b2iANspzQ8Xxp9EcJgg0R1UnaIFsrgpW
U8uVw9REFVs5EhexkPd964/hW5ATqcLL7/SVfSp78yMtlTnmh7On+gko84UadVC1S9u6vGeIrETL
MBh+K88+9zldSC8Lq9MY6zYBcqFKJsAspG7vi0BpgpAeRsLW4QyOXQa/QjZdFG7O9j+23KOZtp67
/i4sFVH/EbfAQ4a26QYtuIxxs31QeTc1sqeKJea6e45nReRyGb1nyNxw6jh9mttzuJaqSmb5WHk/
ZvIDyBPtqhiqYX226/lXlsBxAtz2yqhVeM/Grn0VTOT9yfDlZOdZ51iaVVM/Aqu7vl/Ddzw5Qppj
63ZtvY8lY6nV0Vn72j8cA+M3PjMrjOvtE1WJcJ2Lo/8CCkhTWM2zdzZB9SlXuyc33TTHSMNLxNbx
qCikVKSLgZauc7/zjj8DJWLP/oIwUKsE4nqHm2oviDkyMeZAgq6jM+4jcLNvek/oPclNyL20OesH
eQ31GXtpYcoEJU6E79pF/lPhUVN9jZPUsvCSsQzMYhhfAsrDoucmjleOgPcHmY5kWwzNV9OouYCe
SHPQ/UAuS1W7pqlKWeDwtTlV8q6Q+09W4go7l5w7Dp608brirC3EWA8eLef0KnqBOqvqa4Maknmh
Uoeut6u2s9sbf1yXG/Ip2aP+NDFhYUUGCZHsxXMpCIEb65A4zkp7OfjcSFxr4jwNVSsugr0H08Ih
BX/8yhFmbUmQGiDmN4XK3lTvGM/7HlVUahgTy0LiMlBF/njO8/2CgjP4EsVYfTRiYWxPGFCxTjQC
599Fuccc2yFqxHCMBMG1PZf1cHrNBN+9iJ0gfbmjaCS36tk0LYXWr8ueoiY3Rteahy7H+vqGUXXW
hRVcDI3Cn313bY19bDAXxakJZHtb4APmLYOiGACzA44hgUbUEQTYan9BRyh/+jJMCvkumw/f/w2g
oWMAB5mBlkQMGiykjht8eJphuhpyz/XwR5DL760psiQwZhJlVZU9I6js5RnJuZRgApaKi0a84yco
shAanjtd6sE2jZk/KnkSCV0RjRxh9jk4d2cJt47hn7abrAXEVPbX24sTvfvb2GxUcvBRUziziqGh
TYIBen6HQXVNOKD8TYj8YXubty9L09ZipC4UCn3aKz7tCQG4qvbN/oEVJA3xS2g2nJM0Hj976CaI
9X/1DHkHp2G2nmIZ6NQ2cc8/rQBp2ijO6G5KzhHVuK98B87m8jkmHygnwDFXNlUOwOVnDjcWEr9V
Iqj9DI4C1FXyjQ7bSAZV/yu2Uzo5mtiqTAv4WTP+Mo8Hq0RYA2vj6RdtmibT5ZcsR2+j66uNLtHX
gc+6R0BU/KL5awKqgsBQ6BJzDaAKMQDzex9hxJ6Hc0WLB6LLQSzCDbYULUjcHaLAeeIgcjNG7168
DG1RSR03fz4DofWbw4l9+UxhM28O1MXiT9yFvlzW4P3uyoq8UOqL/nl/fetqLVyx7G+K4FIcnolm
nPJEj/5wIko/m9v0rE3HjxukGAq1LUpwcICR2G2KXZpbcILhzkSzfIPCJ8At+forDiHYV5AzFcDo
oMRfOG/dgbhRGB1sNFyYpQZTZtfNaunxj1dHIrKwEHawKl8ffvRfWlS44g9diRShRLWh+jMxDjG5
gpfxixsJYzdqQXZRlnqcMkP+PfuoSnsZMPmp5yekCVcjfL8qnNnow+sST8CXLvRDF5TDzQFUCLh/
TDn6ewJEyZatSXNymhjVjHLY1A6ZVrrcEXK0FSegkq5LiVhhIRVIKCWnzCxObqz9a+4WckFEyzDG
Kbc6VY8YzHJn+OMIKTFAdJ1I/4y3KBFqEEDovyr2ltWNoG9FHXYoc+Upt18QKOMGg3tjG9ti4sZm
nRXRh9BJuzgaTI5B2tSTyo1WhiPLg3QZbwqDs/N0HGWvIxn7WCKFTzVcziHdQaUyyfk4ULA1etbb
5Ys2MvXH3h5ykXHfBF4kLJgjXVMiDhz4glwJ77OEJowIjLBAwmhRGRk9GVAzJSqf40VLRQVxy/gB
LO08w44O+BF6KxPnsIpwwF+x28TvVOnxroIjOIx1ztuwr23pQrCGc+b30MkOYqnD9c69sQca6qcN
ozya2+67ddTfS3Ic7RvSj1+5r7c+SQHmKfhJ+lv5SEsO077uPzC1imQtOiGhF/TeFRB0sb2jhwr2
YeNwicHbLNEDLihZbyITLcXzoJjHOhnnZSDGclMvOY0/496JZ0pApV6QVv0RSTHN+5zReqWZHFys
T9X+9em7NrURA0q4+nPfcsFAA92lKAzwF+x2K0kitCTeugO7k5Z4n34aQWs/KfEwgv7YzZWuILg+
Y32QZx2E+gBhYQd+lEVSNalYg0zTTCjFjyKAB+PgkHPEtxtVIapRpKWEIFIMAggf+IeXWJWl3Veo
yoBLwovIAIIIvbBwFL2gXoVM+Tjs5d8wJYQ905QNAzBQEBE6oE5s/FubWt1vA78mrDG+M9sqZ3lt
OmgMnN8PRVz4SUUlREGNRBvdfLoR/TwpuqlrpoCnPntts7cg69YEU698V5sOF85VIJwQH11jsC0I
I7kv1VRM/gsxHq84nrBLyN3teAfXRcxux5Ax+9H3gAa/9X1M6qX9jfP/achURdKFS9qPrpaiPTQi
o5N/U0wA22tonmey9D3RMIzRLgF+M7w23ppaew8XsIkJ+R0Cz+BkUZpWyIt2AJ7qTTO6a/Om7BDX
aEg+SpGmVXqUkv7XD/0h7cjmPIWOMgeq6Hzy5CBT7TJMxKoD2ivMsFYtedVL59/MdARE0YFrEb2i
oMzQMo9G3mzEkhwG/LMsLChCOG0HULEn9Avg97lTXyf0bwAJVxhHgbI7/RK/UHVZUoTcwhIeWVfd
VC1BMay6edxDTbd5Vqfj4Emrsens+EKiMWV49Uu9QhaihP4mYbg8MZTGFf6ZnSb1ivl7B9bVjdvx
47FxdihQPxVTPxW0/Mtb9KgVw6hcOET+KnQUwQXNxWWhZLPgfbaFNHXt8ABFXyGbRFNrNekaHW2w
vybiGrPaF2IuiXn3OKOrJEwRUA4gwkoP1LvlbAB61FWsHj+CXmpmTiH1TEYB0uMxlI9/fm/nU7H2
UJFOYIJ+MBLPDGSR6p56bSL8buTh0v34qusYJND6XwhITnyIJVXTkX+ai9tFMB1w48ydJ1BD+K8Z
XmZwr+jSymWpAOHKnV2tIVfxnsOXHlwpNSLpCrfrnAwiQtPhlUjQ1jJDPRRudOKng1vwu/FGRqFM
dsSgZaTd1oAYbG+AC2oFhJn7ZSZQiAuJPo/Ah0Xo1Lqps9NbRU8IVFCuaF5Szs2bZ5/QV6Vt+sZb
HDmWS6+KXYOxfP1uRTsGmJ/xI95WKZdMsi6369rp1DPInK1VqZxyBI03zcf+ZAGaRsxCNSVu2/ts
WpHUADBJCaOQEwUexJSOT9QkqOpE0rG8EgzCISCazS189eimDLzYdvrW8wxqTftoJLhkN/A+70rB
YK6JiMcRkHEFp9X3rMWa6bQsb3wDiY+aM65eW9r057W57SCVRq4+CgihRNmK0JKds7rdd+XRaNsr
4D6lPNd1qCDfJ0UvzcNsYyVhdtlTe29UEx23etnGaIc1RMEgHR+6TdIu4980wOkwuIPKat/AJYH7
/k/m635FdNhWvIxJvE1VjJvLAZL+nFSMe8/e9SAHVR1dGmchoDDpgWcud3YGJweV8gww8CtCt1fO
Hqy/MlHSRdJNRp0/+t7u+8hw8HFI3Uv6Qh8OnQX47WMxekKLaGEZo8s4TZAvIezUvxPGmMGSGgDh
4P7YLtW0rRSzwXws61qMJnIud03ve993zYJDDnREny61peMRCrrlf98RKOELk1+jIjcLQTd/KBOp
Nodp2lKdGfHwD/c94PM9ug6vy9HXpkUueOR0rQOGCDN72p8vqyySQjr8j65n8PeJdBerLNHx8WNE
qP9h0Ioz7G8sYAivdwwQVDBAfJ8JJpT91swdTK1czdooR4E8rolGbDb0i/OB8vWpO3kQdpIZ8buD
stuVPRbT74HVCxaV7yfZfvrhK19c5RPOe12JDAU0p4Rla6tVD5/KA9sJmizWCIsSBjEQ3W44kXGP
+tqwtxnN2kjb8CxX/6i3nEHhRGgypyWMkGuNPVw3i3w0TAXnfpobmxg7KuSQeIpY3bYm+DYOdUw+
qa2H2Sfa6SMmLxXJEjue4O3YHBogNh2rDJu9QcB6N9yqJkqT4o+hiKDFyK8QJVKKC2gSscTy3V4U
X1u8QFe7RltSBLLjTEtVThTv4G5nFuZ95awJf4elgUA6Y0LJ9UnR7cEYqT3+WB1ffwFcq0T5uSV7
1Za74ZOEjBf8oIxQyWEWFhXkby8ZmDhw3AN1VJEM4ko0yBV4RubT4oFd5CQOQ0jdBLdGJuHnaPRf
34OeY022wRYltuTNXfk6KhyYl3dU4Ylc8N46Y2pLDhm63AugB7ISWfEB396qIefUUsQt3ABYcuDD
1FUf9KydWIYCenIBrq/kCTNfZ0aaf6rkUEFrepfQaIEFhZeXFFwoeUck3wl+EgYg3tLQKC28XNmF
Pfr0Aakaz5TYEgCA1jZxVNua0ZgNKGnvCoFdExnOcjgou4/HDFUUCjgDPVMQL8GssP26rQr0hDnT
wUVTHerkLWwL+lQkHWFG75Y2qJbmXeJqoRpOCgDzi95sLBBWDOop8yVXRa782KfgpGiQHidc3fP7
kRZTRAPDtwxigiL0Tw1OrUaQFtKzd5lp6bCu9EyRxdKQTo5T5TnI803cabIrpTRJ8JGOUv3F4xGU
6dYeHjM7xei9fEPGc9TeplAUDeGwECA+v+3vSot1Y9SoyT3wntd+j2DgxiIAYwDiv7PhA9txM0qD
Oto/axM+G4GFT8tHlj782d+pGrKAFh7egYbSzjhdwLiwM003OSePJcZ8ZnWbsTEHfdxG88VPBLuG
XGbMxdlVzHxSjCwtr4uk8iLmXsRAfz83HYndbUprWv5rnnlrYNp5RtR9pgDn2XLWw733mEXXceG9
9Wwnubv7zkQPtwEGNLGoEER601ZBpLK7AqOo8B/O2AKV3IWNOpk2JQkXgR6aR7DzcVzkzfqARF86
andibdN2H2PVTbdoNCqmRVSI4iXSHC9mPRTTEiNcU3vlKd+NjSZrxKrkZKRTodc3pD7TbRJ2HOFc
Y57/I8YHbKlUXcu1+CIze/6FujdMdNY9+bMX49raWVySyiRP66IVEI7Ap+inXjTlYv1vR5AI2scW
jNYgE1nY1Z60a/M6+Tkl/uHe2GWhOUMJX60D/NH2aRBctnmyBcyhGsOP0/NjvcT57gAj/5sCzjo6
ClNWv8wbGkNPa9iHUo9W0EPZQszg8b1Z/mTc+082ko2bnU/k8YrWYzMfLXxzW3wsFLH4nCuXWrRD
t1o8jAiXGcQLf1Wvtwv8MgofTE7cy+GM/DGEcMFcTCY3t2WtT4YfJnaCgAOyNgcsgB99+5FtxscK
ii3fFZVgZltXoHt6D6EMtcYevMEv1Bi/LOgXTqVEahu6s8XZa3C16jL5YwdEmRnI/LUb0/SHdtUB
EV2REidSueg+LcDWq5SN1MwLe6fKYKx/1qfTrbu8dpDJc7v3zPRFRvCE1YB894wezE44GDGAiwMo
Jauymf7RGeOwRl/OmjhEBBMeCpES2OuISQNOYPqZe+5zYqXytS5uvxbCuYgQffMmXxoJ7FpTNwKO
3mM+x9ilRCTnETdSk63wiT3Qx0NLuG+9PqkyJmt01NAtWACigz323LNN1zSGlvxgVE75/pPpzh9R
zamugsLt3PoOmonlNm9+CXCW+SjNS1pl6n9IvHaQ0vwqlGqQr2PfbPT4dKZmt55Ed8ExAkK+E6QF
nVqIeYDoCnRR3+dDR/awGCqYlnBvcW6Puf/K/E5NSGMYxjYLSBrTud6GqzEM3/7KNPFx1xIHvysK
HAmxNYOeO256InlcAaLl9Acpbm6bnmBQBcUMMPnYrKo1WfBhw+5SMBBHw+GpMqjagXZ658UbhB9i
0YL3C0tC2/o+mfnseWAGhjYQHq8Gh5Y986Pm0kcDSJbU1izPpBGtHhgbZqTo7Ik4OG4XElIv2k9o
Cnme+QzMOG9yywlIYk3mk0QV3iH1NNgggjVYBofRL1bFsWhAMYNRjOwEQaXFnn+43aQwvgpfFeNB
laRLm2KUpHSB2hhuK4fBoPvYipfsLHPDV1v159leGgJV7f2dY93DT4lVnk+1OIVjfRXs2bBuA4SJ
WtnNpct0qmu5VMUY6S36FrLwW6xDJmlQsnfD0WDmgT4DoNFhSK3tcdNQ0CAJLNd1CHN7H48WWmBW
56enS+mnP8srdLABT/FEZl46/TicWm1pywGmjp/kq/1lPGke/IFHJa6ImgTViCxK3aR/Io5Vk0xu
0qnM0zPjjVK2dj6xZq3ndI2eEQL4lOKiqZmLxfZsUVXI0HNHWYXVto8N7X7ExYrZipwQ5SmrQJoT
Y2W8p1g3F7HotNo2HCfVcpo4xkP0aDrWSBOOpg+5iGZGUvAjmbK0Ks83/Ytz6Oh27LfokiT29Q5N
2Lb8mdVtPMuIYPK2Lrop/Xi4X4qwvfUvWc/E2yORmSuswM0RvJEupYTU4dT63wu/ZcPg1WDsjvab
z/g/jHS/5xxwU5H9Jsk3vk4qpKqvE/l8+pHqmMEBS2jBaRhR+6N+x07iksEckXNARPB2cNyb41nl
eJ8jwSR4Mn0DqlCIpiQ2I7JoY9bOCq6UCiicsw6oavDtwsmlBD2k0yAOTFG2HTAHgx2IzEwqE/p2
UNZwaRswWUzg4db7CMBC9LgmZfwbBrRHuA6DDy524MGkZM0aYcKoW5rd7mg5UAcv4kHmvFxjaae4
SKiImnttK8Pj8q9ms1BAzEHlHtWJhJgcQEQKMa2haMugVD8zI0nml04PlnMv3+DcSUa5WzpnCCzZ
7WhptpgUeGUr2/PisOtA2wUVoqLOmhka30omAQrH1nq2jsFAMGhT6nRsQfozZvyCik570npGm7fZ
Y18WmZWUtCLpHxSnDf6IT3HJkE+ihyhLWFAfEslluUQMU33pu8CeL1jSJrUShlb+j7EClDEALoA5
sVUHqX47kZ8S64sZreUcCRF5jpcKjuICuu2i+qvDtDH2/fE1ixqaptg3jGrXfG1P3eL8o8FZaFhC
A2HzyU3wB6cVKDpx3CUcCfHSetCvByveo2Crwn7h0S/Nl4NDBOwh+PltwU1H2daXIYsrzruDSNkU
VmYzy9HOtxYm+aiaszoL2n4HObyq+3h/HE8CGxDNxH5YgUI3SdFzwkSYzsgxokfI/Z9j7IDCgUHF
d6YXOuwTgSlz2PEg5DzNlTPWzOeqeB2Sg6JYaIEMaQ2pkThRr0ATp9FcuFrW4ZkcsFtd2RY6OnES
rOvBfG9rVlkvdbugE/r3JV50bsO0eODNJ66FCuBLLbR+ps83YsoG+XsZt+J9Kx3HXLz1DpCnogLk
ZsSP2oQNSMSU0hJkjH8sChvNxbcHbmNT65TAvIoEf4x7gpozycYLuZc+SUTgk2T6D3ZE6vHT1JsP
Ks60cvHAV+yAdpOus25hQunaPHhENo5jQqNvaSQ3efArRxLnMl7Iy5m0fUX/OFEYUJLtrUNGGMSy
mgDrlXX3eUHWyte1pRtYMRFdnV5/nSOvvAB6bHqeu4kd6Wu1hhG8RykHvUbbwHCaaDK13tiMwdD2
L53FHjChndd1ssV0H3hlaCAn6IVcsH+nxCIAzZH9vKJM6fTM5EZYNjcs9uHQkpuGsbf7FC8w3HA3
ZDGhj6W3aOADuBtJ4LSQDfeTFYbP8pbT7/pzScY0vuRwXqc+fd35nGLtd+vPAqHfjneGMpT4hri+
dGBW07tZbl53HjzFzJKnm8OirvE1og74oStWWxwADCEJdTkWEmasnF13fS7owC38acOpb3PaVtAT
xNedXTnI4fCMfzs6WX9kJkmWcAfdRGsBZnjNnOVeExDLM+93DQPtC2RLo227jkuEOoDpltnWCcnq
4BdP2NBW67Vd74M570kA4irMIIrZp7GJg+9BjixZ+jpn8599caMlF32SxvHW6OTBr7JLlIf+xZdK
ApftJvgDCA9O9OWSv8UP8QZyixj216iUfHED6HAvszX6aoMphLD60nFwX/RlcTSbtZ64VZBCV6bx
a9mL04vqEg7FfTPqpkOmi+Oc/j1sVJxau+a1PUZ9DAK9TXbl1MZpM0F8C+TFxJPyIlifykMvKonw
sp06BleBb3vd+tVQxlu6Qbcq2nnmLKf7kFhrx63x0rUXUfMzs2knZJ/7wCVI/QemJJmUgekJmY8Z
RO2HVqVWorOKnSXCIIlgOOQRlqB5nYcaHQdmPjE7j/OxhzKys4VdO9OoZK5KpCVLjPVbuBfkfLIp
pCXDOLui17BoMX2jlgwLS1qN/alg0b+wp7fRKiLqSMM/B7fILprWUASkHhqGeZTjkgveP3o1b4ua
+DVoG2ROb9FmDR/vdWf8QGtJsnVG5mkGEk21EVx3SMpVNHKGtZUY76toyuzMlDAzebcoBLd5TqOt
n+cindyNHZr/DvIN3oTWNfI0ugjn4DsGaicsKyxGfIgGzZmMjEMlEwxMqTwmzRLq6l5wlY7X0pVd
Tr1sEcneC03uTe8AWo70ri1RFmiyWfN/In0xQZTg4PKmvms+ighPqzccDiBm5ms1t3mSZe/kqVkN
/3soAAQj4lqjWoj/JjTYh8ItmHlYIQGTM9fSPuPxDzxfkVIZh5iyZUPggaBQPQD0gnQX1YRsVWb0
PnROAL4rOkoXlg+MF2x8tnwmoOYlEtTUbeU9Yhuo/AaZlokW4z4C8zSl0bQTWukQJgWMqzYtHhfE
CjoV5AMuKQTGSIu3YjVF9HyQb64/X4HdRjKRSXBTu1sMLlR32/5f9U58mJ94QYVuLENOz3MmoWDA
zF2KNlyzrIYtZ4uFnYvUQTNwRjoUvPKnbXfcAgBQBN/ITyCo4bNsHW44G25b63/M8welhrgYUUwA
sy1+kq5pAuLVgPQbUWUREKoc2Gpls53w9J8CRUPfDztFC4gYgATa2NiLgsJa4m6+70QNuraoRF3T
mI4f32A4fp54PKz9O9lg2Nw0UsyPffjer+G47Cj0HEHIm2p3ztohN6wJXTSlnmRhddIROYWasjMb
YJHNP3bVKK/p63MF7Bt29JuBMJL5p9x5HFGTyiXROMyZrveBxedkJj6J/bja16hwzv5K/+0kJYNJ
ir05L+oTs0i4naanwcg633uoCcd2YZLzJv+cW9+2Md7Tj8C+Dzb6Xzq0pUiDTKuFM4heTZTWkFw4
eEQAe8zcP3gYI10m9hdiCTvjnST5xx1XPI7NMOlIyn2fYXWLzrRQ/WCOMtUWF+nngEIyxmCLsdOp
f89Ub1q/vbGXykNdtKAjKBxs3hjVy7gEPVwGFhfn9WZb7Hin0yQuYKbnFfONCDWkBSq+i3jM/NK6
ZpPN8iMRxA21OnahOaObzaERUXttoBylcLmdV/eIgco2eC2oz7tWK3jAUddQRCqwl5j+EJd+zEgf
fHC8XxjzyrFLNSyltz4d20qRTdcbVULYQ4nHg/Y85Oc10suZmjAcSgtLeg7tqJDO+6hdC/wvn294
L1w1WUom8IDYPMlEB4/Ns/fsOw2TMNQkhpzZj3KZp1MqvkQu8PgVrB7v+fe/a/BstNFn7nLQlPqe
Oqg2yHN6sQS8snkijm+0HZhsnjSrrR3IlNfw4fwuH1nJ2Z2gno52JL1lUJ7gLfUkdAFK7WkNvezx
Pqqqg+ix4v7Cc1osAcCiQcUjfMWzdQw7781wjnWiR3EXahvEe7LgX0mfpQ4q+QDXRtczJvVOSzN6
GhhwGdyF+rSjiNCwrkRtkalQ9XscrM9WP74dYuHKk60UtduPqQQY0Ye7bXA0hvRnqKrxNG1fFZ7t
zvlJG6kVccvSUGvW9xCvQ99tH8ZMm+Bas6dPQFncMQdbX/uerKuvNf3aoU8Zi//7qghptzLOnFVQ
0PKbaQyF3ew0k6NRkdnEge/XXwTGU1L+S3pKexPPGnjhgokCt+GMvbOQ4z8OSAXyo5qRlN5GcL8f
JHAh8FMpXPULGCHejQVIIDYOcovwjkkUjXJIKqyt7tOG9rYnrpogkHXV0q4rwZ6cYw+dbsrbVwrc
gKnyYcw1VLNaASCXO05XmB/xU5nQbb84rIi//LwVVCXOGxUhkH4ydjR7t9BjxyPfVcsGZsOfXqxL
umFP4EYybSQfx4MCVbe/o1f5qA3a58AREGvkCGjdktEijTjhgv3jk96s7z9lZBEderSyxZ+NJriz
xJ5l3UXoe9/gVbT+T90d74cZ3Gf4HWcctoRqhgvBw9bBs0oIWVm1llwh4rn/gf9WtPplOguFX8PJ
dFWEq4hOkxrXoLIzMjUPaiIivKyFcbmVB8W6oW3fPDl/itQOIiaOcz4CnYK/Mef9OVXgcCvaURyG
w7zzeVvWNYL54GwviR4IKEwunCiJorhYbl9uw1AwxhUI4uNqHmbeMR/CZoJ1rpiO+5Gm3N92ZAGg
QNVZNlluZ1q3i3nNoNqbqnWi7Q5/hXVRYeivW9HFcUU54BaG0U6d5OPISDqxR5XOhDj5CnV1PXB6
SRRUKqYqe1Cx58GFAfT6nZB7BGn3lNxm0XHoLvLxPM6KcSUDZwO70l359+lo2e5uDHmo79YNN5mo
2zabGJ5YHVq6Jo2syxvBlmI6mOBmjHW5/zYBJ3weHKFbcyyUDhT7Q9AGgB8LlDfxjF7CpHnX+wM+
70J8pbWHGHfNufPEOR9xkEL4KWvlkOjqWYxdDc8UWlhVLcofQDRrqDUnmkpx+L5UU6jTLayZRcTc
M2YLuTjrl94u+EA2fJvt/G9wD8r2zksGTpOkm0X8PRdU8Ere4HFagcxezZHfcriaTwfKh/MryPyg
Gfse1Q6JZqsPyYfDUh3h8qOk3Mx3bQKFxbQ8EMkxAj/UjQM8TkjnV/lTb83Q8XtxxwKUHVMiiMqD
HzTRZr5O6rPlO46wUzPeiVMoZfG4ze7O2or0TsNCMo5zTTKmXrUtrCgURzy4CHTpI0QYP25uuPcC
Jo7U+Te9o8Wlp73KG1YasWc9VxnJR1DsTh0i5dHBF2dER1YEbDL0gz7O6Ted2F6pCjuKRnbotler
x3Vg1v9HzaJkDL01vgyK82zneH490hwHSky+Av8qrm8lu/Vf8NrrwA73cCIIbMKBVI2ON53s3/r6
U4zvb9RWrx8jRnE2N10tCtXYbq8FO0aKxYjLkxxJY+wTQSx0cSvWo56A/PLH1zoASfRUhp/K+la7
ZX3+POEdLtesjOg0txWZxuWFZYPJIcqQcfrQ8yKJSmY+jk6PpmAvjbJ6hlQec3YrWfHVgQMHkbWt
T6EmSlu9cwDsJxm74XDLAsnhANowo4S/9pVjzmsBuoRR38SE+BF6xjTtPcQphiO2tyzLPV+p+Syv
w928S/YoSvXxaWOBAwg4l4bv/nY3zjHHYcPmogg7yPC0GSm3hcUGKN+VHCA5z0ga5KH0tUqTHF8q
ZMKlvaqpdKypzejtF6W96+4S8oqOYkuhEsU8lGCNyRuQg0xihQok1AfTCEuLeD1AXhx/qmtjgUne
y1wOAYJIKKXKtzA2eKz6s9A9DSPSKV87HOGif8ddCfM6+N2i4dQA1Pu6UpZDsuVPBjGlRrTOoeJm
p3kZHrkSWis1oRYP9l1htHfP37cQBWoVviXGLav51PvIge3ZpAIIeofWWUCL1vlLRue3MxdOgkIO
3dnZOdwJ3oMZVqTFSl2L7A+VTb4uhSlFUViV05MJEaMUlVTJJoHuheVOs7VHaQFuoLrKEJZSW/Sq
ClNWB8GcVdQDnsCXk2IaXmtcbex13WImsEhkHfLmej7LLcjWNGjQP9Jp34dyM5t22PHdJX3xXHlC
fvpTCbpJMQewjYtF8uGzPJg5pJ+80THpzzpCPTCF8rCHcwuzp+pb/LCcajCKHb83TSjuBYAd6iGD
46VDgHlCAK+icanw6/jr7Qg97nt1TXnk2pVUTCAPVqYvJB7JiEz/yTPC/xrd0PYQsWFlh1tQ9Gq5
cz5+qSWtyjm/7niho+/pENpSqVMkAg1mI6UMdr6rwgVYlC4Bm0Y9tkuwCCx+M4qjhsbE0tH09FVm
hafF0taHOCE4K2yjbTOTErl6MKovnvjNkGbWBnxlLrdOGT6TapzwUJ0HiqOYiSOhGqFWkmOl2VZO
8Ga5yM+AXE2gJ4wnB3CmwV/xqBKk8jr5h7BffMGaA0bxihhJ1TdW6ppw8BpuiBuZea4rpf3HrBWf
FXUPLnXi0JAG6jbK+p/JFwhj6jpF2cnU3GzCpOb1qjDVEtT42VEnkbe9OV19LB30voeAyyk6DKbt
2dml+7u+hkoQNon2o2SIJFqYVi9+c6mau1uTHfKDnvQ6Wc+LkXbiE7mgpEsfz1vuC6hNcztzLfb6
slqNfoUmxium2CDABt77Qk71aoDGLigGcvEE+yGqLGVciX58EApUdCKVvXUg7Fn5YtKyWKW/kadF
oWy1QlO4mk/lv+1o5jEqC9xldeeHSebzR8z6jeQZVisp4Tj1cJOscNgOunZbO/bpCteAacsuLig8
M5/11bWCsHNt+U9mrT/I8KzvvlSIDYoXq8Zx11fXhDTRz3iWH9o9E2SZYi73KKA8qRD3Umr7eI/1
eGL5w4OGDoZhuBZrxgZe9Wf12EzTFyR1CJjW+GmHVrQ4A6UCdgmfybTg0UnfMbd7AySlN4jr8gFX
Rf3tFWN/Mxeya87CWR8JNclYrfbXDAi/RigyYyXFMZ673LCmWpeofkiflW6ob/unXlnTRVLjlMVK
R9mx8yHMYna4C4NYYas8v2LbXJOQY9NqeTvqsuHCF6XTwbB6qUMIKjEzOY7ueKO5dHyCIwC4HXiD
M9GF/8GGUwzbB/P3b/ZLRzTpbXpbEbmaxLdLNvTUHu02ml64c0ifnvYXLTqR63S/7Bo7ODQAgQvj
yb/05E+HnY1UiX+oMyAc1ccri9p+AVUXiAe0+L8mggrRfDP3RmQ/lJW4Yp+O6Pvz3ladqzEvlRnz
TxRiadQC3yfJ9c+cZHi/Wm2Vy3NwW9lbuGR7/DKpuEFV3kCTs9fMxGjJaJTn1KVcbhKVZhbOv67Q
Xb6op/toZEwICCVbCQyn4gtas7SEq+uICky/tbVWNa3BrG67n3At4gja09SdKQjEcOnblBjk7oe2
l7OlvlOs35j6IySxJwUN+tGk4e/wwKmt7EjQwdA+3SqNIYdAD+rklzX+vr7gMSU9SgMZMqTFQRhY
LgPp1P/Bvz9tp+AWb4mTmhdD5LqyAGx7s9cTP+mScZUZSXAaHhGWfhgh7Ye8FJ+NU77r17vywOMA
xQWcTmD/F/23zuAJ896qBEWCCM6hAq0uNzTQ3zsuSLTtY7v8mQs1Bzs8gkQQhq/3ijTqSzrho3XU
XQVbTwwsqZ6ZTAsZI6MwcjA/QIe8C1xBJP1SvRZmNAtsAaTnCPYqIfICzBJxLWgRFidE1Mthngso
qMNN0qY8vurPf4McrJPACiMJKqh1C9UZjLWzNOuyrlOKPC1v0ITK4PpPRTgx8UJ2aHRHFn7+mN+A
3rvJzDa5pHW3TMYW2t6j4JMAKkRnKb1WFr4/zftS8yh9Lz5AEzn9AvZN3w0BV1bfudvV2XZTXYlG
EVoFHzQW7M46HYEBZ0w2R0PAqD9XSEsWd7cJv8vRzq1XW+SBpKW5XUyfzG4dGK7gkNwNDN7rkRzX
W+srtkI6x9DYEYDLjMu9xZRc8tGNB3Uw/lWdsLFtZp1XUCoCSi2HzQn3X/tIls/6JFgBmQ4nhOAt
HQ1/aivXhDJvbD5OoU+lIIHD9de3HXFs69eEdYSbfs9vtiP9tpKRMd73XgoCx9mm1zjR+uVQzRvI
js5nkJxbZ78N1Cc6eEGZ9T9LqHS5UMTSUbUPaf0C3av7Rupd8pUr9wa6e2xRLUwna/Cp5wU36B49
5dAecj93EQ8nz48I/SkQg26v+1BFhw+e+qxALMHi9uXdCHEfWcCJjun7SWTIXIGWMEi0/sofTvjJ
9fR7dwG+a7WFEIsc6xxJH8H2ZrkOPndHnkxaIkqN06mR8tkjGJCFSjaYii5HnTRQ51ZCzt1senMJ
SGySvSizT7rxcYiKk+6kWxW8yj7rE5Rjp5uRalFTPSGvLbudA6YoyA6i3ou93cv4ZF1POI58BcoO
ztbJgmRL5IXX3NwdXAqLEBK4xOZUnf4cKOGyAt9tM9uhS5hHkuzOGOLuxl1Yyp3uU/SDFbT3Bd8t
Wpy1N+Ro06qFVykm5y9Lo0H0Uk4akTaEW+3q6qhhU/Bq11v0UjiebEQMl4/GJE1f1zLygSVuzYhm
mMuFon1bIvR0mxDPT80lBcNKE6hpqY/I0SybwaVFvHA2KtwInj0cwSS7LFIDXkea9tVXX3tM1cAS
TKFa6V7+pfknb+OGkSfB0Zucz32fLMDzSbbF6FiXkrc0u0QWn4Rpz5/KbCeAMvSpVYKebIkd8+xK
LKOQdx2flRbIipk+PfE2hcdDr2vNhZ0a1eMPat7e15iSXttxFzsO+BEGJyMf7ek8KLrtdch8r6Q1
ZqW3WeMnH2ZmTL51WvlwOhtCmVBQm/fPk9ZaDrVcQcruDUuojz76TsrlMfhgjc7zIkzoxUO+OdND
v3XL1Yt5Tex4nzVxugCsUQfO6uJ5Lcyc6zu6OR9CetrBFerlzLkhfrYbYWfubXRHI5I4OMG/WYDY
qBpbd1mZVGuyc1xJ3VzSbU92gfddzWxyJrGg2dR4Ttwb3TwGfuiLx7yxGwBPB9gkaJK7j0uk5w3f
sST0dDSbv3rxp1AbS2/WFatdbPhvIExkIQZh4tzQ7seiHSCGuOcVKHECUmDNKQRr2tPHs1XOVFdk
3YRVgwg8I42Azd4yiExIiMHFOR2tgHYxMHskvBzSfXW+j961fe6ViTcEsBqcTp8SWBkZSfSFIZJ7
Zt+74YM8PU61ACdZhFGcBtROCQGJoSdLHC7jg6cz83Kni9tuTfnkvqY5RxSEJp+kFR18cK4L32VK
ywWKeI4C8ksZSFKgPIQHUvkqXVNQWLd+KxOs+mZCpQzvK0qMlSHOnBMJDNOvka2FcAKgtnF9kFTb
73to7aJaVd/KW99gQydCUvtppPbG0odE6SkItSJcmqEXffMREuAqlX1BEe6cXqmaG+37iK6ImQCq
JPT/Xfv0bsbgmD3ZrxbVNFLe9UoaIpQfrEe41Sm0nALK+rQwA20+3rs6RyDdbBww0WlhN/qcr9Si
hWoYN7LvNAv7sBPubH41uRBkLCCFqZLCpyryYcnXSbeacil0rrt0N3HblqbV8yUDmzZ6jCUtu70G
QLuXObSM7lWAF3s8Fn89hyHPsW1066zUL0qVKgbFXRUMSarUy5xzTTcGmon+WTTRo0xA2XSgsDAK
FLe6vOyVX2jjJ5XbJkwsCF+klyXA8TB1LIQRUTiSoowTvirsobfVxvRGrr2vJhMgCKtPqSSlhiWM
TW+UU86Lt86ednWI6YPNpPw7QhUvjHeT7m6Y6ITEORsQvZWgmbuGySeAdcZ2gXUsUz9ZuDU5f2ox
qktOXCt1YF3ODh+JE7NfLn1WhlcaGNtkpXCWfSDIPNiOBmPKaCfprulXXrYQ6Tk32GSI/5ZsXTy3
N3b+ZgiphEkJaoA1AIycjRVQI2fOT/NarsiaYnGGBoZvy8FxlOB/DGdqvIpISLBNoWr4+KFs5OKw
TDRxV4FRxrEkSxYwXPyhaEa9drBtiXbgjY+k2ckaF50TiLIBAcmtN90azQYP2cDDEYnzDythiXil
14s/xLjQyWAWkd3QyIfOYqJ/zusofiFLB3WRiapowC0/oRufMp6NbIKX2Y8yW75/rWXOB+0XUDAg
Au0VQOKkUfj627Mb6W8D5NuAh2bHrMhc0YY/V1V3G2T+0+JugYvFppa8vsW8ufTm2aDC1kd1ZIw9
j7w37nWRkH6DL8+IDVR1sI2qgpBg7a+U3beHcFdL3csA3VuOY6Oh778oimJB1u289uITBM6rsTzr
SfVPeUnZRw9sa6HViXN7r90Di6ew7NoKrax/M7OLNb4hz3wluhl9Z6gXZbQR/UuwrLu16QIzHFVD
PcPqWsFp/2Qj3BFIxhK/NLOfongVKjkaatjTdI/cNBwjuWmSyWx5LsAhctUTqhnC1/T++3AsyBNl
1+QUphg23il9pZhPlspw+qFaIG7eI0RwT7lobMuaPASDAtdKPmPFYqotk6vhgoIZayloZbHK1BeO
2BXi+I6KXcL+Q6duLn6Px/7Pm9vaaa/dXFhp+ao4XKyGyfuDYROJM56mbpVB6997lze+K8KKfJ1Q
rlGYLAugXeT+KNLg3xGHklXZfJdP02sqQOSeBznTbkQzxkVtpqOfsNcgM8sIXiyTeMuXjE4CL7fl
RsQHVOhQFZe+AZYZqVZEKqn2IpXDZ9Pf2rFi1D5inLN6G880tG6UYlloC1pIdpF4CujOkWVkrAr9
ScmH9I/9O1WKzrEpqUJ7EkU6YWIOaQ7x9aYj7mKNO0Lq936LqzBMaAnjABWJwqutH+pBeFn+zAR7
NtjZDAn2uka8dSEOxkdENq85cnqrl2JDZAzWPYr+veCjCwGMjXRPbgcgaldLbo5Xc6TOq0H9pHhZ
wRJi+Gshf8jHNkkIofbclp0hi36uXEmXbnVeMbmfKhvCaKiVKHYIoCIyeNFwkUHOxh4nrUpUvSGv
oG+F6ITDNk1aax9SBxb2eZyFovYlE2Pij6vZwLyBeO80egi+yLiBSMJz74PeBp6clvuCqpLlvAD/
CCWx40YGZr/zlW6ze9UQDCsPHlYFS96MKqJnlQR2ECrCIryKVwD6GxkA7xF8BmuzgGkWiMWduZ3S
OKFAjkXQPzkpSwbNRbvTKSFEHxJbVUk0hGI5EPFZEDG6aVwwQ7A+Sd+bTsaRcdUlodW828T2356D
9TAx4OA5gEL+KHF9/Mm+fU1KFRzM+uzFM9EcP2T7qHz/Tg1+Fq8cpRNwtudB6geP7CPWs5QInAE8
cbGMTZop+6WSQVqhAlk4eju6X5+ojdth8nUIvxr24+rMIhQLXvY5DEWQaYCtRITTkgRMazGqgn+H
n+xKzDl1sL6iNZ+Tgr9M9XcGlTx4Wdb7AnQunxKqlAddJGHwLXe93HTr9TLv+3ThMH5y1oh+EYT1
av2BLb01a6yrW2ZChKII8zZ4bFFLIezSdjeq781wsTp1HMo8CP+Cui7w6+zsQrOuMwz1uUhtMWJ8
VKtxwRG2Vxo6KDOJjOKLfYF2WEgzo74c672TyiaqBOJb8kl4Z4wJKSiA1xuGknsPnT4gbddf+gSR
wchaHRW5m0AOskSF6Isy9zFhHBUYBpobM3Sqx11HND2iZ0CJ57vmrlVhe/Eildujvel7eyGZAQIv
LVaijxtt1pSpDcHscfHDNnNetBSQzZEG5KLCwokjCmEx9V0WIHaDbNaVWOUUsVgJ7suRKT+B58rp
K44gCHChoTTs7dC6QZsxpcCSj2hH2JDgF0Wl4KUQC9coJRzY27VsTy6HLr7bSZE9xqfNShMBrofb
WzbezBIs4gRnT/e+wko9T4lNeYMHLWS4gDJnFEq7d0qetsghD4NQ6CFa+Zj3aLP0Gm7bNLry8bm4
1+lj4DZDJ/Woqw7kdPZDy4IM0GKCuNs/6rGvu+KtTEnbO0KJ9CNf62DBDhql83o6gM7zAbUHQWsk
n5WG1CMel3bQ/GIszaQjx1urrH7KFGqXExVjm5oGpssR9IhTYrse3ipoKYWKlu38/iGVIF080Fpd
naxpXtI+jkBM9zZn7f3Ha7TD4N+9E7Ie3VfO6YwGLpHfLKV1/Rn9XNa9uCv7Pq8FeUVQqQfnFEf2
30TXa87sY63CmwtLGVmv3ZAdl98IJx8YOJWAVXpa2yQ1YWxyzPGrU2ChLyTbveVFl1jLJwAavyqK
s3ID9Am7MMlTGWqfgvRcGK89nZJpYIiIt9LBWZ1wSy22HlfXLRW0w3IkLgusijKx4NdxLgkLJBd7
63ICTLEA7BvPrBmi6MDohBvt3iKKWCWXNtWFWZSn/Cu/zia907aiTq0uMGZIvvTEm2sBRsLirbhP
8vCTrSvfT8ErI4SEHHuMDKOUXFKEj6sr6ETz/BesIvDd7io/9ODIgggXYmliaczXXgMi8QPD3/kj
GlPnyN3849NRvQNmPX66mvIAYb4UfN5Do7bfynq23weYQ+7QUZ3+cfwE2UdwkRhKMNpXH8L5nJd5
+A2C07YwGMQzWD2H31nfRFR5wVzhju6GKW03cTUBvtU264ObgeDsKJsEBNIwG9HmteNVPf+atZe4
c9tVCp3aJYUmaunLH4SniBf7bDmasqT6HtwwHsC/O9LHDRPEeFlJvp912FT1NNUn0sZtdmcGD3sn
tMuUOH8qQsF5tZEtUvN5X84Xr4x91N0cPjcQ23+r0SWbQvWdkL75km1TNv5E9er4oTF7wZMuQaHE
rpy2tSUcM7WkoJFBwv4hNH8/NJqcwlj2fxBv+BEaPzDY1A04scIIEnYPGSn2qeDeIQKjD+bAhHbb
5v2ncX4NlSniRq6SCClDVAWNLl9u6TAaz8Gblx3Ri6bFVB0LFv3+wy4KcZ7Le2NWr2Jq+wPYnjxH
TmnQFJta5Qe/Cqq5cnJMe7sc79dfm+tDeM3bioyuXrHf3bPKHfpn7Q2UmUNPhaovHFZH5lSvbPWb
y6qehwDNIdfLQ2jhY7yDX9loaqwhVJEt45GA9XyEQxQqHlKnMPs2JQ9Y3PsJOcvIv1W2c4ai+PR5
z8CCzCTE9GOR+pAYuYd49JF1t50jNgYpLoKtVtl1tS8PFbhBBVPwUWH7AIWiwhMfmNJBssVr2p8f
9YHDREn4bCtmxQPoMKvRwf4LPbhUeeEspRzNNpwCBU5noabixi69APUMlRiHq7yN270HdX6Stpa9
wKlTdwQBtEdb2P9hqTzLTXFTgnv7e1a3bx1jAcnr+NM1EOjApe7CffZtmURrPRHO13c+QVdIVxpE
ipIpY1HVlV9Lv0/kq0DHI7L3Pg7YwCgV6PaWnah5B/PlSwdvKxKsESJDo/D5qOA98DdyBF/TBdZ0
Jhah3SkaoyJjm5C2p+v2cyEuKm8PA0KLKWXCNTyz2mqBvv4kAMqk4enJzf8++Cvl+clyGzSnG9X9
9RgEziou1FO4Dtz8JvMfqOsrSaLQc0VdWHLLFRCnG3C/8ayCwsisoHpXLRR6lJbcIY+ZzJtTzNbB
9klphsNJPwoHsPRY20+S5fLyM/QJEr80PGV0A50FWEMUJcO7rzO1ctyEr6nOUhGYDQtA8XgSvmsT
90K/zD29jUormOnSmuWy2ydNlaJ1YUgHqsK1+t3VxDvBFtbGzNacSjTkvlFwyBBn0y3xYAwqgN0C
JY3i1Uj6O62mInor86xarXfguQPBcm2l/5jClgLoGgOLmTdOIwHmuqfDQz4QcWUmHW+Ab+VgkKLm
Hryb3/03JgYHFycSAbM/dWb27DN3RAhdhsWmcltMi+NqkI2ufvNLckenfAq7/a6St7Z1hrxwGWGl
92V3nQK/TvbkwcXqkkQJmn4j6VMXuTSsgmAHQbtuqIgGT/IQS8KL4WMY7Ci0oOFTpAZTh48z/H1Y
Ggc3p+caLBdqNYlllafQoQnj4PIXnyGLgBz9hr0sEO+zKQDheF6GxB9vsLL1mA2PhUH/Tp9sIsyi
lHMQXlKUMW4YXvCVSci+6z4CCY6O0Milg3SQlq+yHH4lPRvXyFI0VB4N/0axXf8/4qZAQHc18N4x
28SWAOh/sXI5do8pn83G55cUA+WKtdNkHL4gOEaU0yAc+koLfaJCUwZRG6zmkmInA4mKu1spZFra
qroPWOQ9PaDbUMNvKbfPCznLDb9sjK3UkVjHPw+556sjs8dQRnBapMVW6x3bM9M2wIN/c4CiVWqo
MAbAFnvYcOd5alXvwsPscTRMwAlVJXaMqsULTqraQrZd5dEEHyeVxHby2fbU/gT4FwC9QaQa8wh9
21aho8EMMMkYqi0pL01e+qDRpBGp29sF4b9PceUGxIL1nY893tqQufZPfL08ChAhw9byKFC8CAO6
OPZXxR5bv9VHBK3Z/s3fDpcKb5kzMexd+P3IvCMen1UVb+9D18OPRWPbizvjjLc7kmpNX+btcvwc
w55V6w4GqYXPtV63elMmaO/nIF3J4rrHJ98+2Hh1n5Tg5g/A6NLKG7p4sktpOiEkLjB+Cap1UFK0
cDxyw+fnO2D6mvMiPtRvsDWzsB2nvLjJuPWV1VMaVvCCTJ1SjE/Cf9kR7XxVFa7QZt5jX7jpY/Wo
lk1xGZDwJoJC8iczCKST6dQsMp+SRpNujNclEWywZmeDYyVbb+949tG2IOjulloa4XCD/9zC97bH
TAtgJDNzZ9EpCfDkRb/jSuyiqwdcFxbsYzw6r+azGHydxIDnMitkz6JbdZ2VsICEHwY3q/gM9nsF
qOseEUGL2reZWJBGY8a8BR4mPgM55eIKpKNBFxo7+B4F0xnOW2pdHlIkdgira8vi5QGLam/DPMsw
OvXdKfRM9QTsKgR4uefU2eUkAO8BBxIkBW5SKBXU8/VftKk6YF/89BXJt/Rukd0ngC4WYGm8JKXP
iINJMzM1Wqn3ENMb8wqN3Wnxor/SE+ai28ObnVIl3e5l5raHsMiD2qKc9e6tCttdIvSxpxGf5C+U
rsecQ2k19McszuetyojoQYEjWL5mhLEBmSpceJJmTqGBf6tDLRUTmfOaRCWc41u2/KaunYed9iPN
/W9V24+6CXbjo96EgZzbu0PDGxxuWHSjVCqkudAApiaXuiNBiZ6OOHHG0FnVJXzMGfd3aw+03iA3
s6aHC5kHrcQwYDSTjG4DblJjwgyCgNq7s0SDvQryn2ehu5/CFoBLUbLJp61rVSwpzjGR5In11rJG
fxnldQfEOI1yI/J3ebJJaZTCU+avmPmXCkZ9gTB5q0J7nGDkFF5Ph9ITq+dzeLfQZGFpc8ifW/t7
9EiNn0yewnZSsCjgV6/Gc9uhmIn4Jj3L1NBerZJH3sEpXoC+yALR8iURGt1CjXRBkSFxrvL/w7pH
gxQKvPML1Vhy8bT5f5mIE7fOewM9k+H34FD67xvMipEY8rhj3rSyi4cDakfVEBHWLJtaJrrtO0k5
3yfjhY7GjGEW13d/v1ZTPtrXvvBYNzQmRojRc2AkPK5x6WXlXlV5LgiQV2MXFO88jrrJ+l2eeB3q
rRGLRUDu3jrmQAj4lB5xRllx53QmwrSVMu0v5ikw1HYjhobwv4iu421Oc9vgTwGD0OT/k7lp15zx
0mz+mtrwRNMmnWfoSQRo447PB4CBWSn8TgrXH3aCcAEAlh/hYBGIxsY6EcjS2z4htzzgnSWhtajE
yjO9JP7T/tc0aawGMuGF8dWbaq/hjmreZm01duwLXoK2Em6304gdh7P/yonEfcNCoOjcXMu3dQek
kddSCLTbMPiCUxWkTtXQ5wviTeNR4TYzoEIluDETjzZadxb1V94qibDVzreU6IeJLAoxB1Fx63AU
i/ZoE94FSxNqkewxp178WrgacAUJww58qNmivLV11HjY7OG3q7w4xXq5tFJPf7HbVkkPBRwU+O4B
D8pgxVgK9uRHAlT6Y5gY8AXzJOY18SIjlqlFgl+0iIP2TbYvo9KqM0aulwcGzdw/r7Qi++HsJHHQ
BPgm7Ag3KVZ9dFByRgyoZfTxZffX0x+NwTksJnnf7DY+myx0tK3eRCFz/DpsYF4Z+ZnaZdn7bWMU
SMDSi8YvYKZiX0tRAbid9EokZCMo/MLE8dfG7odKkhKiZfajXxheu5WGgfOsO3dvV3BltmtXpur0
lToRGo4cquNvIYmIX9zUFAS0TbJ0B7joF4oPUwd6mVqLLZj31AN2fElGgmoa76W0djcixDHIbK4+
NINjP69gglyVxUVWSEBe3QxRiCquvKC+uPghbIOXmHksDjS+6eoUnwioVuS4AucxBaEPnE+tsJpg
oAVwDfi/uk8B8+URKZU0bwP7Xn4yhWVL2sJKTKPNAJpf9VopJrA9t0TOXsP88dLRKoECoRAVX4nR
XGb3b8h7ONMS4t+WiRpVgY+lwiysoBuQz8FhynoaxUDfT3nm626f6Uxp0/EvU4lJlxPRtwpyH4v8
krg4zB1oERUDgI0OCy3FGF/j7uRIvGYgmZGGsJ/HrgaFh2iqivt7DVRcOaUbuDTzVooic1INbw3S
4BFQ+9nMWcc/s2Ngo4tUHAbGkDXTX5Tb2ibS82Bd9h2QZBU6GJgkAlngl2C3+FBHo61vMZZZYINC
SxZDPjYzeR3ApSznLVyvggfhIWp+Z5JwavLLXGB82rsoXdh1P8oTugj/JS3j31vggPDpS/KzZVo0
uAvRrsNkuuvRphgR27oM73WC3LV9e9By5XazMX0FOTgtkPXXtzIpZISujb1WrL0n+G4dK64VoBPf
OtHgNgrfTJlJIs0/9XNkQIVIXtTZ0bKHT6XW2nLWOqks7NKEechSRshz81FmUt2zl4eVetMTjD9S
Q6CTm7CCgEBN9HxGfh0jbOeL0Bxf6N0Y9CKMmGYLjC6jhbQW2jiv0JvsKF2Drd9YBjT/dLTuGIFf
369eEc3isAb/qPDgnpb3gg20x+HrdZvmsu01Wx7paFLSPtj9bbd09sFBuxxNO17fvnX2nV35sag2
M6dfkI/L48oqjb31cYxTIpc4J27UavO/j0++k81VqPBHpjIe57iKQo4rp5SbD1A9ohnqXgfk4+wk
8twqv4tMAehjRgoKaNqTUJPptwbTfkUvwRIZMOaJ1UiiY/6HuCY+h+hYGVFdbHn3Jk8XI77eMnsa
M+7LBgZePNWND20C4B6bJyK1v/kN6dIItt9+4EjOZr0I4tRSbU53i9MX6v2hDrDeOy4o4iWszUOp
DkyYV5zkGXWRbeBxtYsWia+/RS8iNqXnRjznCxvEU1tsomtjQDlPYaIg1TOvIzhZRN6eZbNgNpp5
7YEP9ai8nktgoeynmCZ+nVmD/xx0saEn7q6r8T7YyWUm2sR1Lz7HdrfsOgpsBo8WxyEt2c9Do+GH
XWTEffhLjO0IYtmHb/gXz/QYwxggpuiT7+iur1/4sSu9m+d1NOIX+wXAfNEblJhEOKgtqCSQSNlw
+HWphpv2Xexah+7cCEN8jmoXaXmA35+t9gBYMYtyTBG0UtrCrJhhUN5eYTgi5q8XFDURJjQBIDnr
x3bh5IsHt5j8drUl3riSNno4Kl7HxtaCwjmv5AUHRcsnmMRS+E/P//9Ux1fv8kz21Rs2n9JaKrHa
Iw+esB1WlNCdj9EWqdZk0cBNO58hLoTbA7RAPNoCPgq2vt2nb2ZujJ8ZzulcxWaVf0r539UwkHwg
+quIWh3yLzATF97Wrfjuk+GShm8AWqLeqL6jo2dAX9sHnazawzTr0M5ESo7QK/2AD4YHAVhUPBGM
qBs1lRrhxmzDenuQLzrmT+kZLoQCTQYNuW/UmeM1MWV3qe+8TNcT75n9pwfEvsniZovXNJnRaJBY
wpMRSLBsTKZ0/HsVevUFvDiF0BdRM//kFqV6xDSfv+mtubLslS7R6N5IZv8Uf+5xPXxj8refCWR7
wNFOPjbaKeUbrUaISNuLSu4im97taQQrotnHE7Eg57/Fn+iD8nLBTp7DDUNCIghjg3oopaUvJc3l
bnl/eyDu3WQzSr9xWnOxT156ODbWPTmHPkCJuEDudBPUB7HSQKPSShauwMBhnfvOTtnU0HCIRqqh
Sh8nd82ZL37ENy9en1ynmFSHAHBPr1Ojw1h0tyCkEuT9NmZV4Xqz3CXgvDKjr4csozHERkhT86pl
opVJhoBfxyIFsXXgWxg90lGpra+xsnhiPvYpS86KBXmCZseMSs4x5pyV5m4glEyrczMDEleT3LH8
RYjnVFrrYh6gbjuJaUqZpm1HJDSInsqwHHo9pEYnqrjWjCjW1BZVtoa/RlRUUi88w08g9y3HkXmR
/QAEHCK8GWpwLLTAnji42iFVVZo+ogkCV3zGe20oFHrEKIzPoeORPfZwOF3KqyqIh+zxhc3YCVHx
Px8cPxak1ezqEJEl1j2EM3ndtoXqdAkBgTlr5XnwmRDgOwS7ANlmMqFlV2ON4rRRctVtAKeFsKYo
0AK0ZA1+irjlKOhFKAlhwWl06k+kJ4ydByZF4CjcLJTFWykRy3oXuYs9WBToTptGLNIQCygW0MP3
/SQRL6a7IGHBSWSZMOpnknbmiwTk62HQUlKWGsMtEit+J3TfYmeawBRMv22lsWCZA+RMJVeWQLWB
WJmfH/oPbS2XeEl/g7tt/8Ontl3+VQbs2+pODmwruK+rEXAzWq4dGByiGyj9/+EMNPJ75MGyu0p8
AydUd3FfqZ7XPk5C2tkdItkA8/13ikqSZpnecfZESU64gt746GJbn++KyHVl8LIRV/EDz4UeSjds
rnIgI+c9E9DlfZD1EGqZI46Yhe/ts6a+EdN1fnZHcAu1sleNlFy1/fNPBtJctQY2XOuXF3eNEEVM
2D0/mrkAaH8sj3UDHGjvXETmfkV8Cyk1jG/TIiutF53Ia2jp4RLddmvJBNv81EhjUTMOuj9Vl/cK
N7BoPTlMvhZnqnzkIOlSEBMfkRhi0Aoj5u2yXh8yd8uMJiHwyKw/ElVc08zWfQpzzas+c47ULWLI
+5itUV2WvonCwyjSBRe0mlImL5WpfooQctPeg3Uwb4roegol7vFfiy/EJDTjdXH11ghPJM/rE7lQ
YkGLBaE6rTASWSo2Dq5rWsBa/BWHDfK8c5+PGLKRiILDitrpBi+/jLpTAoEBynUAumIB0AAxtFqk
ztA9njRxIfKKYRdS/AY432GQ8zrQcrUzd3x09E/BcMOxA5JdMUgJ3yqkD65HrGDuoV3i5n1d4wGn
6cjm+9MMO09B13yrB4aGTRQWe70KMRgdAhw+QzGnlzjyIHAwfhk1TF/ggenvwV0/kEbVT99ojnEE
aI8Ds+dRqIxkqh3dqMfeXs6chZN0ZsOIjMzlLkn8xtAbI46wjv+lV0xK7erxKKQYE4Com8quCxZ3
LK/CzmfS/O8rSq9H9Q+rJcjO0Z0tpDmTj+GJ1cInyoFCGZ/Rf4eO6dmf7VbCzr5xJCWnnpFxz3CB
MnAGRelsvabgU2G5SqD75NsLdFYvQDUtmzlv3Wdzr+6KmYUS1euBgvV+G0zcdI5+LQl1bZ/QP4MC
F9spaH/xclPmQZi4qgJnA4MpOcZbWY4QUAMbFOiPQOdZz6FlLOAyBUob/rTrClqp52PulkrHwDme
lCWywpP/VegSSbyn3gmVSPdmxZPPYtt9r7Rtt5fyqiNzrZDlEwas06hOZYM2VeleWNRe2Xq1Mn+C
ije7V5OHsuYfNY+egTYBDG78eNLWwDMrqGEkDSZ+kECoqcDpxhWpy8AxL7Wwprdjqwe8pxh/C2Ex
i1Le6qVmiGsIBrnew7rITAXMrT9qLe2xvTkZ3a3cb9ZDbwxIeELynbBSywmWUy/bstELM4uirK3o
VB32bXGQF/4Zk04E26ou+ZEcGi2H/VtpmN1Bvi77h6ZtOB2/BFlypdtOOm+IRZulpQ+gPvn66qsF
Juk2j7SYJgj5P9eTMzXnautANsy+8b1syiSJqLL7YxjKhCEPxVujXB+Uzv8G18BtYQtVlUGSj2Ab
1ycE+IB4Y118rNVxFxjWhS/Pq0VPi3TA5uK8FvAGLtoJQU+ZnrF+wmiy9nFWiJouFzzEMnHDpz+f
QkwRrrYSsMD1EzIJIpx/yLf5Jkp4MAAnhjhJKFK8S9Uy+0I5CzsrtRagrqy9ILJdQxAfWGtZZF/g
HgO0sBUSzjdWwIgFqSfAnmvaxL658UWCT2+ubO80iaFJZq+6w8tM5o7qa58ruRAeDzcEd8xUrBjH
nunbWlTu/2lUW/wmB9YaTjep6wDnXucMIyMnKm8IEL6D7GjhLF8WCuTOqslTf2kho+m6AcHrjF6w
5xNhpuyqrUfUgth0cvbMBJsqzM5COB98AGPyLQAdvrLJPdgXtj+ev5nYOwv7wkoaPY+FiHo6WI0u
uBn9ZB5fbcF32CKTYJCa4yaQiIFqrQH/7tvsYgf40to4z8lcK/wMiuALltSbHX5SfziEgJMRpclo
vhjGEfMtvg9Kz7Up+S/LmleTuzXQ5Qapfro6uAwg5lGBx45jpXKxsXVAkXlglHUmkgnLM0PPiekN
iMWSubPdk2vRc5ysiK+oSmCTE3pKcvtFZ5kMAXIPRtvWoZVJ2yMMSUJSpdJCL1ZCISQiaX535iBb
aW6AirgnU20dHgARMglRStYZStp0Pl+t8aayS2J7XMuLXFHkxckXG+bdNB7jO01AD1dkhbXSz2rX
Br7tHjHI9JzD35d7HMeZnBziIaiA2IhNLKNwOD22d5gBu3VmTuviVPOMgSsPTpJr6DAQucZkXB2S
wIXfmvI5h+Ju8IonWb6abSBjP0SfGJfYtNYtwm2b0fr4JwHiaz2e+r3+aj7TV6OUZ/rJbYzp5DwL
xa/7XYFTnlRNJKMj+T56YxUPbSSGHe3Jmyq6K7835121cb2a3q7lORrGFRz8X9FWUNzPXXj6uI1S
3CjV/DjYdcHA+Ot3d3brY+jTOJkPJoPBhcp4llmNPWLDuY3hIYEs7hLuHpFb4QSH+uwowLvUoZ9/
wV5/llml18XJ3Ghm8T/NRGMHE7ysDKC1e1nl3Z1AgY6hdnIPXuTUOWG7Nju1S0MPXJvXZN9Ym1Tt
8hfhAcrWuOtr6wErkLxFbeJbfzEnw7jYDJUAHduG84iiNr4CU1PuO1JSPgswK2Afi3Qzf/mbgpaT
LYSnLAr4T1VoTm9xMH21CIUbSNBDz44QkZMDgvpHObdDRvPWBwSocYRvz/3O4RltZxWyaZfy2uce
H1zLaH5miGtHCnhCSPOLmErT0LHSUssEVPMIrBD34iGaJOozwrhSkszqRCmo2LMeZb/fJBQXRK/V
/QXDmskQK/7MsUG9sFOKefBae6yVgc2U9qLxN+TwbHtAAuuQxhYPh+RYCE7oqBQa49CddGAp4L/1
BGgHbFzBvMPitFEMJlIa3+xYe72AfbBA/tef4An9CIwfDoHSXXafXZ3M80fUxncP+lbDFJ7X6+fr
9WnE6xfgF2QZTg+pQXaJ3/fTOodC7JP4uKeWSkSAUS/TMD4qR4RD7sJ8+P3uF+IAY+fMs/uEOFs4
gTZ4SRRoffsdgXdJiszUDAqBUzsI9wxL5FUqWLnaMil2+XRrU6p0kAub1aAXHo7D0raaoH0P1Y1p
FEyW+mYtJehhpKRF8SbAvjwilkMs46vriwjlcVGhkVhL+tjPNqnzPoIrHCUzGfQjksuYV/ercyys
LlNan600bqXPDXt3o3r94L+geZ+0UxUWMMPXLs6Z8cXYtB7qoonh5hRKkv5Mam9PbFSInUQWXLZX
hNUgUvsxNmhmKtK9Q7tcfjYGc6RED6Jrp1w3yodyuumdaNtBgsADX+aLVioPuKz79c/D7o895lCt
YST2vME5Qd7t/47dmPOv4Au2n4dlVLQIvM/IABouAPmSKuL1hXLjBrBwZHHtxjQ/VXVB86nTh2As
TeFjvpXau+27A65tDMlV9rvrJFI+1Syz/kgBL1j2ng0QYXsNd3iPiYSskD3DK2+XW2eEsd23e5PX
YWp+SP/NNsb1pkIT0Xp3IcsI0dEg63zJxkLM0ZYQT227hP9ix7y/WK2OlDXnC0NCmUBXGw/diFmb
b37jYHdfVrAINNQtvmozws/qh5J73Mjz6Hq4zZKFeeoPKgwy16vW/1v7Lu7CeOpI9qGJJZW3buPb
pBhPoOwCuLHbdAoTi6dDHbaG2EJ1Uua7MljI6QlB0pesQmzBMOxD+DCKpoLb5RQsDADO/B5kRrXc
Kf5gYPalqcbzxE5nH16hopVl4TdK/LWFZKsXSyRpGabgPQpfzPo14D+1CAXMELJ8OgEUjOem3HBT
ep1Hhom00smi9xsaxy89Bgp3wXm8CknlGtxRWBYgMNs9qb5mHoq+2/ngKRLsvEKqOal+ZsSf44S4
/L7GPJWeN6YYWhY+uhiq/KopPpwI6AH5vKOgMECmJuhlLlt93jTZqqBKPNzR5BXJRnf4NBA3ql0/
lBNiQhhzx8E0i2F+ghvagtPwMACMvK26e2eGf9dZvx8iKARB7pIYx5ZB9lyJ3qD6EFkHGnH6cYIU
VByxXdPHm6x23xxqXan+6UNoBRr0WadNq6xi5JTDo6p+FH5CCLBJacUfxRWjtUYquid3aMfKEBGv
Pzw0CxGDt2AsrLpwhliAEsGRBo/wV8a4R1Efii+726ruSi4JDdL3XwzBBXiqUV8tmQuSXqd+PWhy
WrUBHdt5vKKeDg+daNMYT0evhKwpapcVdgOHNbhkkNjR2nV9mL4rALezkC6fvw/y3JZr+u/e05Ee
7QXF9J7XE0OWLKmk+P8F1PVr2k/kr55XomHQP7RaVQGBY9vnUTBc8wSCJc2lwm4l6PZ5ajOx9YJH
GXLux0fAUHjYQFmzhlHWmIFlL3KzqhKOp3cFcVccHTW4fN29YROSz5GDHhk0nw2i7VvnITWh1Dha
wfBVZ1mGC17QoIBJx9lrTuAR66huKXZ/qlT0zEQfMFhZVj2TBMalEQwv9UzbWTwJeOfjKU82x+PW
P41ypYfrQNc2Rj0np8rM/fovk5T4mC3cuB9BDIg4cia6M3/oPk1RUNutRbTqtCyqHFOzbtQKgJ7D
6rAJD3XlMkje3s2YT/nwMZzHMtAgyZ83m5JPq5oWisBc5a3IWCioPzJSSt8OkYh/Vimex0JaCZxd
3iEIgggn7wjwryLrV9V8fto54K77BQ4HwpbL+/hUkoYArRT+q93IAc5FhnMEosuB/h7TDnVpnR3g
noGUpm02jsqogD6YmSjbNhLppol1h03bY+9iewj3kM78F70rpLM9irOkr7OBVOU/zK7hseW4L/XA
zavgUzMuoH/AmVzHzg3YmK3dHvgJ8Klnq5ZPM7j4f5N7t8WywQJw6v2sZVrlVM6eWRgyfmfdZ5uj
oOicum1wesNUpP+CQjEIbP9dtaJY3NiQbqwuR4QPvyOnWmgjJzgcdK2CJa4QzNUiAtHOIBClzQqs
a/Rb93DvChDaEItf1vy9lnTosFHnw2gCRqohVeJdVT+h/KJwGTQ5Xnr4UDajnJsVJQuk6kUgAMIt
d+BcvwJt9ubswcjiKwiRStjSbiCozIb3wQOSiKk8BSmFTmu3ID58wnrWYSZi3zwnaFTnnreEFNvw
IofP2CLMvVt0W4GvQ289xxZFAyAQ5FM5GI0KowtZFbvdL00eD9G1LFNFYRf7KYtsIcuv9h/hGvoY
HaeOTQPLOUkGtsPOrh/TYIEXiViqgVAE3gKnDy0PFgF/I/ko3koiGeqqFiDilMNAK0togFjS8OPc
8+zj/F0po+TjsORGFQpjhBGg5fy8btdE8Q+vXRynE1VICpB1A0LwvSbKlcEMA16veLSxqCZmgfSk
DfeWUWGW0vfWiFCVUVojToKWzbuX7jaIXIUVWYVlCExSg1bGeHi6UpDY7u/uOdgo10/u9agw/Uzd
57RbGtB1kVmyshUAW/WDqEoy9IDq6ck8CyIjz1QN1d87roO1EGpCk8Kc7kuff3/dHIdVvS1tEl8x
5l87zGO76V0M4vLY9yG9BGWcGpFQPi+jA+Xm7r5ij9ZlArLd2NJ7GzKE9YeZvrzIE1lukit6sQE9
ra9WPdLIPCy7axcN9y7fgVNPTlmqxBd1B4QSeLaIMHZ2KGAd51FE3Uh2elmQ/bYj/L2cdwwOO7Y6
q4asXE1BWf2OAQBzpgzsKUj59a1ob4ZS0HfutxcZ8Ou491hoNjkZOi6jfBlMup90RZg6eV5JIS5A
bmYQfl/zzYShX/bd55nU9xyU7ss99uN+6YtfCaHBu9HuiqZwyvHtwu1zwGxHlTgdtkA9rqzicbWa
/SBvVIw9MUfkIxHduZ6UzV6pgg0W2KdFeXo39ZBtZ6Po1IQ/62oopNP2NDETbq0JycWzKIvrVrLN
T0uEzayY1gXqPpzjeosaKT/sYJT59C78OmWY6KAJTgaHUpIA/rByFmXmhhfUNJCRvTROzLV+UAEc
V6EtnVbuVJtdsPXWpAFcJ7B3RTms3L23xPZJkCRKHS8hkVbT8cP7F/sWt4gmGB6NIZWbz56APiz3
2rUkfQWiUCCj+GeeM1sUTWRbrjmFM0re6Q+e6f8C0sTYcI0VsUnOKz8s2fqCCEdTIChoEXQApe97
9Xtx5ldVN/e4DYuveUgDo9p03792zyVGz7DDY4jQv0hQ85Q0Qxt9wW1bx1bLWW7+ZX7h07nlZSAj
1NfpzOkbc8ioTuPLv6BS83eU3VhTMf7nTFqh7NbitXJnia3XQ7Tybj60tIO+fcA5dD03jUaoAlD2
zbQAMu1laVBsneQMPpnzhoGsJHyGtlr77TIEG/ZfsKjUaDRHiCtmU1IgTMwUBULIpQh4xIdNuv8N
CH+fX3A4Mzn7P1FHviLlwk/ARbuyP0NMJI2ur3635h2z+fOuw/8Lhr7/50dm44puTFsT18MiBleF
INvU6RjrnqWudojCwP3slvXPENydQvq+S4DHUFpOr0cj5+ggHcS3tTwxt2G/MdRku0F09nb3Alxk
YySSirRj/8IxSFUmL9aNcz33ErsPCFHEwuVFCIFFd19YBUUSaBd8NGmAaFFqLB1GLYNFzd0iWPF5
ddOHg7UmTSRQgDVD93JLMKUPxuXYSiipGnMjHwGFtTMeb45vqwgh3sOF4f9Hg0fskCYIUSTaAXG/
l/9pS3GIQDgK4x4EdEL32Ks3JH1LzXwn8kBXTHSatuBC+PSNLbMPFymcQzXb+vAQLGzpvbUAqo/T
qqbkvZ6fI5fzmPpoPqYMK/MxpcEX/TH+lpzF0+wcNjQAa0GS/eW2NDCh7Rv/Zmyffh10bm/TRTSK
7VJsw9nmz9dKpM9W2X7Q9AgD5gB73KqCN+4022Eu3uIj0pMvJB0eFivoYbXRlhTOiyZAFIrFb73o
rQrCc4zhzd4OBe7HNTtC2fYmRplb8YcOlmHiLkwjKO0dNCTSs23d4W86M3/8e3jjONScGm9L/wpt
e3dGC/AynmhsfsuOoAEji8Cf6oD+Fmvjguc8XkgVL1YVopkv5ExvbCRDsJ31mz1+tK92dOxj/FlT
GxutkdAduA+52KKKoWMhr+E3Mz0cAlPqPXZcWTOGk17iCHAjvYFUOI/MPApdhVXOzgT1p5oLcyLd
JB3c/+RJSRYtAwz+D09/RrD5M5D7YEpkLl6+vd0y+a5x0Qr8s6fRLl4eLoEmbcgo4Sg5dtnA172h
H3GpFWTTDURw+Vx8AAodm4JUYIjeUA009ir9TXqheWIavUj9qflNZ/V+AtehIMShXlOtA0nBLwQ5
7lcuTWuPtdAn+n0G+Pa9PQafLBi9xZ2Nsidp3BDZMMg4fGRqfO23kPkoOgKBkOQlVi7F4Oi/ldqu
EPKj0P2XCGD+/3Jx4UCfe8iljEP9pF7cKBgxBt+LLy0Ve8m2WwTkTHxrhW3bPXbd8bsTl5iXowla
etlSs/Dz95Of7kn3vE2unZ8nbOtelWdZXDlNl8q/avQWrA5K3U6PAxIMCnloTT0qko7vcbDM4lVc
AoczfPfbfTWxneew2rCacEDusc7XBLjSqtYR37CROvrcirNVbEIZN5en3oJOBgRNqEq3PaXAxhQ3
0ztB35YdvGHtFOTyqB5/oi7bIiBSNzGRLptea0LYFb86Roait+zGSIzZqEJDgHQ1ivD/xiZ145uE
Yq7P7c2h736NA9t0omh/5Pi12GUP0TcUOAnZT5WyWghVG9N+iC9eT8Z7Dhix6/6rqIkeJZCmd3ay
3StaORC/xE/YvpVi1uTMQrzwR+HyYhIkWpgyAJ33kzvfJpPPVk9IAI9+rVC8REzSipK3nN0zNeAf
UF1zkzCMYYcseq9KtO8xcRGw4JMVqIE9cdZaJRQ8j056kpI/kAzsppIaWHLqP4JhKrHasXN/Q9wt
X2cQWvr2BlQ4v6SGG9ynr8G1cBWREga3isPPubdc/YyTBPypgJ4HAVnmtrKLEa4Uv/3QhwtXauXP
sUMKkB2qQAWAV9SlQQmUCYA3skNOXYgtA6vqjc3LC+1NSGn/F28P3jCMefz9YdZ5vKQI23roriBK
V/ryjqfcndrZPvAJY8artJ/hshzTS9jDlyI30ciuFjIceUDc+YT2fSsaoYTWYTJoF9p5ThmFBL7e
A9pPkYG3A2E/X7CyeH86GsntKc4MtPB60TQhycH0MlEzBj87JUqp9Xv8ZZEIU7hStPjqwfsBOldE
IPX03Vka+Y9iOFF5BMq2dBPTJOaN+N0sENEID6zy1q1X+NtTtxb9Yu4wsKJY41lWJoOCPPrR8KNa
C5/mI3rkQA+aC7UW/tOw807O9HADzrdDM2Y4tOZnBOpi7qetGSdWraWf0kmMr2mF9sZdpzl51vsX
TgHnZz6MOVxew252Xu0CgkQq6pljp1dEJwztoaHbwJQ485HfNaen2kUz10gmKQjoZ0CSIuJlah/T
k3smb5I0wuoet0aNzdmwkvbCkjbUWhbe6tprK1oBMO2u3pB/8oWULy2YZlUWO+pU/JtQMzD5JuQq
CC+WfxD/shyKJ5rUIjAlmlkBLNv1Y2oOsOeGtJaoe/5ZRNQosNklN5sV5wyeFBr7f6awoizdqJJ5
f2IRjVeI5apSkodwp4rO+sYxawx4lPVIe3v++KjazVd7s52PhYEpxEB01j+ekIeRAO19mAd0C8+x
5b7qbzUb/ztTj3/ImYRAtBM5SF9FnUvN+kULILimU8Y6ac3FLWUE2jjDq+gG6ambSaANa0ZJnHxW
U2oe4iykukP/b5eB5tOGfGnkNhwT4z0KmzalbTkvHRwneZHEfPbL2ZHLXK1MzhMDWwUMGss6dDSi
HRAd6rKCQAWcGuCyi2FZwBGo+PCQnIq/yavWrLARAumSvRIowqjARyR+P/wcG0vN0hIEmS2tT83Z
ZHh85omEGNi6iFdOQru6wGKIwQmFVx6t1MXjT1G32q0z8YTQ5A6qy+9PdDsEiDWds+iymv+7WlIE
64j3hd4UI6XkkQrtfv57hVge0bPTJXtEL7kE2Z175oEbfGlqqOeHmq9MOhR/Rz6bqLoEHbaVsFRM
T/2xJ0gWsMtERuWtPCk2GkTkwhS9aOul+0qlv+8VD2vInDMkbm4q1P5joWKooADSNKQHOPQPk3kN
YtuphfeUihH23ZVGEc//rSWwhRoDLbXjtmYm/LPtWjIETkmw/EHLBhFpKCUM3rGpNncDUpun8qPq
snTv1u2WrZKYlbxsumrB4FDP+mCkgEb9FuGQm1yh6El4oJdNziq8DsD9CYuAFcHWcPmKbUPZlJhK
8640h74MHa0JyPGrE0gw+fuQHyiMT7QzYpcDrqnopWh5nH1pDwYjytbXPvUhjC03sXuvsBBSxqeH
jQOj4bub8g+xup2ShRL3tzRNqDakgYmYIGV6EltfN8NBJALys6hLUNV6D3vGhfgf0AxRUTRm/pEu
WeuefndwLlVbrX7OY2UMAhYxN/di7VMBXY0AbMco2sGoag+JqrmiUZO8W3C7qJqiX4P3l2UBkOv8
EpoGG6ikvOoG9Z/jA54KiUjnO3nnqCP31icD2xL+o8NpRuijMf3I4sDjRSmRVeWOjWWSMjSy9iXP
/UiN+hVOo3v+PYWq9iN/h3qrZre/daU87HN+TDgjur1Lll2W+z+E69rKeqJza+nyOk1T4cRBQIfK
8db7JKtaGcei1JDEubNtuJckOtyvfpzL3wYmZvNGMBdUJrHdtwDZcLI3H3Nmlo1RstrBmktPC4X6
D+DGRenp5/NGHGAvtxZ8QsGMsgi8KX02c0DXVCeSGREbJA4Pp5HXCP9jSWpZ/qm3Df3wfX/FcTCT
lDSENFSTKw2f3AT+JamR1xJ/O7iCr4mcuCXg313QDmHvf4YuOoEgXLSuSqtAAaBVTSyc5kXqxstr
614Mn/dcwEk+Xhgt9FTfoCn5VAPW/rlS7Hq8g5hHuDbREw1SHohktGghzsXbu4K+XHNjlikmPVd7
ayO6Vyxtpu9IUvS9uT+inu+HjFntqiwwiD3usHlCxtL9ippaieWDmoVEjEE/TkXHort6ILzt814H
qREYyqt5hI9GW0YUZ5uhtTbZf16k1d5K97DDYwsYcoVM5o3vvKW13hgMIBb1iOMSJba27ZKLs3yr
pX6qbKLKy8qSuPd17yj7FGLX+uhOmUvSnicSnkaq9w/aGUNeBHEJ90pSx1Fy7XTe49C022jLR+6N
Ds9obOdUakUBS5MGzwhVbMnjbcFxHOJJbATzyt95ODZJtsX6WqocmbF0qSwtFYbF3xZBh7Fl76i4
y72uIYHZL/mPd5Rsi42V1XBq/mBrshPgfMDMqz79PLcKtsOVgJd2RacV3na9EUcSoDKcoLwfcu/q
fBaX4dsLZh+LcKJ/g4KMjHfFOtrlHPwYyBXG4PHd7/DrWPHtcIChXxK8mfr6F9EXEHn/4xy8bQES
0dLFImHudOfgajQYpXTm51lXDKaDurdm+vi/v3jMZD3Ar5LvQsnrZM58FENT/7H578LYzO24bLun
rPiO9hEBpZoxHtqEi8NJn46xr4Gvu9XORiX4UbzIW9ZOsXcoO+Q5b60bpQns4G93KWw4LEYAw10d
WM7KdXst/ddCkCrils7B+2ozBldoxp0Gr1dwxczHFmsUwLxYFTyczqGjnM5Jt2OI0ZPult2uB2b1
4kbVIMjGUIau/TDRVdSMNk77OyOV/kgxQMk/ePCVUT2Ul5aqiWODCopeJmx/4bH5A9SxO8Ilp+DM
JceVd0Ry3k+po4Sk5RnO+iRbWJg4dxqfwnuC7MoyMKkr8MxPqmlxPwM3EpHzFqTmDSdufSzhzDpU
aVpooLDIjbZ8Fi1NTT25gzK87YgKZJ3Rz2SsL/x/ZjM9TGEvkXpoNLlYO95GPERGTvTrQAfeF4pz
uJAIJiTknRfMVfftW/ffbw9lPyeTBPnzSLvmxX1qpipce9nNvv7h+gQeji/GU50txoUI/nk/Z7Xe
C9r+ze9tnz7BZoZVrIRECH08iASNV7Bspu7b/ARcvqNWqDbdaqc2ZNhJCmWDGmfr97Y3Ne42jFma
0p4U2mAjFrwvkBPHVYoXUCOnXVR1A1+WbCdmolsSCFkDgEVNcJbNJ7x1LbWj0qc6c698Ze6VeqIF
cao2I+HkDzCkEYv+HSmo+ON2AIGbgp0LXUGA6f9+u3Zwu997KgviSQ/RFiWBugyekWVNDBLScIV9
6dgrawGN1tVKLiKa+ynYVwkwmnLSTWFf6ULCZXHVmcjIxyScUbWEJqYMW4jmFK4JDdIUKtR1nvns
gr2rfRjN6X7qsA67lryq/SkZJHBol28OaDCE+MNdGRdIHEIes/jpbTfDe3Gwzw8NVFgXBcie9iDR
GBzcpoRjG4IaTnJptrYXGTM5vUiUUwI22kbYy/d0woFswXCSJdU/cZbYpW66yjGGtVxWAXUa58KY
oNMHPzN3GOl3ho61OtN0+U/HuLHt/NEVhE0dSlPdCDi/D4997yCL+l+h8JvI8uH4Y8Tgq4IxfM9a
rriWaYJFktAMkxJT5Ed0NmBTPeutn/yTmkbx0BTMlDSur3LrTDwxI4zVyEFiZGJrWxWvKe7IHJIp
okiEd6YUd89+1E0G3W5tMv4tYTtwXqz2r+pMjS0lDB9gUIm2aTztoq5cqNO3dkxx/UD26JRnQ93b
0lPD5lNklK+gD3fu90KMCFkyW+HKMLRPD7oW9MjLBiNOVGEYtDrYCWveM44BMOQ5ekPUgxDk8m9o
0+pZ9BZrCc309QKgrtKGz01L67WXxDS87Y6otZm855RDqc3vdag18C6Y6Iw8CfrY/7jTc9mYczVV
oD7VHEo0Wtos3pcB58BF6kU3eEnl/5r6SVoZzfOTerwIrMWTW3ALJufoiIl2RehRc11oAdygLGtA
2jLE3hIsvw6iAwzj23CuRqpCGTqTesuX2Xj9gVx+vWNxegKB69qzGnuIjw9doru4M5H6SQ6rLVcc
wcglgKQnGps0iSTUFxqKbNBYEL6qnWUYFlZSGFagOroqvOclnQnnsomwE52SVdc3YsCs9otJoAnt
VRxnOVITGpiRPdOEK4JyhZ4YUdzVgJHlrNPHECpeqLLkQwl8a9oAt0i6riuBpD6C1BBmDtijZJot
/E+2SzJb9GFoF6bvEl8Y1hoXP813SjpL/TKoLbbZ71SnTOBQEe0Np/3ZQm1v99qANwMjNSLQaOEG
AoibCXIBSeJLsUrfcR6+eADnYtsygzhj2X8TPYBQfBcUWxALwcY/zGDyDw62O7W489ML/Q5MsFcK
8t588TuTdwKmAHTtQqZPnSlD4XME0qHl4Tu9vPCY8aGzkoWi+6Zy6uOGFLq60O7mxk01tdPLc6cS
dx2/ZlfZe6XX1ZZ76HxAKLw8u94tfD8pe7MRSDIzQQ5fXusaJBqL+zMdYazdSlh55ymA1PnAE3QE
EbvaxUchp5OKgzy2WW9mPy6lDpT76YZj0Iuaq+iuOnK4zzpHYlT8z3m+ZY5Iq7CTSpz3yNsaupGK
Jf0TvDCJ7pZaEn17KXnrgy5ZuVctvmrepTAjInLkUy86vY4HfTryA8uQ1+6VZndEj0V57kluboIs
fV5erEOsM3blZvkj7348tZVHJ9Iem7AQCwYfxkUIHxVcLUSvAszPwdhPaFfxpvAv2mhYv9sk0UPy
tF0XbMb52W8O6GNmQgTrycWUxyKKnFgztSUmD+nfsg3B92soO3hqwbPuJQ26NoCUzuMesymbt7T2
UDgPXN9s2xVkYaX9qq5EO0clIoWV77pTZC0g4WuvIA8GtFfmdAr+xkenHZY0GJ/b+mGqYSonQ9JD
4StHwK1aE2czx2c9krXjmBJYNLD7DRFLiLjGnmjYIbu9pqBJf4TVXIMoIpEfpU8rb+RyvT+s5LRe
GdxyXPxbhXZSxQNt2uALQDUxqzinFLSlFsoQ+ARMV9IbT3XLW5Ub8mQfXKHADr6UNvpcT1sC3Ze1
jnh5l6lpbo2FOTenjyavfxjD+1vDy6iDdZvkDk5AinRey7cdRzo+OoouSDS4P+UO408EgcMfmU9e
FcLx9Yidfnwy8ZgUVD/Ga1PPwjSYZ9OA4rErWlS+GuIe+8gFzeJrQmcD05mGNDRWmRBDGrq7X3Ta
BD9TNWsQEAkkemd9cf4fnewfPhuVTlWCA/59N6pZifwzqHm8ZeSQ0YXM830y3IDcqj3/tLPXpBW0
tCn0lAw7HXyD6VXVkxqF7dqPwdXwOci/ZC5rD8NuJ7qYBeoMvSDvx0sEGFYSGJWuBQzUOlr+BFgB
7y+z0xrfUbwcu/k7LKs+Lv1hIxwtWDHO4oxShealsSd5MwSf/8F3LBVlwFLor51pQhyH7/tCAITc
gBoLxJx0eAsCJVcq3QP1eU7nL0R4BDTbPZo7XSq1Szx71D/Fui/PkZRMMX0UdOz89ZpYEUgT6Dst
ZZCzq5EILI9yi3ATIMyhF05ed0ekrY1eWwsKHvhEmBZdYkyuDVI5TAVcLe++OhUWVxIxO1Zh8GuJ
iNd3Pbjpq5zupHkzU05U7NshwkcvojgrwFzWzCPWagmMLEXQECNwYQfA9New9z2YRncKkQfVgF/L
V0OhyNcDwO4eoP5o473zME1lscl0I2oanz6Ms83w0VS9VFzTH7+z0chq4cAUNPQwullgK9LsE16a
Al/6vGaHlcCzSrINszToM+9zhOxQpYMkJX2aT7fCygk3GVk8wTnlU/PQqQLlvf0A//o+YSKW5hXp
GdLppoOkstEbs4xEaU1KK3RDp6+eFTf+aSkoh+WuuBlxW0tHHEMVBpd/xiv21j4Inm4zXzJhFmmb
bf0Ea2WtXP45Iqs0fKjQnvPUbkIrFt7DAUy1FADJ3tTvVDgc1F2mOBgG5VbQe5RxhRYcR3067aN8
wxk0lr8QGS5dotSW17Cx1/6bAhdl0wIip9DyXqSnWqYkKyOEZ7d/ZvqRAuUhpcdydZmNepLcdCDY
ijQMXNdZyb8BjpyIQTX6NLp+jL8W6AyDYLaLxGqPyGutrm9QOtrzdt1uqRXXMGPXGo/RaYyrcy5s
tIsXfU+tueKtoxJZhsxakNtPHyqfD9IyQ37ToVfIGyDxVqb8f+1HmTnit/vG/zL9v4JIhJu0kTRy
6nF+nvYC1NWuRxlr84ne2go7gQveSTQ3UCg2zgFeP2/+5TdY8dOiM+lKZ3MO3DCvL25eNDppz2Ri
NjNPnU4y/yzriLoCN0tpAqw3WAEvZv+eV9Reb1btWfFZcj2XNIExLwkBjy3tdfOCE1EAHvsttbDe
jJRvVDRb8GmqYq0Pxk9OVlh7xst5Wrq82bYnNnofjZD2Tau7hl/gILe6pXkfThj2LHY+77UCqywS
OC1nhCxBUAQAZ5r0Oz4zb6kSEiwJEhP4D9QpjueGfYKOG9vhw36RdPHojSc/dIq/cwcfsVm7kfFs
7jDmNgSFQtCcPBhv6WglzxjbOjUXw/BHfPEGeOUW2CplR3RWF0bZ38NY+2lRRQ6/whB4BRRYeflb
3366hKpfsi9iEc2KyMOZo5bB+7LH/sZ2KpdH3lx21zKYE+HqyGlYbYbhASV+rmmBlYLHUtfs4ypc
Y+8nxkHxRauPTJOWvmc2vmvEE0ZxXibUPRFEXlTC50eVCE23Nd9n0Vxr7XbYDmAQHbEOyhFXDjf7
tK+3wu44mVgctT+NTnvnxo0huiTlysDBsoc051leDMsNg6Gu9wbTgHTMTIGPzcF1II+P0g9jElY2
AYi/x0gog/yvuLHy/+6L0CJHbtUST69IIhxANRkSGqSVaPfvuHfxYiD63qgIquPRru8RMLuZAfi5
bDsC9MDA3F+cV3YUnM/NQs6DMImvu4e7KLkaN1/YLfADtTIPr1Pwfba34bp2ZkE0qKCqqqbquRq1
XCaDAdAQzXSUHKXifAjq4eM+nBXP/n561EdT/1v5FwmW36v48PRas9xtisKioXfxjOrQCg8bo10M
pVRXdIZ0iv7UuZ0kiMH1yBrbRKT3S9E3LNzzmwXHeACzhW11ZbwMuyBTJ1H10xkThcjBllRbdbZt
PindT0OTwpDaCJk1z3IPcBWYItWND76YbvA0dHbdcZXWN9kIx2zB9+Oqfy1wzTLKKXw29D7OmxdU
7xYfHldWdCCKJEdjZPdf++ZNKWgzxUAp2YKU/34QfhaohAM6S13l0y+2PLmCIaTmrlz4XuzCcJ6i
X4YAWmAIXmVNMMUg8zn0fCgWH/U3s8cINlfbBfc5ZRNlzgpbzgeyNgVs7D9SoxxyjpzcfCK1op1R
k0krtin0hxceHzUvRP34dnIwzOLn3MbgbTAinyXiYwjE7+TzCT8z+S0g9VIQM7NW7iK78q9GdxZ+
zFmj0ZrQMZk7sV4VmRw0x9pRxY4YUb2m8RqK06Ebb8Qas5HkwfMt2ydwR8wsZtGjctaxV/sDhgSA
XyEu5aMfmQOjpDKj13aHqdiIMk3tx/84/ZuYOlDYxAufqkbPmwUunGCsnsLGp6mlRX51bPSAZUAo
859hbdDfwTnkRY2i3Vo91VcLFE8aSLEbZIuoInGQSwjcp2mtXJmJ7+8r6c/3BY3WK1urrSk5MAGr
0tr+a3oMZxS/mQhDLFXQ2Ub2duKbEqBDYOGM8s7qgktDKcTbfhAgs6jp2rdpq4Z00/GBWOdEZ7TG
voHcjJa7yzNpWxPhHwDpcyMFoLF9usj6Hu61s5Kd1tZ2nQNMDGBW8DaDf4CMB9fpzZ0Eqx/O544N
hWdHYSfNFpCo4FH1HyXFHfufwIDOFMDCq1an9v294ybJ7U5ORou+MP4E+zVHZSYw8J+JCSeZy4ah
g8oq4llukDxlkqv/WFL+Y1h91TJtSlrflpsnTRjNEa6nnohfhOOlOsjfI7SrsOTSaqgwoY2X/tXW
j+l3f33DaGxkujXJlBC9sQL/l7yWLhTakcQjT/j30DYUgfaJ4RUPR/uu7i+IqPDhngOeuwBBbgld
L07fNmWMry0roQSgNZ2SlDJrDKm9Zl5Q0C22YI+E4fRl7/pbXZOlTK2gHX0BKsQqIHUGIHcZueSc
e30V6IucevyPSTM20eocUamoxwmJSVLCl73NUemTMs0rpiELxmZAW23oHPUBFX1s10Tg18tM2pSz
3KmA/zeyzRT8FSRByTUR/qmBUmCfNVYkHmynBCK0HcZYOXcjT+Un6xY8ncdve27cVXWVISKHX0e5
25qegUQvGbW0Sd3bNT/hNpeIBZmcyPd7MwDZmbDwkuL/JLYH35tXBkHavXQKN/knvbepZYSla794
KlIhbjWJd3OPFYjhoI1MU7Bu18yBmxxDUAlUYA/vowkbBRbeByCK083u5A7dfjDyf3Qo6MZF15U/
pfAJ+3ppXWrKbSN0BPuryOx29kESeCioS1GItG1IGDJgmXhk7I59KVvRd1EyeUEYx1gn3+cKfci/
ClrttJgkx81usz96NkkFWB0eb49DpOT8cf2GmNuPfg9TfmheOthL2RMxSOzvnX2z0pXlU5UYWGO+
nq2xJRr0GYH7eqyTfi0lbtIBpq/Ug1W3OhDQ4eXhKOT5nIk8E+b59o00ByzxqL8dqkrcocXrxEna
sOIjbHiR6aG0wXC4ZT1seYh3+blSG6LQfRGOfbTNBn+k0ZCIt9b5i7lcqtd98YH++nLo9R7X+HWq
m8LRvo1tH8aIukTPyqdmCbnxRa0uU9x393k2pdL0Uir/7sgdlLJV4jerUDJ84aGTQIm8dpGeo9MM
v0Frcjshxok1wEuy/PUSPvRW68dyPdqs21LpNTbj2N1SYRpWkrvkMv2IdA7ijQlvWXliEEg4Bs/g
s/bZ0L3OZziUlRftIY63N/DIAlHtgiMMqdYgGIHj0aNm1mDxnb/p/z0L13ay64sfTFuMeZedlQh2
jN4s7jrpXZ8cjNOf0HOcVo9jQLSDbzQTo1EOu7gE5Bxq70NpTgX/zRbAcCNk6llDgJ6kcX8oBeTE
vVa4ten8bUary0z+I17Yn4q6P018XgnSh30HV4rOf9Qbqx2cn8qiYLBrR4rUoTQn9J97xj/6GkPG
4c57zEgU3Cp3bFmaTNLtXrvjeNwKv19vNZ1dntxjt2aBiyFTEVqalKDde4O9X1zQ0BSeqBfAUkaG
ORBDr8BXX4D97C0bJ2KQGtZOFYtWKUS7upzmLl8tyMyrHOM0MVgHz3StOI9Bq44XvV0qatWHVPDt
UAsVREhcWpekf9wkeqXMaaKXa75ANjYSpz5xOdJuD5DabWp6+T7XyraARpZyCG+J2zqtNf8vH4RI
27NLwtmq3J8Hp6hoVGpH5FB/kX/mDS53sJIaniwPeNBDGWXBbkASI5anBZD0ZRjmXv7aflcYBCY/
0WxpVTOXyJk6M6Y39KRIS3eNV/D+/gf6LNZIW+gIV78KayzXFqxQGOUnD3Q8+xp+dTPCCGdkaNjE
fDmr7p5+ZeOuEQRsonxU9jKL8jkzmKhsJp+DiTdt5xV48ywK0ptH7P1r6aCTyThEUGMGMy8gs/VK
eFnNDiNJmRn3Zjn0Rq+LclOT5hddP/8UHcr6cN8HMd2APyj7d9zlTsV6BTAnkHK88ZwDDoWf5ZEE
Z8h/Zfz3Cx3GyKKgsO0goagWRhQ2ejDmw7+bmXkYwDvpJzuOSXYJqGqVBO3dNLaL9vIH9gdY5D0w
TDKqpJ0XPekaJKCF/X9a669tnpY1FYkWRdMa0fjtpk1FHHZ21g6H8WRaJzp311OKhYKB2Yv8jpSq
q7G5HjnqVaWfoP9pOmhdPYF/9d9RbT2DZOeGyrVuWaP2X2XUbiYoJXApUuMwVpJNBYn/fnPBy1xs
MxLdGURC60IOendXO+jAuUQQUHHZm6SoXUOMaY+5ivJiF6AFMLiP6Iff+YyRVuMd4rpkdgpfzjOI
Ugf2hAPF/yDg8KOF8Y7lQAOAlRoit973g/BlQJEuU8gxG9fsBPuD7P+ZtOcLa9nxUWVAsnxUQdAV
iiCF/pMohmqvWeury3lrSsd3ERRVQM60XXe5Abnd4ayUZ0Vu3arCX1ZAaKBFSpOyN2YEueEsFlkL
4n4oR74+2FCLQrbYJuidY1hiCfgSGCiLR/poyt/PC2Mro8ymXh9gbcxczyPhLunTnQiu7cWVz4QA
J2cw4rIDhNkhrExFMvRa2heJv/qNX/zFfDoztVWOQdVOq4SxSn5r3cbOO+piLMYLMhynjVnWRkuz
T1foqOtIgSwhBWhX6WUcdklEmW4TCMqhfveNAqYvUgCHIHrQZpqbB967JRiso8MR8ms3oH7e4MrJ
6EiSGvQDLXTt8VfFv8+3/sunSgwhmWDo5WPmTspdGmYoBcN/QUBw6JKoFM69yCNGPsPtbWbZUg4S
3Tgn0Rm7U/MhEi8kistgouIOFO6DJvnhPzR6kwn1NxbML12wFXO4Eezzz/tXnL4GPGq/jqAdqnjV
vnYfb/i5LJNLUV1dgGabnjWrKBh8Ak6DtmKFn/VPhw4liQ9vH42Ja1qLfWLE/QBmIOHMO5vH//PA
ZdCXEcY5fNRbXbi97NWvTus8kGpDF4HblPHCYyuTFB5G/+ChrpRUtWnuoorUO28Iv2txxHuflifn
k845KltD11G1EaIGlyzsFxw4JOS2rxFWqmIJQ/htWQXiJ2BRPgn6GtqzQqrR03+QJ8ApsgOTeC5W
xMAZ0Gah/DvY0XwCzEKxMjh+gOWupotOOjtlvY0AaR7UgzZP0cpc69Cg5dTxBAoONPyqkS7z9Kth
NmL49UL6fqgY7eL/ogkhhDTbXYI5iz/EVMWhavvX+qQa4rasp8u5EBF1R95b7Gj/rkpOVyc+KivK
xu4NAAMqipfNcENq2HQM4mVpvxlq4gPILDkE32Ic2YBuFqL2SDd5UhLHwfFX/nL3tJuWO6/1ZI3i
OVaUpS/OfQl0Zfk8StoIX9GBjPH9ueAnwFQjVaPOfgs/5qzS6kBtF2r4NPCach05aC7qr2RS94L0
lsuM5o6P1S5nXD6KEmymxjWLV0XeXPfFOv0n2/gcDvri0ddS1UU2LLQdFPfmogAUGFApKjLg9zpP
Lbat6XE5gjwO7MbHHIKo6oSZJXHQYmiMpK6I1CoxUUublLXQKxnc1iFu6/TcDJs+736VNR+NwNVJ
1mYljo6QpjE5WnYBUpm/TXA46tjoSYMgSPYUl9w0bPS+o/80D/E9Pvic2zffULbBXHiZ7EN1wbyE
ZCmVs9qn8y9/uNgHJUETwsXQ6O78Yx9AmY770d7fecIRVlHm+iFHAsm0rx/pg51xCjZDbaoYaaQf
WZ9Mj/oWP5eM10na5LVrBTk9nasiBAhvPcPJNDvmtKMT9+nId10I8xDj5vMwBun8Vy38OWh32dYA
81nfDyvUWCBtc+mw4vmDZadv0EQzfg+DQtDypXtbu5eufZb8ADV639vi4s2LN1fFA/KC0xQXewdT
beSgB5i/vWzXpUyYOhOTrL+Iq0LZ8iTsCmqw+7dL/DFQSnk8unzsv7nsm2hJdsdSQCm46YcoziK9
yIVGExD44tXqqCnlmqDlxcfJwlXgMMxFxhReGahO0RzW916I6w2YBIeMEH5rsGwFsEkJYKdHSruW
qVNg8b2wNU5ijFbok8LDwBA/vfnFnMYsEynZjYZ5YPtji3hDYui66iPR4t2Iki5K3IGLD79oJZyh
sbEF+v/XiWjCxwNj8RamE8CMyeMZtrWKeAtVgKRzjVpoOWpja9rDKON3feU+lX2ppKQvnZfCIuug
dw1ShHyGYMZByU7LVn0LygE7GVuDzwanYVtmaIoKC/A/DtGpyCA52/pqun4sWMUzhBoRJOwognrO
ij4vwvoLnn3i+AIgtDsX2G5R1Fh5WEuad68OKQ4c/8w1ynGiTj4C9t/Mu1YKoyc93TVrYAzdWh6P
DczQRK5mqgn8d+I4cgEgU17tHyZEmQA50VLA7iQlSBB45p6o5z1FAxCS+9Q9YOyTQ9Mj5Ko1UJlh
GMXgoW/Adegv9CDmm2gfYwYWtIPzu0CpKSPp3RZPGcARRH8ZAKlZBfhBKZJaKTxyNOewG1J71y6m
qGAVck0LsyFNbwrOfvFMaw4/9PZ/MVn1PE+aCEcTNBeaAzs9HAyDbSufp5dz8bl1ilu+MGpcsncE
Ezy8W0Y32/marvKzxT8SIN6a7LPla9YfAIHkQNApaSJMNp7os+sXeSydfTj2rurge/9X4gi17WGj
MCnzx8q4nvvOnAk081/KQOx2jvoU2puavXI000ktKFHBG/QmgLB76YufrvKhGsMLc7ibcgGF7AE8
Z/v4JxwzZ6HqKJY3RT/RdWqtnnaOe9tHr0I9OapZYPaBD6jzBdmH6SHa7VzlXmJSTth8AKl6DGni
geJMCVmHXFTGQPGIqxBoiOcEiKwnq97yVw3loiV/PaDHI1u6JPbC7aBnfrt6Z0USQzY4/R/GoKJs
ZLz/dabBkFqLC5Uyc6+exfhmNRusiEqwBOf314neyIFbd3RvUIHEHiKgnmErYyoaC3hP2Zq4YV5w
Lf7g9jmlAzexggMo8+nT/CSFC1JL+pJPWJGh+6dhXGMC3L7+O5qNUiswHzkuBB6DOYkv1X+TU27C
AFSTqIlKr2r4qZKI1MPZNxArfhquS7JNAtKiridIzm8RFVeyJcIeY++KX5HgRLXfSNdNa5MWuvxz
0pCF+Wk8E3C6JvEHdmuC/Qmq0knqQMwz2mV/4HPROoqgYA4lG3dv23thvJDJHzwge0OJfIa9Akoz
dXzRFBjWWBjxjuox6EAFtx5e89zaS2S5tKWrJedJ8rLA5vCBiPhOVqDyyy8b0RnkQ8EbP694BCM+
NDP2FaxR5LaF69Cc8qs6iY3UOXodUUCcrUbu6RDIS0Aij46RSDjUtg1B0rSLZkzJAV+8wh/Sm3q/
9aZzA+kEwTkZnOdAnS3dE90oFzxlQ0twLSKJ0Va4VkIwfcFz6KkHwLpXhybkgLasrPtDgPO77W4a
Htnll1K2bFMnNMc22M/B23AdWdXy7Gjjt/K2WpRQYbP2WJqmY5lmhQHsnE3b+5H+jPPNFSbBvAKG
XpyqR22JJ6dLnCmirjuTmhP/4IDwB3FIDPPP6FGRn/oN3fLoq65EoFQ6ydVlbArxUyrrx5ohF428
Kpspso/+lhJCzqp8oBISzj2Le2IQNJCYvfN6AN+ocGTi1xkFtlKPv4ZLNexKX1YqDS9v+wNPSLtM
N3tdxD/k8RYN2LUhKV436GFJ39KBKd+XWT++l+yDHqiFgk08Mi3iV8NE7caygvGklLUacIJ0iKtJ
bSZtQwCuubCxXUPmeGhNzVYgffegz4P5LYQ6UpbKyFQl7gd2hIVTlnnsI6eShyCfm38+UcWIuhgk
Q8MKdCiTDOg9a1q63HeBkuvAE15HQfnbfnzBRe88ddO/UGR2W6kFG0DUCX3v+rR514OnLTRuxDzh
9tqVPSeIFRIjAOfIUBRwQ6gW1eWMVd7rRTAC5Ly34r8XWiqpZJ2KCP6YtqlQ41TiBO57srzQOAmO
JanuNUjeKIETK4RVSgt2On9X3swAlWpDIggY3yyQ77an94iZ6lMXZ4c0Mpas8bzObyfCnSv7OxHX
jgMZxpBKV4PcmZo1kdwwWEI7TSXJw+xU4/cmtkRUZg3VM5i3W2t6E0baJ4ItOwxJ87LaUC0sw0bB
2U70dSD1nUeU20F+SkbKqRA0KFet5hdridfegwHLYdJ+otRjxOsR2Qi1kVia+7jbYCPaPX8XoTKe
vi6wcveXaQGfqzbMzDxqCZtoWI0ZXTBc9AMnO76LQCOoYIqSDUUeWZzI3ZNCcPE66PP/nhvK1P8/
VZkJRZulfxMTk0xGG3tNBxq4TwAoOHzOTVEa3qLnqj0oCVlcdokHfSCqFbN3H9WC5NAJOZmGf8Kh
ng29SHlRndL7rP8pAi+eVL11i22vXGZCFw8tq0S9d8mz94uRRjbbOL4y15bnrhr+7pNY6AGdd2KD
ZRp05xPh45nkEkqSomevkYfinu8WvPQnVhxcDav9yYc9IByg3ZxnoQWhnCgK7u8IgYefLQxXxwvr
n4auG3P60G7RIqmrnFG+aPTc9CHjGfylPfGjOlcVsLFtaFjG6qisEjUEQz6xaRoXcuDC3du415nz
F3/2v2j38prJocRdbUtC+EyljUufM2VXEJX2parXNmWf3aoKczBnXAOfXZtaw6RhT63HhR9QMPZk
cTtpi8hOuOLUvG7LB/kuAW0Eqf88S2sW/qTTz9Q0om3SHRUt78TIEWV+Dsj88OQ/++gOcsxMLb3v
CksScXTdt4EcuZSdZt0KjIkJtdxBimfb2bqPjtfaUoJdh6/QIkDtOuwhAVg19pDOMcpn+OAFYtLa
iyrAcjE2ft3f5hIQ/3twR3Tbc0uYeWEcFHWW9M9rX6smRku662vQTlZiHbpbXjs4Y2VjsV8jfxEY
TmnI/FlDw5wYKAQCmhlgTYiRdfcvbos4fUDUnYcQPTZMLjMuDRktcDS8LfnB88MfLyOsXgsKu/UB
sUkXfVfOcc9lYmi41g+RuDQhLUV7Yiwdrl5v7z7ztEy954mT5syPVrxvqWQUWBx2K6nZ/Aqlh8xR
klTXNHSxsPVK6Zr+rNZXdrCIdGo9ucCAGHLBO/uMEqjWb+S5g5++Zq0qoI8aMx7HyOBlezkw1PEg
AcbRSDFpojbRYhMY2mAzryoNTl6SV73x4WNxRvuk18nX4jGuoO64bLjtDRhWGSvaqqIVyg4SqyDz
eO8BoxIOLyPd776FFQPcE9oZVG7D1bQfrbCY99xBYA0Q6PuG1edlqnQdT4Lpu99cnblzEv+yQ+y2
SkoTSETf+Gq9OmeofYNQH3Ryv7aCdP3SENdL2IrAAmRP/j+M9sp+YVldlh6K04vFMShCg1BjhNZn
ABcYttj7rkNC8qwfoSrv4dcyZm2lW1Qq0VsJIK51okwpwF13mgN1YB7Cwh3WGaWlOh/Sa9+n59D5
pYPJaasse6maZsFWW2YEqXPU5ZnTfnXLw7d2yUL5XBIbe5e2mIyHeHXh2skmM7ZpcBtC3NbCEVol
UvdiMPEYlXs4J5Ry/btk5g+V8WC7F3KSkmtXbpt5JeJ0U4bzkCJq83A1DyU/l1+RWxN7kR2veXfM
L0WfnbtsEwvVyP2koe6rm7APMj0dqOb0ub3Ze25zkOce+8xZeYTCK8qafo889ouvPRlMS6xMYYXy
zRt3S2+6gzkCfSF2VFLoMMdoV1soAzERgTXpFQUKZTf0MuUs4Ryyggbdpaxjzq5YcI9FEsthBScA
/0lRXgVpUxEnjZ+hDkgSTfBfjZKTzzVqmNIaVQXMm1Ov/LUd6fHzXjUEaVoB0Yz5RK8lnxQsadld
+ojjS0SRrGY1Iu7CKKKKZdZ5FGzg3mqDpwRC1O/oKc1rwjkA8VD+1n1GIfxl6cnxWGpdoaNQnfdY
PMIk+SdchwZ+VBrJMs6pb5WQMPR+lDQejdI=
`pragma protect end_protected

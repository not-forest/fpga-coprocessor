`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
M1CpNfzXaqex/nZ8BfnsvjpJzITgW5BoZLmH5rskah50rUAqwcrzlY8mDAKJJ+B1
os9/NCSvqtoF3rRiGrJcPuIUdcEZGn1HQX0Um3OJDv2CQppmFeBetHcuomU/1KNT
lPGWI5XfK2dFWzqohFYOqsU3xSmQL/Kc8xy0z9MNfBM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 31392)
dPhS42AVd5qvzu12Af964n2XTkYFbnxHSc60BcrzrLD+AIVawIJzsmRH4YpWjT2t
UBD3gw3+3gHiIU+9bxBxxp0TObqhguk+4Os5xK7kAT0nIwMACD0kl55hRJQKvlJY
jFjBE5QCQbchWAxfGtQaBCC/talLasIwxdX9DpQRuZFj+WNW/tkwuXO90+d0p8jK
F1y06ih6x/Qa9Vr/MjsCEE6IP0BOt1LBbLGJtjHKvAHadMxCT2e0fuUcuS/9R28h
vZ+GY0mzouP84Fk/5t/fFBT989P+9mdbE1DTEK+WasbdAzGpZ6EDWgrq1OGVtSkL
5k5rTfPEElcVP/zAjSP0lVGS0h/eJ4jfeQL2Dww1m0LnpXzuGctlmfWoX49aTF4I
oEGhAj0ev+DW2fw3QSci6krbZ9sI9mtl/6JQeurKBO66xqiS8ALKGJ17HNubeRIC
pET74+poO6FXwVtba7IQBqiXXw5ux8+z5aKi1xn6o0DCGE5krboBxY7jHdW0Rzt/
nEuQ1X7MHWo4WhhvFHiAXaBZ5cERdSfvi4TLmDsj1HZcIIHcdULnT6TD1hrH67CC
mJ5C87dwrsjOxHPPxvkWBDn8RCBFSboO9gvtztRG3ozV00/mssbx3AHwAGuLOJkn
ThZEoe8A3c55BLrGTZ2Xlxn7fAAEGCWt0Z5rB7GaIW0MGOTPUZ6lTyFBF91Rtb+y
5lQ29a8LZ2xb/Pg+0k8t3iKTLq7bdUTui2CsKVjehX5nZwzF5HDJKK1UNo/B/AjP
U9q9jhHO4UL9qgHd8moePlWily5DIu0iyClFhfZA5n2NWE8TL5l7p741fMSjz724
9KeJz2aqjJpiFiYKja0UR8fXIsG5Pa0+gaK3s6dh/rQUX+zqQ7N3FC/T3Ky4m2zA
TSwMPPCV0wIpuHArDCHBIR6aQH3rmPa4nHoLgXq1L2nIUeXwakB4vQPib1JWqC8X
zWpPWNRDkqJA2AN7HdQpvc4/1XrvJI7LPS3bC39rwrZ8tc4bmyMErZAoDzChj1/J
sBHI3C/O/M6FGvcWQ7tvavmRA+RlEUMP1/KmNQQ0qZnS2GomU/bG54vJTytm4c2p
CDAGzz7se771knmwj/x40C/I9JcIP+YPEsdn4flSxi9b8P/oVTnRoVi63Cj7x8qn
9+EPIL74tx8A0J1TlAlcuQOKfN0fG0nH0JbNEH68sLOjB4iGhHxa+EsLrQWDRkep
Hh7pCbg6w6p8cg+Ut38B7JhSnaF1X/aK8quYqyfP05OLSuMFjeJpxSmVY2FrCSRf
2CetAiBwJwlccoFmrNI3ulwK8FdUocd2vLFXI9Ig8t01spEOkU+Sa5ImJwGpaEpx
ZzjBaGH94+Hf3EzrnHd4Q7KVgv47xPNdS6ueF/kO1KYCdpBPfQadULrzxmRbV+uc
zCX2h/jt8B+heIrHKb3vtDIUnS6SxY7fM0jixrV1D+N5ohSDECopYWIKfWb8x26x
h9NS1Ab+RtIJMqPP1LibvbqzsUlFrZxhQX+m8c1XY2yRV3Vef6Lz6Way8sTEp/MJ
7a1jcXF7JGlYF5MktIELQfDtn4k5xQh37YMqG/DFXLjHe8TzKA6vPxC1bY0nBVzM
n6ehccxMKD5ee7Ae5JVF6uhSdEULkwHknCkcxj7v6yCs1PLN4DtqhFAAHrmgpfF7
h8ufRwErH5C30D5cNvA4nI4j9aTU0iH6CaujadXOjzs8S/ADZ+XctAWToZdrfQjw
C9NRfQZTEXzgI9z0Op2CY6W3zX1brC0OaPPF3ZlBWr/Fa84ejJkXBIRYmaAcQ3+c
D7LkDwaKgTxejCsDsULYq8VwXcCzp0cvdqLmC3mnhzhdwvS1sabKQDWr/G1GqSE9
4zmW9gTNdLbojJjP3vc2Uo7vSwcGlbkf5P1eKhj24DHWk5sSdEHXPPoco+sWH/qk
KJcxQ9pHbBmAXmskaXTEL2l0TckCoX6IiwlA3ZzpeZ+wgwkuOjZPlCjqPMu6G7NX
swG2D7jlDcTZZpJ1UM1GpvRh850qTTBpx5Btn/HCwW0KPeISSXD1bSGryhMlYe7g
DwGG2sVzOpB7FcfQAhuJXca3sWS3fE7P0b+CMx6ILqvILihLNhEp4zltBA8utnOw
AtxNssXa2kVcuYkIDlf1aL+jgoyZT7zDGKYzpCg9SxcRYTi20Gm6d7+ALC8dyshU
JTtJBW4M7aeUVO95dX3A3bAKd5BEil+cEzmxQJLQA/e/oNLj74VZIWB2bXQ4agUC
vTWXwL17IwWcI1i5iwlUjSS1f+lcFzwq1HfILiEGZ6K8iRMJfDRAMlnB/A4A3084
Tgoj2YnSjR+c1sQ2xkuQeY4udR1EyHb1AoTPh0G7kx6J2PngnKK1/fU5N2KnX+xA
VuQYq/7FIE5eLEzNmFSkMEMbcONDkuzwDGnJR4P1bCDRXqDyDYBIbptKOtSv75WS
3Sai0wd9g3Hhu7+42gp/sm1rogHwS0UTZ6IbHcp+2ottK0LgrrqG0Ib9GtpgHyxz
DVnyKM8qPMb4cZZJNK+R9Jk/GJt6aoBKsNmzX7b9GXYZrwgAww3aeMFmnf6Sfj1g
yLpmxH9d7RDuE1UVq6DBY2qJZjdpSIPoqGO9AkCWd2BUmQpig8moQxltTMk6r7b4
P0Jh8ZvmYJmis07NWv9eK3aQoplPExVjdzUZ5yMs2qmTFNCGJA18RuWGSBspxFaN
rAk0IW72ONXNZHxY4AOmuDsAWnJJ3HgakcQVrHP5SO60fs7VKrqrf3Knsq3GhbJA
lze7eyhFaRH1IFSXfnCS3OeOko2FeeAcPdCbF7Usmr5/I0ZPv/DZ1jlDaEP2Xo2c
a0NXZ8AppKjqplhLfprhmV5A+PuL0GmpCbkG5elcWFbzEHxmo7+VChAZmvw4Orh7
yBboH6sqJqFXl11qV/2vWEEk2RBHel7AJHr66tb8zsVx8wbxboWvDjDP/iMmCobI
pICeVZNyo0d6AVEDjlLxGt8IeDpj4bZU5/89/xt/XvjL3JU4Ynbs+DHtLipOvlE/
YDrHA8ZN9d0Mb9GToM/tbOzgEB6Pthb/A6Gtzk0BQWD+wMONm4+dmC4AmILEETbO
MXMwK6dbLhKatRIlCPrqidp2E6j9hrkVLmSvbmdeJ6oEEEg2WRgD51l9iKWf6lCy
chZ+0w+03OnDAnr4YFYRmeovL5PbfOKF3QAGNYzhlfSXPgVdruTuhqNg9j1sHrwe
9v0e12I+YgqKeOfp5959tBSnGn7TilgQ2lY4ddizl4exym39TGTqEqIl7B0XX1jo
lZqdYuSBfTuGtWEfPX5y7RkSyrXw/P1gg2rKn5nfqmcsiCVy5DjdToETB9LEvSVU
PBNMJ/zn5ejeym1Y9v4p92+JMSOHuxMMALoANFfY9vcMAy64J4/TW3/eP+LxzlcP
GhorG06YiLsfkoWJP40hqDZK/Z+pUagCZZ3RzMhdovjmpaz5rYL+zmOmyFfHqNx0
hkXLnuiSN5c8j99WqzyoBH3MZe4XTaxQZh+PeoPeYhBjva5m+KfTPyP8dYOgH441
K1pWxA5GbxhGLoc+VyQ6iMB7nR10aRn50EGwMuGemt+1HwFvfXrzASo1mc8XwWDd
dlyvarBMrQp5kqO9cAJNtesWHgXN+qS/N1vLyIjgx2lSAku3hVu630s5BEsQvxYk
VAgx7tMRtkYVYB7/ixhWGexEA60eZobjgORmXtKAU8weT9Q1OqRUloLii+jQJHjI
T9WCl6odH+MD37iI0A+pGVTNNQhCC8/HK+7XO0N4s3QfMZWwg0/8S2BYaDp7L4cx
3NMBxGKhJAxzusJDQF4D3Ku+EjooK4ne1QMXEY22uapV9gFS7U76NAwi2ejwJliw
YjCOrvmgafWmL/i2bwh5LLzAFiLJVAqhB0SzRvGEtdC+9T05Ii9OmSHzcXVSRjh8
+pfr2LQ+tKGsy6QR4QqX2vJyosv0CMfAt1DGrn7Xk7AuskaXQarjzrK0A/Ed29ji
r8+gfLoc7xXxQirRkdpkV2a8PnbJKxjbtWxpSUUUpTnewUv5ufwhfzXXxZoFIpmH
CQbbNPm/fanGqgr+hUcb6dI7h3DRX/66szlPgVzDiheU6r6opgStTUTXxgvJrcQs
WHjJOA+Dj8q3TSKx5JbZgkDkta0XV+44V8DZw8lLxpJHC3RfFK4QD3oFaQKpXQAO
Yn/TUP3wfe69Ez5H4mjrBhYdNTFVYgJO4G/uwh6Kgpe8kRZFohgQNDNUGzkSiRsw
5pWCPL3XmSxfVMWrL2KxN1FrQaeIU9R0S5Qkw79QRXG416AQvi0xrcOEglRkB1er
JwL/HW/wIF7vQ6Qs4+Zc7chYOADghKzwiIXP9RldXacE6NzoMoKN+KkUn+VtHrxB
7Kmb/2fcq9jSQyBzVMTLn4LFkl3ppu3NxH+UDQ+6JyoXCltu3NMBnWyUKVI043kJ
q3MacppK4CqrUx87t+gAs0RIkTBY955fMWnkxjrhlNIjjYSYLuUfepV9EiEBXq08
9RLO2cT1r89iZ7kF2+TeDmce/Hd+iZByY2Mhy4Cs+70yqnANPWLQdgDuFDERLHc1
4Z4WIgYb2EYvsukQEbw0bqKMWHaXN4nZCN70vI/9qXRKEGrJCljZ+vWwh+n/af2Z
NKY71qHCkWbtEIgVA0IcrmU+5Zsmhq641EznXnISDXoGKZOIMkKAYe2r3dXYbQ6m
E/MxbaCMzbyHvy7PGDMZbQXsCNs7EIBN9O8atFQlD+FDJriTd2Z0dyPxhQKtiSXg
z1Pi4GlN40+4DHmlmr9UvCdXRZqcr2kMT9yujYX1BV5Krq4R0vsQKhIN2kQ28ohY
jPKGj/lKjNaDdu0fIECHtT1OAMCnK4sCTfW2rTK8TaIf5CUUPBOnHT6y/X9sGMfs
8fqEi0ayMQlVLOAeUsU7L32BOPDGRyZc09WagmdKMBP8B6GiCVXhq/FUSn6uj5Yi
mLVEnJGPQlbLVU/xPmfmhZTa9nNIxX0FlMDhtPvjELG/iSmemSC4RATRLvxcyuJ8
cltOiwJeidcumpfBseFg4Sc33HcMUP5S3PYcaew/5qIdoYEp1rcbYwzX5Df4kNue
sQW7bMoFc3+M7G9FW1+G1LPMXDyU1wB9lhx4DaT//Tk+E48MdiRGBT+umrcZcYTA
sYqFcHf6AyYPiLtaMhUZgE1meM2O8SE9pZQecvm2jih9/35HM0rOEzhjVZ1QtO97
i/J6betFHc2wBUIjxeOp41Vf/pZTEfvtqYDQ0cd7UoN+jVNpLVgjJnUmiXiAlr3p
ANcVJC1spaULPs+lzrs5In2KoTks7s0D1AtKoPx8FkD56+YHJltxDKVBcshVn9N7
Dz5JVchNAod6YBKUNFNyVZ0I34xhhBzgm+HWkprr5HTNJxkcE0Sy2zroBubS3AjX
9k8bK0nbnSLOPP3we4/yFHsGdTTACK31HzdqatRdTTg7PAALbC3rY7FslmGcHMRJ
m0D6eQLFXlqGEKtp+F81U1JzNDCzIhfO2ANglMeJ/xYUHDWS0SAxIjjlGdTZyHKz
S/eahoYw37ABwpQUsH5cGrj6CF8wzYIXhxBjSCXgsJKv27ljwyZ5hpi/AryIB5ru
1Npw6SKKJoKpsNrGUJyDoRHSlTIAEIlA4DpMbHcD9Sulup/1BCm+jg2QK12ajIGI
zBLhCZK9EUe32LHSyNkRpoetpJlT59hnMghj1J1+WA5fg7BRx5sTxOQehGavkaTY
DydXOy2SKQRV0/yiidlIWMLRHnHcAOF0HMF8KfxB/XqQsgbfO5o9QhoiPviP9acG
M8490Y5v8S8CewT8SbHs5CaNW6aviM7kVCZbJvfUkC4wnimVBciWHYXkFRh4uVSw
Q7ZUZhS5JlR0F9udUyvVRqVhIpoX46T6z+AwJ6T//cvl8dDiooZOxt5cMgT7xX3x
gJdy0oyDpLYlZBcgOoKEoTa19SaPDQhKaF9sYwTELcMtE7RQysszFo+brgwGmGHs
5bvW0WP8tZYVg1QJAzbZUNJtT2Eyc5dk/bdbMoOcvydwG1G0IQ1eMsvtFIcL4GKw
cK7aUfrUHyGzvmMpGx+TQeYVf6hCGcbN+uxTHY7y9jHy49s9Z51jFAoNTFhA82ME
snftcpccoF+k42cIQYxYnUtLozB5ylH2t8aCuoltdoaYz2YdBlr0ceIErxzZLkI/
gwUmd5cqcgfDiPpQeBQLRJZHHzxIZnp+jbIA+RMJgim4sZ87wUWozKIpwjWO9UXr
F3aYcF88dwJinsFTlornMafF2W5r5EP8OcCPtAOIWpbY/6ZI/xzXh6Y/roCy/FpQ
BIdExl6RxHJ9Ws4v840kIAhqJMTQCIEhXUqojlB5SUuWJxdPtUeeCxFvwBMnNZig
viGnbTHLPWoFYtNId3erQGLHFV945YVhdFXpV42uHPWnycJuNGWqL1Apn8Vttye/
gjmH+/ACttt1pYlRVwilWtZfcKiiEi234YcnpD+n9BDBwBf0YQ9n51a/ntF5Ef3W
vS/wCcvdtkLjzBLPVC/UOy8eQ8L7cJHjI8JOxTKkEYCAyIN6Yc0zJFDmWAPwYt/H
KJdGj5bgX4e+pgmx0ON2nDre5JMh8RZ5Wshjk+33ozJlv6bGB3jISqN7mxkP27dN
k6E7DswnufRg956jBIhZnJZiKg37LpW/5lHeC6BxTxHQ7j3Pvz1nDVKMnY28pLe0
FEEVcldcZbc6xmZ9H1Pmte9MqgxivYlED3XLMti8Y98WhpQqGVNHZKb7F0XJ3mbJ
wiHg8NY8xWtOWDGMZJCt7mV4+xxrRaDV22NfMU8y10ej7LgaVE0F/0a0l9UrPWAy
lolK01HDaUgCBdPkDTTNDm+EG3cOnG+enSxtnxWqhuPXL2i/Ox0jTHkGgVotvJ8A
8RrcfHMaaAoty0W01RGhpcjgyNErZK6iNbG6ls1+f+i+YOn5Wx3A1iRytNLlDtYt
7D1S1Y79EsxZvphIlqMxjrkDtHGihpZNB1P9o8HkBoc1K/huJQim0ury5Tn2Tyk/
cS1ir6d+SXhAAM2I5doL+q4Pcfa6umqN4uAzn9QJ6qDQacqXUctjU8SoKLRGVwD6
YkcJEFPjAF0Vor6I1e1EwVFpS1hdswXo/4oOgEWNsjLRb2NSh1nm/+kJmT+BvCdW
RST1DBIM4r1iv/RopZ0gPlzK3XGEv6ZfyfsX1ISjg279W2UoH7gea7nJnKKGJWoC
VxR2Ixce8qyyucUG5/bAQUmTMWcLaKCwyTt+6yHBVdGk3JxtXqKP7NotEVkKSJ1O
6+1h06z06ftY0/fM9q7VP4rdcBl9LbmPSSqX7JVj82WPXmsQAZOhQMBrVycbd24J
GXAvcqVssrXoeTZF889gtgTAeD3bgOk6Gz6CcL6vm0GexIWIgL/prZ1DXlFogGgH
b8J6FJoVks1bAW0CYajcHAFxy4iaUHQSNJDFmWTtz7mgMJRYpws537CxVD5FOlH8
eQTjkzmdwnyUEV+RfV8gTYSnlh23/akPuavXEvlduY9iWomhPihWu11CZLx3PX0k
J/+cL3e8/oeVJp4NQHSz6kdm4dmnOZ8iZkIUytSWV1A9tez+K2coy5twtWyxNeCV
656IL/84whqlZO8j7kmGej0YgtXRV8qVAjGjfv6biM1H6sr3wMyLOV11ea0PYRYY
EOPsPABS+cyN65JDJa7ojiathhfU5W89L8KokAN9tjuwHjP4dCK4lj93GUHDxcU3
GkY16SSmhnnIKGmkXISMpKXt3Jy/QEGlT27ikppN1ajbdoDHGGO0Nyzn0KU9Cihs
nCEOSNJgSeoFxS+RvUSGYxy/XldbXlOZkJsC9oKf9gHQJzmJlAK5mCzt51EMTven
4hByN+hAca68lz/saCFbJwSZli6BAM2z+HykraCXMXHX3DirbhzIyuty8p7owFee
WB4VENasX4Ye15G5O7P/MFhVcUnKLd1jH85syM8sxTfsaTKdRQNaQNmi5jctgPCb
Hgh/O8DrjVUjz4d2N2V1dCNk+gtSsdjyKJypqEvbAHrzEK/P1+isPx7vk3Vxy1S4
gQMseibploEradsW1rtfLGFgRqjlyzRN7jbCrguvMg4ML7M1Ae/ZIbFDdSo1Ub5d
Hau7QoIfj6YU61TOk0aD+nJeT/D/vnufNJm9sXgpJc+f8qNfxx8izbPR/NnimciT
oHpEx2L0ELBdSfSgoElwT1Ll21jigOYuFBYwwKxU4RceHH7/JOmw27EPOa7vJ6zC
LjOKhPyOcRACfLkCXS3pf6j5gRT4eKq1DIJuAoNN0t5XPgXjhTDqFBrZ7vq31FuO
7iGQCs96fXakgnYXCXtMSpD2uRu6dASCZPK+twS639Viug4hhFmtyQG3Hbs8Fill
UKlA79Kqsz9D3s9EW9OsrwSF1hlJn1+IK01tuzkCOaaYOFfOy+pQ0o4ykMf72kFR
DRyD20dhXtkqER9VoZQw188T170kck1IoRrLnK3WEQ8iWbs7lSy8bdRHq+ya0KvC
kxa4GljhENwh9jWKdhbvaEAgj/kshEdvDf9lnKFPTbqgqnvIHXCPBOuwZLgtsQay
v1AupamCa+esJjZJqYk4M3536gIHxXrGmzXnGzQzsQJhWx+H6GhSXcrGg50JknZL
TBZ22JK/JOTeafwqUP/vRT0V4/2+bFUAVepXVTVzyjXp86b37Z2Pd7PyPUQmpCCf
KnGznab/RarjgvJL097Uw2KFhq/QSuW2AE5YZfT7XLVUemXc4Dt9k3v8T4g7WtiP
iwcPZ0SZ+YP3PEB8lskS3RDDQBjryqPeZRld3hOXyzjPjrnO4DI4vmbZCDg7zj2c
TdISB7dXy6ZqaIWZw24Tll+rMaTaNpHTiQM6+X6p17RqpqOTdavvWltCbgYNRXe4
rWgfL0nfiNC+kDtrIu2pIoAPM+ME3hfj/RHjaNO/m1c5xV3wZiuJ0aYhwxNVCBOD
r2w6pr4CS4Uv6BlSTG9N5mCJZWGv7U4Z8eG76Ht6kS1IbtRXs5PNcFJp3afLOTn8
t4l5rQ6QEdUGWgIfA9lW3TSLb7aulZ2rE+gz/RTCU13dxysDxxp3dB7X2z7VEuGU
ZRG611gVtqc/fT6Bvt1T6Z22JBi422QwaKCkItGDRy8HF5yUg1Pgfjwyh2x5m6Lt
lMxFUUdGNO12Q1VDU1cLtKgesrkhDJF2hpxs3FEHTGCRNyVugxsFWHbA5ulS9zf1
XQl57lwGD8u/Vb4Bkpa39pcqlRZOkjXN2anIZqcX39xFBeQmKeIvEfpoq134brOw
A3dPTTJ0TbfQiMuh0kG+WSOJbra2yghq+JQ9nDR5XemYJU6i9OUCq02mJZvq25wI
rqjSDVpOqcrdGpC8aSyyvod5e8tpYfjHoijcqX+VatpJx5oXsXsgrK6iL344XOOL
xXjVjDULnpv9+m2dgP4to50Uy41zZ4k4Sx6/TygdKCY06EVUvY0CIwMw15lk6VsM
fV4Y9Bwvng9uEkmTr81dlhDn7kZQT+ZKvQwymVj6vA8W3tpJGmHrxUkrOjeoD/TF
k8+DcQE6IB+aQhVLRuTG8URYsHJo8DCiaomHubLD/4dKZZ+/5wvHX5T4DL9bA18X
+trJYxwQAb7sBYEqFXaDm+3LsCSEp/WPjKPewfOPgZdqtCIHWhGVNqsdWxny5AG2
ivhI84rxbaK1aDAUpwKVNC7nmyQNo6yZuhOOU1URCHSPwJ/4F6nMjR8mU75gXkmZ
V51QIHVXKjmLhvuQjl0hMzR4OBnKEjBf8sOIIMPpV/Y5cTs9ZKeR7kMkfAu9g0Gd
8e/sHZ6+wyNYmxGyVpS4WEoFAwH0lPrtqpjxCEfzerkYlTHEuJrDyqEiNqZ3PEje
8V3sgPg/xi3mCuWKuxLcT/n9FLUZd02tISndpOXIpM6E1n1x5FDwqbaOlFe84OqW
EobrUZ/Px/2Y8SmaNLENQjK66sNFz6tV/eoYghPkQtpW2CHYgLqolL9hN8BHyLs2
SAkz3F+g7+ry6Dnwnl3eK5IyOVuzQZVUuDdFq8YtOb9OXdZunSakvsS940wv4Oes
0ZdXplO6GOTkI2TEcwC1yu63/hyJ0Ci42QxDGTD8PhYNdKGMj/XSeQfRFFxVUFpe
vWTu1LCnla3YI4gvTsD+WTF2DU/qTwMG3gZGEhbK9N+fE8Tnpknucq04BDac2mIr
+V7H61Dd0++AtUCCB7IeYXxGkjJ4d6rGGM1AW2ovGSWMVwI5uekbRUDfdv2ZmT1r
K1YgueaqNm8nFMfIkNBSPyYOsH8+tVdJyaUPDf5d7HNMKs0sslduCmsrWOPb63st
HMsrm9tqUdq60GqOIpcPCDX+vFImfxzjSLLmTes15KhTSOW3gJ1j3Zl9KmDfbLb8
oOVi9GXkdUP6QRa7VDBiRjMeLmP/4yUwP5DXUykleJcrLNIA1wOZT3QlDE77ctVo
plJ7gePhyuM+7mkV9XH0hJz4T3kUBvbIWwcebn0IIDQ23dyT1iVhzaRciDCHYNe/
elEHVPTZ0GrGJiVRXt9WW1qbgaWx57PaubUjy44MqsyxdvFFSUYB2pjtOvlxEmCU
zefwgx/oP0E/6xf/NQqbthk/0td9qXNfImJSy43J5eqqkHjPVJ4EJi1jN0YYNInO
jfuPLs5SP7/A0XVsqPDl9YgGBV/7QcjBwRDAgQg2HEfWUXf443O28o5vxGCv/RuP
enAbGhiF4fL5tlqtEjDYqKM/Rcbw795yRKu9MyVDIJnGd+KPwsjZoN5p2d2I+jvs
7Ec+SPxH3nzLVrste/vf424v3bcFFn8jFrGbmlssR6cnKNMPLn1x3Jm/BnTK43gD
OWMuqtupqvvAZ+iTJnxT/xfC2EBO0201e6ZwDVFVYczJGyhzGiYM15Tnvd3/yIcD
xypcoPfYAGP55OC3Mmvqq85k8/uhtw+LxedDxfHGZmAhnocQNHSd9ck7xzQszpQ6
k1wTi2cpDWeSJRIMjmh1r+a9I8cuRF7IoS038KSpChQGo+qyyTYssocDIxuC99iS
I2r/iJ5IogN2VIb+/owfwOtZmhgjRoXYWEHb0yzqs7N+dXbPOo6aGDyDtxJQgv7J
+DJZf65O970VGg4SKoTxApPgRg6htPCgup1s6yjM/BKtjHmPMSrhzjq01JJ1YGOl
HWrz4XBh5cvRlH6G3dJd3puHhT4FccT3qq7CrrZDPVfIqEbxGdwKakFkHOUB8Vco
9oPbn3pzetNx8KaPszRKIM54sagH1r4FAijvjgibSxuuSDdA5WRbYBfcV9mFzMR4
GNAdhHLcHn9CCt7zEGEIylGM/fGNXcYzt8+hDSk0Qrb/SNGl0kPhDTnXAsWrtlYw
ltgsvVclZeW0o/kbMfP5cIc1P9/PsXNVAzwzXtqHovme955g6nSaGVSxz7K5fCxa
pIXCHRiYQx422o29/GdyurVjN/EbqJLiWZH5m34Bh2EiBSwr25BQfCZTT0h5dD3w
IeCWRXAQrWB5UbhTqP5/iBbDd3kD8k7Y0cdyhHh215dAWgIyqPIAcdnrzPlwq/YX
9horYWSMKLzKzEkHQcWSD75jmZb4WDVTbfK85Ha7/GDyT0vWmqSG25LPoUUwKmY1
E522AlYMHIepm8wTpE3h0KMZjz0GHGCnh5U0E8zPdjQtSLfl6rdQHuwOI1OpoLB0
AVMMpgw9a3pKjeLrGIbKdUz6VGIGhkg0sKQNVGVOVaJdN3tmZ5jv/mNuOKPEBeF9
9CPnPnxFLpTnTVfK2QtRJjCZqze5PahI7tsX0MTdDt3W5vjZ5svwM940pYgzsf4m
xU9M682Sr+Wa14SGo9KIIm/gYbSOrpiqOOl6CRoQsVb7c1WW1kl7cpiy/UP0KWM1
58aHJpPVl31Sy0Zr8YYnRtdP+h1IRDqxRNcPClY7pP1iHTOiyvZz/ffc+z+/xnVL
ql+a6g4UQ573sBS0M/pZzJtOEeqjjcS09Avin31T5+VxDLZs83raOt7wLiXcZYI4
KMYsgVI8MZetyFDd7a6Eh6csrrezkp/eM7H5cBKfj2NwwD5h3/E75GWaMboZ12AP
xocub4blX2c+FG7AaH3jD2igEVx3TIt5LMy41a52hebJJmhoxTP+www/HHLSAjmy
me+DVSIP3Q6OqfOiAdyCK1sxSTvG141odPNPJPipqVewAXHfa4eBbuHA5m3VaQub
8qKhryh4VbjXnbcN60wdLLQfdZrEp2wETh1TaP5SHmurNZAD7TwPLHkP10536NQW
FvqrX77zOvL5vKK+HZQpSUFPifnv4aEar3o9YYreUTn9TtIfwKRX10xelLPxmZ87
yQ6N262iaxAdjPw+T+G31pdTMIqYJJeB961Yljxfqi54LKOEw8Awb97qe/OEYXHu
i6yTpNOHQ3JGm5q4bLzaVcA66+SqHUUM16WgrM8S/XUOazhbtTO9br79setxDu27
CrsiZBBOgxKV+DWLEuq8ZeF53EsOXtgr1Z3MeLUKwg3LepVIZ9bBoQTWYVDQR1cz
93Il480Wr7oWLQF/lNVzUgsOmUn7A0ao4pCia3SQrub5AlD2JsDo5n4aVvBOO98k
n9ykIa4jhj2h+gQTaHixBgIW8YIppkk7BFyFdPfAi5TzMh8BaAU1/Zf+rpSKJUL0
DCHCHpa4U+zpN0ux90rCXKOnBg/VwtabDQDbjgDTaepUU4AgAtQTC8cKjjSGnctz
8QY+qMvWKsygfH7m9RKmwSXbKZX19NPbgZUz5YvCrwcPFRPd0ilpeHfNe3vIgZFF
XnacQ8gY1qTC7wvsSNP/+9nlM8Ag2iC5sn6zRg0YeOZhItbWMorm9f4nUW+hcGhA
X6NQylJyyX03zxM3K6LiARr3p4D32kWRelKLbCeXESlEXlrBuTb5VIx2JuCD1Jwe
kbRQqPOXH6VTCTBGhGhWfMmz4pAGI5BYK6fsaFfAfi93sVnM+JS6EFOSvEwOi4w5
dpgk1sE4BJggvQzGfvkj8R6tIoQVSIBHr7ZlEJfYIE6sdZNhDdj75xm0yYdWRz4f
hwSIbtSGWL1OLwUAyb7Jg1ZkN4NXGNhxQZJXynk+o8sw4Kq3HlVz7SMwG8m+HFCf
0y7Xoq7EhIfW7BogJeOIY8T+PkAFJkFchqS1hGQ032sKKqXiBsToYvulIRnKeP79
z+nqECqwNYXpinJx8AvALwPVlFmZLYe1D7PLdGUh7evSby+vBf4zJv1MsXKXxi0e
3VQYNUUuYjacDtzwTuAKeIJQhPbn5qULX7tj2NkxpNOLnL4LDK/H68k5b/lL81c+
3f5gX5jWwvk6sSF0h/IzX831PRBrzcDhRQHlD1GdnTJudV8CeIcbm3W36I1we+Wk
9gEn/JTyIpgH2i8uQN46nB/Nm5fyeRg1WgUyT3tBfgLWiV9fuAJO9/3dW4YCqhNa
kNI6UwMdiJXcexSSvPLY5LiwPXoh9ti531aCJ8n0SAdWeeH3zGZidi77oMtned0A
4apC9GWjhVbkGv24p9LHLTDhv9uGHhay2eB42+TBXYp/0LPpBvb6GVVM0NFcFDaq
ZQBB51UdqmCgQ54o2xOBLxxKpN1tAwPebWsPu8ZgYuyXrTAC1sgN9pq5gWHF//xM
yrJ4bOZ1TUe+ajXBqkWb2ozuV+nHBpj8xV3h2D6jipG/sSmE7VbZAYQpHrX/nfZl
YoSwZMDqqkbcZk3fz/jUrBRIcknOqkwftx6p3coffyIRNLZj6TzYvyY4f3phImt4
KiFAE/nyGdVRMd7I+xdWUH43Ui1iTih5bo2EK+XJGu9lKk406Mcm1NRBq14fpB5y
ov0gd/QWZquOy4Rg9LV1bMwAwfzYw6MQ6YCFtxvdtlOevEwlgxNdBNRS133QFVxm
naQsPvIf27BRH1efL/xmQY9L3FH0uDW9IfYuTWytvDbA48L5BVRKZ/EWD64TZvWb
641k23IUxdmbUQCc4TB8dUQii+wzBSv10QLXjIYXEJucsCEhtTbAKA6pYGtU7L7b
CO2jUTN+XjOQXYDLn4LcVaKYO/u9h+y98aFYgNdFoCKgMbJ7xQhCo5rjDety+d0v
u6pVIgswqgx/aAlXq3GNoYnJLMb6jfZqkIaZB546fVa4QcvFur/tTypa5desQpPC
42Z24b+r/qHR9w98BfBr1FHNmOD3pHqZSf5wI83OhU9VdxAZ1oJQCISiAYQ+qzF8
fNOuMempnYLJRidSD3butjmtUAE93XHuPeHIelmdxJ5w38LFE2Kb4BtERz6by7by
rO/97WFV3+yGmd6jXisUHb/VsOXFZ5jsssKyQQb/QwCvjz6+BatHK+yTr5wG218g
11GvLWaw0OPs0sMT7cxg7SUJWmlGm3gTKvcAx+/wSq6sUidF9SPFeE64BPy5gVcW
QZn5dB3KWrz+G+E4+qk7ZAyiN2ZuNlSFAbu0IcbY/pFZQ/hGZu3XsJs5IwykiZh6
TFihhKdnWCD+B4+0Wvgj+0X4pMHqI4U3tSiMYcQ8Steox25lqAeLIfNT+6NzQ0WI
Yi/r1Nnoehl/D0K8P9bh8E+QwUgCe6i6NN4Rl2WJFbjIYfCa+EhxGPnCT70SO4AQ
wjOGu1KFHvr0Znvuurkt2Lc+6V4imcv75OCK4j5dhOObmfJynkn2HpRNQAajrN7D
3q3KUPJAfqBPo/heQqNFMfJYD0Px8ZeR1j9hPVBb9jc66N6e5I5TqXJoQIkECpe0
IwuG4AxXeNb4YmKLM2N+Ost79g4c9WHkksq0Z21nz3UD942VAeW6lmbTPWM1jnr1
wpRTgxNQanB1GaxKOgEOVRiQKtdGqfpAkCdqk5sW+l/XG9HXR5uX/gzTue7JvGEI
70cXMWZ4CHIAAXBnn4pSzO/fxtGztWaxZn3BLUyWC3N9K0Z8ZfOlrAh6ZLlbdR1t
ENAcXIQxpgfvX7D+AojiFukB9XjRiNi/609rNHNdkP7ruRyfrzWqakYGsOzR81/h
h0hg/fQk4qaq1cu9wOGYlzhUS+rvHISbh/qWKeP7/dK52b1M0Xl0+SF5nenYXER9
NcYPuIqznDq4Ez9iMGcTZw5rSM5lE2RAazjNvmD7hA6UWMTOcAbrbMvHRSUKW8IK
6UqRa8F4awGOur1EnU5N7t/LiHOavnV5NveksPz3PVoOlt3aT4TGcuh4eTNKhbpt
GJoshWrpY59tOOolCeNtHMNw6ptV8Ac/zGLs1m4spqEd2C2BinZnDxCQtOtf6oMy
cPCQSVgtbvwwoLBLS4E2Ta34JlmkbceAPxZpDcm4oTvfVS33aH7AIgrbgsqzp6NO
mAzDZUs9ssGW4InH1U5hlz/IeKwUgU6132IjdV3tELAdjFmDySEI+PdfckQ6ln+s
WKQl2EVinlDMQs/pAwrYePNKG5B9Fe+8dmdCQYWAlMjrz76+TyQ/rgQ37mJbtvvk
/KPdYVzz4Wg99loFPMLdYEupv18/Tm+YDm1prCh7LMvDSKOi2BLyGF4MDZaAReHB
2bT3+/pG+NsayW+BSP+TY3/tRznw9b2TlchhbrdN4vGF0j9/pcJsmIv8tf10R1r9
lQHBx6uIF16Z1xq0EULJputHzXI0HmH0k2jJC8UFbs207fzgN7sOLQZ3Ow62wPfH
SGnBpHZx/B+J5V3RQq4kWEP4ZDELYF1j3CR2uTBTAu4ndIhM+HVp4xh7biAKYmgP
eaEP9FbANcYQC7BV+2TStxxXMdRqRNgUA1RPEl2KyZsTJhYlnd8UqeE1FjcFJe6T
vVdOFwbhjSWikOgMPGkkIqzCLdY5qAkeN2rzsEpSM1pfEnjK4whSZLfwC2YrMt6D
Uy7RwUH4yjf2PmgAjeDBWNUq/9EsKF+uSPwP0N3ds2rt6Wxe8sFLi/1Dgdstcp24
IHEvIdNFVIV1fh9FVDfmXKCw8b5iJs1SIC1XheYhJdY3lahlbZuGw+zFbV/uYakz
oBAhGAsTAPh9M9CmFqhJappwhbR06PcDkVq86akC7wAMybjPW1IOVmHbuFbKfDzk
GYmFiArgt4P0/WbSTLil3OenDFO96sVSkRyIFUX08NmtykLZTAdEwcGJpbq9lpLI
NH84G/Fu2SyrDQrJuoUP9TSHRS7Aycw7zR51wSQAEVUNhpzHQvBfbeh4DGcnVXQ7
a84V+iBfWQRRY9d2pC0Vu0HnIx9tyN+U+TS+VXr9i4W5SWp3pCJcIpPQmFTRNG2R
Lv3fqTBbh9crTYUir2vKyoaKyNmUMnW2zlDUvPQ00kNzFvs1kbRjyn3Y+YVoZ08D
or9VeHDNPiKHOh4AWufeBCOvfRl9eAodteeN+itwVC03K84aMPUc7JhBl+UXzs6h
g8Jw0aWnCSE9Q8a8gJGBcCQuWaFJVJkEzeue1Pzwe0pMWuT2e0Eb5h5bjtovIROj
zJJ2sjuNoIj3ChWCd1+wPzOTM8flexFYBPoev5UDqYFmFkrGW9yL0PgBFEu3+VHQ
ZwzXzglExNuG3rMiTbPUaeUwYQKRJeJFtB9hf2ibdmOCv9amjAvWmdCQxDQYg4/e
GgjkxB0tha3dVD+6j8L5LxrrIJ9TfsFbR02f2r3JARMmhKupAaQplWXrxRecCCdi
tM5Os06DQTgXos8fnImYZR+JJy8nKOLUxpk/nNof1NSBieV+vJmZSZtXUOnOv8+T
QOs3sCbKyzZKR19LFFs5NkqlcV/8PRxRLYZ+ByO7a2yfb+QDeanPZBUUMh6Zhlqk
PJspTb4aqEq9y6yZpVWpiWrL0tiFl7dvouDdrRHqV1NXlGTMWHeuyzjkW+93BN/P
CgnNwCYTZf+8cCklYwspixznUGx4Ygzz8EEFfHwXqWgPH0DrHvZUqAnxUphxl4Qv
IPyiVY0dZfA2QMyDKfkfqD4yDvhD469Cv55EdQtto3gpf0RV2zi9SysTsIWhGZGy
gjgH3XiKMZaRqyjzlYF1XW8+6lCOwygtVEFNrOI4QRa8eAqBmX2zCLsnDfpnVDCU
LG55G81pyrS7we2lQ2vbFxj3OXYFXO+6D1UHzuE6qwjRRoZSj/97ZTQV9775ApdL
O8MS/Fn1RA7kpz6JJSiVQO2GINbLa19PQeFZIsJbHlsQ+/boLTI3S852VnFADAOy
vfaWMxkx3+1L6s2ZGD9/mHUAVKwQzK2AOa54k7rAMXzYUbc9MX8gftZzf4ZUZwVh
zOkIxsugAWjZnga8C89DlWfj7N1MLfXkH0dWFCPY1d38DTfhWAOyrjKFUQofTyI2
Ru9HXIm04t3IdCt2X3wQiENoszxbfDcLnRuVgLD1agbGIVOeYLAyAlaIWR4YgpCt
fZ00UwF9mLPuMjBNpJs4r5i4cUc9gvRncIgULen9aCfeKj7Q6QvLEw0bdmNN4moI
cld301On7jqdrmtCJcKGpUrjA902IQ6GJWCegEARzje1YMld2mfIMxomob8ZWLUq
c1+9ynIYb+MDN/LkAL2uge4tA17bc6R5sv1aID6gc4h5gnRjO9I+1/zh9Ir8WxSj
UufZjsvNoW+ErHPvXlocNwM7RN9jc0hfbDJaermeQysfNLSEjlLLMhrxZZ5S4ZO0
OEyTdLWf2EWGjgUn/akHYkqM2V0/Mmj+2B7zDlw1qXwidsNfhRhw5J4a7MmX2HvF
vaWewmbPSXplVPrkJQ14hfXAM5V6PB4EASAz+pFu4SF0tIL3oNYSphvtRTzo4yjN
8iv4rDBrjOEaX/M9RtzpBbmDB6ub6kTc/vJuTVyFzSECpuo/ICDxF212XIPlqp37
P2wfSC8dBzdl4VCLdVVRch/Hlv/sbfOAazcMyUhxKqm67H6O9LUSQBqNFy1DypUV
4kdFMgL0J0pF7BXvI0yj0/MWfWmIYIE11465siUKU6O+GAsaiyqlBi5jyha3zG3S
eF5ohRS+qymkG0GmH1VdgJbLRagmqF4xsFBepPpnbgyDL6lsCwKEYHDdooq2Ml81
KaoJTYsWsLZGPW+7RenuF3ffAfkdtOZe8RISAV5x57r7dv8i5LnBN20ftkH/iIcZ
cgfbnP38qJ4KXMRXCSP6Cf3xisxfrB9I9st0SileMdcahVBsTKba0N4N+snJAjwT
N1B9GvXeNW9XneuTmn19axCG6jtquimdmgx3lErdhWmNdkUjf+SOiIasjTPoDbso
wePBbZUf8RoM904cf+cJs8ZRIuodsWNFJVFCVMyNU4xHO9UhN0RS9kGBgWdDbPUX
r6hJeU5wqyrxkVmYcthRCe+AJtIRGbFd8cTjY/J0DttVcYJ0wCEz5sLEEUT7u31A
mmG2076iN2LUMQzUUigWoyhcc1aYwWP6cRH2mWpL5jOVkovzkM5OaYtdvudLwJzz
EkxBSD5gd6cwcdzwY9kravJBsVO5yB1c7hnIQDl6/fA1/EkB4EO8VJcGWRh5jqsS
V+zuFTScjLW9MmmuIy71NhAmOHmQ+vPareeP9nIQ+oWYOT1SF/8b7fypUdNGDcAu
GOOisUtIkaeFdEicpzSey/yGZw+12Pe1v5Uj2AGjpzRRjUgvSNs0biOFo+DBcRmx
EYuOuA1ZysTLSsRm8XKDU1speyO5A3oQ/WQPqT2ceRKejl6iraZNgip9FLOY+E5l
nbvNVeglcxj6ckjvAxJ9rm0N51g0cDo1HBd/UF1FMNkVpjbJtMpdNFkscZOEgtqr
+Fl0uxHrbjTEHJhYP7sUH+lgAJvbzXpwvvrD+9ocL4ULdzeVvLEtpR0qbbs8Zb9B
Xb6JRhuFlxDN9p5feGnorotG68qeg0X7tVbzG0lEqm867WbAFwcTj7mo8dNfa0zB
aOOWRtxbwmR9xLnYwkE98DpFXXQv6+WwYqbEBerILGvg5rl3jTTT/Iyo6TWTBrgv
ica/e7mg2wTiz7wc44qDBKy9z51aOtOjjDrKr99dK7jPbNLfEVGwsVd2rIRj1xA5
vYGEaFHqsxFfuwpdn+KwR9IAg8iRmzJ66fvrsE6Qcdd38KaJvz3sz6IrRMaDAnzL
+3bOhPCOkqGJkHAEAGxazuwTFLtVb51qRQ3AgHAjXwgkRqaTQf81GE60RVc4iUTD
deCQf60zGF0EkrCgA1OaJJtB5gwiMXwpRtxN3hrbdjqSZUFuGlZW26JaQKq+Hgk/
6yacWGOAE/AQZX89dnhZ6YOGroC+EPcwgabZIchYFdLQvx67TD3QMLVkaAu0sFDs
LPpsUfoxMeYD7MlDnIR8lIgTwtRXrSoYAA5Ca5nc3It4bVFI/0C7oPpfHHTOcWXn
hCCeOtRvQyNE1yBJUj5lVTD5Hb5ng2OwNlH5uOpvM9qM3pHdcndNxn3xyAUI6Y6T
0clqVYCGGxRbJkbMlNCB6UrP9qxpzywBunmWZETePuLwIeUuV7wY5chxzk698njh
I16oMrVxFkFGFYhLBi8HgTySUJptyjk/QIL2hYG1E8NnkpCgYkyo4TVotb96SASY
H+f+YYQnunVo7sANY07ZgqoFVA4qJZT+U3Gi7fdukZaHviztLbL5skuwwMbKaLnS
TAZZVkTpFVceWsMrM/I+XSpjuvTLylf/WghhR6ciTYDSmq42G2a1VcyIVXZpBeCn
XIGTa9l2ChvT5IEjj/AvZKCQwZkYh0cY2vWihZqzg77gAGU4nCXV4fxXl8hKzWxf
yzVliMHmmUsu1FEPCEbLkdMSxL7oDTQN6P6ihqMHog9jW/i4GNWYYiybUz3OFOzC
3DNSzM0cu94tqMZTvF7ipLf+2K+yYu5lOQX+LGZKs7CHaNdWLDZHFIxiBGxfcaNI
eWqMS0OAA7A+YQrwuj/0oxK5EPWi+Tj96T7aacKcC864Jfjr/R8BTv1cUFOHj8WS
HuGRrFKzOIEvNml/sVf2ztuP9aJDPTHmqkhHWTUpUgvohityPHgWctOeXq2vDwd8
EfF0ze6aD1ApjoRio3+luE35claiKbZsXllYFRMan8WhVZc6MiMAUdsceBBkISLK
Pwccbx4sGn71xjnBQgVbM3r2TIP0wNcZOjs+M1aEtba/h8/pbRXzE/+xFgyQB7nt
U4B+Zpe8fh18kwOHFthzFoaoVg056Xm27Of69QansQalY+kSITebHothwsj6ckQh
aq3Wh5liF80EDFDp52Op88nJbrC27BW2Gqp9XdnhCVHj2PIUZbk+W4KdD2riLebs
YEnegL1WjkfdRtJEVrkpaF9S3KSrqdzWFmMfSXtnt8wPcJgcGGIHQg6//qxSezjj
aKbMpCzg25Cd0arR4KJfuDdXKwWxTjx9gqr4J4uWSB728fd75oGxOJ5fw91s1wHY
MgHbqGt2px3C/f/Ofc8yPNydXn+w8iqQNeUJVT9Ru7BacPsYLyirpDaPHgB9rz89
Wlx+31i7ErLdZaHaoJt6xLgl37cWBcpa6AXqta3f7ubbs/yS3b5Z2/7LYu/pJWn0
TXSQlQ+8/fIuRmbJm/Sw2PsyNkrTwPnxlNpaXNCB7IYyXig98VHCB5xDNkzbHrPu
pDXIIJOLsChwsfV+Hz1fAvOZOv291T0wYun49r4KuT4QWkZ8uC/SIFzVTzPDTkWj
jsRyIr6H6mU+RVLcufTVo+p1h04iQlO6fpuRUMtcU4ov429ivZpGMMeG6JuCAce6
S30DIlyE9E1L26QuVu33Dnkv9d1SIfLhr+QF0UcjVtMPXKnjQG269s30SCIxnps7
YYl3+hNxr6Pp9O5hooq23QXAdC2g11EvLuXKegsfPMLY4R5Omgf9CgnM/AYmwX+a
sBTz3qot86Jw2XgkWLhnk68gWv8nwe2hGH4pvfnsj9J90wmMN7Pvs3BMQAx71nRE
MCo7vKkXtL1R6BPgbAyC+PBMTz9T25wiuKN1Gh0iaXXIZbwkauo74aFvy/80PMpN
n5kfSfLQatLreiSB9NeLWGjGHRuRpoQUhHrY9OhT+zAfCvDdhN7hqKvVdsbQ6DOD
Ix39wTFIy9mayJgJcuQn/RHRF2JAVm8PPgOOLi7sVVdJILt81D9CqoLwbSDTxPI1
XE+GVxje1FY6CGCNNLzLJTtoh6qXtVzEvn4ZrG+Piyou+IbRQvTSnqYpIvpdrsDE
otLWovElzoO4EdPFwGn2hmIClXzZQHQcwuYvw8JnBqchfL2rgSNLh9wY6MrG9fvd
/zaZFs4PnVWI71l+OEL2R0N6Kh+9JR3q6CnStTbTeY3WGZOHThNRr87xV6CODlrH
zR1az2HO0yoMlWaIZF5AGQbi0KmIpa25R3GiJRbMz3LKXUiV8a5z1y/aA41+0p3t
ZX+4ivLAdJTpUqxMSd8n4YK8RziXx2eL3fQocdAoFdtQ07mRWRxKfzwMftdzfR/x
AcDDNmL8HTxVnuDsculDdAAbshDH2yOZ4IOcMJ07JXMn9Gd7AupsW2PhVFYZLxL4
IYSQ7nX2eXrS6RBFIlVILfbuk23M2td97UyrRuwPHyhWuRVRIQOhO0EF853N6deC
k7FnIRqrQ6JOykUJvd8iunIzB8NEZLqowvNx02d1blVW53+rYPxYEYw1EmkEUE4s
HPXww2ipZLAuj8A4fh8K5Ew5vxbpnPDqahvTVWp1VRe4G7B3nB7bpW1eupToQ2jP
GQssFER/Kp1cuDHIp2HuzBIYqlz3PDzCaT/UwE8x9fmOP2WXt+XIUtJYy7nwarxn
LxlBdIU2VfyChxRd6Zz+d++1+eT1BTfx41ykEscutWWJzJsv/AJXp5q+LbEczI9P
C8hmlYIaYKj/EVc7tQRvQaodxgVkoqK1S2YK/9H4CUfNVCBW2xY/sOeaS6+dxmbB
tJYISW9i8A3sSMuioN9x86uE7xziiP8cLhFH6hJ6BOWhKzrrlM6jBo40JqL2Y/X+
pMozEooMTOf5BkGyydkfSygh44IJCRWIKi1ATLw98cQjzVcVJY0olv46PtJVSLbk
+XGhJRTHm618McMMoysDgIML/ALXZf0O/HJ00nl4QE0m/HnMW0syr9Z0T6Ee5PeU
3ru162kkmp0zBhRJ95gZ8fFSF2EQzGhDNyeq5ZRF3ODiT87OgMVCt1khCN6ZoNN5
DUAdKUEKB48Xa1hPbfuQUcPXQEtwWzjrltT8CgdiTVksNWOpQ+XobR/qpyAS1X+h
zCd/ZKB/mWVX7TAuHeuMEJCMijUJjAcprmGbmrLjgrtQqUOW/8ucAhZkdJPCHu0X
t9kvQy9oqoL8yl12bf8veZTOA5q2keaVr+J3gt0CxsVt3QhSN+1VDq9609iNGQ6p
z6skuipQRF9rDK9UlOEb37nXGmibixsaM3G5LkdlLYiImziariVV0tCt35IAB1aB
XeiRI869TUQb6LPqRTmDI5k4QAP6DTV21HX8h6wkMY/apg8QBUOxVUWUctkE01W1
fXo4vT+sRGw1qC9idlrW2n6RNy73CQvlZZ0XQ7T3jzInQLd76yJnce2EI8er9NSp
s5e+RIxescj6sLWwB58wo6HFPqMxUA9Qla5s2dsFYHsjwQdhd8iYt657uvYFCK2c
PeD3VLtmWIdSEMxTdDumDrbGbuv/eo1vsQS6IYntMFp4xQ8Cj4LBe0NjEBd1g0kH
kJecsoRGbG3rDNizEXnOJsexEBRUrJFIlVjEvlI88rUicx+2+pTwy79CmVLJkskk
fgtfKBzsT+KxmRwzUGu62U/DA1qm2PfBJvp61TrQ99Rqeo3ARYm7m12NyJiDWayc
KOv3hbszhUaiGetzYkF5epQmcVVNLDcLfpNzU5JKrGn1kMy5c+94krEZdJjnEAb2
ntKRDSgEqKXj4z50gnGs/Pymy0TvfKRjzIovK8PbvF/3jUmld1jrhfGKJbyF+E4m
hTwY9yeUU09Z0NSuTfmX3FUU8ThzMcj4ecTuudmcAYrnKXyE86shKFx/uJbPXYqt
eJJwF9untopx4+3fA8W2UsqruyH4Ks3TD2jqWrE4fRhxCO8a/ETS3LzyT+v2RMCw
wcYHFDMFxhhsShhTGxSnXfz4Fv/4la01J780g5Zfae1qRrwO8NU6MCzcqJ+avuN4
RAsfZAvVJf5xKin4t+Z05mfglo0NFucwpwKGC7G4k5HNg356ZGHb1lz15kygMntw
1c+7ylC3cEOaKAcDSVX0PkuB8am+8/3y3lJ9RtpIC40h3lLPFveQ9Jmq3B1VaaGg
B8lGzA4nPsFaNlv8pESF+YVd2cjfyLHb0zq2I64OiSrMcznbokRs6816t1l8LuBa
iIMevy9+q/0phvt1up3ciGoiuKRADpzZrOG2+4S0fBsF7US3VG9y2hdKxlM1/XbS
ZkfwYZb5UxrnhteQSeuX6XXtu+vAT3etBi/3/bZl9+brIQe+SNv/Ji6aeJuzJwEO
XOHbpzn5uXBxmW61KzlzdjDtgwFKMd2vxgfk+q5mr3Lfd2fA3gQoWaf1e2be4sM0
AbAPjdMAd8Vkhwfi3IQsOXnZUlZgFWBehxqQp8Psj2o6Q/Vaay2kmC/yot8RJlT9
jn0iPMPxzAG1Du0mUGeTsq5HlOWxYuOf6KyeLWCdkymQcn1TBOSyCEW3Rpgr3aHU
vSRoiOZfA47vEL8VOIbP+9rFDNJc1wAb1KIpoM29IRsB8zkBukj6yYKgo5w75lMU
iqbH08IglP9/pi8sYXjr0BQYchDQkIDZ5OPYHvBZBXHNeC0wjHra1CKQwsMlg6N8
xo7T8FJQe8W/pQ8J7mKxnIicXuC6xBP/Nca9RTJzBEOjhHE9uFQeLeJRMFjJihWP
Bwim2YctadRMQsoQG2dklfTTRVGUKhxVcYRIkyLj+mmKqbXDM+9fAWfZI1jrhWX4
msA73nSkXQG+DTchBvCDmhgmeJEOApEjkxkFa7SdU4omb+wAdKkb9Icvojt5tKVt
KLHTQ7jaAQXFnTXn7ltMV7wDrT/UqyPCMx1ucOIaT+jHvIET+tbPwVVOQmx61ZTh
afS0h+OjR6gezbtMs9eaKrPIZb1lHfBmUWWSUq/khBpT6rWTJFoS5zo19PZPckCq
PeaMdgfTZEa2I02mGC4O+KEvUKRBoGSKpvYfhZa/+Ea3Xxg0CnLmM1M707E0isMc
6WCciuogahwAOW28OXDlrukoXk1vZ4XgNLkSN1diP2jFoZd/Lf/S42dCFsSyGTM+
xguiz8MQyPpVYycb7qU7LMp1eTxIP4HAu6gAbED7GefA3cLwOWqPdYy6B6ZKQNMa
IhngequDMO0oPhnISumR6OihK5og3vX4/SxdEO04i56N3+xjvLaB/njeJ3V7AI8M
WOEcRXgQQEwt1htHVDvbiWyj1xViT4XlboLqRTCCke0jmpfPZOXTkreOPXy9pIWA
q9vC8/jKX7hfeLtA4UB052EtLw/AYz0ZBSjUEAXB0Bu7UmkmYQMm067jVhxii57Z
01SyMhSfpsirsSkuIhRTtSnv/zxdiPnrjcCdf/2725M39+t4Nnm94C8IPowB7wvB
MvbB238MO8gBzNgOWgACN2e5aJxDJ+QW1UP4XD//DIFVgDS0ajvLTWoqu8jVG0oj
ug30xj12D/vEfR7uUgSabQAMCCfySqEKM6IMz8y8XxuY05wgeOwxpor0DV+TjPM0
mRZU44ZHURcvXXi2T+d/DJUmKJLKFNM6QJxDPyDz4DEsvaHylE1RguAaXR/JVrEC
TpnL03mUzKevkBFpXPq8hCi+mad4cnrhZ1gzuIvmAq9F79Et73HWIJf5y3ni2m9Z
e1CgOy2TlKG+287a58J3JbFcUD+TKFnHKEDicoa7nNLNdbj0yNI3+ojmukcrTvn2
k6eWevChOIdaCN5mDCivf9NcFB2efWkkWLIHtmcWmbd0rJgEDzuMg7P4QhEAvb72
XgepSGSuHPo+CXXbjgz9C6Cjx59EFce/V5WWkDSMpigtiKyLXLxSF/EVL8oEmBce
VEhKK0dEAuKNRvjC6B+lNDwovnvYci6kugiPcJgNjPn/AnLC7tKVgt/Rb6/fEImQ
KTrO+Be3/44muK7KzAbPshoc6rDyUJMQuiuupdHobcR9TmBkf+uIhLCQ0IdkLa/X
fov0Wsrd/PUydjxdkhoadaa8/16AjohrROFR3dDRl2qGjnimcmR7tdL6vdxQM5Zg
rt0xWLWInHeE4yRyYwcvvrlgCZxXZkpRfq1L4Lf756HLat7SKPXn++7YHHXrOoze
sSmJDdFenIkZ1pl/8TszDc5W0v/c24V7Cteb8LwowUqLuj9t8o24KZuBIC/xJ6rx
vZoiI9DDwGIixpq2DVfsFY4E6V5E2xV8uCRPU0GmXMXMbh2T/jBk7X5JcYW+c6nu
su0L77o3xE3YIVYR703o8hz0BTqzNMrSU2uMD7DQywsNPWsHxRgjuZHMijT6AVy7
jXxXsjFN15ISO9aSB9+zAOostXWVVFhVt16p6TNdK8lgN+e3QQ7vObXvnqch1ygB
rfC9kl5u6gHbSJ9yiEU4hlbx3fNKlBAFnVqBmSCfcMJW5psM3czHpS29yDGmyP7U
iiXi/zJelWEdS6Oh/tBAVQF4ve9m77ysCLADCaTm1Aiq5JfSM7jrQRBKXC3oDqcr
inDlVyOP4PEq3V4LEJlTrmvn+IuawDQ4E1pFb9ppY69pzKpkRodw9GvD7ZvHL6Xo
8JFG3WqKoMwovWQhpnXcgEP1lRe6YWrsMqCezIqG32JYM74ud9v9ou45YJq/gTBU
p/EhAaF3EBaOXXIRmWLCVABjdj35XU7RR652bIRy9HFJZR0dTPH9g4/dbhsluB0M
ahPedgndm3w8SJEsV4u7SFTpCzBPUaHsr0wYjodBpT2FJvfXJHTAv/Bg7eab5CVx
qtGSH/FjUYjhAZJlAbYU1xc8NDYamH2bcTCLXjFE2GwGjl+TBsn8VKoJ8X1Usbk2
WMIoUCXf3DF/38ClYHXQDISyFONzf2Mt4J+JZLW/sv//p5cuaCXpThbuSsBxGxSH
fsSXxM78KDnTH4kTafX4ROCX8UcGfoO2hbu3UxXFB+8bwIBekmx6uobukh+9ATE9
uWvjcfou2bnem4bfOT30U+IhHRYCpRQTtom5HZzimpj/ppuYTAQtsRD+XVNazI/Y
29fv0JA5z/OHug5H0dex3m/bm2w0dVikW1KD4Sh2Fr+uOrIOV4suyIDs4JEkwCqX
1IQeRghCnkFvMHzPb56/sD324O/mVsZxRc+ruoOQMCRd6aL5Kxzq2EZgNlxJsBrI
HnHv92pADhacPqp+oy46QOF+CetniKGGpHSJwkcWkkONLMpJD0WzPh3kuvpYLWwh
EVGqX6YRkLCDUQwbzhOGXFQe7LBRVU4zlaQAkeY5nEwfzeT0q4+R0sieRWAT9hmB
MA+BfyvbxxjpllbWKP7jaqAUg2ScLdwYbqCE3ryYC67Er8DvrpgGXBd0gn7jBvrS
H9PzxJGrLnJOgU3fKNcVkKV6AtJM5ypB7ohum0ROUMBxn3YOdG89lkbWNJK9hTh1
87TxDjgGA+EYRlB85sc0fyorB1KOHwDzomS2YDAKOxSFRxzdQTKXKmghE2p4ZPX0
caJqDMS05coVDWs1I8ZY7PSCP4OT4ilTKXH7G418N4ym+paaVNdgl/6LfoiPDWO4
93XYs/CnckvBvgLAK170c+yvnf1jLkqda5/I9DODbG3UrXPg6Szwr69ZvYCa6bIJ
gpmmBW8/C4OAxBaN1Jspcp+0PtNsLi4evwkLUDFK7m/6B7PVJK5pIFHLlR4lgoOu
AEUAcl7t2hu+v1iwc4zctLI6SY/TwoY+mK1b0qvmXvYG0TsBVdX0f+jA/IcXtusF
pkTEoslk5U1kYqOhj84IOGBOuiJhoAna57NEDviK+8qkqeaFztO8JNSsj1GNpmtX
N3GeWs9wY1+Cl+bbDM4w+8/br2y0O+09OzzENXqe8TrqbIAYXcky+wf53F1G/VeJ
v9O3NgYbgMiXzQtNLfHQDsaV4HgvNNGryKEeu8i3ZMPMHa7TT9gYD+18Ro3hPU3M
UcyTC0UfXVNDcctsaSJVl7zNSHmZdUtNh94R8ZsBdgsplfBqYeStdU/RpdWYOhbU
ZT29JAnZvhutNNiC4DGASrvHYdeQgQR2cenIqbBl3Yb8Y/8ByNpdgYsekTPrQHiJ
l28VQyubxbUvBngoYljzxtwrIK5E1TnotqlapC4Yav0NUu8wV2hedcL1j1w7YzHb
7EWQYi6UuH9XfFr5EXXcexjBnEHLG3bGu43MnXs02jMszsVdL8joJXr7XHFw1Lyi
OZZ2LG51/dM+13JQUXqFh7JETMpGBVtWdUuq7u2clQ6sTM+pmijQRoLxmXm+Dj7Q
yj+ljj39/0rr1TaR7+Lq21r3BHtjcrxJMCxKtdYPU7EYUSmjJ6kINiOaPv39+jRf
RtQriFacUPVfvv2DGPLQCt/J7+5W6S+R4vSEzQYL0neIEE9hpKyJvMIru6cxRMqM
fwNFmL4H1dMWcbKq4tSzcP2zj+YhQN7nwdhxbuJS46uD31FK4mixlkC5WjHQUbIv
67XE/GHe1BRcmRej2lkL4AYQx4g7wLvL3FysYaSFomQDAr0JFXyJ9WIPJ0BUcoVP
g5ORmXR6Kt9MIx/RyIvHbQU3Lc9qHlnB1OVlxj654waMqxFtOXYzn6ZnKmWt5kRI
RadA/Z1qtU8bKKCAhuIURyRYRDbkqakAO1C23/OSKM37itCoBeQzwQ2IVm1jpy0Y
bRd+GKw2RGluZ70fLbgbrl6FeNKA1a7WE1U64aEapDvENbUvUgsZ/gAJxkqyXOz/
dZNp6SND5r+QVEPEJMRE5Bq9IkPAzMzM0CEctBZY8QHsl7/nQNF0IMC51riiMs/3
zwRDzvvTJDJb2fQZjEo37kVO7wsT2Mh8XYTuKgGFWooq1P27gsU6fft/xDqIXQAX
4RQLUaQwBf5ABJutRdoEW2+yhgmRu/831zZ0F9JI5jULbJUVu+mL5MqggcifSTXu
ws8535IN72WDCSPjGOaS/NjwgnmRpvqjnvlOQSBeaWWreK/NSvLLh1lXSBlCdGut
a6fThBkjLGbLY1bTdXb0ONitQMF9qsf8sgUFJT4T4rKRB9fsFbnonlCXYdcE755M
1DE9DHKmjRj871xGzEkd6KKBtuHItEUBumVg0NqiWBiw74n8+5ydamDvVKQw4SWf
NN9Kj1xUOt4helODkHev0MIezUkSUyiDTW9Jsy3uE9VlVxCWRIeKY7LFSvaeZUKD
m3i/elHeRc9KJZH8ShtBXnEXsNcCilcaoBBTZLLbTK3SEUwxURqqOwhhYvViodaa
l0Zy1BiDNZPA/UsrJQOT2guFtFSAjFo8kLipy8N/y1B60xjFXWIy254ZGq7Q+6QJ
WkcILirYXg/q5spvcYIku2hIvt2BA89GD4qgez9JuWpSaW6KcYmg4HPY/eOyX314
3Bjmxhh0jy7dRIlBr7kYtPk7t0RKdCpoxPUVdPrkBnO61avezs97oi6fb9mEUFAE
D8vPuZ2cwPhLzoo4ZLW9RvXHbgHXJqkTvjv1hqhn1nhQCoL0vhxP1DPN+3sGmEWS
bsoDJqobZJPUUz84WLVaLzp9JO2xNNPIjZCvBIkvI1bFJwEqnwMba1TiLKtywpab
8ioB2Koo+cqXZ9ZqHmAifeCvqweOSmeSUYTMqWfrMDZXNNnoypw2PeDLEa/1ZQ2P
ETTle5nxa3s8VzvhIgj9ccQZRWQIjQNU0IxSvuI7Q99W79Jjkrez13ZGbDlLYZ5D
Ir8ezdL5OOnv+36Q8IUKMnlLLdzeyGHHOmGuu+lgkpaAhtPhTPDE72l1mTgsfwH6
xN7CwwQ7kL2KzXQL3q1KU7rZBI4Mjoyh+CYZ42sTUesJKl84gx6N7u+wa1KBAXLZ
K5ee5KXMnQ1BGBLMZT0JkaP8+xI4M1OzKLz4Pch5pIDD+cgdaMm/YR0AKHglMd7c
18/fidx/VbYJqLKJruhrPfDkhGkVqX8B9zrhf5PVf2JrasSEP3vJ6DYLbqP5r2jx
alm4Wd5U6xJhDJY26D2FacmzM99i5dYc7nlWTo3h/WzyJruE6eWsovctTeY64TWg
E6gfGy+Zk23pwH21dOuz5tcnKxthLeOv9K/t7dSyqK+UUnkOCEYgQK03FP5NVKUw
JCKhhndfnEOgrrR19fuSSkKBN/HQ27q9q0+3LVK8TAcvGBd1QSDcS8EU5KauG9H6
CNNkq8sKt7v5EPLDH2JNnsS7U42R9+3BEtIz4VZeD4D+CwoWgZhu0+nyVMPRbYsJ
FnMkJOAzA9B8IfMnIzXtVI4rizRYrbEUzLd5Frl7SAozEVLGzNkDZ7l320cWrEXB
+8yaEP3Snd5N4NmKtPqZQ/FBWrZFsp2Fqpi54rTZRB9I5MKGqsX9uhIGEVS2FGJE
7Gplv9VCcV+6EtFVfuxhIBZpfNNTA7Tq3jVwesQH3yBExVDyIkjyEIZq8ee3F6Iv
TxmDyFoYoTVg4tIUGL48RoGWItw7ENNLcT3kmha/PuklnkMvJcXiYJhjU4EceJKx
g6APMWKAOsdg4jeVQiL0PsEMn0q1GWAGzG3vXGWWqKYcmAadCaiA7SUWL5gGttr4
r/MFL7Pqgm/tS1zoz98V9PtojiSwXewfD8Bz0sjJHFL3uojBLN7+63RANM3o8YcY
bNSzeqQSUzdFKM7B/MuEn8/YCVsaJ/sH2D+EXfe7iBunwj8ZKEfxmd+wxj4KVM+g
bwUmq6tA+PqNyJA9RjKu/LPa8sk+ZV0HXlvbKx63MnDpN1jbT8s/QUmdbRGpJrvV
CG1RPSaYVs69GftphIokKjoxB16KrjlKIbD0KNebhZEC5sAm1WID7PJsCL4p6cWE
V7P4l21hL0K9TNxA+AM/rwIDxPGgJ5p2DquqlP82c03/6N91vykjq1Ug5dflIIno
8+SPwd9vI2erv/tZ8V7cG/sYgPXDt7PPilhkceLUZrbB/f9yIsx+u3J/3U0/PUYJ
Amfv8vrjRBuL3L+CzPWv3XlpWN+SHPL+loxHU3WXe7UxfvncIo6cvUrPkkY96peh
pHsKWuR7U6mCGPLwkKiap1aR7bhgBeKuja7suq/4Snr56It0uXcyvshY/+Sym5kJ
kDz4HF2YC0jc52XpoNPKQ2CC5pfXP2s1bw2bWQLrpbuJJqsjWQ9moPIPemnFXELE
T/Qj9978ylY95KmVOGIKq/KrRQR3c80YuvsLc9z1T5Th0rnFbQS7bKZQWBgxXYip
KSCPSFP99CBhXKvvdEgqmbhFdUSdjXLFwMW1aj/ZwlRGJ1AYheu16eZwx0WImW1c
0C6WxcNVv8ightgfrPm3XL0u1V8kCp76Mns31GTydzH+eyN/MjW44e736lZ/I/gk
9s5aNF6AeeAakdEEDA53UNqNZHzNMkLBzVitrMcxdBN3bKep3TBHudNAjyOcC0L6
dhqooOYyGA4bJ6dQCEBQ5JwC86Vw+2mw1I0mYyG/O08fcWptFUYIusNberDI/Q3w
AKJneiay0eeRs0Fz9bnKw2NEuJn+W4yftFa31iEnsJCmI9e84IkqpUsJl853wJ8f
orGgLTVInLysPydWpilfoYDX9CNuGwUq1OMij4kOW8wsm7Lhdj4EBT+6W47A2Ndi
MQ5qblLFnoMHFibmD+yOmQByTKPPIepiKco1mSbA2Pj8/H+a6wy+x/CcS1ztsZYt
v0tloHtaLQeH73SR+RJawUh9q8q0sIRndMLjpONv1jIoeSaagdB7sDP6tWocJt+N
mVlYe8oag8pmBHM/1mEgzl9Cukfsb+MbEkLg/oIsGR6EQ0KjduWLrgVCxsJAX3Zf
kR1Y4Z75yPCA3MtY0O1XMrtdhGeccQYxS/6hK1mRm+Hbs1/x+Jsv45NnBeT/XrEj
BZmS654MY50A5U1Uh0yroEyoFftXoiLvr/nOj02u/4T73y7rpHnme4iSO0IDvQmi
XI/FMB7H3i8hN1DBUX/zXR1wm1cLUzu6q2iebFvYmsjnFHG5gI8dxBUPnST1R5pI
WRVAbWCM0M8G+AtMR1QMF55MMOMSY3JL4A3zs18e7IyrlP/Ixgjs6FPMgnK8qZiR
5rfMbmfWz1a2npZVx6toZOFX66FS9ap3quwWwmd63ruw4+bVULC3okgERpJa6fyb
KwU1r9PlgQIYAVCvCqaFdp11O9XRPDDq+8HlrQyHQcN8+ZSGv2eqaqsiNeHWtxXA
6o24z+kZvxgSbWIzh5XM2lajBedG2U0ut7Xl8jbWH+TUh/azRvzh9M64aaVLdw2f
yZp7l3jKpUeLJ9ASS6pvj9+qk1o3dtUttdq0FwzgSaZuEdaMrX9yCAelrW8KiS7f
tHIb/+wSHxFmty1etjtE7AGFVteTY8LmvMKvvHB+v3RqDzvA3u2lnMKap+GmRJFJ
d5AgdqyZ0JsT2B0flHrnXwzAW5dsovMD6Kywvqe1SmcQygRqpgMZAOrbnVahL8O9
IvatZNBd/VkF7Wp/iSWqqevArYJZmIJxwYKFWTpzmfGbvRuBJOEj32klDvsOa3a5
9KcmeDLmGz10X2Fd5aexfLQd899EokBB3ewRQ/KF0VKSWIAnE7AjfC1ancK92EQU
T0fNg1v5nSxA3N/Fp388Pwj6A1gmR0AFwi/SXcPTjDkZNEzxOeS03RR8Q+IwHaJo
1f75K8qvjBUKjKbaC0UyU0dK8qqiKE0UoTez/aybvEuWAkiA9PQPKBZEXWDjxA1S
gGLmZNjt/woKSA4+Rl3ceVs3kK6GIh4bleHpRuLWcXDVR7JkFFYy7Jvf5HDYGM1C
gjaAIa7EW+/BaC54B4RpgGwPZL7opB42JZoI3xeBp1lQeNbZE8IyG2terZ6k+SFu
QVNA+A9QbFY/o5TZpiOXkQNsg/aVDjJiGU5KsEecehvghAX5jxuEOII9XRr1d9zT
4kxJWlTFHk4roNL7iuhkn9FU1jlMA6ZdE4TQ4IzVVihfdonndQabWgFRiNza3VC8
JGo00tyVSpYUCNz4QoLqYQy7/m+a0Rl/3/GTP+W6mM+JCI7eTiKxPgccKX8Y0TQw
JEh/ep3clZY2pKK2pQVlB03HPmcIaT7z5E2At56hl+Dw8DeoB3REBxJhZal3ifZL
xOMTzgTe2SKFPl+4orlese6PConZYrg+mBDcpL7MVLXdFVbQ+Oe+0V8hDYkyzZBE
XEx1J/bQ/Qf7W5u4stc/AQMNMl/RxLfGvXIf4SQL9X3q3l2bqpm0zkD84DOv6Ook
ydhTJBfdThvKJWX1+OhBfn7wv9fWhbllE4jlbRJhLidmEtztq4H7kTJNg8dXYDhF
RX2Ff1uJaELOYdT0FWwqI5G0suUPWT6ajJsxP6c5MtzycexOERZ61f1K+HVn164g
16RT7Z/7iq4YDIBCCIu5dfhYN50VDcbxl4EM7eKK9laJ3f3lEDhZ4hVNs1CBJm0Y
XCsGzJPhpStmLzjHgUfgJlUyif7QxfvWBuTUPBPCwDsr1bluLFroM1DlkQWLGUmd
Oeu/jtnGJgbz6Vco3Gzu4faXtYNI4Ihpxe6M9HeXXiZ9VibCadBHKXppx7SU4ojv
4iTSg4B/1E58xaQiEF5CisbHYhcGXH9NmjMg712Bu2M2PgXSrynbjSLeAEkUwJiG
3XIR/oEgOsYPFkzI5FTytU4KSHw3rMzZHfzfLA78C7EWBphIbFrSTYgaahknADlA
Ywo07XlnqqfxvD8oPDjpv7TMTkYFaXT8q1+aul/YHXP58Ct19KkpeSd/OtKqLN72
uTk5WDVr7RZBoP69e/8YpWydP+WsXI1rgIouBFvVOogaP/sGHSTYHKlQ5suCAEJR
ixO/GxxJPkbjMO9sH3BSchyeD7KYlip+hLmhGvrGUU7Ne86LnWdoPhBrDCsxrF9a
hwXkYlQ5Z05jMwlM4uTo8l8vYp9FTGVsQDeHQ/JyL1ZI2t/vD1HeSLLJGXQIOdjc
XSfLo1cEwdlkQdWKmnfWbQlJ93/FgyE0VA+tUz+0eYSiGJR6ikFn97Zc1/kAaDQy
LredBZ12A1GMeNKkhq86yfVdvPQ6x1QMJ5hARr9yVcS44xnPS/OXVgDjGt3YQ5pN
XcFKBbah8NbHamZMx8vxNzQ3EBfRU0bq0V4dGq9iOgwsro4EDQnIlTClybTuSNx8
7T8oxNqTUMiS3dHq6Uvpn4t6D8nzZ9njXFS17hqpdVY1/33q+7u4dgyfPXaBid5B
GyDpzhOqUPJZn+vjKcTKur1exKviChKtEuwcMurjuO1h2kE1aQZpposuDKu637SM
PPKztzxG3ErTuDNjpyMpXh6v+nHwZobl55zs78Aord9Nc2+NS4JribXLzs+hgmEs
qgoyh7jP4dpvmRe+bp6SGcNCFAYpP/OcbZSt2T1A4O72scpjpJWuxvFxp4oV0Lef
t9JMlLz47GeWu96c7Vns3IL4R3qIX1z2CsM3Xh2hen6yB3ZFZMyRqT8myGXtoGqW
EhR/9eTqIJ66sYhTtH8hfbtVeAC4+25MSkJ4uagR3X/nLyI00nwPD/9AyVyYHBQn
hGqobHb8OhnuEoh+xqD5etgXExxoOnqyGPPeew9rsDFUVKUUWcSpzZxdIHJ65nc9
N1SeoWwCUQsLyQV+Kc/RCJ7DOZw0+NShJF8V2oWbaozFPfW5DyjpouL1q3pUNXuK
mKo9pwBKpZ6FkrdjHfpeM4xbXw027iWw3KnSr+6hoO32VruJsvIX2DjcJjPJqtda
jDEJHbZ2D6lLeHGUrIkxiNs2gpNJxhr+MjOTEj+/bfYM1YiJxScZQSFev/BNDfrH
iOX8QKZODnVim7bQJlaUEXuS5CljZQ6owBtilXQvr6BRJ0xlJieZYYIVIJmasuni
uZP1y5uB5CaWtJe1OGE9+FZiNdDB1gatYJhf9jOtykIrEE2WfVUABjBh0oQZtMjh
TJ7ZlwOd9P3Bq79+0ScZMS72djJsTMufIwAwRlqpDemm1WKem4qeKc5NmZiQO40z
ES8aWvnDZrpl2Y7on7pCoXUfwfXMcPnG9jW1/8kEQ8l0x4OZyEUsMcO/NT7lDVr7
Nt50A5ciKvDqp3+6ZQ4PTQN0lFDE+65huQUetUvrdXWnhB3W6A1erK3nsOooqNLc
hyrO7g7uTqwERsus/MvV4hdPe3ec1f1D5R9eQP2N2b1KymJOSyZ6/2TXC+aPno5u
SrhkRcApFzOONtDqLluotH0A0jQyCrKplALnAUL8W2hL/sgrCndjBeEBVBRQZzhx
Qo8eUxA9Ms36KYEpfcz+P0emR1JPe+xE+auUVeW/lAzsi37SX/RCvMyE/LybepFH
p0W3zOhPycSFc2P+9F04SZXd50SoDOutvVDlDsqpSPE5SKSNG6FsI31kKkDWDl8H
QiYv523RyWTYryMadlT8XmW4iOWxCYf7vr8Ea6Ozqiz7rQnAwGJ6loL1SHUV7qD+
CgqYpF4uk6wTAeXOoE4QdvbzYVI1+Czo385dVUgHs0qzMeA5diiOaYlP8h0zaU7W
c0ZFbTRGghPGnvya+UMi24EiOFrqrYWNlSF6ekeN1cs6b5soYKO8LFWIrv1yd0Vr
DPR3styo9rZE1Z+FFVbAgtl7F1U7t/4OnBUrDM1TNHdnpTrkY7jDeJlyozfWzyzD
83QUNEQJXl18UeBy9gcz7AFdUsuFX4u6lAcYPU+FqorYfwSSD2QyJK9ThFwS3ohO
zg4bNO/0cpcutfu7o0xVsgZd4Q0cZuCDM0ExV3DfkJMKSYgAn5v7bUnTcnSFvl/8
6K2WgSSUCILFT9nwATVVcY1Mzrj2071SbhKPQkhqnzhNWZefbAffLDWjeF/YSzcZ
9dCgF1raVgi/kn74AvW52bO16XTRivGxd8I0qDF05pU3volQ732kvF6XYH4Jws6V
vnPGbkjhkmrerE4J3kTtal80F7ymXiTQl8wcdel3fACSDnx1z0gQ7n1qk0i0lH19
HPTHJp411zWNWUbFq7Mq/egdNcXQbbwsrPHy5O2b8UbphTQeVNujXe0Z7E6A5Wqz
mfmYI9nWnLitnnEmfiw6IAw2AyYT40Yw7TynEn7SyW2E0/FkHajiaZAQzmTTOj9T
td38nPEHK+tu4Mvla4XerEvk4KIcr10v0jJzFYy7hAuElUQmP9/T1CUpxGJjv7zw
auKzVG2Wh121BYrMtmbOiYmjKYH6+pDDNwrOgBRS/oUrqJ9quR9/ynLAETLtP/7F
cXDWzg7Hl6J+Gdgh1iXFdLLXnwMbx03cONWrnBgFZv8qD1xyK2gjL1bImcVYPTVW
AFIEPSzd9BxHVIbID8+lXSWLNxtmaw54GYyUkvcuRp/cc4pwKvyWV5jGI6NE9Xw6
hJTWQY6JHyUZIGlvDsd/szxpxsFCSwvd826PZT9PNYz+K4f+cb2ejjfdw3YyolRq
tHL6RNoqba00Lb/76asqlGuWnKLFGSr2h9QPmsB4x8CfZhwonUrlCqnoVo7fKr6v
95N3VnblgY7oL3WIGrZsi0McsjMGhepcGL97s3vNkFMwujOmYvIOEINJRvQ0DrwC
wWwfpm87NjuqflJZKbKH7J3q6pimbrD7/05GiHIpYoqYyKZHtmAQtMwWoDpQAx4o
E2JEXehdYXdDE5b3xvGwlcIO5cmACZiXhhTzh6iu7VL46tSikYi7k198hR5eo0Ra
TMRH6hPYs33gGf3KINMy/jHborqF39Q33qll9wVa40c+z0xiKKuqzlPTQ1tS/bv9
DzgtiQ+PBS1KTE+2qxIh6TbZvoySnDoTmwd5aXkXO9kINGGvZG1ltXR11mclhUO6
qz7qg+7B4U2ICnLPRmnud20bCAj0P9SgQqRWRMpUbTAcsgBsW/NBOz5LkOdUi/3p
VA6DCe/G471zNCRrfvWeL21t9mFs1QQTUO850lMKA/O2xhiIKZcUkyxrUO6kNczD
yRTixvp6lF0CrJqxmd5wPDYVCApGj3SXp4aT7HBpO0kvDuj+SJ11quSXRgQKTLk9
POPY9XFdHpzMeKNOVc/HF3xisWCUFauvghYlJ5AZoK2faAk59oP2xbp2OryuVvBN
9nYE/FwMPFcc7c1VnT6VbM0o52hF1PAlZFSFZglbMoFEG4qoCVV/5arfdulikHxb
jZ6c+dHd0CRgLPiTByRDrppSeBerws2B0msx1lMuHXT0Bl4RVxMEe0lqgWTiLX1a
DPkMffypzlFe/afv1y1XmjBnbKFUmM538XMKbIXKBfa/DvJGugaKWhM4GGxMfjjY
+BoEnDmlR2mdcdhnDIbdTfIfTY3SJeDUtj34b4q4a2c9Tzvv11ZSL7iKghOusDSA
nbACkZxwGbjr0E6vtN7kvH/qfMib5WDjr9P47KTbBLKKZGJW6UqIXoqrbWTmdt3v
ArU5bJ594bMZOLiUMT6SmVKlYu39D1cxSSDeV4jv6HjU/VVoKQQFsydAkuvKXi39
bNe3ueSaajQQ/xvOlSKDAx2HKYCg7ObsjJ2h7t1a7lgyhe3yofyuQmMxAmGoeu2c
nsRrmpDD8tMISTb8K5fAolVFtgzcf0AGDSf0y6YTjFicDQipboAZlLdypYLIN+rd
4TUkaB1NsexOVkAsd4USPW3E7l6eO5Q1h6uW7eqHUpzpzrQR8lE3QiKA1JfjF1MN
C7fNEtxMXTKa/rmAGx4nuMArfTd1CHaM+qTr1BCxaZIRLsN/UnhzRf4IOiEjzOFB
yhK6qrlPcsFNk8SIy7QhuAA7FW/YEq2vZj2ZecOPHRoGUMJL4vdkmjEFyE9ZlFvJ
K9jWrT70UUab3gnEykWWyEauD1C/q1I5nhrPvhvXgq557wVuen9iREgF8kf68Db4
OHG8EwS87MzIGrkLhzoEsJrtwOJKOLYPZ/7D502mthO4FDWeeXpCNWJgRSeH1ptU
ESrEhMwE7oifcRfxtcV2IEbwGYCHcWuSGwpFrpDw89KlVuq0NnelJFP6uPAoOlQa
xtzGXo3mw28lRccfoj+vz0Swqs3BrEV3tDy42A2dVBoo45vgXe5WhFh7lwcQoI4u
XynIzCpPl+97Q8d5RZxOtVJ8o4n7qh059vwVxnLsfNaxW5qtZTdSR35notOgIZE8
6v9M1fwc9EVI/ZXnosOXzdPGJU+4Ra3YxMdHjE/vZhWB26lLwSA0sc+PJ8yj41xO
lI2blkUfbt17NQJTtHCSmGuqhVwSTaZUVvMXmQ6BV6YytVtmRhvRV4ktOwePQtH+
yXuY/sATBr/F8Sp2BlhXfEF0C0oJ698nNJXcJCXNVSwif/ttlRuSC4452RIukKuI
3IJ/GL+BRyHViRDWKRsD2NB1j0lFmr8brvPxYJNfmXXJcm378nwvgY0UGH7+mFXE
ULl0UxYFW3VqW8en14VZdFPE/T+M3fXtrdkOhdcoLbgUlOlBUsJC/xAoOmwxIw+U
D9tTnoXRrzxc31GJ8xI+tE69MpJMSIa9cyIUPIt+HmCPafh5OvyVGNzJ/e5D4tsf
UpwZXcV11b+E7WqpQH3k+FNyN99rasTQMcwpH+C5m8C3zQ0muK1yyYMhptT4umIi
1BJHaa5WCwwFQEJlN2kJhmL3Rtb954qMalq29adoxhCj3DFuQ8TP685DHkZ723RX
NJZKLcmSjWFC1DfWyiNyUiVRZf099NERnVcfuzJwgkZ67BIIM8nJlBs56OkM9lkz
1YIM7oRCCyfX9gOqmGgYvaYr0TuYRFkafMzb8KY2P4rtYvEmlhfZIP3bzjnT1kZz
C3RmWUNAusZJlAkIZ1zDhXQbApBKI62wFYbZFgmWu3edPCwmfXzgVsYC+lxuNwhR
AYOZuyInzFs5G9bd8pipcAGVcfETtErSZZbKwibhGxcFUKGMY2ZL8FieM8HqsTj4
Xs0H8+lo0xAWg8EpD4+BJLsf7A/qtnXTv+qOqCRKVj0t7NqI7uHHd23ttTugvOQK
B6stPO3lZb+sVvAtDve5wzKFPgbIVgORBOQu1jgX0xz3/P2TBc9dKuTzV07p0qcO
TkyEry8vPcHSrnYzbXCAn3lW1vCsbHnUvnMYV4iOuG3C9ubKJvIobWw12Ldq3hJL
cQ7cZxyhU1Mv/JFMJWH/YEtYGwdrDEAU70AT9+5AqzskZizMawlw1KIgTCmlgdnx
/5idzBQDUJOuuaD/QH/udBHHaxkJ8EbsZaOrITnj7hSnDm9lFRYkS3V27HzFNj65
ONHiIy16+UPwjFeslfRFodyeeoIpYJZ/Bbrpd2s8XJ1Eu7mR7oXSYlDKjujwA7tZ
EwX4Ygw4zg1R3gStg+Mo5ZVMbY0DTN4Ki+OiOSIQrmgCYp0cO5xtCZmcKpofp6I3
fZfd/Sbk8TCS8tJbihHUHgnnteXvs4CIn6/LFvznAOWIPoTW1ZGbPyrNVd1s54z3
ZLU+c9OArKAtlT0KXugGg1qOaB/F9U4R7tvXYaNef7eMiSRhIHbKY62JYKxZEVjn
vMNWJh/C1NQzY/DxoE5SBlwaJDIQxMZNMz8Lsqyb+20mVE2kqKYd4i/o0F1CXoW1
AS5KJ4vQRYjr9TaTob/1f06oa554UiOV7w7ViCWkYoMf07KECTm14OwiflT4kafh
bIXvkLT0xxazySI8sjN4Wy11ln79t6X/XZyZYnYIHEnH5I8TzrjTJ5WJaWGhEHBI
cCo11uztHe+n+uL6t48Nw3Snr5/4v7VszYofz1l0aOJkeLVdEMpy2SHoUGhGKzzc
N2YEXFtBmPikL4rslL8BPoXdIJkQOdq4L0DyjuwOm3cqvaQ225YIy/T6+44MvmP5
lEMnIcY1SQOIbQ8yHsW8NSxG0G1E3eBwcEz22mj9AdSKvJA9KFCGn3enV1zExk6r
HtdnP4LTwM/fLdS1mxm4N8Bol23ycPosouJfy5Un3SuNRdVF49Avq2AqQeueEZVP
cq6RbsalyX1AdkZ2dEZYoAt1JbPzbMbnSl9ixi9l6Wfmbxwn+gZDAOS47yeEXifj
x9qn/lR+X2E2lv0uVYaMn2rA3PvuB/RVbvkqx7aGjK6Q+7iMpFVBDFwlTXJ68bpG
7Dhdy7slzKlh4PU1IhXX/RYr0mQXBxtHW5B6BpmhBG/Dj2RJY2fWQSeQqjZU1HOR
XhH/XnUdLQyAZyZt6o11ijbfyVqoeDW5t9AiVWAJTMdpk5ejwu27kUQL3eqap7lb
+g1moL7TPUwDE9af/6VKsiK8cwaCDb+/BCgz75AeT9MmkDQAhD4LZE0Mf0kmDVVZ
5cpCatDNF+a4HV2dglFqL9xmoe+KXD81jGrp1nePQr1Fidy06jcKdbE+AZPkwOm0
OrlUEgOhSGxdQqHKmbF3/hhcebQiNHPFvJLy57QXue4nVtsItJ901BrXIxsdC96G
lTB4u300aVJ0t64KFpa7COyPUM55i+ODpvvrTKdqKDVIGBAMfF62gBnQFWUiBYGX
btwcYYNhp3eLUI0anEZYbJ9wG4NtyS3WNjgrVqHoJUyczsk+vBSNvdqL08rKPx5r
SKUGvNIDbPjecp3MJauisovPZsfHfgdepaP13ZD1EWwu4WpgHWrGOr6EAstCQlZb
MP7trXBPytiINPAf4M+Ld1H9+HEAr24eR1j/NxilBhf52eU2svgB1huxMpyBYVfo
h3YkyjBrS/F5VOGJ8T+G7ymhHMDUcahtiazgcRgHY9FUiVyHq1tCKtJlG7pWgfUC
jpu1KgvGx7JinqwdooXs3jRFNUJQu88ENQL/WN3Scf+rhaEC5KxXEFhCmugnJJ2Y
Iy5D755WKZ64xGzzfpPvo54IUyIlFOSHg/BsIOmTl+PiBmBh/LLoVOiPIfSiOcRU
FdM8kxsgIwg0iiUnw1VVKLTKmznCCmtiy1DOlGj7bZNrEWg9FbZLv23HYQObaDyV
Je4RcTGA/QzUTjxK6NI1xmBxxgjEA9Roh+REYXJHEC9Wluk7XOKXcvT6R5Jqd8YE
J+H4UVA7mu3wcgf/7X3fqmFa79mHSOQFuHuAKIbRnNLdQKHlQd+irIWCkBKarkyS
8SFi+fwu49blsFgTse5D+q0lWruzHS9WohVOQU5RTQmw5Nz6pCVSErNsXpe5/zkg
N9WjrWoOFVgZFTXi18vv3YP/FFdN5t61fi7LeBFEPtYoLa3wAx/mdvyvOJKInarM
BlseuY7jjpxKFWIAetps4tg+pdrr00AYuzDfaVN5O89DxCnAm9lRXS6lrsaLgLVj
EsuO5UK6ikDikGAP4twmetG+F9dn/gSs42Lc4IZhgXERmUuXB1aNPuE/iXEpK+gS
tGfAZoklw0k0c/8s+MjqwXgR4ZvxU6czsMG3OfENUscvx1rpb9c3WgGMStJUZ0GT
XpTZzjOkvP2dEywR7u1Y9/6Jcf6jqkLbGnUoe+LQqYcEgYOu/IV1rAfhVUDgqMFg
IT0Flys1Gn3LV4lrqe04nWZh6kcgdG80rWk6OjFuqpheSxoVaXbazyA8vK8VVRCA
st9Y78DXn8ncCrrjTp6ntCTHvIxe24zu/QEp/NNvp2BTJMngLb51qcP4RHLwsGsb
T9cVJc4oiPV2D5iF5m1ChXIYGW8VbWLPcjs9Si4vYoW304vDRfV9IUKsWwWKwoRx
br6aW3wy2I1N+xtVsIt1PtJtU3AFTQjs8I+8q8/zmLkkMmI740f9eYQ2yO97XsHU
jxkVLcvAuoee5xrSgcdyXzqiIK0kmrUMJqYqiYFwrewy65j/Ck+LRQelmztq0IIO
2lirP57XZ72Kxh+HL/VlMuI1V2g1AqSYtAajMqhHgSlRd6sJi9Zc6Z1qMk84d68b
sLZ/bF65DQVMPwF0njrfVIeJGMc+FwqEV1NfCUcyFrMyxym8c0U3GJ0ZA4pN6u3O
nQLxXcqm65Sola5R/jWQHE0IXyGActkqCue4XeqMDCE8QOoEzB8We5fBv6iU+w/9
Bjz4FxAZdS1q90KTUI+Nr2qpQTzKK040tRWKkxNTSvFwIr2FwayBoexvqKDHnuy/
6xRrkTFTqSI7aSNJxmfY+H/p5cRqx198tpAxNYpN75r01xcVVPAfR6P9UPUzqB43
ksMwJJCOKy18UxBwPj7CJeqp4BpGtKN8okRSIiBxRUy5ejKFw9LE914yYNEgJDiv
hezjv409Dfg6fWbaRXhyGx5ZNWKFmnbwsQFwqEwUpB1zZ18/jfHPnSlIGshVns32
wIJ0MoOSzOThuPbVJJ/VM+/EmychFgjzxsc1FykljHpbokSjii1sY/dXLslvv55B
eGABb9aqU9/CAT3uZ/aFx0aYCyjqC619nS0jqVlWqBsDyEw8Q2MWNGGttxpSdFm8
/Z5/tYG4Rg0g0ArzcZc4ThOjRpSERlGO+o3QD2ppnlBiaaRKh5cVmdDDUWLV78Ny
Lei/TdKA6ph77AzvDwnIWLUMAMkdwX/sl7hPGGygKUdZ9gBdT+DPLjtZ7+39s9Pq
iip3oN/I90u2JnkA/YAWhmeLZbf2VTAytLKmgcKBK8CKC1L+Rb54+7iObhLvqS4k
hkUVYx3xRT7s4g/zBELvftms5XFojwi6XP8uYQtCQmmC5BgIs2g+KqWZVqmuUwoO
3fOAqbzqSXSXzh1w8w73BiN1IS5jkp3q5aDabmmnDGv9D4BL8OAsmI34djBkkEoP
KqQeIzqyU9e7aj8oDJjXF8f6HOe0lrqoldfYsM+JWHHIM4q/NaK0qCaCQ77t+ecT
0uD1lzdXwuKMhVf1F9gckUEmFE82ZnacalfWcZdgGAupvhVv6b2Zft94eGCAz5a7
kSImt3RUTI47pZ3qRKyY/QcsF7svL4D62HjIJ1tBslJ59diLCJkvFnc7Qg5E84jX
YChNZnbfnv1EWYIHuY54x8lMNA4W2scYutthPJANk1IcIYQXgcxZkq55TGCcD/6D
TlZ+Ly+MLHnYT73PuqAo9jMab/gf6hyjeTJScxsCAMtmTpMx4kIgxJxMai0X0Mdo
Y7pUdrHFYaokHhn2K3VMgz2bRKGDdT0WxPvUmMfhfE2GKXxsRrQ3gVlrYgRTfLI9
lKsJN4s7v/H4UPFqG3Rzt37JO1Z1ZAlOpDci8s7WlhwVKz3pp6PQOUmN6HRepP14
q5JwSnENZXeOPvXaQRFUZQQYG/ynytY2py+li0RizDel313/zywax+d0axqlQsay
jBu5w1EPLjl/sVmcBLm9SHgXrdrBP8/Fn8QlpyEUWh44LDykjVrnNVNdbC7vLEkg
+E0Q9ae8YFovjIoUr+HT8V0azHtk4+BETRnRO7c8pNLUGHIXRgsasFRHGih2JsnS
xwjpGdXuQKRsn54iWN6ai4rMivExgtTrTE3LrMvR0icBiUcjyKymZLi58oQRwzZh
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
iMvtaGNAtrpjf/QgcUMDLpk6BRMbxkMZ9zm4YP27BTpEhVZsTtrBZ+TcVt/RBEBO
3bmF5ELDR9f2+UnSIHDEfOZEnyqYiwXMXdXhy8A1s9AiC35YjyQBEF9d3dDcH0Gs
DN9R0vBHTt6i70JvAfq8eqgo0Y/C6sAqXjuqlT+KQeM=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 6400 )
`pragma protect data_block
GWbID9iWmNHbVrzLbxd6RpsGwf5YX84FDYpTT2e+JcdozJw/3KiWRWEp7NbIauW7
8TzX8eaeLqaP7aofIyuRhZb6s/A3MM/lE/iZTYhz3vDNhjOgQK7U9P92GCPgcGHk
6xpkMCO4p0+AIiyImgKdZyFEHy+uCRF0y0L6aXBRCD1BmFB6HjZ4V8KM87400O5Y
92W/jtDoWcVTRSVXhA+wdTSM+shsLtj7BWSH1DA6BuKEOU6YEfPbac3yIhi+Ce+0
/6BV8lZ+0x5E7vrxvrlqqYDPIfHsrgRb5dA479Z2N36TQCzJmvRYu2mjHn5xSiUV
WC16aZzHWkK2AyjJ9Xt7KJS79w48o+JxfHH2kldPCxHfz4VHCCgGxZaB8LVm+wNS
ZshXbJj247E3jaa9VeaS+8zTAc1d2uD89CWJGkgaoGE+HOSqEI64mxke962Gvcyj
6ySJC5DBbP3X7DdVfdrYlDC8kW3aEzN8ofju9IZWw42w2bj0+xJ7Qd6wdAyBGNvq
EyAIlKTQ+K4c/UP/h2TLMntk9L4/W4QHth8AZtMh96w3r95er053b9ek3iKX/DxC
nBEnNLLrrT8NA2kWQ83HNteKXLV1zFedyYvM2LR8v5cYngx1CwHoJKK/7pm7kST8
hWIYNancmWSkSjepAdESrf845DoA3gEZ6f5K1RZRK62vnEp/Uxm3KmNHwyrrjpE8
RmnlIl6GgYleegley2+PvmGMuzfUBeYOrRS+h1CdEQerVo0VMjY5EGLtL91Iy7Y+
K5xQqOgtDPNzzh8DYBVtcLm5ztYQYtAAPx8z1l502SWHGr8d/MpY2lPksZqKSZQr
mey6i0TFiMqWZcVHM0NsjBx3+4C/ESsU/EyF+OkxyVHOe2tA02EO3V5jktyqSWb2
ZrzgTD9YnxQfAg95ecQSdMT82TxjSgHMEsS734hvDjXdhsRmNq0Q/2xp62Q9ZJSS
X83f0KHdr86uVcPe4j/XPNywSOI+a0dsqLsCROHIEmYv+Yad2zzKH1bSBriXsuJf
Ibkp864KfK+zLWYRbuHjOTjb6EObB3twl++wl0g//OGwMys34mxwJbVeHZKQm5dv
rvAj7kzIQJp1J6/P+geOzDloYIZubnPvbpCvx+Ex08oCaD/lyNgKRx3WMuM3LkAg
3zJWSSiXBW+/5TVF3mBGKVxhniuXfu2dX93N4F9i3BWtRdeY3cpgxNQ8tU6CRSDC
Sh4IN0tAZCw83ewL6o5dEg6VBcogNJq0/KNG6QvzMOQ2TOISnkeOmu1tDGbhTz9S
nFiAhxRfUBU90wZIrDJpQNmcST/BN4bvPMYrV9ZODiq0SLwUbD2JwgDHPZq2b5zo
2rHM9qAKQ6nxtWThXw0iqhnGbhHr4M0E7EHXAZMW+GXcqHNA2e0TpeWLoAkm6YJ6
93+dDF1pxXpk1k42h7joGvQ5AqD3QhkSUUbHgszve3JrSTk8CFgq5FO5UDPK4cnn
s0nbuNUpJFEvRWHOHIXAI8sKB8IAgP+3bq07uFG23CzCY1UCThKZGVfR5BsuLzCY
/XAXuXvUXMmDVwI1yKNoa0hANEDYNfQTY+AYv1mlVdrv9Lkk8H2bG+h6bYiv9pV4
ZSg5VERSfVzAklhd/7/ExBJo4ydZKIaGBn8j+Pr4Was0aAlotRz6lLk7MrfDc8JK
+jWMtzBtbGFj7WBeiWk1G3ulc7+mamwmGIctUaO8nFc70z9W3CT1r1m67TMap9YI
pAT/DkYR9wD02BjbIFYfiO8V0PNidQldeWaSjxwFoYNTgvzEBUXnDeppo2rbL8re
5aImC2tFsHqHL0wbDayVbTHiiFjYHdYSdz3xTBDdMQqNpcMFiWxKNWSnUD3XQ4s0
Qnr0uk3lRDpCIA5Y4OgIOiB0wZHg9svjFRnNZuNzvEhdO76dHvrG/ymeqHABblI2
q1tRswkEdmg9GSgelB+0ejSUuGHKCrdRQ2H78DcaUMmT3XlS1z0K7OzgyAhMXfMe
LN6BVeqgDgB4lE2suINh0IbhPtRudHgN1EyLr0obhnfZaMJ5bPTMnTWCa736ZNWM
914T22WseSuKz9TTyHrblWC4HfRhyOJ2nTncJ7sClcTFCE5dhXBXLz86wQ67PTWX
OtOivyFzOyutbJlKiOW7boKh2B0D1kBE5J55JpoHjPiHxBQbMLtX/YLThHbg4NAF
cFstsvqSH4x/0b/2+vDUZ+ec0T9yAQ3kIVXnJqOzJP7pmI18PkBGpnS0uK5Aqta+
VpASewYz6T9K1KGjllVT4wD+3mCwHAMKwRMyYuJu3k4UtN8PSp1lIVIdL4LbF6gf
R2Jmdy8XfGCAAMSOYAEcZ7+17fP2+rWG0SlwvMvy8FOMuAPAt/YWwBcFtG2vCfKu
FQl7SpNBIGDq0XyN16d4K7Im51SupZx4JuOJ2fKsDw5D/lV4S7VTPhnvf4EAccox
aqfmUN+IWSpdZdD19gxxrzILwAeTbvDWlsyuN/uX4scxXTf6z7qmpTR7NFc4c7+2
EYmPd//5Owk49+iqRaJdUMVUIl3iNvC3KvfGwcecFcLv9pIrDAqLdElrIRkWXQ08
pj4+fJpRggMLwZMH01aVq7sWHqE0m7Rssfyg49fDwd98i/o2XH7RUwGvTxZJou9T
RBfZPmScpqAJasQ9x94tFk95EAk3SEcbJPcDyeu5qGt2R3/0zfixLoL6itjeSHsc
p0beJrYG/EAi6hI0XU6E6M4SiMF6Tt9fk01S++TloOyVyPAgJH8AbBXoy7tt5d8r
jSWRl9CF7RpqpbgN2N2qwTQXOu4rYpMNwKPEVwSwEUQpVvHTeOJMPTGd+7yY6Wc5
/B9vGYVPijAORARwnrDTYlDPEkX7u7ucIIB6c6pwlUfJTB5VZvGi3fNyBsgY5pdc
NGbavb5uD5O8xpZS2c+KyCdNBMpQzFA9ebk5nZVoltPasX5upw0cAo8fBZt6G4iZ
NWjrnoWSTSFRRSIPHW+6Xv9+Jyvw3oHuHDrZqHJ6q4S8woFG30GnSpljCmCYEp4m
qgd2lUSQBiy+vt3f+mwD+QwTufIjAM/5w48gRa3JjyjD2SMtMd4xg2ZiIORVW0vl
qgHCrVBv8Sfeb5AlWzM+nAamu6WjUfmlCRCKWs6eOTAgzDZpd3rIhfidRLrBK12n
VH2SeIZOYINPtagE+vXexQOJmLTQMG5+4AY727IC9NNil7euegBr4EhUm2vZt/wQ
k22ta2RNyGg+2tJafrHZSLgRIHhB8EbetWWUXVHkdLCpsH+yot2DS3478+nvna2y
ohiTCXOs5Sjiq+Brkls9HqQWr8saPrZDjUfysDRLfOL6owFvEQ2oTCbQ9SG22COz
Hs91D4v4trmIJPVwjX/UxvA5Zg+TXJ1EtR1ZizpwbsWGI3XKKza/3zUWZsJQGzt6
GKenSBMFVv9jTZl+L2pJoET37BbX8d8ngHbC+86XSxuUylE7nUtagRr4lR3WEHqd
8ox7skUdRDyDJ2N4957zZayQtOuoNLc6H3U7FIHzZfSWVryC9nDjgLaC/TrTNAOH
Oj68tspQKJc9flgUE9ZpWKmZwt4Y9C5n/A9H90ENDnXVhrXrdA1L0dJ6d2x9ZOou
1/mqbAwR6lSMeTRGR/DsFQDLDmqP+wB2GKOGnGvoHQuF6+cYG/ZcojwkIg5HyEHg
s+BWKPVF4C7IbjZhvqiMUwlKWXZdc6n5gL5lgx9E5LInvtUu4W3829tgVnmKKM5w
zF0ymdMtfqtgo8kD6Re0/FsD/Xf1btCFsZ5fGsIlgrIEVNHqYMqys+o/kb0d0dPL
kRoDdTW0BSalcKntHEkhzwBH8iyVNm1H5CAd5U9BoPlqMfrGVQ65bnXHg/2ZcZXO
kN/vy2ZjcjYrHNvsY0tPs9xrwHsmLsP6FRTKThbe6Jc9qnSu+nfN6UwmcjHZv9o0
Q2+ml9P8EJ3NM7jKkk7FLjZRRLpVStXjhoQ0dzYg483f4UdP+u1WXpXfN2etl8hr
TOEMA62U/hDJpzgEjXo9nyalMKYKxU9wvfF0FOQwjSMibikEeGy0LaX3k6T6gn4i
Up834Vbhu/6RT0AmqNXM1L+ajUYVaUw0sIUb7lW42xBGCTeMZm4tDe1CyH0M3Rkj
f23HlQm99KyZqpAFN28gC+xcRO8brACAJmpivpQAhaO9t8eHzSP1P5Xr/2MN0mme
cMmIVFsKA/q+Sg9IATi9bRUQY1BJa7m8WVpvL/YZqKRoB4ETaNPqfI7kxKfzv6+W
eqEwF9ctYAx1UbHlX7RnuR7QfDfIamnf9QknMgMb2qrwrar5UFiaI1pZfxssd12i
Yd03zCR0zbT3lpfcVj/9s3dGJJ5WtEcbnmIoRlxYbblF4hblZ+XT0LZN1kXnVvAe
rDKaIJBbCGQAbJpSTSL/m8dkzcrW0z9gsJpF0MEXRjS74BYKajyvXNyUiaoI9mRo
oD1wph4/Uw53rSkDIJGJVGoPKrmemaZ0kEpiYUs7O/TRz5qXdtd6vWM/xnXRkp4f
JdmYHxI9RrNXfUEe8+fLvF+fpqvJpWcaVj8aqDstFwm/c+VGJVwrMCo5f9Hh/xch
pmqJUjDIYb1WW8c8fpj/JbK+4XrWfzCMhPg+Uw70k8+T+w3In3caeKVbb4QEw/fl
h6ZC8RmnlZ2hl/e9A6xdv+hWRjIEGuKwVbAh6AciW+ldKzLQ23BlwiXLL+zaR2Z2
bZFoLx7wLL5UNPnXlej7lV1v27WKW7coIW5+9/gS+eOSu8FzN57LBcK8mdU51uS3
qVJ/9PIvvqg9qOqUAf4/Psh5cSAiN9zFvQXF4tdNzE6v7gM7BmNqhfzbJpavXMlm
PNJuTououwHCb2YR+aHAoZAxibYbsaEEbmssV+eDo0lj7vsF83EmMDPQcZT+idfs
kyBkvKggdFV1od3mHrIpAG8Xma3/VrArxFttKIdh1z5u/7a2DYIZj8MJ10WH1NJK
p6bmikO6WZt4uwH/5t2BFLtwWoCII13jS7rgiBA0Atp+hzmBNt3Q8hZ/HQ77uEKK
TMPYsW1Eocya9bixqoWhUrpSDi/cRXu2GIGJmd2elwlDe0P1ZDbUjMOa/4GqJ1db
Eng7EqLTeSWhuq3rVgmSUWjqEjfKoqbUPtydY3oiDTsn4VxKoEXVBL2DNDh25NeG
7szCV5Ojej3HhZ4Ih8YkzqTmE8zU5mqjoFGYJSH8+kUHN/BbsnFmArMccinB7AUS
jae1P2Rlyf/bfXa9pIf+9NmbYV9DC0piV0I2UnjcYJfm8DOrdDNZNENRqKh4FWHJ
COxuNkaWf6vDDhPLQM2Z1cRwkPzEtGaNzdcs7Nnb8RoxCU/C9JoPMsfgmbxX3QmP
rI1O3vE0UFce4x22CmoFXp6Ajpc6tapIF0lHGKLD4vj5nlMd2FHckachikA1gUKU
Ym3bUVMDEsG1ETmYkFkPQMekK6oH+pfXCK7EgQ3sqAKSDc9MSpGEKuxCQ3QeAErY
QypmTmA6xjFLWp0Q1ttQDyA9ldYaZ0bmSF5p9fwivAOLa+5Vk/IFwjtO1iTFN1vU
hRSLJyQWFhO9kIBeI7q3m/iGEFZjNpghlyYyF3x6nkIyLlpVuMUYwtY7SYGxbThb
xhR6SrVS8vjLPnLtWIoBQc4zb4/WzTXaAdiGh68AvuHjZ0dd/RSMqAgPZWBzpYvS
bUYCK0jnhJIxFqPM3aAMB7hLSTQo+Lwumoqoinw5hCG98kixUVc4kLuX31+uMi+v
9o7ZT/Yuk3NLN5W1YuZ5+AW1ikCPmFXpTpam+f5RZAjEJecIssGOs7f48EQUVUas
7hgbKDEuNFDBuNWQTNPsfkD78VSkE1Q9hjTz+LY171YQhJhggIj5xJ0x6emLuuvF
Hc/KZAWkFNTkR9c9IRG3xF5nsUDma9QEKfMyMzCsSp+dPWBcLyTIsJK5ezVKVL8N
R51fXAVfheeKsiq6I6h9NC17CX70+2HJv1w3tFEZ8E4Gd1CuBbeh0FQufkthnGYb
7UtVEHp3g27eXKspkmSpve9k2my5fxBktN4eJTNXQBEbpq8VuJMunr10XGvUBCyO
NsV0lcawejRXNdImTHyuNSCIvYMMoucI5puKE3ORcGWkbERTR9BWWEc1BQMvazcc
6TwdqQ2JUhpC+A216r023JBAZMHoT4rCWBNpM3e2i2RsSXECBP//cH+0hC3uWOQR
51j6InfMODgf8D0xQBPMySsk7OW7vr2PToPlPFckLybdX9/mBzslKtISBCIIMEH2
KKuF7beob9Di+ykCEVIasGOBS2znS0W3YeaPSqBiHJbZYq/J4Vqgkt8WoLNhJZtP
cUdh+F297Za/M0Al7omL2cPuN/485DFooCq6wp15zFv96+2Bc04iUarL4TQaSFiy
QegA4EHGRxVfxapH8FIBDytQpkIGgF3TKnhHbs5rUbr1S0LWaUMQt4cJtr+mexwE
Wcsw1DLrc7q81GelXFw8nVoqe3oJD5MVwh8ACbUODy6CxUIhCehq0Nx2FvKqlqZG
59CmIE4qOj5QHiGGx5ghtC2uJ7iW7xc57teG3abk3OXvPUebEYkVfT7ZxpfQc2hN
h4ErjxRSf0E42YSJVXe2YChefbTEc30JmbJ2mzf4IJpO5ZV7r16daMjlkfgwi+fL
IH6wHs+qVcIR+br1u0GW5nfFOIndfuAsrqXm0oTuDhL3cMZPnuhoY2mkfPOX0YOE
XeFEDUDay/K/q9jyKtukI9nvlNpyIQOc0kw6TXhqIUdtv78wilGcdknIQdtad5oc
gmTLgv/Ae7TWZiS5QtZV3KItoY51dKRfrWlwnycJmjDcrv6UOstoMYFuLbOX7h0H
3n0U6UGGlOTREf1cmaR9phP+MytN4subwGfaA39i8ydolHFC8cCvIVC8suM+r1RE
sxqkdypafCYGN/jEEq+qItqJSLme8wjTd4ZQmDmeBFsvWxq4yBPcpndTWggPXBqO
pL0KsNleO6lMnpVeLDNQ4XW4jT7FwVkkvC/34eweL00VOsml2FAlv8IebFN7CKgV
NSJ4FBS7jJiU7t/EkD97S9BFGhoyiCHIW8/tDdEH3aCK/Unqyb7eN3h33N3aTv23
+3rm7NQyXHN7l809zjMq2HSYS+qBf575427V6O4f8Vq1A9WJCz2KIRaRUpU95Q56
KxC/eWHiLKTjqKLLX8iAXo7YKJpgCvgQ1o9nYYYdrOyOyGn0zdxyuc4T1LLCnw4A
rcIiKZPA8tv34fBzJE+cgPiTlJ+XgkudC0K/39dqKwT4jXIusx+cOdAHEHCvU8J8
kBMeoGVY0bUSF70JlrQdgD/x/kytMnKly9eXqvytYAmKZ2IE+lmOeJDNZjrm1SeK
rqzvWNRmymQ6B/NA6rdkkH+TwcQFat+cqztWLevgLXBaVxIQrqg7exfqip/gbwXn
FYJ853fh1uwHPllp16viO1fqAPfVJ9qfOiQ0kILmZTuAehKiYOyoV/9lHMJ9WcZk
g4kwvFyo4wN5hCG2b1eUkc7BwcIhbejSK+iDvA8mo0J0N3SRHOuvBHX0/fqY3/C7
P6oVYiJwptaET5tmSKPhqcj/gNxYPbOzjEjdCsaOdJh/SDICJUOj3peQNssFHAO7
rWeirucBx7zvRkIRCAGfTN4nyf4WIVRxOqOCpMpEivNsagChdIiDx+A/iW1aZ6Li
QG1HiSOub9woGHYq2d9PcnSs0zSWa7COwJntwaTSygx+Jx9wR/IJNaLUDnM5nhay
f2YQ+3sj9SGb04jkAETkpGmpq1ATR6wHOkjRL44/XgCwoSRA5PQXMSN0E0gq0VIo
Ci8TXEfopXMlqe9gjq1r9EUWiI9Yw+yDnP9vQYdXGDIB0VksqvwAnfWipBvPkZe/
mkDmU8vG8HMxFZup7c0aAEFgLEc4V4q/gcGyzNUApLI3GFYQDt9DIbtRED915qEe
y0TKBEFvr+RyhhqbpH5kKtrEuO3Uq6+mh6BXHbsV56LS+Q2ADLHFp4gEo2uglynL
UyKNqlE/bkwp3vfDkeamoHE+3Pe6aNc1F314XczCDf1g/4h/vWcEZ6dHi1Q71tIo
1L7jImjPOh97dP0Pt5B04Q9p5cPgeShr4DH37TtHe2mNAD8NxZhosaLMWzAhWicL
6TqGQyNfJAa8tTC8858DoVsu00fMvi1AzXlx+MI1LU3oldjio4Hcq3106Ly5O5Hr
hnAf1m6oibRGivJIU4K/WYTn0u0R4hk0eV29XtvUAzyyOpk9XAb7EeqjFdDwUxp0
S+E3Y9eZ4sEVD/n+LrhdZmq+o/zCZ26GPOenyizwqdGjeScNwVSrKx9Yy5HUDExo
E45OJiONOVuvoJvyNvbzreh+uf4bc3rkno7LLpW3ALp7qk5powF5WbKdeoNx9tu0
GCq1P0YHOMWXZ9r5rkvL1o7fU75Xmnv3iCnPVeb2RT9SPqZ1GdVG/OKNEr3WpAt/
tivc4Ff29skphGFL6WdW5Hiu7UKWW5J3GZsUwbm6+zpEJDgCl4ygyqOeshnidoHg
2B2dqstDB3Q/r+BQst1gBjB4R/F0HS7PwSWHnR55ySKKxl23PwSCkj3j5OpoiYJ+
ra+ZlxquWHJeaafb+jzoqQ==

`pragma protect end_protected

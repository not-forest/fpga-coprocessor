`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bEfUSD7v54Aqz9jHXOKP+ddRUoKCowCki6okHI4laIFSgFxAARWjGggLR2GwH/VP
bZmrbQoQfB5XKs/EEAovp7bWanPip5Uy6yBVKY8lRUS/X/Dul9zo2zLbJV01hm5j
KTmXPXzHRwB3FX0MHHVLtftcPjVVtAgBJHXPkO5ZjmU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11696)
6mL1pFDnbeI2b3Xu0yjK8NmpZUZUB8OGIVdN83JA4puUXrNl2TgDykfW7JLGAt92
ypMb0GTNusx7WtmyokVekP2uH0opPvZJN9lxcXnHLA0WR+bLjbmW48VwIztxMe/A
mE+HKMb4CCHW3huqkkKfr3KpO3qU+OL16AiORPb1MwLIVtYEgtoz6uf6Hu5yBxgM
rNmHRt+sVqqZfGy8c6nGMDox8dvbSHpWLqH12ssMY5GmLKcgd9/wySyY0CD0d5A6
0aY7al53dFWM3iJXNQ2LugprzqW4tFgfC3Y/b/uErr2eLRruAR8oncpAhT8UdDyZ
El+hBgOMnBWx84Els2mLzzSewjll8ZmzqFUyG0ZOz6Pa2CMnavUSh1vBnjoS1ppU
4Vxm2GFaXEZJLHwy6xmt+DiMIt7lnlB7b7mFP3Q9kphoSFfoZYOKfD/jS8GomK3U
KWTC3P2p7cToer5cBCzrk027Ilaw+3tsZf0NE+9K1FU1M2q+VGq5VtcUB173vIST
9SuQEwew4PX9ZG3rsMtflOPP/nsPwBSpvgn9Z7hUlOiOinNY5BGyrxcIX1sFOhx5
/7r1VC/2Rmkq1jwmb/mOksK9JZl8Lvd1VSc+G/KHWkWtDkLryZfO7R49jVRYRSqH
kuQhOIlBBIDOCUztmWp5rRp4T5IMO+yxI5nZrWrLwugomiRogzSUezpi3NGCj6/w
LA8A8Cda6tK4HJLwX9lbginhHc3P/ITYoBN7GRmdNP+In3f6ugUY4MwWD7jlQ5qm
8fnZo1W8t7mezlAsVYS66IpDDQtfMo/QeUGlgMe+nkn675OiYaRqxbzc12zzVIQe
fWub5GW/LibQXi8MZ84KycCrGN7FR+t45e2iY3LE6EP5n12+SURRvAmO32Bztl1w
aSiSJWE7RFBUVcCHaCar6pPju56y3khUv1PwGzq4x/Uu+rmUVNq5z8C8EFtKWjZf
AsOiGPuz31WXHHZvMhqujWYbR09eiejGZIjR7lNimIsw5s9jjmZz5+YO5T4sIoPv
FrV88GmwiF8b3qu/edJLm1D1Sz+FLTVDtZkz5EC7Ferz9jDG+keYnSQRTEsFnpwU
UnS4s2+nPCmuizdjdW9G5nQQNEKdPxg4ug1hMNLphmdsscVoMsH2FGgY2sQSgdkM
9R3fdq7azvUu6eMIRqV8pi4lVMWZMlj4CYrMum1aucqGXuJ1a0nifHbSWzjdtXRC
sw9zTnNkxkLM7cQwOo3iTX8Ha7DQpxJv7MAzSMi6EJyWhgicf3u1YhPJJyURkutx
e6PTszoPpUFjjbfBsIQKikYzqiL+JPEdaIv9hgqq3sbpHLCATe0zZQj1ffAAkHEi
/c05WS3xyCYc8ypjTsCk/l3MeQe4V37qfHkYWxM3W4f3HOpIv1Eng2i460QtqiN1
4eqhQdH3y4xElIfFt2n+N52lHL2YcwzpX+W7cj9fRiIzzzw/IVJOQQYdawDOZPsU
Lbwdx1tHQpdVFVfXJ5qfGjnJNAmjESfQhM/KyPfl9IWWIhbRn9Eo+0rk367PhGtB
YxUaerdiT4tnF1Ry706iZHYcMSfx5rmsSFVSE16ZdfsP7hM8FuMC3771hVO08DU6
hz7ih1Zhr0BIT6JCjIHh0TqZCYtnBC8Q2Qh6wh2gtyiVFR7ce2LlTbgMjpOzUEVW
wv17YqCMWhWAlFCCeLrmYthrmZib3in5e1Q5yIcnfUIqhHdsfZytM47M8SB9mQQQ
epmCQ82kl9NNz4eaRgWARB2GfNXAPcwXG3BffiFwRk8mu1Cp5OkATrCM3HvGNBUY
4t+gwTq3ohXXRjJVWp/xTcqls7HA8klgR4qd3MjgBrrYFPhW46tfgei6SXNl7d1q
uQRCdc+ZtPLUP7kGNU2tjtzhIzNKxQu2ijHJ175PzBUSYErVv6TlkGAVnNX88TtX
/u8N+se1mNeYznN4dKTsWRy4UVtwH95Wxds/neR6YHtrADHBGJfSgBRRhBk0biEr
UwkCjjGLGfdRZbd5K4C3MkVx+5hj3ABXETijvOamWtSsAyXUBMBOF28A8m1mYo4n
2KSUlIgu0JOb6zf/jk+u6u/lGj55dOd8d8dCiaPg4no9O6uhETp3rBOytoxu+JvQ
E1A87RCj6tgyFYM1cuYIg4VUpcjIHTT7P9Jzubd1BdS13obqXzJsNCIeBC3mCeGA
uKZ5uY9+7Ihf0JpchEbwyLvgJO+ATGECzBrwdVVUUVCEIoFwEhhVP2PfPBsCKq6m
N3QftKqXB/yjHzn32uTSoZVInc0eJyvcl4/hWv70n1YzWM6CDDPuRds0ioIDLbf8
XRuEQPg9RpULOG595uHIiuLmZ6/tDigoB5OoSNO+5/Nf17sU4QYQ/etYTUcs8ZhA
i5tq29J5uuWDzKJ4J4Hele3Q4idGAouJlSdqcp59nyp8568B4werZvr7u34d6aTX
1Stywxb8Ua4a9D1SkERbkelLXfoD+W2MXBue3bC+zVQtlNUJ1PYHdBURKXAG/2Yk
0wj5WZDBT11JcQnEdkkJRGWNFmAOmA5xFGyCn0gUdvtMoiHP83YaEgysK4CBizDH
hIi0fHOJE1cbnsDCbmCb18Kadf8Y0Sy1wwUtO77ipGGoP4AEz8TWac1Q3sWj0KB3
0gVwIBfT34tsfB13kvCOcYKBGOe9fL2etzzYRBzU3EIkuNV5g+EZpgu6UOr8lFbx
FI6b9vdyNgSHXNmbqdKLW0ZBStJRqzZ7SAFG1fd2qHkQwxyD8Xv0u8bYwIFrGoXR
xStEUBdDVDMn//b0y0IVOJOBp1DHZKWYKPfAJIqlfsV2qFZ33rJcVUacY2hjs4pr
zQahguG81VJd0O6uZ2hhAdDEh4Mny9fe0Br3NoBNjVYiKju6G83n5fUjbOAYKA2b
YTY/tircbFUj3Uy+SVS6lUJm/8xwDvQVCHP7J6MbGKWinKnzPriw9cFTdjv2qbRT
PZI7DI8uBsJlKS6N+YfJG2Oor3ZcHRgBgbCBsk/s7Hkj1QMDZryuyBMtJgCovrUu
i4JjM8QJq1imluYXGeFpcTAYLJT9BN53fpYcMBfCiVNWZiuUT074UlqG92NBGqMo
1SS5zqeY1+afKuhcFE/obPy4OVOaq8PbQKXqR4ECV4/FEmQkPriHwpMIWmyjEuR6
84XDEOY6yPapOewoBprDkHoCqMRHhs7AhjZzfVFyYOsJ/5T6qYPrwIuvkTPk0NEu
qzXZq5Y6AKZEumAC43z2XjR6TJ+35qLsPQLVWxIeWl9WQynw+CMfrtHJdl7iUPpX
hWuwURJZ68k7ZxdkXNwuYInoIgrrwJBTHRGblFQyiTQ6r1pIheoQpBOT6IjEJ2Js
68f4vM4yjHRP/lstdekOatZMDF2+o4s3Ww7tzS0z69komg19McoyWtP1NVXhXSCL
S3Ce9o4C2tXN2NeQfUDEfYoApfsAGWSyy0r2xRT3dMt4ncsa0gVaYif07c8fzQpP
tSV37RwOqHRkqKox++aVzRwW2IigtWZUxlWewjjCYHGtKUJJe1YfjfftG8VPgGmn
eJHcvL4wjU9HQKBlj3Nl3vmoseNb8EKWK+9W3xBLxVBBqpwgDbHhzsf1zZBPjul+
IBRFl1dGKBeUorDFDmxmnQj/PLnuplwdxR+xKzM0B3ap3DofwFEjjumOv/MGyuJg
EE4Agd59Ug9eR3yrAs9CofB9sitht/e+/oRkxGizJNU4WNmNPu8FV1K4bKoo8bIX
ZPnkT5iffBDZM9GSrNcH2/V26BlQUJ0A1+1Wt9Jlj9BXflftxlR20H2MEGgg/wPH
oyxOrwcG420pcnBXZQtLMWyNI+671xejpcCeEj0F6IgGdHwIOqxR2jp+UEVlvrO/
H3B09BcmmMJymXTSisHWz8lXyj/iU0KlyDfo2uM6lyC+vJCYqS6BUM5tC6k3z9NA
Zv2Pg077yce85cNMGXyc/mckGftKB1hS4b1+tH6nThZ7cZNctbiwSxbos+aRtAGT
MCMqUhpJsPsCQJP/wOWVxw+PbdHzMunruP3J9d9Zl7BcxW1aLaoUoyCd3r0i5852
UZTFvc9xV+IrwjZQxnExX94iUjNGQM9HvoN43M1r8NtHyBg7bhcecpChJUsv/57L
u8ZKhSjLMIEg4MlkMwXaIoGUbEBBqiDuV+EcA7vfnNymINxWizughOnBGTcw++BT
45/yuccmK8mOITsATBoBUNMTGZy73PxyoiSdyAn7i33Y9DZz977dBdV/57q8E6vJ
bog5PoerPrMK74+w3UbGJtIdKZc67BHuQdUcdjA92sLKdqT7/xD4pH7Ag6lTDiIl
z32dTsgvhxiGwJlO6JTeDPJe3p2aqcRy77RujOd2AGcOzmf0s/ndMt482hvRDwjk
71KZ4YHVvPEoB6pVmZj2Ly0mWpUZYGpmVwaE9QltesV1E/nGcO+YZ+tfbCM7w2+C
/Bq4dysYYuzA1/nJMjhKuFux+fzyb5Z0BG8eczFzYNaRTSWgoDbVRe8O/2Fumcl/
l+hvMNvB4pf+IPShD+W04jBXPBWYX3MFCl8nJzTCyaCk2XGO3LeC6VmduJqYHF3N
a2yr5Tj8BI533zbZ+oQB2pj5mQutjG7qk36PfHE6wap8tSDUU1k7QdZmXLpD98vt
KhaquKU8K2S5tMN6euiCB/tgU9M+4+DNu1EAWanDAHRWPMIKbV1I2SxJurHEK9+s
mb5fgG0RLFYP5wOhBd79PXW0eHcNSwl7sdMXh7XFmWNOquSQu8CvNXi3MPdR1583
M5GgBXDx6tlGY2Akb7jZAaH0ZBVeVNNPDSq6qy6a4EmROtyFzsDTeI03n1cXGEQC
/iiuNu/L+Lzyy59q+1AT5iQc7wkM4TtzIxbumy39Ji9VbygPLJc962we82r8Zh71
hIFPPo/cm6jRnn7KAUTJebMuIh0kUYSmYtYMhMeVGWn43hz0/MTWVACsQsVzg8bo
2sDvUdy5G4SXN9HJDtYI2AQfy6UEN/OQv3BxZX0MlynT9uqR4d8f2kLq2UszT+TA
z4uawCjbNPz1fEoQ2lUZw5F+JiQ4/PCMp7feiT+PUINEnsioXdTQzUH3FpVvjsQN
zP0dGmbwRR3YcNVTe8EEV1YMLM6ct5Rok74GsF2gt9oiSQFhpq1SFZAizpMo4Tsi
uVLwBJVFkAfc6la3eh8rK9LmnmcvMvtzVGdWbhAsENZUav7bqbIZrPRGkbUmJtrM
7mEgMDpcMI7L81bt74lqrMp93UY7879m71xR/rEJh2T/Ni/OCIfm4KEXOgf6/1/w
2+roTemsc+QO2OEHh8J5K+fDP58tekDx73hAevbnAyJpz9jk/XWtxgIjt5BMBb3C
YgViqLAn7hC9S525WxtJoGvyLTQPdD9h/ZaoS2LLhe+rfomyM/Xaog6JV+6fK/at
GWyDCWsDKcLVjSQeq/pjnODx5iTekYu6f9SVzuLX0b2Ur/q7lW0r7gA12OqE9DX2
I1Kx2aniog/H8fAxWHz4zBXjqHMK7OoDoBRSJJH5bL2zAvj0Uo20ICm1NwY8jEyS
6oVQop8Z2D0KurR/G/ekL3xhcoCRcqE/xdvNXVg/uysYHUGufPxcpE7NL9qeS+XG
2uayyFgIkq72JprF874cVYoMZJt0o3Ub0w8bWJYYvh4gToc1p4wXbfYTUH3lgUX8
g4gKd4IpQ030NuAquOSjxd9LkahxTpuxkgF/NM6PgqzD/bGrPU4bMmdk6sJf3w3h
f4T3iZBqusLoNYRzT189e5aEoiMdg4RXN3tUy55z0D4KlKbbCtiJiymqlK0BmCoz
J0LX4u+v2cDBJEnzhCxQ7CsLvTOrzDWGpf0C6806i32aChr0yhXwVz7oGgE8SdEx
jCli1Yv04xRVOcyF0bGBB5OmmecaeNBw3wBZYdPntF6FGzlr3n3ohAQTU+WiwcyA
CVoONsul0vm1mU6U5Kc1ELqq/ECgIMkjTTONqiL9LaCNw5ugxHsfz8zRB/OnN1Pi
x3DO2AaRF+obcGbBAAYq0T77L7uTHj2FiXOPC0YlgX8Z4sqvN2KOOq7bzD+pohnx
vH+OLdSINKGihENXOEIQPTXrzjGjMf1V64WwMtCu3mmNC7Dr67ZKCZZR2vXZewDg
WONEtAJSc7cNEBv2wzCGNpj5qB+/i2hK5UsYsLVwcGuMZsMZstAzTflIiQbaVWjb
LqRqkSlZ1SVNeS0w478yizzXaovyoOvFNVqnUeuUTH4z20GyoOPTl6o5WtNeB8dO
DzJzq/JELISh4TjJFnaigCxTCInL7ZG2f37/d7EhttNEVfvukih8iWSBuaOxlQuO
Zhj0wxfye/uY5vSjXaeG34wld1p72sWAlRRl7x/nJCGbUbNWkP2AjQ6d86aHlsoC
cUCGSC1lWQZn9AFSWKhHZ+qjcuigUlM2viUVxw2W1lkhZf2dlhmr8sVFgO6TK6Ke
2sNj6WkDcN1zV0IX0emjEJvz8ChlXu/pgcWotXHcNzcZcE3vX/xZ8ymN4bV7tUSq
VDqgIqFeEa5r/GjqoDUZUbxfgK7IJSqmox372Lusq8EWT/bjtPxGmqJdMt9QaeZX
sElpVUOkSgA3Wzc65oP7Ocq7B/sl+BKF9/z6WzeJF7fJKn+76srzoEpIsAgGm14q
goseYfPP8UShushGDYjGlXvk3ywfKxQ0aemVbH9JbxbQ9V1fZjR5exWbbzOjqW7f
FKl+u5Z5ckoOcZR5s0Go4VxFq6ePLIDbtrunvI3bc+oTy/to5VCqHWAH82E38k49
T4FCtMpnQeSxpvOlyZgI+J/97OlH0QL7fs51nvJ6A99aG/HwxHkqZFI1wd6lGGG/
lqwJ0Phqiw1pAyQ0xIry6donuYE8v/HWkQApumbwVmCqdrMSxscGBB9T4g8l4w9V
BK6+dGWi8qWmQf/7HYLWAKhluTHabRZsnNaVEWLuPxxRgbj/xMYA3vVbjnswE3I/
s9XSnz0+IVR6ILL0LL2fX83Hp9JI789Ws6aEDyowY09Q6NLhp9G3fJc7PdMkwsuF
j20Pn4fqqMl7iAVdpKtZA07I0TgWAjDwidy0I6w4PVFF5/3fr9gWqAR+4Qzb6Rbz
FSZJS6ydujKuiIEBNv07f5+7w+7irZ/M7Gf3znwOUXuZdTqF8i1WaQ+iXJsVQ4G1
5zp8M8YaRtysdYwcebg5IPBIGxQ4BkER4NAZYmCX/ttAkSrWx9UHETuMpfWoYJaM
0jQ47ln5Jpf7qGBUbaaUysbyb2+Ox4uYFuNZ/RF7ituK64SmDLJrBs36vyG33jYu
W5InUSb5b0nTKpjcgw2wHpapeEjXfqnnAYlCoX4PhMAEzy0Su+/2jDWR9ifw79rV
29F9bmSeG6BBPbQNSs+TWBIDxBoZJcUYBZT9mb8A9PEdmWGoCNJJBnJgJrRqui8J
8wEKQUdUxe4DAq2qWDY/PV+A5qQFDB+5Z5V8y1byzES7BVoDq1715ws3Ub/JOVga
AwOoAcyStuSKcD2bgq9FKN3h23h4jpyjmcFTPjcbq++3f+tFFa0UqJl0uKCrjQ4L
0t41FarhtK3IclGnYQxzsEKYDnbk/NjVcDMvuv3sjqSzDbBVdgxAG6PfXlp0jmC7
QaQKbBTzERC/BcdsfMxUJjs9B6r/CjbsQv/DTvPM3p/bHnSB5kwEgol+eUuobd+T
AqnotuuefTIOXDGYbIW42r2o+wtAe1QfJ54KPe0sq+CYZSuN2Hg4awuOBaf1dAG/
wsRKkiwT7djDwHg6GhQYpZtzNJm8L5MNgFi+xSRr9kUQWDXLcYz8WdpeRAW5rQ6a
lBnRe/Vn9u03K/2Y5kM4YjpxJja1Lc2y3n9g3YWQXYgYCZe04uIv8N+V5WTT7yui
UpzVgaYQzvPdFyW+Z8N2kbum5Nbok+TfVIBsxPo91uakCdBkaHLj/VyQuQftOGLE
8Yw340rjfm3W49nr7gx4Ho3m5nZAoOXRw4t19HsX8GnERUIWwvwmRvC15LMWvocl
wdUQr+SpICYXXWSVqfflC8Fu/w8MaTn8zEzwYg1KdPsXGPk+hbxv1Sml3+iKhpaV
wjDzE9DU+SNN9eaLPMF7X1FmW5bSlRbGPbxtVAz2dp/cR1Bht2v/W87usVEBX05s
w3KYmViEXWK9DoF42V/l2lJ+sIID6szsouC0kiO/NrWGtB8kcMc2ze9CV7KCjj1+
PFL1mjAx/foBwkGhjaBefGvyzGNJJSF5ZVC63WkNRwiIrqnBPkuHt/dj2mYin0HH
+d1QXiY3/lqfxGzMVsg1bl5SPnKMAXpJZDRVavaQlQIo2tEdJSx9bnY7lSQ5LGuO
J4ZDdb9m6Y2NjjNiv3xn9z37AF1V2IUhTLQlxjCKOGVL6fvGFnNywyjsdD711Nk3
r3bso1OBjIBrdrKBAUAQAF5WgPYZTkNlc6cnwgqFvZ05vvKAg+ScXOvEgiPuOWUw
aYQC68ylaKyylKNr+FKB8hnVeo3RrGsZ76/7ue9iBaVxh3bsAHX6P6SzY8qzxSja
kkI4uoK9Rw6zDbDLRly7RUi6btia2vUp08PQh9d2n8PavNIwH+/JoVhTpxdZkZnS
86ldgQ7qrOs6f8N7q4LrLbTR9p+fFtuRY+GTlbuWRzgsh50LIbnrptL/PF74a4jf
VK7Z/Rkj5lTAyHbAIQeBMG5mTkoElckqoRAW7rW/N1YRfYP5Fh9+MoaPKq25NDID
l3X55TmnS0rOuXE6s4pPSEUehQGbZiXrqKNwTM+EPKtmGh+D/WmU5RCfNM3E4oJk
DXFAcPCbVml2rOpSSxaoSny4z0IYTsXeI+dtH/yAOgs+UbgGqfIIp0vDLT9O8pFw
hS8+8LJA9FNkbMbeleGHIRZuPC2L4MYeDRnOFayaHdJxsgN1hoWKg1nr6JlaDsF5
2LsCjmHIgn4CZA6sb4rWGcQI3vKxAvr/gbcCiYCgwcGfapEbLx71bG+Molj3EnOS
Fu6n+OjYzopHiL0MCBmc73qN0bxdfGSEZe/3YtG8kjU/RzXmIR0Jmf+xrlSp64/s
jO5aVHZ9vR0OtS6RsnYvncwYVEVPGdHvFhjuqyXLaxX7Pds62k8VP5di0FAoawjU
xGPTuKmUpPoaiJqgZRd8oDOaPiiecTQUbtwqmEG4IJ3PIO6nyujwim28c59nBpcD
+ySiBqIIfz/9AALUt8pNkVSwBUFWUQqiOAxZeAS88hS0HQzZ0J+ZvQTBgvp+OaCq
KR/gWOMOe7afhmGhti3pX9bt+P/o0no/Gf6sUtMPto9xTXIp65gkQUpjbw+3Drjy
gEOsuWC7K/OD5uMOWmC7lg3NimiQTKXhQk0cbCZlQyvvKpLPvTf3/oJ4WWzmrHWz
UeoL/aNaJy+luZW00xnuEhqfEKIiSpdBSUlT8cAJJkA8MxjEOVREQpzItBQrVDsi
IMFAsYBo9YGX5IIrvJgDaSNnalyv8HXRBofaHsqM7n4bDO3M+HCYemmMx4hJB9oQ
MIgAWIIc+196T/QHBD4IgkZw3beW8kqeGuV9UnAgnbUNNHdad8KYB3Rz71b0v5Hb
jTfPpYoY1PNSQbjWJIkihB9Xs4R61K69FeFgwILuLG437h21QcSz+4woEUNsIHTp
/GI+BCz4UoRJz1bwf7WzuBzxBRk/fTyq4QUOA+KYWE8SvIEv5qRNwLs0xTE87NVB
39PyE5r9ZDanaxGUt5EB/Ew3Hmsv0Uupv3+ft13yHh2mcfpknWr7fI8swFZ02bvB
UgkuUBjq7KmUxncPXWFYUhOU841DihDGx1IeblnTkGE13HHESdnYuUGqfUQ5H95S
7lNJT6QuD18bSPyN0YR/k74ohXahHrcYqUzOwp2KrfJgqGqmmV9qmiG1QL4UTLKd
D7Mx/LFuv74Sr1S9w4XWqnFPhAnuKt+W64uV79yf6GpKLrSfWwqkyTViwkLtxKtO
DlY/pE2II5CRe/TfAznVZsK+FZH2GzqjRkO/CLA4akHa1GFjAiVbDivuVCE/WJEL
Fy6noJVA2ZZ2F0ilmJU3VuTDkdzFaLa2yqV/V1XLh6X8kzBycxaKmexVB1JE7yP1
zTFQV+ccdBcNoCJUtfUBIQ+4URB483x/rlEl/okmmoEciUWkIj4riS8pcqGQTmUr
9H5LDvsMnxElWpz1ZuacmCJpC8E5JfvqRoxG5xZbNeEmkgBrqF6/4lWMMIWOjboj
XzTILwFpZlA+MRnEI4ZKsmvCuLD+HbOLNqVGo240Rpi8uC0EvC6ZyBLVqqrOgn9J
T44EbZw91YnRz5Jo6qIdAI4bxZKalJ0VC8LPmwFi3f4Jd5+7LFfWFmgZEYoJFydP
2NF525PaMiPhgw6Zg+1ginY6DyNzbwEgeNnzvdgQZX8692QNug5hdkiXeqX5X2Hf
8vAZIH7cTa3brp16H9FdBUy66mtGZK/oHEX0AQS5N2kLX2TGlsixnBGOkN26AvMR
njR57LjG7L9fDaO+enkghpThhPKCX4MhHVrN3JN2zhLZbDhxWry9ytJ0Xia0SsMy
wIMyp31gJk/xo41UCr2ypzIx8m8pOITBRdfqWiqBLmoYPCBwET6aldhXkNen9KxQ
kqPt5AZyviRxbur60SUFQiDNnk0EKTmoUULQJycNZprKlHKFz7scus9b7oj5Ihbx
ozK32DX+1jkCStKvoEM5dzCbkeAtTg9m9LOoaQxbZqsE8bePqgzWbnrq+VHRWTE5
NERZFjAUVhthV1JYaAoSVNl7sfGtJ6DmmlhmfwoQvjDbwZ2bN4JsZ3cdu77LSy7I
4K+PMdgHwbNe/Ro/9NU756S1rOrIySyChAbia5tMFbHf8cDZqBE0HRsjHGMTnFjW
4MwEZm9p3uFEAEWIFaO6JIfnrbUdoVe36n5j4njz4xbC9el4eusWEIcUw4nUKV4t
ulAEFYI5ASaUec1Vf+eFeV40a+Gp07awtldomCDlg8YOhBW+02Dxtdg6wpMUvxJR
Vx4j9q2QFq4pUYbglN51L1ITtteBKIIPensYCNPWhoMVw4ZfFgDsSCSVHnuHRAes
6K9Ox7jwfgKg+OMSAzdlsTwUhH2u6dKSaL1jqoAeVt/egePoKilLcIsVZOLnprP4
RDrzoUZ3/k8aaQYjXdxi129gQrl59vM4MyGV5RltNu/R5FFGgOanZ0j38CgmgfvR
qeL5eHtD1B7ZYRPVMjV+4KrVAnsalygIiED04TXNqsd6iK++bgMA8ou4iWewaP5X
jHWs5pbTWN/TJSp9OdfwgXKUj3zgKBSoORrVjejeFT9AC2fKbWh1dJxWmzaKLVD+
ByyqtHwRByPXdt1Yc9MAf6bjYOFcBhTq3DQNucBzoQmLWxZiKmHKqjicHHjZs7TZ
Bj0ZTfT/pRtms3Jvd7agGC+IIHoKXf5+cILQzEXvDhYzo4M/AjD3v8iqhJ5BuzZi
2+7lYrne9kJMr7r4kiBm/MGcahX/HZ5bTo9skV+/+PK/7kXV2+pww2KFGl14GFpJ
TjW87dk273bTMZytfx5c4j5RFuX6dm+h8kWFkVSQ945y7pyM75lbJb9jSoTqSW0y
9GI3fbIlr7O0tQTAaUNBqmFKM4bzEeH0g3S/1QPeIaySaDFfgS/9hqTcTcF05joI
esZAhtiQyUxh9roJ3f5plJCzNepVJ51PNJcGPQ6AixL5auEUGlMOxQFkqQtW9Wkt
rHcJouD6rPmOyl0amsOH+oj2Lqz+wb79xOSw7H5BirB7Qyyrg8VwzlragXVm/q1A
ysd1F8QWYOYp+RzyjO8JhONxfVmjnRirNugEr1z3HW6KiRDaHCqwSNRdKAe/W7Ru
lqRY3cYDFHixrKDbCCrV8kB5Zdyc5vrCBSv8KbxRdSXFxuOP3BSInQs34XGkuGBz
nMBAE65g81QHQCqm7zJEiFOBENjSP+ebQxC2BN+DXopFlhN7T9FaUQjbuxmgNGSh
orA4EDvg5NNlRYHQgRR0kaQDOYkyMHS89L8Hv+ppd9cRXPT3aGcmIAeZ4nx3We8X
pzzu5gNDtx2xJ+ZIDSuExIe0Wpu8Uzm2Yc3yvxoJeJP1Egzg0Vn8Z4aTr8LBmCJw
qfzBrMnysmJXG+h1Wb6slk8gPV4Rz2+TYpMCNejYGuVP1DOO81Rnjb4MCX17xoEI
/0AmAhAKFZ105xod3WicJX3HHZ9UEX5NzvYoIyGM39JTKnaHfBAbOz+0eRjLTlwT
dccNHOY+n5Uz3PHP2ZloexoJlgoLtlkmBsoxKwfE2NBqNWagcnTuWcHT0YF40RYt
3WkeYDbK2k+S8ZyXgdiFa0x1rjWxN4MMNE2/QHPl9Lz90forFEc+vTVi5PazyGJD
zqi3z1332Xnct9JMdVzh3HHL8gyEszX343Ua4qPviOvyfaWkUtgw8TVpnd3I+u7m
AOA3XpMGLd0LylO74ITHkssgorYiAV7elD0rqATnLdo+6f6IAEl5G/wbibJ7CeAV
cl/9ZHbEquUKEp08nQdYDeFqgsR4PJE8K0ArgYafzDMTea5cjv17g7wCYi/DWqZY
OPGj3dy2Zwmm8aDR0H7GYDyKIAmXoFspZYkfIZReis5D7naAuFHcLNTPOgPmI28Y
qCbE7Jj/dYOskyz01pC0MEGSHxjVtAn0r9lbwS1+WAV+WE9jvDJl1zvLnt2v5Kqw
EhJ4JnwpE4FRffRJU/pk7PknN1z7mgvqGIJ7xxVAZyG15+1QQ5z+ZuN2//O++bme
wTX5WzzcIxKPXD1mxBdzYlk7cHizD7A5ylpv9UQf5pGK71AalGiJY3e/ROIcSNDZ
CXDMVxY4l/hBcTa4gBGVRrFrEsZNv8+Gjvf+OFuMCi6odmmhI1yUHA2h53bkwfGZ
LG19VsjYSwCcth8Mws0P9ZN5BWijMvMXEHKHX/Iun0zKc83ymBa9qgr1WDSvGzNO
FF+SxRjD4baeptW5PageV7PRhrMXSrlssR/U6eJAhE7MSujO3BH449vciuD85eil
gHztTTj5VFVYjegLFG+I7cgBxoGm62eKWLQSh3Kzb43UJL3VenkoGXGy0On2BXdZ
ZSbPCOfBzDIuEFOATCPHfX8mID6O83QpZebAjtXykCJqsguHjSRWjtTVUpVhBT6A
OmTL3FKsQeBRnY+jZBLCStBcyInQiOXQ0aKmULq4Hsyr8vmY2gXqZpGf7VKeHSun
+6MQsQstKiuhG/LUxjY7w5sTN6XMtdNzV3tDoYG2n6qrVxUaz1aeqYRi96r2fsO6
Ar/X2rux4kdFQJc54Y5FpXJnyoYdUj7Pr5ZyjEn7qItrURXTgBsWNJTkmRYriAVS
n4vWi0ey9lZphJdNI932goEGSLkzqwDMp/GXi7WFB5/cpbm4JEqtM+g3l7xwVbn9
Wq9gLnRCAjrZ0g1a3HlbYDqqKfzY9AIp89HWz6GMwE1w5ffcsBaTLOYDYrLXXYTA
68P3E0PchhhYHKZM56w9ntds/3EFD0On45na5b/mnylHM/g5sR47UC+3xDbeSuQz
Xaov9hBIlLO0Ju1moetSsrqZ+uC9W83o6e2C7MVCvNIwOvCAfLCogaAfGLDzotJY
auDVBDEwP+/Ed0Bwl703Q64usX9l/ZXtkFP4x0m9+Ak6LVdIIxeI2C7y256kBdmT
7UNiJaj68xFtPLazX3lTaQTC4o/q4E4GB9UeDtKfwzqWaJDvCpbUQ64xY1H0tgGn
/mghcQf8WOuUIp7iPffP/CZR+ZoRRSnVGK1pDFFJUbiCwtCX1jSg+8sT5hzhUoK+
M6rmUPm5lWPfVDXLfv5v6oC2XAxfPVE87r1UGzpO48TS084o8MrlbJ8cXgWGh8mR
/6AyNCyM5dKNsqWoh9Lbzt2NFh3uAOjbMD6YdeXyP+id00gJrFkF5ZJoPWcCcMsB
Gc9rTTS0Z88WzJjn+3h0lvbwc6mLfunlYB4uivO5Zm2S8OHVjW33dH6PDJYD2MGf
SkahvNtMVLzMLrmzSiEuXsBV1yjtEZN2g6FH3/b5MWzXfDbhV+TDbcMfI66d9Zme
+JONH4gFbUs++lbnzt4yL72sYOTcYkQdp3RqG+3sei3BTan2kuRRIbVWOB1/7uG1
VrRfX7RJmlUcK+q0Ug9UCxKB1KIaWDysNNDnYvTyH15HIHUb/ojvmsVxAU9JXZwi
rA6tHZfJBro0HZ1xg3U7SQThrRC2WzvqRcKPeL97GVIR2wHaVx1s4+OptLipUtGF
xdAkwb7CP+gj8RiCz88T+1UlwtqCKNFpcPgqhKVFr7Xcpa70ArOu/TkHYWoN4ok7
zMlOin11iYQG7cZpjA7xdSSV5cfPtBAbRxMYUqH0gJzHBUWs9F3vW5UXqTxjkY+S
XfMEJB9ivEy5gI2pX5P17iRhP+TUhGn/9sRj9FpBoTtqH4nkhXXTYd4NcjZgUKYx
3NRWL8LmOKD74dHxUGoY/TfPri+8ig8ZljmU3QB5B2N9rfBK20uPYGUHuKPdCCi9
GC5lLeU8mWImDM/O76I5uRwL/86w4lK1ndUrnQHytj2jStaPQ0UP5GA7/GJxeXOf
TPIBqd0wfBzIa3QALaRK+jc8YTyv/7mlfi2R8ehganGfjkFIC1hHxe4836Y2ED5O
ESSto7kZ3biMGg/eVY/mskIGFjCozA1rZqOnlj9zhxdTYANnJopO4LuWBY1g5xMz
9Dh+XEAymsd29PddNX4v9FmGzV3nM0ymN7/PjUcXmrszqrp5KgWb1e6GJEbQWd43
D1UFRAghXoZetmY+A01Q8VMp1SlJcHduwGwfntayjvI/WuDd1AT1yFj9nhEEfqVb
ufRg1OD4+vWlYv7wPh34D5ncRW3duFz+96KURYqo8HFBmczd41kR1FnHZojNKkLw
wUUaUohfSZ0IhFOierNu4+46bELA14pU4GjlAfYspuTCV4vzWcTflCeYl/XAvAKm
RCVbg9h5jo80fPxca7C86tVvODxI0nusPofVkzcte99r6hc5IqesTxfsZX7apl+U
IQuQ8m43qdFIcAh5eSGMFTAEe/6e9gwjulOsOCxfcKbwKiDwISkIyTRNuy/jbpDc
XzCpSA6bJ954ytjCQjZy4XaArBeeZNF02XmP3cr3cJSXUdov3YACnGteFdb/XDSQ
f24yswO+A1OWmW1w6YGON679ouCLsoaTY/b6iv11yv8bjeFtNZ5eH/5SjoMU6Bi6
rBjxGvGsaPCmz1hVdLVyl2jK228yzjADFXfPffrzpjEivH6mLw1kPi1kMSyrLg09
UahhYz7O1tYPcF5Dz/bTbOQMMyaLtTlVKlwrZf0NCRuDpPs4RhXbwvwsvYouDFe+
6t2IL5djANZdLsd3cQhjQWXGRKJJH1fqG+qpi2zPk1PdbkOrCmjjiryNI6Js8IKj
ne4+NSfpULb/OHZvpR8CZt3v3/CyjGyEAmdJh7ykCYNGE9U/d89vEfplciymiLFU
P2oZd5YHHrdaER45J8CKT+Cf9oevXM66e/VR3dq/sT9il3NT2xbYKmwbpqFedDSK
x5s3fnAA3QUCCW1FKI45KjcwoO6YAbFyq46YDuuB9vpyCrA4jqYumz1PCIHKl0Jy
wtqdllgOxOUmUq5VxNn9XDF5kE+ff45hOdFM13+hA01t7EpRHv5KIY7LIzWkXenJ
OHpbbhGGGUGsBml1z39RNiSnT4p2w1VyJVO96Id+d6owKVwV3JxLbzoJQXmT3bG0
I7h4k3qndVUSmEUU/0KvdpxFV4mUB2zAMhTdKBsjVcM=
`pragma protect end_protected

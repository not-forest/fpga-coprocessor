// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
PU/psFFkjDAxwo1xACNLrS6RPgpS2lN/1Rym9Nvv0tBft/slx++Ffg4/l4JqUo4U
ezMaOqFIhk71fZjmQYFz113Z26JtEcKCtwQU1x7eA+t1G8+yAnDQuBtGAKuwr5Iz
tG0RPWZyMIA6DLgf5hmC2mBBBdKYJwzZ/hXbwuGXPaOAWgKAGyPTvAcGuF37skxD
YNOxNuCw69KEehnEH4kPUUJnvLvOM/Ox0myZ+0lBDFNYYQQHVFjd04Lssqm8RsZW
1amdd9XHxhs8rAxAV4SyULPOo4vvVG7Bl5oNoE7bxHiRuShU75B26VojN5GFOH20
1aUOh3GZw6R9g6rMbX/vIQ==
//pragma protect end_key_block
//pragma protect digest_block
3GBNphn7fwJ2A+60gVG9MGqay+Y=
//pragma protect end_digest_block
//pragma protect data_block
CUQScaWYfHdC7bjEfiefGaKHOsDT/PyNyXYaIpySLVLHc2AD23m1RHmObTIXpjsC
gXpifZ+o60BLZ+YMUYBq0S7PMamI0xMcDg7Lun9D3Nf68vqIa1jalybr6l/ke0sY
z3Hwi5w0ifw4mcKbDTqhuIkpmhhZvhUVAj5Uxsh/kE4/kABxi2NRVZV5oGTgvdMY
q6S5LIo9Gj0+pwxI9r7/zkKrHX1lxu+ugRuH24B6UqE001TH2dGNXqX9SefGON+S
/sAlauvldP7RKgIKlwNnQdvyAYmSH2+/P9UEXwaWPBLnkfz4ITzocb2l3lO/Ta8O
h1zDN6nWYtErlujzFQYGMcKLX7aFsGiCetDziuixMPtbg8KxePPtG3lHzn0zr2V5
pxHucdiBbJBGVmGlI7kQjycVWR/vEezs/AWAWLUwCQy9RZY+GrZFc4GOJL7MU2og
nPHVr2PL+15QbkxiFnWKCkDVEzJ73RBeThm4o3wkWlHCFaqjWZ+dBKlP6ADdPDoe
AnfHOG39VzYw0l0LFeEp4yur4M7Zt/23u/YAkwGVW/0kvszzGiYb5LrZdZ0jgWp/
ABjnyOOr51AUDGAtcaXSOC1JE00my0WclDSFWgtZlaSAmpOc2HcCpxwZpdR+hzJH
Vc4B98MK+xCgwz/tlpXNPRLL7WI3JDGEGYoYfqxNAUjoa2eySAqVFHl4NWYSwHx8
SRzhA22TaoAOI7Ew8uyf8LeOx/6jKslr4O3sQFDsijACwuHXW1OUroMfx7XtbtE8
m/QGkCsgTn8KuiGbzEfzzdjp3PfqhJVaQD9zCjPkgVKK1UymBnkbZCCPUbub6IJ5
RZk7YEV+MwoSj3DVFPyaDEAG7gHDnvzP+mxRecYJdZgXWePftGOb1PEfWssc1znp
v5IS7frUbFrBIz0zD84+y1HYz3k7evZUvw+UddsC6oAj7bRMkarWS4zPaZCdBjLU
/VVWZlPf5a1/kpeItGay4nDalQE7hfNXoaNGsNJL0mC8p3VIWUbKDqWWjPbVZ2F2
YrXeiV9bbINYRSQ82eAUV1t8W0BQe8noZGDQWMx7ve59xeD4elXpP43ToVYR3CAS
2mhDNNZVlG4wHyRjti2DGkKN/p2seKJfBbYcAa+AzzVmw1fyFx8lbN/8rnt/6IUS
PllhNzInH8CRf4TVHfBUjqGY9D3CBMmau9phSE5Zwn4X4yzqH5iOghzzY3fsg038
1gGqzbSDUJWAwXuDc6sgZdhCgiMeythKQquqkAAoEyMSTEPqGM0kzs9tghtQH0Dx
FF5XQwvz+ynXRKbMyIp5lpbYfr91WBcstKh0L8a4GPK01L6kbNzhLGgXrHirC7xL
uM2tjklE3nWOcWPbNiuTr1jEUjJ8/uhzgJZI8j08V70dyfdD0xuZCyVcLuTVawcB
WRfShmCRUnv3YHe4w9Y3ZeLMhL89k6I1Ubl+YydfEcSwMuWnGoKhhGZZ59724bcq
t83vYVCAMqG6Gs/vfbZ2Clxdmk2DaOyKxclO2kLiinlEUYoUysv+mychWN6HwRBI
syQiBQHhBPeiQZgD6iPdPC6zJlegz/KEOuLvXKLNZB4BmK8ONX7AOE67kO1iM/vY
oerPc1HM7Rm1OjtoC4Ot6uiT70w1MR+fvTgZA6HVXLHZeqYfdupfnUSP1SOudSnd
77vfQqKpTY/UGx+EsunHa0QSw/8ho4Fs2BOiMLitOmPRWXaB/NZBq26zNBDRz1ui
thUbzPFiBTWW3UM/Ot8Jn+MnXb+g3sY7oUQhU+Tx9oqoAsxmhVii3Di2DNEql8Ij
9TmoQaVWeqt2+Fbk9/mFNipnh5hnnmNTCAlVAXKAfPz6BAcbdcYzZAMSAxMjDSzB
fOMZUDJqFO/q1f+Ojnue4TQzAz3nxDPYl4VpbVEPsL/MCuNCuyRBkJSu4NXFR/ln
jyHa2uAYO5plAYgjaSSwWviVwFoM7GDrr8TDWCJCO7wODDhnauVeGwNA9zmHDBBS
kJJyfjiYqDtsIZrnWrbBH43StX2g1yDdjeN8lbGWA8qHo5jncdEbC6QJaUv1+A+B
cAaLnvSpX4C/je2Q6xinB6gs5qMWYLv6CPwqYc4BcwziPNnKHo3lnAvTCBKxl/jd
n2CBp8xhtUZkqFRc6qn3kDT5duC7DhadC+atu1oLXWBMLHIJB+hGWmYsOdC8h4NN
/C4lQI4hc5D1OfC9+ePpd5WiN1wMAV8NmQqul6vzi2SIUs3BBkEje732Oeg05Mvv
akLYfPAQn1SulKl/K9TWMQef5btibIKoLpxkEWTJ8LaIWrU4YXCTb4Lgu2CQchXN
ddIuyWGAPZ9BNfRckI9tWkvO4Oa67iu8ZFqIPP8pp/ULZbTkKtdBp2Li1eOnzSqX
p3s4xwyH70yy9S9mon2sTQWwMPjntyIQmlQY+u4gMzHs9IGexm0o3tntfQVzxcee
SJs/RlkWEgPMgTF4WfXE87b/KzaT/MkLVOxR5E6d9XDYFVf+AXsMbNY27xNs2muu
+bf75CVULxzcCwd8OYu+vKoS/f/LOT+f1kSrV17SYFbmNWXVIFvsqpmX3DOCW53q
yvWA23YHNKl5j23irJJHjXGq9MBk10a8Qu6zrwfSUEF0QBmtdAONmAHCb6amW12D
nwSm91HogS9ESMhtDFQUaqUA05AwF7iWQyEplItSM/cgGnOt7Uf1kIZ26XxxiTBo
wl6pTvN4ojVNnZe0YIdsLytcfnABvaLaTtR9aUVqL0pDD5k9RvlWqyW9NwZ3H+ai
2oBnNQfW9MzIKYiPrI0KiK7PFcv23SC09c+NX7Q9CkNHFLWFQXG307JXZu8VK4VF
obF5uarjf5ueO+5Pmm4yG3uojA+Qsx7IwkZuuOtJEmh5hDOZ/2CL2rpFM+Vqx83p
puAYmNtbZjXBlI0Mag8mPe7N5laBM/U7mpF0FVtnfNqrEPa2IIsa7CgKMpPzIx5D
dXIS1qZcdRKiBXmhGnyBViIuEqsqY7cW0J1wZDKaJ5fK3Wn6nFAr0pNeyRQWQiBG
ljgHA5lPeSusCndLsSGMm76SXl30U2pLSmQSfKsAWmX7AgVUAwAe/Ocr+FTp2VLV
+V/FRMB8vdxzcDxv9bG9tJyaxYxtMAKp2Ox9W4Fn/QBaFYUxuw3n9s/af86z8j0l
ai1qGBmv8VdBKPEOhUmjqAMQJStwFZ3KuXRmp5MSCW0T+oTPus2NV9r0FP3+xXsp
FisgN/2wuHJY2NipVZ2zLtAFiuA3Us77+jk30ER2albV0nUDeK/tmBnNSkFuueuR
ebeCNuA8Xpq9mroBX/k2gb0uZ8RT/NKRTsAnOGbfI6F1SXSmp+xoHATE3fDvWHj4
bhX85BMZo4epiiOQBSixUx6HB6rTx9zSkka7PuUYmVLhKQjz76YLtEtD01wxcJSs
mJVZ8CmRf8YMQOfgyqClVk8koj1ig3NEgBM5R6sOcjZ4mCvafw34gCziBoCLm8Xo
rGkhmWnoOt1w134PQ17gTtR/vPW5U4xAr0LOgeum1B1dORradETaN266c0Q4HlLt
RaMtkPvv6MXYVshYlJ2rB8b/FUfyPjidZL4StQQhgl6gvjFuijHhVE4e06Q+3CJL
HZOJQhgEMmykjfpmUlGWY5sa59fkY+EVDNT29yrySA4TnPMns+ULNH8F1oeZbvUM
7AeLHI4N9T78Rr7TtKybtJjFltYpDefcniusgDCY5oof1nV9UauztKfyoIGuZfd2
OKmlM7ZD6ageOhfvsKP5PcLUp6Eaz6NRyYN2J61ZoQUYI8yVzOAWIMo+1bpdQR30
+KP09y6rOiGB7l0MOZTypNicBZaAsSqbLnBGiTGaTzh6Q4NZxaBzfv9GxHZKdtEp
nnIWO53xgGC9Z8JUC3+FkZmnqSLOdis3qLC3PcLdRySn27NaLtIdutkN//hAou8P
Ms9lXbHrwZN9ATfEzyTzzwaCq5tjGLkBNmyH8FG3VU+a3e0bjl6ZSZg6hFapdya1
3gh/YSCjLjHsmBWy11sCLEXM3sqpPpGUdibNV+OP5C4dbQWQSio9xAnL1ducaMnN
fCZ1Lzn9bKNEcW5PylvVQGqvEJQZHGxtipiqVHc9qDGCGi6DGdLpqakhskH5AYl/
kHSluhwdLTmulJMcTiZ3qOl/YEc+kcyvdOBrrJkxdEfDRVmY9POfBDDmRkFH8HCv
kYRJgYEEwjZT+gbRjMLqbQP/PkORdWtw52p9bfxlEuDqk/+i6q/LRWaSA7pRxaBJ
1Wf6b0fkRBOCkYOSYBO1eA9zU/hl/8EIQV+azAqO3zA5wJAzKFl3XfqYLbVqRIhx
Mwni0MBOMWhUzLXVPuFkPcWdwx9T2hV7+qRJNAahGVD7vE48L8wrYfpcXoJa5t43
zbNAff5LpIXy+qCMBM7b+77CyDDTvqUs8sRSSoWTy25GR2Rem2z1GZANmi1EYxXW
K4NbBPqYjgTsqnft86y2Iu5FGUy325WwCzhhjMCZbCLAvQN7GHpqbOsDyvxyOO45
ApABi+vSpYccXIOV63C21nA9/nMKVdcHnrURcMo6+vrUMhuhwFFm82BP/zZ6IJHj
1Q8ehPUAUrpip31xHjGtSCVd+L1Ha5QrGWTHGIWJWDa5Dew0F0kawUKPiPs1P37Y
Iihnv2BuHOwLyuvLIYubiGMp3sf4Valt7pjrBzB0FCguzpSqlYMZ/TYzU4EyyMPn
ieDhWoMrO+2kaUpoCM5Wmdam52mEx8q02weasnx18YQBCPR3fQyJWeuuA1HrshdK
f+/kdGYEvmA0f1I/3/iY8VcAQOIXeFfN7DDmlOW/57EXCWeUTuJsoZkoCDdjtC3a
bbn6QmLepkEJQ2DBfYsr4TSt0wsqO9uopvsU04RokbYARmsyd7EH2NGs2JSoyuQd
dt0+q0df4Pk9wESS/YQD0HlYpQ/VHU6+ZX9ZOhDWavhTOrun3VwxpXNQbfRseUPD
mHFMyadRHn2Bku5SlcEBaKyZ8aBt1mCDqRxyvGcTwD/UMaUHAoOXXtgBE+43EbeO
f6nynogqyPCNtTVo/VtN3LoEIC64STcc0f5hKqkI7q+IUQYOBQGbfBR6+eUes2V7
yZOHBSETWH/DOioWZfuUQIgeD85zsJXwu2D4I9hbPBog1xhF7evrjU2kykjq/S+Y
Wh9b+WOsBiI4OC5xztfojRrz1XsaXpMuKD/KGArmGWheMDLDOpmbDrnQAwxedKxk
PZt2ACcTAW4Kcv6A5JIdBxO+iVc9+jPmT7wJyclezzdSTHmkqZdmd3dUvkTQ/kor
XUHP5IIPs4fcQBll4PgeTsuqdf76bjsjuQV+BrafpHnZWi0clwMKub1HN28bgIy3
jGi519h0deGx+DAf2lQ8CmIdxVsZxx58wFtOEG0fh2TJ/ax20NbghU5basffNOV4
pjSEwA608xNtCgVIEKsK5QLaTrcSXD7Fw1fu3nB7TOO83LTugKiffQ3bfcav6Uom
CJv0hhSAoBxjNed7ZKARBOJ3l/KNnFa2o++WUrLD2H1SHvt6zcX5A57cZDRmISig
XtfOVNMJz8LonSaf3wzcsiNbNaTn/PunFKkwgm4pX1w2G64VQhgdrBWX8a0C7lR0
qZoTK/xEAEwRqZgIYTV5HqwIPHP/4o5oliqTUGSL7DDrwoxvoNsJivWNbAJqSSk6
OchfgyMS6a2OKChYdxeeF0HbCywEi0FoJQsaojj+UeZVorNIiF11C2XbLqdgYVtI
ohNE1Ik8PeHrkUbSofv66huWSh3BajiI6D8ej2EOHQVw7OYL+CTz12ghI4RZP0vo
78hmhP8N5jcjXs5So6yrY9t+LXFtoLkZstOhzEerX6o0ncAfzrXIEo6w9v87Qweo
8L0RUQM1GxDQYg8zi3fxqEhcpc4ahZ2m7dYqfc6I9jSZpUUEvcCPOmw4J4R1fIjl
5HOI1uPgrFpiAGgFVyguUbDoqb1EVFESqOiCF4HseJmGO3ReQVAZ94uQ23H9vvvs
6EoeNkEybkouQaQKvNd6LJQpZvNyr/XGTfo+iFnzsTxkYwkkxext+c0ARTYFYZg1
tVF0+PRHsFJOkwBfUPJxSXaQnnbYwfqL30wFtyQv2LHYk3OcLnTjzCupEBLW2NR7
rVCiPCoxJOe9udar5q+BIQd8B1HlAVzADPM969ZeaMHm+jQ+xHzbfWC3Kr+Eh7YJ
4858+2T57t61j+q0/S6J/T5hGAITdxfiaButSINcZWwKvhp762wDES4zcGjY7S4t
ZTHlUYSkjVDcPyT1VRnDGzP3cRb4XgqQgxssgdpMvI/xxn5als5RRbsJSk6+Eibc
LJY7LFoWwMEfbX0eYrdlxVEYLs0XIph1UR9pLbG0rZ+XZmg8mh5PDz8DoE0QfFBk
qVRrNiHHmTS052X3PttUNKz72jv/ADVyvIPqaUovh8m0Gon+4Dg+tbrJFO0djO3M
TL+35Im0eD5o5lyhSuUa12LSh8BNPG73YKPiGHHOcZdIaZIjue0X47pqGXvz4dXx
P1e/DJGlUUX8knBaa5fTLVjxAMTk7i1rOKWsV9PFbX7eRHQrTVQzuShoid4bkegp
3t8Z1oYBO/UI6qLMvAFOCyymn9rUip5VmL4+Wp3ICP0H+5pG06DzyXv7aOCCcgSR
rRa/5kkVhQH3uRPgqW9V/vWUqU8wmB6+V7eAJVL5WTT40u0Ukl001kh1oYDexbfz
m1bhrTks2wmn3MwkpD2rjzbj7lpT8J1wdaiRYWnkxKQfOzuu3CPXue1a5OdI/Gv6
FetQYZ59frXyCmor2PJ70H+cg5GoXBK9J6KgM0p1aIooQ+zzOfyByocIR5s1NGrn
0nFAbmdJVrA8S6HlHidvulNRSUCE4dNEdRGCHi+So7zZt3mPgk8DEldWWBTOEEW/
zgFZkp05KMJ0/cl6Np4D9dLp3nlbQMPOhzvWmTITRrSUuMuyKQSRn5kOzMsGJ7WX
G10fQyA+7XW2Iv70CWw5BcEbY50SXp9+NOqtz3MnuSwh2WAX2Ci+ocpwZT5o+gC7
yC+4uR+TKdgsZ1wA9zhrlK6aRLGAmn+g+xFrapolsuH40lPHWU+eW8gwW1ILnBYf
sofaq+zWFlCfiEQ1DeI6ti9XqVbvDn5EPft/y8IXB4/5kdttcFKRi6m/ko2kOfZ3
SnmAbV3itI0jZKVCUOcTHYY1a+a3zBlVH+c9D3pfj2vVHqkRvJXU+1VWsNMX8w72
0IT1UKFgzd5IJxJsE0FMpsDMynGgTAjNRWwQND4UACzoJcvfMoD65p5Lxs2ZIEye
FfyPvOmfQLsF2NeohnX9alAbYi6aUWqh9pw6yTO6f898/TmBnPvYLnmOYmgUZciy
n9QrrbP8+CAWVzGJJ8VGs7DiujoSNEnSmBgeq9Afw20kKyi5j8mKITaEIE9ZBtKY
o91J72Eo8xs95L2hDxAL//WAXltzkGTTN6LSnslXuRjuRmJqd5uBOxXWtkDSPuaN
7H/wKXsa+5SFjlCqYQ2tsBhrilxRBp5RUFqy0OMdoHAO/648zYIErBdDR92hfPdC
zWG7y6ayDdU8gMc0/l6NqOfCArZC7SbgR/HOOUyLzaIv4cMPn1oaIrW/gCiZkA8m
Lu+DRzfCWDlrfwPcNGC8QKg8tc0DvKeuAw/3QI+Bp603vgnL8N4Ec7wCh+a47LC1
Dm7edm0eX/l1z7tcmrmkf4DHFcnGLauv5EC89fhlTzccPh9GNnoNpJrIsx7y7KOz
+S80GwIq1lH/Fsh5pb1TmDCPzh17kQBTc7TWq9BInLwy8CPydZ+fr0lXjOOpRwLk
Xp5/Qq8g1vqRxQ5JQii8+Vmb5YYeJ1I8UiK1EpvXOU0pGAumYuJjg0gYlZhlA5mf
A6veTybq4X9wovC7yW57LiAAIuCbyA07iPIyWL/F65Gi0DX9fAI/YwYl7oRJe+zV
eWBp+FKqtwc/hZAT2aFppwfdcmXqhXr5opYESjCmdjVyIEvoXqNG2hMBjlf97b5x
0arsWsSprUQukGyFNEa3EQWR83UwU5JJsgNOJ035hg8XXJKOXm8Xcn8F4XgaFuYl
dSEqfpj0i2gBxCxZwTOMsYGj8hUmNUPqgWUG6Om4xzIjZ/0JrfQSRnY4StUrv6go
Vafe6G+9pMFxHvHqvNGQK1qLvR2DWiLWY8aTghW2E8kWFDi8Rt10Wb9hQwspG1Hx
5WRhPYzz8Ydbw55g5yNr6OUTnz0bs5/KH2f+gvJ5ZcHJJKeWVCIgNKk5OMSXGELJ
L+sn7qCecaAv4VmQX/H+7y0Sl2tnNSA8N+RQpHm94yN8k1N85iof+zoPz4PwPJcL
fuMYC9xYlMuKmQarGAvvMsz9Jx/8Dt14z26SmsY2sNxabYre+eH16CkLcqdL69mb
dCCoJtg5zeHdlhW8ZHrctzkQVEo7DSvXWyKtdn0ltOdUyeXW3kYgZPQSYdnWO0qV
D/NsMm5Imrjs8Dx8Z+Z8RdDqYVQeivoHhhy1cwQ2tyftO2QjVDVDyuwnVzg+WAJT
mX/kJDF7MP09b418cBEyPsO0Lj3HOltGlzOz54ka9biTZXGxejbYb1pfHRhBAtdt
zDIpPJE7ba8M3yVGubrQKdxydK8QjzpZMpR+t600r7MXKn0ENiVQCpSs3MreboR1
ELUEokEJRkLeMVpizMed931YZoEMzx04eFnq7q3oB41Gm6/bfuO2DnR2bHzIZbUC
05cgBMBxSJc6XqBNkihIiNXvEzAcdtMtjsNxvoC+9pDBjsujD/RBi6c7GXaJeTZF
8pAdjyQte9DsVdo9apqAAr8muY6ylzLTLP1YHgciWX+H/qFewjLAxK31q5ngILBl
+0fUnK1ws5X/BFi1BkbGYYm0w+f9tVaCeAso7VHgim70u4SWEktOn8F2IGf9qwws
FibNtf5tZO638H5XO4XkuySTrYAsnEeK/jB8HB6Fyeg2F7nkiLSYcwpvF4oL8c2Y
4QLRzo818S/l2ElyQKIZVnfTEJjnd2oktOft2ihKsreNCFb7yzzr54tSxTZqknyE
gbQzToJNQtsbzW76K+JU+78TTb6RFb2dD8oZHWiEZk0ZOTq7Uc5JGPn75/4db71Y
wdgqLNb5iDr3WvvP1HkiTqGpGoCGYOJ649l0j/iGfkmXhwqzStdupnYSnQGEPorC
7XUOjcqykO3jTgjEmD+MBHFtc3oPZtvDocCoxbqBEtvG+4WqbAd/PLu6HLyQYDbF
hICmSUReHds7GDzocXywYIE4duAgWkrd0s/lMXa5bVJ61zU0SVHm0oXoLHboKQoe
gKl0NkKzyxgmCFcKo87NsxW0Lj+gZ3pQMmKmUW8E/FiUiHC/p0IXnVuVUYnAK7Tb
gIYfHD3t5reMqP7b9eB0HdAN/2x5LvWHtvJB34e38+ST3Jv51S8D+iTB2Mh9dcXm
eAxr/DKGMsPOnnri219bKxi92oXUgfibbVBKACzyuo9HSnG3WGMKLrrVDSEl14to
Ac4jr4lXMF9TdjfYyrOCvQU9nktNkVobLt4MhsDxkA+Fb+fZFO3HFUYbQmzGFSew
3hCK9GypE2Ss+ZzQBcs7I0Hbt67VWH68pDsK+56J4r1wbGebgtpS+5uzp1iLgKVf
NAnoufEnCsPbWUZwlozbJiDk/h+1WS6D6NJ/SOG0OxPgyMBsr5AcRdxrEY5VI+/W
PVRdB2xjNsq5f/xXMezeT25K21+UnxEkDKaOfAt/EB+WbLIjFGju1aPeo4/ov2PW
Kuyf+r6DVq6yav/kW6zz0jxCIz5iTb/47fwyRoP62RuyoyntAm9NSJfJv8Sp4sWb
sE7hWwUg+TtO8Douo96K6RnHAv+cZivr1RNtMHwGeOcPQYB6p8EGIe04EzYVrcIC
EIvXyTC/riB21pvtYe80KjCQTPcbSn409RD1exN0rG0amPUiWoF7999Hk+OFHmN4
oHwEkfNf2YleQ1Lz6oGI4v2zzjp/HNpcR0GkXrmURy0vqycllQeNlYvN/x5dikgy
9/MZ/TTVWRbuh6B+fVKBSGJcMx0rADxfIpiYIzblbzBP4gnQsVHxcZypnCRYCa3y
lgVpBKqPqRQEeLN5aWgmHDRyH2fUtRvkO4ncKLK9LbhwXsdWLmt/+B12X1Q3LCO5
TbbmudG6GYiLnFeCFenTL2xlp1YflX1QQXKBHkrofYHPV4DWFBjmse5MqkU7iSBU
LNmaRyRaX10E1q82FHlYdeho34nI4VwUXBY1dAxJpKk0IDaLkIP8zwshdvGgg3ip
MH4NZuLYPfwx4QVNXZNqDvl0pDzG0qg5aDG1f79XNVdGeSN5JWdhJK3aWiLWrGCE
h4e3D3EKLF8/nb/A5byBKUTIM/homPY+fpYmpNL3Gmto+Ne40UsQ1p/RA8ACCFSo
geVg5PrWdD9O7RjUj9LkQpi7lenametT08Okucx6mQ1j6VDL7WrGZ8mYYHMH7dPn
MzPpCwzbivpESNfe7LQV04TFq25T3RBFke0yfWwNUueYbtx/4uNQGWWSWwnzCFjD
QLT0dkHknkBQxrjfLeP0DW1RL5Vaqi2RZyNtlSFKwNoC8iK27Ee3ducRIqG79K7c
jY4apzPjILisOgLfbOSffDWyqruDz1s6spT0AYxaRFMZQGliL/XH1Gaz7etE/sWb
1ebpU3RcvCNUhE07cH0RRBJ8Mmma0YULHvzznBekPoQE/K7HJA7F6rItFGAgrISs
AOtjkIOjjRd0REVpz9eG/TT8EAnQYpipjwb6f+Hn6dP4DRos+BwyjEUvwCpN1w0L
Dlc6X+wS238D6PbKoKurJbiC438o+/mhqmUXXCheBwcVOBkOdJEIhtmX1DJlkJxy
bx08zhWyLvdnM2k0dQrrGVk0uXPMykol7YfqibUBqu2gDCOCQ2ed7FpTTteVPlXr
2A5bZeCzyvspZHI8hKYrAGL1VK3vxfruI2EBADpO4rvqY4kjt+rRl0wieR6K/6hP
481fUM59hQCQNRXrG+YhnTdAX58lSPA9P6SJNnqbCc/a9hOGpgPA3LpEErrithU4
/+bJrNLJXDQPsa0OADkjGdebAEYLjlnyvnYqbj0Mp0Y9Fm0OlNcrrV7zct/JAjzM
nfhjcA9Kw4xXoGNG9xEgUTSG6QvfCHCOaIed0sHJdLKhZwu3+ztudEWuuvWLcSLm
FeVSW55Gd2ks4mH7nGXDgGkv57CxjbW51FojAnrguhlyCGvf984wC+mGDx28CCIH
Kwu20JBdZGO+o0bCBH43AgLSqV6JlWkCMktuWxm8bA8alsTCDm4EqShR4izA6Wjb
ENG/ObO9RHOiM5Bh6M7Qz1qhIUkEqaeSnyTzSUZIxKrNXk8Vw3EKHwfXnEx9Bjlz
LunB9rDA5TvRvE5KXXb8N5DY1DsKQAfjOUrQ+37OGX1Hpo0yM6FeWzvMrSLoTHXz
/o6A+MTEWFQAQ0KtzE9rYOs4MjgO3ZcEuEWS8GDo6PFmOXZqaDM7hKG0wpfxH2Zk
dShbzlx7yFLaFmD3nelk9bW02V8WEJBHaE/npV2mjveC7pMyli9uwXbMr0eNCyrZ
OfXjropZdf9HD2XjJPqxSkridAV2GGZ/6Iio08/SLXIAP3wkldpUca8QOMfNSe1R
5u8rUJlnSg+6YmnWbjO051YpeSxEKbLbsE0/BRMh0F+mEGrRl7SV5DxBmQdJernG
x5PQssRUlJ/CgK0Dvn1rscKoTSSb5LGUdpJ1K+dZiZ4XWu8XJo0iwYBBVPmtmMBA
A8kMysNuvgaQCUTbIm/7HSniqav6SsiDObbn/KWcwElHHqpYH2vzf0sR6iaVxgtj
QVUaIrLsaFnnrBJc/M1QN/+RjIPa4UsitIe3JrpaaTP2wgGHfh/fbdvdT36Ju8dC
ypg9JcKSU/A64GuFjRzlcdjftnvzRXkDVp0bBg7sI0ruWh11UX0SGnh0nOE0cx2g
zcSi6yRcE9YWkrPFLsXj9KSO2xNPcOW6C3FFjdU/WjycQaK2l7puLgX6MM4nyojI
oINnbPK5y7SW0x9dfozPNlLJAtf2gW0RMxr3iBrolt8bxr/Xk8wZrOGCGl1W+hUb
mev9GG18wBq2ZrqvkfmCLOX1EBqKcfh23yCDz55KRaQChJH5w/b9wLt0ytwKdDPb
EGxrEO5oi8oCh4X8By5WPgT8HAzd/IX/WBxm1zJdk/YF6OxYtfvdFVOX0CjVJgBM
7FuYOtsQ8T+uOvjIp+FU7hLOJTAd6zxr6ON6piKe5FwSIB72vnaguNH4B+ctmSDH
PLVfA1Vszf154F7OrZ4aswt1rwSOZNIapIBywTfH9QjJgLcPTrNLmxGJTm4ILAXD
Bpx6udDsfIrm9P1CEiys5E5vgWGCzMTlOUp3d6kUyKNLKL0EkP1hEbxYogpaRehK
ICPQrrPPxUNwmORw4Od1H55jk7s8sS08FTrXE6j+PgE95KMuSxUEzTiqyGhaX88S
JjYdqzgcvgEvp6H+dlXfY5QHJ5SoqNc5pfymh6Z5i3RHOxuMvH9IPe+1/cT+uGiR
C2r4Ga6ZkKbZyjfz2NPjJeDbmXjdE7Wb3oJ8g9cHcEl7QwZIB7CxMlZSqmI1lVs8
LxSU4HrDZ8JnhJxaaHNBsgHjpu5Xs6WB7KMR4BN9/KjEvIzPUTIbvAJBQi6iSgGe
KHWf6lBZeKqoAq3zx9/hmcilV0w8I//v0HNE8HqYp+PK7Wva++adIse9sZmJ7obZ
U+MGccFo0C+ZBtEPpMi9d0y9A0hX0lSmGcu8uwCA0dKmK8QMT+FtsnMzJKwv+yzA
2xAQJ5gLhVxrWzuD+iVFxVXbHEWNw0XHkh8+Zj+sMIO0EU92OU1dHXGnDZXUCqKa
mH90xjB1AfBCz3JcvcDnm2haT7KcdQEi28buMgaIqF2LidC9uIMKYg0Jm/kif1CA
0w/07BTCpBVDCURq5BYGwx6D15VQriAXkFEIpSHlbME/xZGUzRV7KT9fyVwYmRVb
Nz0uwkqiO53jOjmCKvrmQwdny7qtLgthM37kaDZPp8bdoZQQvj3kd51Yqih+kgbX
8QHgv3cHZFaitijbRcgt/QRpSpkK0QIKfuc8bPPFLLKgGrYVePNLiv3OhltXlhfS
EkqDGiCaBscojRXd4kr8+kzRRCK+ioBC55v20I+xvLFSnxO3hv90PCcVwI0RtFXs
6IXpYjoUkU0fv2ctsa9xCigQ+TvEi9PKBgtkGqXwL4CGmj5TcTVF7d2uGPFIOkWw
pRAjKT4FKTvp1PEhZ/blaa4/YcwZ7oCY0u34Wl14gDY3otqNYslFIovg5f1HmQ4z
mEDFYBHQ/k6SMYjP4VwYKHgGZ81tZlILlhj2cTn31NT3NZIoElMr1sB9RRaQBJE/
JiSkADwlr+bhXqF6dGsBQ9f/vya8Dkdxx/gnVTC5J6xp4PmhCY1QqEpIzghbjD+I
+4eTsYzzZktlLOKtze7S+FYyjKJUnjmcKN484U5l0Pu/BQE3+sQG5ABfb3B9t1tr
8h1iLfZ55RwdWTHUMhN8WJodm5CNhZqj+RPrmwi+/SixR9BNjdnB9IrZY21D3pqp
I5IYpSeyH2/122PDFa1voNjuSiizamfjBU8V966a5/3zoD/k7B6/kCFyGdN9aTrA
/RoiebRQwXr2FUipL4cAXLw2TPi9BwXh7UnXCz5cq1zXin1LSM/5SE8pFbNi/2iU
5XyXKyPacM7olM8OS270NRy8vb7pOhLC7OBNXLKiK2pXczT/KPNHOZPvD9YkdA4r
7VI8jS7+VCTZNTtLYVYeqNrXd/xsxRrmrL9PYWcd0OJIvko9JMnbzaMSXERzvy9U
f5vNCpIqPyjnl6QE9pPt7PbGO0tRVDWPgG08c6HtSTfz86HpG/dQeg0eQLJc5MTA
ErdK6cLC7q+LpL2QBjZQRKQh/rvhdXojp8KOsITyuIbfso8XCgUaLn8cFqwDYNoq
0mLsn1s6Q9msePS1AZvc/bKEUVKxUxKeE/nblAsga+s19kJLvVewGznpA6R9pDhr
9ab03VhHN4ga2ASgUrOF35/3vCwzolfc0di11aOtyE+S0gj+8qjBzhvU/uA9hvYM
G1od6K64xd/nkGbva/03YQhylT+MIcgbZPDotX9t0uNDh0r3AQwxS4bsdQxIoVK1
oK+Kf09TqUo3PLiI1LxEzL60flbemwhR2KZfQcq7BAlM1IevcxG1S/d85py8NIJc
GfKO4A6PWCFXGVf0py39J76o9HBYyk5pwAE+C9u8fxz7UALLsE8TpjrkXj+MIvki
QLu/E57oeLt3v1N5BJblUw0OYnkLHLVxZi5dANXlJ+HqOClahpU3CsqiA9+w7k7y
mDI/hmM00uXnjd3ait1me979/5uUXdVHZbn8y0ThjvYHCJsSJjwFpRfxLqhLQVOT
C581w5tiXv4WvGX9hmTjEkr7oD+EzQA1x9o3ysHiAW2SaX9wB+mUWqIrdpXl9Tlk
TVNwUgClSaMhJW6GYL4r5wRU6QRN7/RZMZ4HJj2XbiHBRbI2IJ097UjecIbJozw6
JdUfFaA+uCvCQxbSyZSBFvN5FCG8cI0HbjULLz3a9PPD0etnOcRhHsF0Uvlkcgbb
YrX/3+4ToNWbjVVneiGUnMT/SlrrFBnI/9rjohgyBEE7B3sQjwkcfEvMCnUnQSsw
zUMTCM+9Lj2E9qRY9DjtJ6KrDsV3jUtkKzKUAyYhOdue5tdUP3RzvJog+8OagN7n
EE80Bc1AgyTJ4Ar1gnnJmURrYaM2t0bsNVCky/gBz3dQOHPU7B72MLMFeyc2zTMJ
VQ9hL1Ow1lQDV5wJE+jng1YZPkIcSD4lqhpuPM4UQlWHnM9zETBwz9gQlsdkuEfd
+SWPwz20uA1+XVm2NcFeIslFmERYWvW1FCjANnZjO4KvLcn1rPvClaqxqH50+LqX
4I1ZUVl/FxHDqC6pqg0l5bnFXpED88lAVpqaS5Snyg0+Yqauz5YUYo6ln7xryqAE
2ADzI0r4qYlQPEAQXrFWPsLop/0TD9GYzs98BcdPi6ARURsAkxC+n7kIxu5uS6kU
dKFX8BS1FNBYMd8dd6oJfDM8b14UMMupAocpsvK8p2TGc3kOldfEEVQFSCgw0msW
BR64AYCUmevvkpP+PJvwlyrQHbamSiayi+77Pc6Oy2+wU5UfNn/qeKm2QlcnbWSX
RwMjDL+4zwDMkoKgtt8p+Bh8hoF2CH1i8Pqv+N6nJ8otJiuvOajzjMqHKj/3ofB3
GulVVCQeNGh8QfauRMNlia4Pto63H/JOuq3cXZmxN6ObLKWB2VWnE9VGqZvSAxVw
KsutyGAzGdwrbYgiW48YVVryUIPiIVOa9kJ+jmxq7FD1RyOaSBewMae72TYRl855
Q/9jLkdB96FIynN/8HGh0UHgBI8akYSZwjK0TJDSoxsj+mZb35QHSEkD/FLAm2i3
kuGTWgZAEYJiqaogwKl5Y8ZPKOi+BayjRNgLxZCMhbFydJlrGeFMGqmB4FdlnaPH
upwQdJ8GAjNFlohLepnk+OtL/XxJDaFul/pTAhRR+yYsn4sAhJWV9DMkRVy97U0i
qT/rlSjhLRUsdoS1nRJTrrRTyVip4/Rfonn9pNj8X2JWSmbaoE3v/rv3BmaWlCsY
sKu6QuzGCXqQ33Ifi++/DJ3qMXfdgvf6XQfiM9XuEbg8550/cZJ7nIUxeC0oQEYU
CZKAvNIxR5aZZyZZyUPWrV3orc4vPSr7+wbSkydRDZ642WnZ2T1M6cHIhqz3by9a
FkJ+bMRyPLN/rQjGst5yfk5BWjJ6Y6Fixx3U5/MgLC5wkFlKj/rA9pVybI9BtWlj
Xu+1aKTpjZMra7dAP3IHyA0Z1b6Yvitd63VmO4Up483XPOqa9la1j2fH1m3oUG8v
LlF95bLCHvsn2BIAXQ2R4WW0K1VUVGbiS4183vf2PQIiUkRKD0YpT4CNaJC5BT4Q
m3uJdC3NITNp+pehyJOBTUjCdZhP885XblPPB0q3o3JMVUrpzmIZvy3Ij57Fq9SF
cfEfrGPqy5TVVeiC07HRQAd4Eyd9FUzK4gKSBLHzay8IIbDskX4i05MRz8laUjun
3BMUeZonu7mdDiTzbBj75PciHkPIjhp3kI+PegWUEAX7iDvDSaJXp2lTV6zVnpe2
n+r5KEVYByyK3Q1w6Q6UQjn02wLGs9bnBpZPkEnOb9OCSwJIoQtRTWdEV6Fut6V0
JUWD3oPuBXzqxvGrxuqIgKbxyaAKRE0FIRldLdcNPhhy/vTA19r+xQcUkrj9YKEf
7IS9T7TOfihlNv4iBO9cLy1SeTS+RkrfNtmVkYZA9ek2XsRpk+7DqTeGhxV/28Lf
/6ff3eq2KPXMrBVDaxuFzNqEqIlXf8T5Ll6gl+0Q+DkxsxEPc9OEk50MnmNGABCP
A8vJx7ljWmJUDWXc/+yIvQJTvWGY50V7fNgi0HioxnswFEq9tCA7i1w6Ef1wCV4/
jqKbWdHfIfPbzi6ccWLVpXmUX+7AMHqGS6S4dupU0DONEWyjb6Yl6lV8FWsGz2SI
SRZLa8l3BRo1m+X6R9yhVqbv0/k2rNuq5CmxLfbrOpFaTueidtPjVHAX0CmwiTE8
rMdsHPlZPTOm9edj9NQUAdrflt7rlLnyRyzzThmIJ5VNhlA2UPfQd6wMKGQoG8uq
pej6mLYzNtQW9agEKiNYUxi19C+uYtNInUAIwGegaYfYeTjgZikxiSRaR7pelOIz
BYqiEQtpm0MxMgHmJkju5u54GQ6v74D/KIvh3gdKw05mVfoVy/31yhGnvOlrNhG1
PV+wZgj/NMSJK4Topn1ksdm1ugeOuTlIgGuaX/Us1zn3oWQCkQV7/fhIlNEcMycZ
Kt1OD/yMUBB34ox8M4kqvhRAZj6m1/U8W1EZgPSug9NNR2LnBa6RrRopBSeA3ED7
jUT+sUuJAoMbx2pylexh/ZGez3SGVCi1scw9K7cnSOX7uurfmHrIefv7VKAi8UUZ
IRGPKKj0C54E1e5td6pyyOG9SFtGCDMQfaBi2QGhRHBcJWeU9GZkn0al+O4jIo5J
ZKmLsQYcbEVOP3T0ruf43BM0lxDRkGHfl7BePooxQOULfcWZ/sMYk9c6ohFZGfvd
vfP0GrN7SLRbsi47o47PcmMjr5HtsBa9Hz/P3B2vCNoBVbEq24OLaKKsHizcC85e
I/Wmq5hs5soD0ffP5JyMH6MLe3WU6hbMCjqMONafHmwZNEvJ9vU+lYVt8ZU0n1wD
oCC8gIYR2IxXBcdzIbhtmd0cgOxCOb5fm4uV5cvaN2+oGu+M7GPbFt8rF3CRF/0p
ZnHt4hxlqKsNULDuwRBK8bdpxNT+51/O8SSUVV68fe1371Eno02bqtwLNE0TjmX2
NKrhb3y+ZM5OsvOjhmv4/X/CA+N63KzduFyAJ1GICAHfekZpTj10k/unS1irmNH8
KHQmNpMaJeCUY/EZchiWnuV2KlDJ0o+nHki3xz5mKPUxkEnnaWZUnn3XQrO12qgb
xV20mBKZPqij5YdWrlkFuODMVVDgFUt7eZitMT7bWo+U7Y6GMGfFTavFV7aN3FxM
qc/ygi2FzTViq40mAfOaQeo95WvLHZbYiIITw5lvWdGmdIhmDBbactq9UkZiA8K8
nwNinp/VWCUlpVuoaih7mVD5U+GMraWw6ZSRpCrFMEu63TXeU0FY9B7j/iiB7GQk
IQ39hUoOZClSnYlQWpOO2Ak0F24wOWnVeJIIQh91xVNQTfJfd5zj9OkLFW8Ujo5V
waN8Q0FQdUxnC+VgSS5vMxZRjPCaiMjxrC03XUHCsPYtv3tvepMaiRO+IyvvHdN+
I9dUuVGWZtg5YxYkA3Cn1YgD1lGZ0PJBBakGCga1U0pBmPTGRMTMCPvGamut45up
1psgSGhzgN5Jsokmp4j0AUgm+CdBHvB2Dahp5G5A75MCxA/F85uKVIPKYhoEmyJC
7bIubiptVffiGp+DPoqMqfQcdtt0ZfATipl6Rgj9IBN/0rt78tkvwkmRlhxcyFMt
4cKM3EcnZk2+/nTnF8GUgr4oQARQBvanIwu57RC5tICiRoakKne5HK5Dwk6+mFsp
qvdJVZEX5XBjRVXNGBAj8JIH3XFtTlsg9u0vWoJ3apD8F2WuowcdhyEfkTsne4di
xpJLSHSS9OzDETzTdrlRoC/7tI0qQFSv0NZzoHPsouagjuGBM50O4BaTOxrePtrr
fqXyL1cfl9qkl+imYxDKdIznr4cE/t/g85Ypi7zLJcdoRJ/uQm+L7tJrzHIo4VWn
7pFQfwIVsoqN/jw937pDemKmJpPOZDZ7WP8u8VjuYaPgsin1lRFRClmK457BjQBA
scYURt+LH1tc9xQHqvs/VTkNpyAvH26Ms4QxnpCJLPwUNCj/RrHXytj/u1ld0rkn
kBKZdreUm9Pga26XmhhMPzLVP0saSRJoEZZNIWqr3mlraOoMEf9DH9JeDBSELK+a
pKRQL15HCoTRR3Qd6el/rT+l6+MPK9C/ywIh7vOiLN793kdZb0+HGR6J4jwVrwDO
47P9F/q6MivqzGuSRy3hv/vmkzqaPS2DEG7ohJOdZnvCmvEeeVH7ixf+MQS9we0m
JXSC9WfayjHIS+uO4+asplXLPKfU2i9N18jcFNWklIq5i5803VtvghIG3uG7FpYX
tr/QSMXjXev2gcUxfe9kh9mtehq33s2BTreoIKNIe7/FEc1s22bUbzxCPGIL1DoU
2/um3Kr5jt9Fcdrue3QQj/zR1eqcbrC2769EYEVpn7sUNef3qA/ncImNRJLK4aCq
8RUOeXyUandaybsHtFdX4awVfQ5aboYlKNOaR/nD3tFgwgB076dKNDmLEqRlFW7B
YTXGpS5swYlXvA1ZzwhEUjpDYMJHgrVO3XOWUxiDFcxn/7H/5yegLcz+2u7knPal
BwUAmSxpoaAwuyp5LroFU6p29RJWqRNfEZ2RUBLUhVCC7Rv2vx51pkkM9C7vYg62
97+1Lz2KNAF7T19hi2MjOq2D6P5atJxr0ShEatYmCFW3GGuYviRs8BuVxWqkIIQI
QObzCnvomqs7g/ZCem/gwueAl63IMvVhIsufDKtKKArAwMNe5gN3kvTeqc0cRzRs
FTpgVvAAuSaaZDrtgcezOLs6TrjP3UW4W187kXPlN/hzX5HoK+lpACSltJXpRA4M
3VbBsHIMpeOfsu/HpPvSqDUNnFBtsvxO1Y7N8l7zsHjH8AgIhNL7ZY0Md8bXCHAz
7Dj39exqJXBja9iI75cKARIufzq1nOvC3ChbNMUmvzfOgkT/ox/Fpt54906eni3f
kYUtPj5BWGw5E+xeva8N6afQyrPdcGqfUJT0EZbdiWiAJLW3QdPLfaX+R63bG1LL
8JAeVAv7sueBrO+Gjq/VlcvXb3aOmt6mHteTBlkHm0aGFa3g3J0OrCEfWlLgtsS9
HWdMGcNk8TFJ8rKNKA/xlB9LxrcBsA2RZthK1YkB53tqFAy/HK08lij3r+Kq1pam
t6BUDj2svTrNeAKASXfQWfxUsGxEBccCrWn8y5UX8qF7j0AZuamll57jtEvIGQhU
wqB9WsLiERDUGgryNoRmrsEk2hL32UapWKLP390CfEw2jchwLChWczfDgC/BrXRQ
0evXEiF1VHcVDsIL/hbW/5Q560SDXMqBI6nIiaP1vnZ0G5T2rtfOLCiGw1MeZMWT
GinOSX+VLPLHQ2AitAK36lkL9L3ZMYASHClZAyn6anI9/nbgZztUWd5dvROiPvPp
qejokotSYNGRVtNcr7TOTzXvUGwksM1wuKnfCHe/pzeRQvTdPEEYqu21Yu38/TsO
sdliVtoCLZEZcSLPZARFkBIIvjWmFHe7yjk91eNiDrKKg1gcN51co8v5NRoxVCHc
WwDExSxbtAG/lMGfW4dLP0R+0FoH5YASh9KvwqL0zW5qyw+kfZwWi8VpeJpWKPF0
V/vpXsmSuquoFVoX4LW4yUMgdGYrKoLjnxAQL0nx9/Ixlvn2ATZqrPgK6Bszqi+/
hMb65KRrAz2wRyqSUp3zSSAkPkSDI9Y/FFzdIrTP3JruHciaBqnRGOi5rbhKSYw/
CgKk3jEYpJqc1rfHLpyETL/NA091fKfCiFPeiRwWCAxPj+O6mmjL/FbGRST6JSx+
3ChscNsAQEbZZRBLphJ8RspJqq8vdaT/n7x/1RXUPeoLBvILkeEa+xHuoqZcVsbG
CzkkhGJ6mowK1IafbHPS29nRT9TtVQdV7EhBbRSM+T1aWj4CoLXZvmL5xOnwSOU8
4DqjJLFg3vhxWV9WKtQGOaiZe5nRDB04DWCqsvyuOnZx5zUsztiYF4yf5t/74q7M
/6sCVZaLlnrIJUU89FC1gbaDnn9wciA8rNYX3P8GxiYrgNLiYCTmuFVFHTNahQkV
lEfqG82iOB49RgATMcCZPgoVTmBDTh9bxsK6Mn0s69atYidHcW2vhwcN86FL1ZKn
tPP1x5piN7wAZdAmAG4V9hnDrIhXmBsIR7/Yg2U5tBypkf1YYDuil2pyDt10OW1P
ExM+XKcbSRkxAL5DCQslx5nVe2PEGrIMy04oKTNEE6p3e5CS6LNLGM6JHGKZFpWT
DM4zlrIeQVxYL4eoGh91uqbNh91aXpjMRheCmN+j2+RgpKAV1I6stIX3lQ7GArF0
DYAn++SL9LXLABj4RIaLu7rXz3uul+Z4B+rhZAQPafkF1KHeox6PblVjJSyOb6uM
LLeo7s2Wzp+aOIa2Wmt4bCs/SGA4VlIEv5tsM5jyH3E7SpOGNRF54a0qAKrtZPo2
uXfz9QGD10KW6Y+cfzlc/hYRC05hvn+eSZ8dbZvx2LRKPSrmi65dLj01DJqDAfkb
kdOq55xq8AMEuxRMHsFzSSO58EKPUC5857PJMtoXmA1CcZ/Gg0s879XW2SAtQAHJ
kMCe9tPbK3pd0hxRu7MRg8f1bQY3u8cRm5bSnAmr7D6StuC4AEobis+p2Z8GjtOq
us3yRADTAObQ+BnD9pJyBkfxRf+HAEhX5QRtWxWRzpoXSU+s+gGYfS00Zi3vSYvi
MhIlI9HjmEnjzIBJM9BsLBq9XkEHby87xDGXiWIlAOwCLZ31dxGFu1rDYvTGONU8
dcBdAMwF/HgWUiW4v2ceJcY5ZuU76EPYd7ZcuweMHlOtRik/4lGe25FeocdW7w6U
6wU0ncGmnxREOCBAzTzswjCLm73nUP8UaGYYrZZq5qhMDj/Q/rPZn+8M6e3eIPBx
apvjgErdxLMzqRP6HoqwgznP5YOxt+4nf2yqDxLMJ9dzm3bulCH0wK/1x5Gs2Uhr
/nB+2stpE3fuwwfbXiNokYwuWkN9R8PjIefW5w9kdky3YG8ksveQ5g+vVsJ+qgOV
LH8lCQd+wDge1sHGBy/Z+DKVuUpEuRPuCdl7rsYBmd31rTphd+l6f/0mpTOySiTX
PCKQDeYt+NUEdQ4vdw+6wkMUc7L8v2Hc6pGZ7hT6r09BdPAqXiI1B0wPrtBObNkV
3YBs4yioH6uCpfdrGV0eH6KeQ49oyB9A60oEAEkagvE6QyEqPIEV5f04pjlYOP0k
3J1pT8RKuQaDj9T91fYzCnaU2ldnrpV+q5oATCrRyq+JQjQRX3eLXaPYltuO0Hw7
zDHug2LNm00jHGnzmdyIeCs42xHlMWQrnJC8AdiVXReg9IsW3+sL5o3a0Kn8fljO
reDrozcuNSNG3VmPADXlPH50cQUpF8acbibhtRKVlEqku4Pq/0VN+Vg+H9CkkorD
JIPB8tRiFIYpj+dlTgN7yUXcTps6g1np0KxTxmFDklSIEK2OZ7IG9yglVfIy3E/y
bD3D3qg6ri+BMvL82FczKszZJhm3c4S6j+nVoqDENEfwudbUJk3f6YgyvJl4Cfu2
e/yXlQaqftJ90758oRzPzytB9YQuhjbBuJI7h3Dlzijv2y2M24clociSjs+NU5/c
jT6ftPVt6p0pwoFLVIXSqBMSLNdN8RZf0L3fTAdJIgSJichvfGZ0MysPb7j8rM8r
421XAQgXACUZ5uDxrgy8sc0PaCEnZhOtjbnODXTQPqdTsnPKSfwVatCVLaSUKMh8
4QsEjiKnO6yxe3mvwH481oYr4t8XBC+k10XejfNV59N+wE6TEDbkIKK1HADeK9W5
hJPOk+zyTtrvQpVJPDcOKEJqAvtNVp+PktlCbk5UzQHPyhn8xKC/gHtPd3VdvFZW
r5jAo3HtFucKkYMAOPoalH2tx0XiVXXJYeUuclp/g1of3oyKYBtt69ZS6BxluVPl
J7gV8fyj3KSrbbBAg2+TIPnjIXO4sH2k2Vug4Mp/dhAuVO1k5spBs9vGyLfKqM0D
2sbf0NX0HBRGg2IfJ384/7b4bUg94v2rNA/D1lZ3BU8SmcxMyODgA3b3hJZO4jhl
P1d1v7ILTTZ8tTfc+QsDnYl9KHJZ5DIVHTG2uEVC9yuETmUjjM0PG71UI6bYoYmN
X7kjNwqRvN06Y0trsuc5iAueXaiURKpJZvdSPI3Ff2V/i+uDgWSxaaq5S8t/h/A1
RlC8MVW4euL/ge/JHfwRT49dhxXDff4/+8owCR/iqx6r096NhS6EUn60WGaAMI4p
4viFBrEFowxNZgxtQyfoAjP/dvF+PAjupDwfE2hAn/8Yc05C1hycxBzCeh9zucGq
ks0bNL7xzzu9MRwhtazxQHYoNw3rFmIWliYW2Lz8V4+i006Iy4Bea+Krb8qurhii
sCqxFyqcLr7HXDl+APgSDjEcKLN4MxPbKdXd8bVPWU0mh/S7GQ/8uZC2H+OKbWHr
mPnWzMqLhCQ1IBlal3R8k13LEFoTw4y7l7KbMyD6DSSM4YlkFdygcO6vgphTGoHY
JQE/28U84aJCdnGgiJnnE+SiSw0VPDBDZR9up/Tb1bdjHiw+LykJX1sGRwZCz0iu
b39Ts+syuBPKS50hr+WA2ro+TQusVZNbfPMg5zwvRdClEMGkZ012XVkCQpr/gsF6
BQsjPAXg2z3iy8Us9zntmYPXhVt7Wp/7PIT7dMkCMscTNtNSrtu6pvO/7aagPTQU
uGet+Zn79393KOMayAqVeeu2zLS/oA0Qe89SJVDq7Ps49xOiskgoHl8mEKrFW1u2
/Mh0uo/FdqpjcurrKu8+OnXCEZsmsmJF4KUEewaXR+4yQtmEC4YHkwWMcxrV6hdC
6+okztNpj9qYsa/4xsTWYoWEhZiXILFF7wxcBYKaVb6yUgqQF596x9oAXoSyLKvz
L6jNlhFcTxDjdKp1LRwPRAfCs3N1zr95JCiga/Asg4C/kr11x46+gHUhb769Ys8G
WlvEsyAY//Ch43F+RH4jN1Rg88hEAbVgECLe9ALBCM7/1Ep1ZRap4pUceqwcdK9v
WKjSM4sSQrQ1bl5g9n7ASjkvSBqord1/SSWypiTDwnYQhNMoVHoXWXIuQ9k5B9pU
INnygt2mF7TAb5/GgAPwSxJL0RSvfK6gtfcXoW0Dx9+eZy7ONdV53ZGrXG5+tS56
imxmIg5U7ryJIg749GVfC2SRb1L1d5vKohtYf/DOT8bFjvkY08vtnrPliArSsOns
bRE7lFDzsITx5Cj9Tidj6tJBbmCR6WG5WHpZDUZpKc1h7gu0VKYgXhprur36x+pl
tvAuK1DJGL5+NZiZ9EebG2gLjTaxcIxYZrcZbJ2iHMJJweAqf6/3leIU8nGxinbw
czLw6P8+osgkwAeDrtyVIQxg/Gd1rtHK3PIVOnli4/Z/nmtPHqwwGxq1LPLVY/dL
C/6Cnjv/0pFfmQexWQc46WkS35cOffEMl5sv5otA8NgY5EgjtO4+Tbfj1oa4Cpqt
zQoxEBOp4hOhBAH7a6Qh6GDoBK3Pu3FBOWc4Jrocm9LmbGwSq4ueCmvZeskdHVxC
iUJ2VVcQlocQGiu+Cl5OR8WBLxEW5GouPLzaQ9wbRj+7H+dDEDiaUFulWrwSZ7OJ
oUYqCM+RG0jHbK86SeraFCcz0+ughkNpvjaTVCC1QobM0fXcewVDTQ8kbcFQGGMN
AOgMf9ClcnGs8LWeoUBrhzZJyL2F4UQ4Q7P2BfvnoHwN/ZRyErPIOhptBvTSTeg8
h4W9K0NWbXrokoZHOw/zzsxkywMsx7qGZ01FVTiRuqgyJEWYq89CNLD8NluhNEyK
lVJIc2snQ05GkX1U9iUnma+ffuiFSMVSq15F0IEH2UOA2cLgEaLPQPL+H7PgZX+w
z3Fg64tDjCzrQaFz1GRPbip3ASAOXSb9tBPAlWMg7ZbnyTGW9kivjY3yZSR39fg7
YCQhC3+F2RAQTc/7hTjxBCmpg0zAY67l0LYlISQv2CHQGtTA0JFzf4HKT1mlamed
aWxr8vG04xeY9yEs72B2ucbTBwi4vBN8itOzVxvukhq9aqVwvWgOz2w9jsqTE8Sj
1yn6ekiE1N4wBFwI7mOTOK+5HcQYIkpGY/kiX9mZWZ4tWe2lSv6zzEMlK9wKYGVo
I7jT0SAyqK13zyRnSLVo6LmHPeXYz8VCpwGUwMPrE5Bt6rufh9yQO4tn1Ymsow27
sbMUk2UrxuOm5FIgBCOG6Uz5Wo4N51NNxwswtPE9ohHrgmfUzpwFQ5i7rQr4+l0u
oSJgeL5cfjBIqN0M51r1OrzSgZdHDT+yQ7t/yFKQ0k83+VTQ8PkfdER8iIDDt9oL
1rwMFr8dbXOELGMZswbfE2XzWPUzaMaOZ33cAHgdRi6BY5R+ShrtC246DGssYFHl
f+aVKz9v3ZdQphpKF12AYQsUoPetzwdhxAWGFj5icU2RtTXDXjWN8nFxagzqJaCt
hYt5uRmgMBXnQMIfs6MkUU04UrNsJudGyQEBr9HT6tL+LpeDJkxk23brdmIyDFg9
czGqQblUZfci9FpKlK9GubbmrpFPITddCEgEyPyO2xqZEjB2adD44fkkYIdO36pI
qhvBl2ihIWTsR2BpzJ30ZFCOyurghNxeaeBh+0xOhc46I5vpilq8FkU5RKlu6n+N
9MxwHN3CyBWD1d62Squx9v9pe28Wv2HiZkw+XYIPCUJmHE+BS3AOPBN7J8fFSXti
3oqdcTXdkk3OXEdjw7P5uXxS6AbzcaBGB3heKb0Brhz+BtHX+X8607wWHMpZMiea
0yiPvW00AF5yaq9NhOqxPetccqXxDImxhVYdq5VfrhTS8xVNiF3ahErpUuCe+Fo8
VlQuQPBbl8PduYxoIU0gOeAzc9W43d/ckaY2ZQqOkI+9o8RecJRBxWVEydg5JRKk
8oNCB4m8NqCzZd2zG8LgCzT+tvK6VJ93MZVmeqKFAQIbY+6PK5b5RRan5W6Vd/7p
6oS83HB+yYh3ZDIfcKEkaG1KotGtZoEAB4J4vCNc1nI3vMWDGvCcKyv1BEAnt1hC
8S+FA0pNGBYuMjfcHU+3qIACGbltDFq/LXh8rHieAIJ+9loQoxxRwh7kFvaorUY5
nUp2pT+F72DOgePzwkcNN8AtNzrVeWDJonDZ4iJqdVvOnvSZttTCjQmNIR/W8egU
pL/Iogp0UUZA0f5gyDEFkMxvWHzqGCZMxwhT3IuasA2mrULI7M0By/GDdLZG2l2n
s010OPawXY3YRejy/TO+U/hkcan+6S6PcumMJ7gD2WqXdAsMAbEFYg7WeS6riERy
8Sowc5x5pDoxphfetiSPzhs9G3SP9o+I0g915zIgdKdwbP/QumOl9stRaFrvjl9o
xHOhQXOIC9dPw7HCZhnO/qFQZvdlQzajHEN9QYMlaaiuEUrij2DqtTPw6C9mVEGE
bxaHG7onjMcmMFvtfXDc4n2z3EOt9hzmFOHCXcAqumkifhFBPnuHTsIaC4Fz5/bD
9deunj/HRMoxX5dcQ0N1+22NWMAOe5/XD6Ln0/hh4bF5AQxF719zGvDTrI3PoLYG
Pg5S1HPklD0XB2GD1qH/qAA61/qbO0hg/yU08hdyfCkPGh66NjNEw9mxJSaXxl9M
W02uFNif5nvOuI6LYCN7LqJloJUKLnjF+/6y/GstwrumOrn2KHdRn8f6s40x6OWF
sBPD4dAiN9aArsu1jP7opaDR506NfaJd+A8Zmkdw6OlBVoyql7pvLBiVPqNsgkeC
qxuVAS2WxDX2TWb+kKzCHsIP0jsYJfN0xnb3yPSsTCuIIawLfr7j7fv3lTbpzgcG
8OtfwYnpF6CODP+0w40lJ6VqTCEoBB1M66dessUYYfThTtgeOdC7BetVa3m7dTsm
W+IE9LG4a6Sk1L5pSoP9U1lC2zkFbltABbMS7wIajM3/SBCW5o9JMkwng5Tq8X5r
lbgLv+7S/75AeR7RCZlNJFfTRh62H1/c7XM3CcwNy0QJ2jSQMultSYs3CZXaKy2y
CUVkXtNKwzk4JZXjJSk++lZBThHkz/YVt9kSgfqaPFMjvfBTEZoaV2jjIj3j8vTW
MKQmgEa8OXKjBYCAk5En3uxVxJn7mO8lmCEsSAButU3HdSxgYjwMoWaN/neYY7Xi
QUvpKD3yBgiL/7Vs6Jjr+I4ynGSQJFkSywfK2GEvU2/ZCamYGwZGlBqrHj06Qy7Q
Fp09100rR+gzHpzbC182coHBDp4fv710LT0n18Q/Ny8GI/rm2HOlBoMYB6g204dc
VAYX78HVsZ2rrP7hiUgYBKFntORDldlyKwM4UDfuCDoi3VdcqdHp14yHpdQUn15Q
oVuOE5Jak8EBWVynwP6S+qZXq3gSNyOeTGrhWfanw6HThcsI/VO55UMSk1Hx7qwI
gnHHSO3Wf7Q+eCF6PilxuTHiwUY2BImpr3jD855fIEQT8Iz3RNTcZ3KE05KMnxoT
JpyWGgq7Yr2OEqax3XfMNHmJ9KpqV6OBItXTXUgPvkjSGxa6c0i0LZP/jI9j5gSc
Klb+uh7dsIXIJvfE1ziQOmS5ArsQb/R36R1d2XD+KXPpr4EMiBfXAlkm5e3pCHQT
9e7Y1k2A2Fqi5iQPSh7SvZb80+MKNqwtdI4mwQB1Cv3h4yK/6fosU1q4FYVF5tXa
UkNnxuAYdAnfg/eZbIZuIAm05Dz/elV/yMRMRvTVys+5t+NREYUA/pbZOdWQrw89
jys7dH9KngUpzGZr5unaz1YXRUjrrTC4zM78A8nDcUj8jcCxxhech1MJ9xJAWfdJ
LFXJPYvSHrUjFNPvcUYrr9syVc/VdRvK28nOZlY/Xi9XnjA61J60Rig+qJxHYF7c
Q91hL5rEutlB3VwDxwYViEExagNU9kcUXxBeSq0sPNOs0s302gwNTLZVw0t1zVLt
KJJSv/h99NIxloQQbLJYlIZSddvlUo+frav7CQqlVwVUosER9kNruKI0kNnQWLOG
w8ai+mRmmMaBJa8EL314XBXKjxLNeZiptaRi9kvPIPH/2fYOJGalch4gho9D96+Y
7zInv6VRKhD/N+YP8yXRbXoZwrhbnEJuUgCs6kjdZ7/DQmAfQ1FS41cSKOv3SGKG
brOI/H38ywegbq/CbtXCz97WdiJrB6K9kr4VG12rubYc4nwzCEUtFCDUefmKn3An
0Vi9U4MXKOmMUMbzDzWdzj+0GKuVhIoblI3y6RFEehubDGq6UFvCxOJ7dzY/h2wT
a1bzxSvg7r5wZBSo7boOocojPZG0+3SvfpVVbrxFD6jbPUlySzkGtxZfUOjPXEUG
XtrbyWOyy+0Da1yOc8cvtRunuQSH0o9LVD0yAp0XZodDmn6OgoF7nyH5Gwkv6I2r
3F33nM2CJFew9XCAMa4/MOmL50fGwJIRXtTewiZO8mNEdhTr/rPurgZff0UdU/SI
6iDtpb8FgYa0EBcBnRGYq3s8xVy2bJPkRtVAlS2gNBFv6gSO61ex5MH/85EOe4Bw
Zw6NztXRQzhMBvKrbRpOZPIwg94xEmrmjwy5aDo8Bsit53JKP9KTLfqoQE6IbKXy
RN+QwyhWOxT3+ZCJjLi/9Eus6BO8qDtjmESVgpv+0uWrhpE/F9wSzxCnX5oZV7c7
VOD2wBTHQx/yh/zKzmqxGScNFTc6nBpD/kaidyAfyF+g9owvXTgsqFnuyFwyRG0k
dxmU8/yiCmn3aImTIb1LX5nTReW0MQzT+PPFEGUIzhQTT44eNtjYc7ZpqJwoWm7h
9cTRshunM4GWuQGe6Hh0IH6W/JwLJ4RNBWjJD9SS/lYyvptWyd4cV1LEXEdBxz2O
19M3HpuWoR8hKdKkBtOQPOeAkX50IFDwnaGbN/BhP1BLPvik561DESMLwmhA+zEj
KgByPHLMq8KYmK2+1Hlu7ctbwOnICio0+dwtg5x+j42Yl7f8sg8mxYQ/VLOxAfld
uOQMVKyt02TaCKmVfDaZbF4Xntob25cdHBNw38pMimvJOb67YNpTP+FrLVnVghao
t0A4pPhlHxWgOnEzWuXQfW/LL4wA4OwzVMmAQ5bPKTlIMfR+BB7q2bI1NukC4Q/l
Po1k+tZtJkOI02exbDZMpYLCTXiuAIJqI/GcGV92thHRfilCri3phEy+uBqR94jW
qnkyBcwbP/rU0+msZR6dawY74qU3M7cveUjIjE7zxYdzbJQmYr7I37GgNe6dbMzN
Xn691XLpqz607yaWu3VHrkb/OFoB5owOdFwi37febO5H2E9BnTaMgyM1o4KIcAPK
bKHQmI4qht/+/Df2rsxmxu6E5jBgd6P4leOdnw5Bm+4JtXG8lgxq+Zd8jgvXnNBa
kAOGNvj14jW3ULp/bEF15+P8roSzAYyBAW0aL3rkI6/0sclhdRMs9CP/VS/Ybkra
xXAaVF0VkQSLlov2PmOVgiDJf2qqoT573vVCaoPoGTHgzmZW/dPptUouuEucIpwE
kvJvDAbfsJsLV/npx0UC4Rlaze+u7JiORt3k/OtDvOLEosTB0X77fhSYehAMFHJz
xE+q6MGXfV/oAG0NiSLidjPxBnRZJc6CuA7qWlEA2DQN5vAECvVjzNxnSlZLMkP3
EbRHqFr4puXoF7GKG5l83PbC3xN6FiYiuVocvx+XS6MJ2arRgKJaI6dAJBzwTV3q
ZskUYRpccpbwUH7Z4mtgkib41l3CbMkPbybqkIG//ptrRQH+GPyp2eV0m8k6iLKm
gv0YwoNI+nv/aHd3jv27xF0lO+po2hWEDAMtb4wD3aQaOi8sHBmQDAI87uCKLqrd
TYwLCqNTLc+dnP04YRK4nP343jQ5Y8LLIEGHC3LG0ZSUGCMUfWULDbD7PFu3QAHb
yvbI+AkMp/ugc+8ocjwDbE9OL6aGUxL7Cie78Z28Q8YaBXFeA374s943Os+qjWVa
8t4/BAU18KxwmgZZLvoauUpH9visO6xh/epJlIYWxzcCoqbmjZ3KsHueBsjGnXnS
E76FWFzB9GRv6fv5phep4SRNv0Ef7/K+0zMriNdimBL9/LFpjNrt+g+3FB+WETor
o7lydy62zQ14s0LIJYKLn9xg1peXUbiKoTv/jTjL3lX1ZFDouOoK74F2yKXtB2Z6
THndGzM10GpxdM2dXlrqTo5WcAG/auNnXwqIZrKZN4PwWdj6DPgId7u80HMK3GlU
WPwOU2jRfyFt6dX+WBeC1dXH06xUWu08p9SwnXcuPBp8VES2Atl5UUqs9D4JGKH2
Rn6gy0UYvr4h+vyn6VdcvVbV51E9/nvx49vmPaYlGirQfilEaCJARHoo0F6TChIF
KGgrFpLtbiFxNaJQ23tYQaY0KuFUdkxNx48e3pNeUiZFJGWUPwTtBn8P0oUsDnGU
tx2N1SMO5AYzRbr52TOnq9SNVq/qxpaaOCdGQgz8FKe8iFFtCscoXYGO6Rumy+ZN
33LcNjWgJBr7+goOvPjKFFl7bqTV9yKhrRHrTRsIAhXUU2KQa18KyNYB+kOE1e+z
u2ybvLMBkryuBjnAxJDpHB4PfTnDFQmiI1q4jRWhuTy7KXhcmLt9xqUFQj0zJ39Q
uncw5PimPLWh0Fc7jgGJWJvphZB2PlwmKmgdzs41W95D+VP5p+n2t10RBpsh01Uf
ug3R343Im51vPGUIJ0T+CkgJHHutCYIMZd/u0YKPXYf+N5588c1ICyea9Ck75duL
qsK26tcg4sL6GpfupSk68vnGYYNOVbn8kZORd7O3HEtRnDa6T7591JOZxL3c0D5L
nynf0IXZZYGX/OFz/Hu/ry3T50/qlzQZmieKKBJsX5BMskA0EkEWbTolTXQUjxhl
UNbo6+MYYBGhV8LuDkD7tKzHfktvRvt6EVNIKLUe3qb7eo54mL6tvnD/+Hsr8QxU
9uvGOZhsWvmhbus0q/L7fv2UFCLAl1HAgVWgxm/VIM2Wf4ifjnAqK/kcue8fgZHu
gfsxQK0a5KyelDtinSv2MEUp3A57a5kHVOyuW0bKdtdS+yg+UmC8gIQX8ZTKvr4G
iB9roTK07U5Eui62BfwiWSJveN+HgXlUx8C1KIcyZ8z3TXUJT3Ggp9bOweQkPsLf
8hTT1v3kyBlTzspfhiu/gLHudPAsmNs9ub+2EgkU+bo45233dd/6Qy7sloWr5xsx
U4k3kIUSmwaR8EOPTUIo66OnowJjqzNJQ0SoQnaVtdD2W2Gxxgx4roYlexw4gHaa
W389MNsqTDXJ/dTpG7x257SAUYxhcjUi7rAm9Qoos9EzRolhIn7oyBcxszLJ08td
3yoEp80NlEK5DXJxiyIPE36x605kdKMIPcZki1f6J8rujovfDnXSkHwp0QR2B6he
Fk7G9U4bJE6VAxqytrhg4JIS2GzJFrDgAx5UndDCKL1H9l533IZvrZw9+MtNF7gT
gEi0jzQ3vaDvJJrMpwSeBx80Tta/9V9DBsn+vhHD1uO8tKxl6Kre5EYwhk+dI7c6
yRoU1vxxEoGWpU2Mqnp6Uqz6bbJzihi9vGVxop581E74SO5urZodxwY+ik/qly1z
p9RIsDSVwOlHeSbWl6x1cmeRmm8W7KaQ3xGD1BAD4ocB0oOP0iVPqJ61eW60N5+v
JtxjEUaOeO+8HhUT0ZK3JoV1N/IB+IhNQmGaGP7qDgL5VpC7KEki5Sq+bFlYe9EJ
n9c89j7yWLnBsFDtjScx4mZ/tmlBgD6HelOtkYRcSwFg/fE6scvqA+e+7NtNKtjm
uI6p9tXV55/3X5pysQfviIbASe3KizawlzEDjcQeRq2BawMTlUR0Lvvwt1gFonxY
HVg2vvq1FXCFNPK7od19CDko2HqAFKQHvfQls0X+HaaEP7B+7TTPdsZBA7gp3kJB
JWGH96DNvhTU/MloJOXtvj7gu2W07fX8CXDxFI13OgtKoXIGRQkQysClKUIGsCsy
k3vAo96R/Qjo8xhQGaBNBtMxNUG+iImxTaP6pxgpZ6hnKdf2bWAQoOyXuTMgD0F0
gTLR8KhPmLcXqgCwyoIc9LYf+Gb/qxQoKNFESIiNS7RX9S9UARLfU25+bs8Y6B9S
YObv9aBbdjvB4o1j3VZfxW982ktJFWm0R4PhdXcynvXa7b0uaQSPXDYaP+TccvNq
rcN5ERkwXjcLrlr4wedDfaR/UxGdzpC/lMIikRVR6bejFlH7T/aU/PyNnb0QaLu5
9YG4E66ZlSSj0KtYuttbvUBd8TPadd43tMD23qANeFBJWHUWZbtf4OV6vhIuarxJ
3q132LDQqLmAOt4U4073Sj/oTzkf8Eiu6sjt5rb/enNkqlHL3ShDqlrco3QWqByC
yITW1re9ls5Ng2/KkLjLA6o7FgoD3uAdcQRGFvChd0aFeWQ/nszgePs+N9ldSKYs
J9src9LNNF0rLUKX/kqqmmHF2rjx97owl9FIZ+a64JxCxDG5ypT3xDwxKPulRKbT
osutjc3HwccaFKvwdDXh/6pw1Xlhm5r+tXOVqq5ztI9NAHCYBig3Z0k58YeVb7PI
dKrRY4mA3Uu3ldsob86z+xBJ7p5/q2/ImJ1wkBi2e4IAmb6E6jxlmJGlpeKK7PGd
Ro3YqAsct6sbEvRZXcuALDfJEAjDU62BGln3mS8tB7b/O2351dSZtDyKP7r9C6vH
jQ1NcfDDvwKfS7LssooW4wEOC025yDiNj9hczZueSxFUiFQT6R/gBltOq2dXhb5I
3Sgck/NFxuWN7xk/LYG8wBuhC6mRDPwxolZvt4xD5YfYwaIKFj3VBMkJg8WdaaM+
5zeal6OCx2/SBrIiQGPgAhqSJqdP0t/36ahy9uuY2c4mQbqS+SrHBFh3oHaNxFl1
4y+eHHjfureJmWtGCfhCtDWOLJS+u1RA4EYE5Oof9cCIslUhAHTG73/L12BurGKp
YHynvOcNFHspGVRe6yNWrsgJZRNBC7YetJWbmyibXVDdcntqAdDHijGsbGaUbqSQ
d4H8cy+x/ObhaCk/bWfdc0gVZKd6Zsez7+Dtp/XMa/pvBWoC4sGpP2r9M38TtXHK
Fwrs5+nT18LPMkZYFQOj0+Y0m/EEFrtSZZ1UbZly+KLU/F1PxSdFfY24mxaSfYbe
yUF3qUfX2n+CFbkUXhZADoqMtHUk5/x41+xSeAG9dnaBBrdTRSVQBH0dk7hseYZx
7C0GWjh16pKUXZC6i1ZgRcXcjWse916HhIktUiSy1aYFeg1d9JkRCKxlAr+Z4gUy
C9mkE/8jsn26HcHQzqmk4ZWe2Y9qH9/pimpgs5IwWffFh2E6L7+9WjMJq1ZxWU+0
CQpq5aqvxCzU/PWMli5R1zwq9mDksT3IIoU0Pca1Igo4jo5UNM1371LoNqzCqugs
cQeXmN3KbGmadaGf6EpW/2NM4KgHBks1mlOZLJGPs6HB3E8ETVWFPOJMyeEdEX+9
7YQxzBnV80pqXY6Rw9JPc68NFjtxbBUH1loUlbH6//YC0R8D+wQITDIc+/up9Ml6
wuLDtSqRvEG26bLOu60a5rxiP2eTcJwCP86QVtbtsRrR2IT0GARLAPOmldlPAIXv
Jdmj08nUIwHR88ajbDCVtpQA/q6CwqQouRkvuZtPJFETVSd6t3P0Hbbk3753CORp
zhMQsFJ2Evtb+c06RilDgwlRQqJlGryO7NSz/z+zSMqAiYN1ipqEDq3kC/YqqymW
OV/ojJ4zDF/HgUBCe0cCTXvVWVgb8COzRqE4/ctKStwZ8aqBwUn2+/6Buy9387EE
y6Kq4Jpf7iVaoEnqlrE/wr+JoHCwucU/mwaOkGKxM+Om4M0ohgTtyqu9imHTCjTU
iIeOJOUYc0G9jdhqx2ahteMRNtknB1/50cnCkjDm4a4w8/0Q8LVjc/LjsQn8cmBW
3aFOa7IrNl5vDQLrnAhUhnVVNP9OpHxhzMSnUlbsOlr4piKJCqRj9+4dr3DjjKHa
IRbQyVftKxqMfW0pA3n4lYlD7SWcw+skggKwDbhpz4R3uyIdXoXreXDCq7tLtLjQ
plNC8/KgnfTwGlELU2fouGLRk8QjpflGQTz+e9Y5RY+AvNy2GzneCOMxQ4mBOKRs
O6QwYASQs20LJvWOsoflZjVv/E0xIdKA0OMIK4xtAF7W+4KdP3Gm6dVHyLWDc5iW
O4dxmnkN75W5br3VhWxnHJt5S/g3E5gHnuQVsBlaMq9+Vb2B+eBxK69mITP0CdsK
zPw597BqIjBxZ0IOCUjgYgrnVXfn6Ye2HaJYwlukP1qYJYtrH14tISx8eljc/gLC
y0rIfs+KWWTgJ3aunaGMCvR/7GFXhhnZrCUEKEiWMRvHGG5T44JR5fx3pUWCjcaB
doKEqyaZCu/e0f30JzivV+ATC9rWaf4Qs4+88SH9qap259Lt6vx1TMFcfeD3HCp0
DHsZpPmM4wMwhIRV0x2syj0GzP7M82t7raboaDqHj7GJgr6ZkaojK8Nz2W44j+tg
OTGGh0QICMBqRRWl0NLHkcJ5gx/fil4lUHwKHStSmBLoExzP+Qxd51h5LckG31mw
Bgz/45JhVfzIecCYSK79s2/eBUYoOo7OkRNMwoKMIGmM7v6b1m1XzZ16+ltWqpAo
4dKtKg4EpNSdJFmFDyCTtaWTJnArZo7Z6dOT11W+e+elaZpVFel/MqBgODEA4Z/f
tY2Rlx2qE7Jk411Mq+0Rt3/WM2jJq45Wl+Z5XEjZqtvNghqKd2y4yMQtH755l0bx
D6GIdYFRRV0gI2C/VV74iGO8umFP9htO93wTJLn+GqKKrFPbENAvwDAlR7SYk+bv
stmi3mcEOx7BY0eMHb43RQSnCwzJaMMoyhytHM9LHS7i8vBPXhvKMPxfVW1jKV3E
pf66W7riG4bD27bCFOacUM7uq2ho+Yz4HijDbNZp3pwMQmnUPaUc74S00cRGtrT0
aBcNoDrVCNK8OqEV8zuPnSSqox4r0VnweP8VeV9X5beRxwi57KvmdY1Hl10dRkpS
YGz70C6F1/8xm+JmOKaFasj6a5Bs8Itcxn0Ul8T863VrVA67tlVSInwJHlOnSGHy
5/MFBTiwkSQTQrah3+M7s/MRjRsg/1vSEm1+4ni551ktNKVS6l83/AA0JTHS39xO
0DWmKehAsJ9b3uBDue5wY1xyKH12Njevhqteo39wlRZ443zLTN3J5wX32cQ5Alj6
NppqsIXsyRKOUBiq8m1oMC4tDMx2rbnw/KTRHJsbBL/lMoOLOCVAfhksbMmGedhM
SN3mL4DEFCD1t5VrFJYJXNxUIft2g4Ck6jVDK118H5U1IT6Dx89/BZAjYGslYSVF
Z2oRG5TIKActtFxq7cfB0tCM2NXB86IyPH39f/gNa4Q0WG3J9i/0YFPQaJR3EKsi
wlUVcJ6EFc9uor0LJV8IXVqQGjXjvbidyTieyqy5Y7D7cm2pL3HzFgk9X3y11v3l
4gqtlDPb3MV5ZBpgECt2ygHy9W0PLu5v5xs89JtHTGRUD2p/YpWSGYom6maf3pWO
gnoXoYQqKG5oug8pLqiGHtY7SOmkgoK85kBLy0LqqWoHOAewP6t3sRqBkd/FL85k
NFJK9aFhR9RPnZpR5274YLTpS7Wl/8t5gYcx7B24dglqysMyXlyNzDlgUfF8o9uC
KqV1LVL2JUo0XNDN7m9Wt5PqVUgmHj2RodSpoln9lotrlUyrISDyETurOxDgsIUS
ojgbkgZ86ypSt5rhfqN928r3AbvA/BnwZfaZd+lwMAuc4x8RGAQGeE7BbX8UHRqP
RKjXjsyj/qgYtyk7xzgm9jRSWn2dd9vwoTgdaiwTO/LeplzNasrSPTZCNINXVU4t
OHGa2NVD9mO1GotkPZYUY4KpQ2Xp1YPp5hzO6PwQE5Vh3Cn5KSIL1CIa8Mp7kY/x
MVDG/JlLeorlzCQoOOApFDIog7W04rhbuzozhSdO4/08OKVN3csYErlqjwQOVbqo
F3nVQgCtfu7A8qcXxsy0ejO2xAqlu8dMEwXQtYLvA/KL3pU2gBTWr4rna1JlfqBg
51nRWxovGGDOF+z5w5LmKlE0R7c8wXxngk2yxw8DEx1QUdowS1NZVU8cme7JX7H4
po3Kl1XaTIX175YbR9zDV8Txg7uzvwCD1zKvaVI+kn/T/Rk4lz6969gFPdiXZElp
6eF7kTFXpA3Yi10z0qDoTcLvSocXSB4k7WWSJRUaliorMB0lu1/+o8Y+hWQWypLK
rK1C6mE0pMax2VXNE9U8bCTCYBWLH30PfSuOjWfOzY9wPeD/WCHbDqv/wlwmgZ/B
VS2lrDQrhufxywc7Mtr/RIWI+hqjpgUbJ6Mu+w8XoQ9O3RKXLevCSd26E2JaBWjO
aUC7ptzFJwHVfcyyKBcxPqgf3kFS2HkpIrzQkPGORIEfexocPPbSZ8inTE3uLw4m
cCQokxZtcPaGQsI2kBouSzEGMVBit3f8i7QGhIlfWT4MLda+roQXKvDsdAh7AmZT
wpdn2wRU6zkYTsaJjoN1Fe+IxmjUABuNHVE9DjN4MepYs4rrxQy9wXJ25Qs5XQWr
rh/ZDaXRfo1K8Y1Tx2u1YqhxeLSsvwz18kWd5wS4a7WWaRNQ59cF0rc9a6pENj5b
Q3oV1sBHvOBkZjRYtJXy9alzms1jJG0oB0FPDc0Bfxf9NgILhtf+zKT9IUpTfk5/
aWj+DIkjdb34jiWxq49RAiwTsak3Ssj9UWVft5UNEI6gw8kjd8VacfljDRqr6zOz
g2X0U11s+p37SDEE+hJCTNuVaLE6mxYwhCUzzlCvIpB2VOwHTHpzA4IWqyWlcub5
Hczbqif483+XH2fhtSnEA5Pxbh3Dh5mqqvH9cjovp5XHujKtQhgn1bkWLEozlxb7
fx918+pAUIDo/Cu8FQxWVgiO8/ZpsScW2Anj1z4MFsMjgzx7qwFysnaGW0B7or2W
mU6IGLNmGuBPR/9vj+lVvhl45gnK3iWgnOMJLwPCaGxagmv5VpNIMjWmsOAy21W0
bgtdHeRziGz8oT47YfrKNWaOaY9D1wipVamcI3D6dQMX7c1KXto2lA0pMkSqR7nf
hgKqQSFb3QwFmj5B4p70ZLpRR61FKw0Zezo3Ju7CVPg3CY9y6seIsRL2BCRMgUoG
w/JYfELvBguk1p5Mq0RFNaBkUDICztZYdmSvkNgv53wQnL2K7ZBKviC8DCzOU2hS
X9a5UoFh2tuWMiBDIqc9H26xzXrLZoTHgvH0dBnKNO5bPqKK1ZOFrGgp/Sphly9/
eWRTd2vXrjWKdiJ8qN/0oftolPcZO3V2vn7IP/bAzkir3C2d6Na0TGnDauhDFaSV
lq+cjH+pPTvTOCmaKwrX/iuEpHqgkqI7E0RceNdrTX47N2CMPzpI0tCt81pPU3AY
wqruJRUt+fOM1B3JcWfVff+RRfQnEz9Yo+dGv6XvSdICBQknqygPE9MNn+SuXfqb
slna3/HGCr/MbjhSNzAYf5QUP5NoPbBkImyLyopzrLKYVhDZONWnIbeNZTI4H3FT
v60PPavsnBDYHp7Oe1p4E9Wsx9jnnM/cFDuv0mE9jSuXa8HmexFZxhwTDTu6vw7E
Ac+5WazWxObO9XbR+ZD6ZNPJ9Rt3f3LEm8c0xr0GifkV3vXq9zYwENdyFIypN/NS
NNIITNYfPytUJubfWKcOm/BCoNsFic93Ph+ETPlaukVC/T6ik9RaBghPp79I3L1I
nhV5bEG8k7urK+jSKiLseltwnWzGa42E5ydHJu19SC+M0L21jdi8qBYMTjXmigEK
U7+7DKSdu0u3uYi52cn16icObWijrgZcOqZOLglA1AW6havV1shbwBAUZqW2cGSl
DX8CTNWBPkN0IvtycFmoHwj4twII4vTIAI5hkfWKcKqzDmDSw9Gm+g2kKvTBXsMA
v+OMSImhthnjixbNvNy+15IEsSkjPLyOegaYAcTMmLJDW8H1KBH4ZAv6Zi+++SAR
nkzOWClYvtCtD+WHybUZe1LidmCV0zwmM+lGdCstIDS5L7I5iMztN3/xpk01FxKe
lEDQJpcqFMdrJ2hW4cYHy92bmrU8o+YLsRv9c7rKhO9LqVw8u8IQIE/lZ0w4JJHM
pP7wN/STIQEXVoEiMKyKcTNWOGnk42CulJvD0AsQ28gztMtkNX3XfVxxBvGNb2Nb
K7njQp05HmU9nolwGf42VTGDx3ZAb15i0GAAeOrMB/ymcLoMhSoNUKWt0NwLpt17
8nBt81MMkByJ9jvp/V9HIO8O3C+lrr2hHWV4dof+fLlCSUqmpMdO3HYxPYhu7iEk
/0KZb5feA6VtXjBNc8XHd4wAWpVL2rXTLh9gZBMOEbiCpdqeNrnwDJPQ76+lDF0I
g6GUvdDHofOk+4Hd+32ozY4m/XuM4ZOErj+euGDdNpKD8tI7D7MHoezKbJSOLCRl
AcHaKc5Wfvu4hJIClXG3krfQ/ojFY7DvLzlZY7AQF8rSERxi81kbyDPrPRPYnecL
IjvWw4stsdtbLCqDMpzpaYfYnjtGSPY74P+18ppIfj5fS1bbB6pjcTpCkng9PUcG
yrTTVOs33XekpKZpFb35hzMGEBVJY+jEdwclaL9Np7UGV/PoKTKpnUH3WndhN9Uu
+YcnuyOI67eEEHePOq29Up6BR689WiqE7VkF0HjoVETPRoJ/oQoxOZfVx/Rv+sTj
v/MVFCxyEY5aTvpPE774G9kYRD+fiAWbidfeynWAyqAoufxlZxWOyHoPBf2pje7U
LV60JJp1ajvR6HfJzKv9Scg1OiJrhWrTeB/gk1oE+YM7EFYfGKaOmolg5A3Pej8h
OcAEX7MQD9cz6IZe8KOWkp2ATFhxRbxYfJwBe8RocEaC2WsZAlJppmhMv+H6qhf9
kbP7D1zJA5irqy9WY4SzzhDUssJakRmv0LF1n1kFLRFcdey6IbXPsGvywLFBXlJf
7dE8vdCcQipPj/EsQrwiUQRgeeLSkD8UYRNmtGS/Qi4GDmNGeBEDMv/63fW+OTY+
jHIBXzprqq4jmHVsqDAKao4dfKDhRZAMRoA5tmXGIEBiXS+pid3uKrytvwlVeC2o
S59j7RyPe2llf66+uenPKoJgKMyUq4dlPaqSvC+1OaH6Nxux/f04pDYZOpRybD7j
+lQzLLALjYdnPCy4b4SE8iC18mcJuzesy+iRduBATvfIH/1txrYhOiLP9wAiLcvm
FbZp3xViBTFW1nIVr+xEOC2NF89I/uQTY+uMJkwGtQ0oGciIBjP/BcVb9trRPtWg
n6bOaxI4zmGuPb+5dukPLoLOc9bsEDruA7IYBPYTkMUZIDU1/JDeT5ZboTzl5nGX
+rQO1iPUdnJBiR46BOMxd7nt2/UZ9MtOvVH6CKqxdMoGlgDhfPAO0lZdyEHc8LWV
Z14hH4XW9o5XEQGnc0d1R4uyuYJBwshfW20XBeWnqeJSI/+IelzBnpnE5Zyovoeu
DDLKkjxkWa2VpjZNUSnTfANXb8XIZAxUq33HY+U4KZpndANOor2p7vfRe1OVLr4U
BiwUPVRy+5xUNvXs8/HXyTcGvgtQDZoSO2KNWSy6SS0+CWeD4cpD1BhPv1dLsy+N
Gs/RFb3rnrnOehFKtazzaNWXx6VO1PH4kA4cI18Pv9VBQ7zBTlwCcAesznq47e9y
pPcOD9DYpycirT+zxCfVpdXQGtxSsUeH/tflG02vYsHGefl12a+OublyQ+YsKCpu
7sIP5UuW3uHzK86aeK+z+wS1ia4JqY1OYGDw9CleUmNuJ8b8/6MgPTUT5uuoXKNX
FxGMTB9kd6XPK2ny74EyqB6W+vEXT+GsIJZKz35fAS9BMTKP1mEtzXinmhZPykmY
nb26u70NnrrxkrGLkSL1gObB3TNGm/+W5UVofZKzkBV+5TDHawOPjN3/tWjZmt+b
1a+lxRG8ivYOAkfRG8Z/ygxHiq5g3j0ffiAnxB+DlAHvB2HVr5+uKLKZNOcUICPh
l7ck3KFOJTLm4tW2UYizYIlqHmGxuFQZm+DLjpVHShESMLkwshgsM5i1BP0UiXTW
wh49aEdaO5ktWorR7qol+oEWAf3oCbMCIDCFbH/DoUo06voiF5Ov1oiZ9b7jyZbG
BqHnkzp/RS3eFQg7Pl9oHm31Wgbgi2dgPUia1cZ9KCXzVfgj40dZO67vnyyS/V3e
50uxmD3weEfzZcsq1QYfQnJNFYbzg5V2WCyoTgDxu97phbs/DGTgTiBkGVBBJvJ0
ewDVNfzz5qXS9eEeZRQLrHb99NvsHjhAakxMf0hIJTo/W84FSDG34j2wZcDIaM7W
5cePgjnLZNTjKAKRtHLYQood9uXxoBGiIcJbur5ZAHuJLSd1h1Kyk1O7JknBDwSR
f9g0ghs4LUhMSn6A2kZ6WwC1ab6NNE+B0AUCOrH5HXPowKb9N+1YZtGv4POfsAsQ
eo26NI1t/LmzOywCJMieW/tqnlKj8jhlmL+xxVRUADYNtaxMs+l3N6cjzZDikoeD
MoF05j2ojpgkPdKqb402QcWmEG8j0tLh75ZmOiMNfb6RMzwdwcycXp3GpkXR3tEA
b6zp2xAvZOJwEz1/5pND5Qi/EzfL9LWucdSiGNVDzex/DWnsbcN24neYIe2M09zC
/D0ECdylSfAnu+mG4CFe8L7sNF3y3Qd9lCjOkyK0JYqiPGuCQtloXQD5MIWjAaqk
g+thQNcwx90uEzbVtPQEzzI3OLKGPvoPS+UC/Og1f0qWo+6rsd4sqZ/LaT84Pfju
1dZahwBEsH6CSme0iKZEahETbDx1B1npb1hxvLHxl5UDMxVUdgU77oEpphokWU20
4SxFEGMZy/S8ktRTNp/Bil0eSrFz5qmI1l7dXWyX10z6LRAkIGOR9MKJ+AsW9I3o
rQJHmzAndDgpPwMgM09ja3Rb6S1jbfKZNgcw9uw6CYEl2Kv9imbrP4n77MAJ3Qhb
wGzs3mVVd8LWV/m8EaWETyYo7TGh/EYXBNbnt/4Y93dxw/5NLUVqG0xfEvuOfwXX
OyITavqLsCaVX+lKMw830e29x9tN3W2bUc9t61Gnx1jkD/KsBBah/BZeem93eScN
0WhMyqdnDgCiSY+j12jXWgOWVZYJtC4GJXAnPYgBHBeO/+YmAirP0AYQDj+MCZ+H
60FGP/FAXkglgX7uU72BeRHZaFPDs/V4FH8RK72j3SFZyI9VApie5Lj1yUPVLyG7
hNsXAcCLrF67U+mw0T4CphNGiB4x4UzN1+0DlPWuL+fRbbeabGdKyd1VWXAN8bWi
gFzPtRyQN8sfLWijkqtPtz65WrgMstDIIvsRwxQEYJekXZq5kOcXgwMKJjxA/biq
4B8QBqn6O5rg/aqfwUQ3ka0Y4GpsHWHj5ogLeBP5A13cr7g3YYw6X5CxL47RSFYq
zQNEwp1N/aPhnB3ePTyyxfOa81I6vwVIgKeEBVc7aRcSdPOR/eJnO3cMKTRu3xNq
yORsc3F9aPXzhkXiHiPZ9jHXKzrAnVU+NFp7hB3GT3N6ZFrooS7Ocg1PDFfTHf4l
TGDOIPFddOL8cJgDorCobtOA3Jz57JDQzOnyk+sCRXk0dxr7TPuGJRm0TCW/5JEl
0AWaTrowfCAbt9P0F/5mvDZ20lYksR/tjDwWWaTqmwsn0O50SmHEwEOrWo2tCBSQ
pdoMT+rdmtHSiuvhVT3Q1X9Z7Yego6JybhpnH739bnePFMnDw3lunGtb0DF0yxqF
pomsy0HXCMIeSiTMojpEizRIOKspBfKuDQ8p2DrTQe3C/7sUUR8IHyVfLKiYqAih
RpnNiFETLd2pegRFXACZozVh9VeBfy8EO6uDpjkXpEVtqxVM+6tmAgiwKtOtHaVk
rZi5r3/UlPJTpi1kQpKs2vF84Q648pVTOV4D4LrSBO7JB4FgI7Kh/UJ0CxxLS/fx
I4HJ+1xH+7jxbkakGJERQi4sQY5H0ea94Mwp/F8lbOglUQ/Cn+ETwZbgB+pScyYy
znTM7HuhjFnl2Y4b9yQnaoGlLf9PbF8avpc6KQq65hq7J6X5zDeqirle7AbS/JzN
MCZwsjBWO2buB2YSxSu/DA3+CwHKr8SrSBUAlxbJ+2ypGT1igMuKLxqs9T9RPeTW
9/agYagug1W0eJomp8Ul0uLzOgODXyTc0yw3G9d3BgBKpaSzvg9IFoLKlf7C/ipE
xTwodkLpk5BMLSzz6MEkl985b1STQ4ajZIJUv8Ja2ncM1djYvfXq7hF2tw465rmA
uw3X4mDaPpBFJ7YPzzZ0aoerXFayhxh3e2F5KtDYNBrjUUbwC2sv0AwSn/zjbzTr
zUnpGbtiWp5ACp2xhLbs7uBqsKKQs5lrUVNStPZ50xdHz5IeeRgUcrNlHsc/banm
bb4t56ZG6N4kx9VSgZfkbNipCSGcW5VSgqrmYdsU4c+eZIGITgbnT2I8TD/iyXI7
9cAOWCcI5t20nOYzceEVoGFW65KWhv7QsRm68XKGt3UjdxfLSPGJxJS+nGBIacfW
fJKQstYXq2V57VLUlgvPAYxtEZ39wQWNmWoAG+K0EQgvLDBJQyTxCbeY+U8YGtCc
+YUdj8Ea4dtxiPLbfPOH2FJSHuNQzO+3IfIU0GfNuwubcJA4dx033rxSfb7yZ5AJ
LGX9Kc7FBNal9G3svuKGysfnDeLegrgMV1KXi4ZgvvqqiFUsz5p2K1MrxXV1Z4Zt
CbLnfutRrycjY0CfTeZ3msZeLP3xdLqR6qjOecvxzFF9mtivJwPzOZ8Yj191iC2m
y7qWKQNo3ckjYHZ1C6MJhdQ4mUdtgUSjMVXXJX0mcGXIzH6uJE/+VcCGEfTnCEc6
koOzpu6acp8Gnmuis4w8dxfQrPbZ5eeBD6PmjBH7INDxl4E21l2xAvB6QBzwcwBR
ZjJ68YN++wxqbiX/MsEtGFsmkB+2M0ruEuFtO8AfbTX5jNazvWy/cGe9KowqnfrX
mdEDe2QiFZxksv9tj+54HwkviCfqICbIItgR6+9DJR8p9OjeeIHfjuhZGIVMBHNG
MXSHF1Di+pQassqEOOIvJu+ZuCBVFou0x3MwRwkLDwKK4IZKXhr1ag2NidLLZY4f
nkNT3SWVjhhNUEdFcfS43kt1gycVNddnvyyE+JZobLqQIlLr/dqJEFTMtmB5hRFI
//pragma protect end_data_block
//pragma protect digest_block
Ct8N6R64rUGQ2brO0O/mqbH/i8Q=
//pragma protect end_digest_block
//pragma protect end_protected

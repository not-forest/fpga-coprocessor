// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
Nj9PiuerjJHA+evifalKoxoAwiat+OzjV/MSvTTFo+5fYjhMDkp1LFTJYSGniJa/
E3bdHZaP7NXNf+y2Yd5GHPbSY6gADtKL+a0eh0+PY2pTCbikdV9TdUXWkML043zJ
uRHfyfF6MMTX8UswXxpw33Mpl0G1aid6kzNkNEmr9OkJ+530xSfhgPXXCSN/tq0O
0TCj217gPmkig0DfXpDQLYXWS7bkIE/OJQWdD9qhkziyFBZrcGloh6wzIZNZVJDs
kZlScINT94XF42rQf5wGZhu3IGDPgekp5scamf6j+/T/TaDyhJV4yBlnBMpIvhLc
mYU/NOex1nkFG0rab0areg==
//pragma protect end_key_block
//pragma protect digest_block
xvOuM5HlFCbObN50hWa6mUddZb4=
//pragma protect end_digest_block
//pragma protect data_block
zOJozypwlKs31SRWnfCfoKUsLYtYXw+dtZhPvehc9ZQdYkXnaZgZWQ3pmsQQ5iHU
8qBgQiKFbQFcDemzdH31bK2uN7vk7GsxnxXr0Sdc5Mi0iWD3AHxiEvTrB9LfXWFF
aEqrqkfmMQzuRVeCkYWMvcgbFp/hUrgNGHAsXJ9pjWFmIjHjEz5dBSNYw2/h67n7
s937QvzkO14yP+xYLOu8VKjt4oI6unJkl5Z6HkQmZpqgz1t5ap0jYk9YQAS2OVBj
kEF9i9RQ+fIV1ZzEN0uizSjJvOCx8vF36cfmuRGzctA4ao8QHKeMKJfPb0j3H7Cn
wb91RnIK3luQDWlHP4PL5mJdYO5HBDIJbyC9lIlNVxXgz3yA6h2tk32uOXM+tNON
T5i0rTdouBq0y7HhiijgUUeEBrzXFTQ0GeUeUQO1sc3CSAbBmwFYa6Nae92EbdhW
6Vg0Zizbyb33xS5zH3TNgtqsujGlWRNm5T2GjyNkj8afxcL7L5ysvys3qwYPwkaN
dMbA+WUpdpjgqMNKlA46j4GsVqxqNIxiBM8L4zdL/nQrWEW9OmeaNt5bYHN9GGJk
vYw32GMti3eA2uaQLXIHfrwtt9GygLDXEdQgalUIxJocUtOLcGcooVjGmGKPD/pt
TC4rJDkl+ECM7+Gdnv1KFzrbi8AKZjgfcF/d81fHZFV2pkt71uVuGj8CV8Pij1sr
5svDCg3SqjWhbImcjYF2lJAFqZb51hRgV5RiEEoc7fQ3p6bgHyxvJ5m8PMj2UZ4j
YTiae2L0Iq7DYjMsN6cKage6p0Z+iqUvFWXYE+jHdKh4C9zXkr14do5MdPTnAaU5
W0GqCchf3qSiVMBeGyOJXvE5rEtwReKxAQ1wuNbOZxgaCHgKx4JEzM38bfUJd02x
I+Nb5iKDbD1IHF6SyaRTzEvnRums3a2vbi2QTQm5RBmNhX2hjvJt4qydBkiGVa/+
7sONiXrDCGiBWKDMtK5AJpuy0fWyNfZhzuoi4cfTyX0YrRTX+29g0+D3i2kPA9nT
Ckf0nak1RFBXJWwztqwWLbnSSzU8mcvUT+hzse74hSb6IvoqpT/8t8Ay7TBKgE91
ppqMJDy17poVaJapBcjt13UMWk48GV/0GH8vYgRjBKhwomCJLtGuKvJh+5sOoX48
zFTtZPJA1AuWp7VV1pLbsWwBGs9lIZBrfqxuKzFH0wkEZnL732oRMkUW5b+dVJS9
1knITFNMDTXdZNXJUhXQ6pJzPfpJZzG6fino+FRuNi139U2SYG/FCFO8QLu34YZj
zwedbZd6RVTrY5iDVEgKdft1ThuOYukoIvUFnbMXXVEHZMDABmq6joPFb2GqwbWX
ZvmM5whM4wjIsCD6NrnTQuU9UvqDqmgRDvx6jFR5Mr26Eflhp5CPCkVl1gJEyxra
Ujr29d67b4sUbbZawUsepDtInvZH7NfvApuHK0UFiXnf7UqoSEqFjBAgPE9SF4oK
sGPETLqBRrR1l7qsRwXsblUj02dzWFJNl0C+YMurkgsuT6rb/aqE7lGjG7DsHhx6
EqILZVFqKpYlnkrZGe4+VTKNe3aG0FR2LP15E02QWrIZD2QaF1lb6KFcUHVLTwcA
WAnJjgkERQ3FmBVxZKDJVs7mfhSa9QoA2ampxehKdKKV8NPTwFHSxyyWkRR8QDxC
HVfUOOpuLeb/vpVIhJr4vmrI+RCdebMLaldt3IUBGcdmABukPT+7o+MHECnfS10i
bzyGWudK9psOzNVkplynd1HhHkB9OzBesf0lWlCq+6R1ARfmMAmOZkxiFpFW7Ttq
TsuVh6VaF5BqCXQitDhTfZrP0aJ09SCyriswBslyCOyYnux5f+GGkU6KA4P3xNrz
DVOUyrg1ZKHGtmKJCoaQkofK2zQZcu43h4DxCX8+FVHkE5/DgplIe1IpviEL4g42
miuVPF7hKwW3kCvxakB8LMsKhNJMHZDTj8v6LZTZXo/9L3B9Bh7VwQXw+9PuQr8g
+u82JuoOKoiGnx7kDv3ZFGWvzwaxInWepTKXrUzOBTsuzS5UTmUalin+zTuW2zB+
ZXlkmxFrJoxLz8V9i97fu9gmXN6rP1wbIYz69UsCSr0ntnT/tg/Vk8IJ21zK4l0u
3Me4nIq1ZD97B6SGMuZzgEvjPxrQrnqH4IHbYbcKDoPV4Z2u/sW8DOQ1txvmCIeG
cViZtTZ1p/lloHIj1X8byM63H2+HkmuMnchOgGqRZTipc0uujx81EHKSkmNtjqQa
DnurSTA4ZqlCk2dTe10o8ODMj5tJzThUvw5w+UR5xfSvuuY+6tHGvtubq+ZUjyZz
oIs2EYuOcRA4N0I+INwzb2P2eTdbIGAdZ4SKeG2e6xSao4+7Ck2fK6Hk9LayI3QS
NAKa5onGSJyiMe6eQTOSOMsqa1BAORtjieJCN6CvGjEpzyZUwePopmO4YaDzXV1f
655DjP6mmOovRGmIcKRvo7V05Wgvoo10IX+qlmEOqga8oef9orLypW+D5tSIrrmz
7XvyzSGoyB4vvgv5g/xv9y2Crbz+s85PFx1s8foTgzL5byqqZdPbhq9jw5Xqq8L5
maW7sa6j2fX3Zod7qvBk4evsXkeypPVTYXjaDvCqiUeIqlZtqcTGEDgqdwuZlwKG
63iIG5LSHWzaBh1UdsA/NU3I60bpk3TdRt5Z0pBU4xUqosscjJY8P2lJn7GbgZB4
SIKwdNha0w4bAHsMIGYJimHqAboXdWCtr9JxBqSSZkAI1Pfhl9TB7nte8KD7MR9g
xrPsr0GMd4ENa6OMc9vdeGL9ZLjrRrBb/B7892bluRyeYZNWRvnUt3jMAkuhRiuu
NGi9YPDUsPDW4SUL03OYwJz4p3HuZm8GDulA1L28V8nOBPOvZsznpiq/mavjpCLu
5fchrJ/eA6yjvHTTkgJTDqARQ6w2JZvI3Whs3QSWxIiPj6LziU0XmR2Sn9UtOW9S
tV63Ibp/H1Crjzl+SajdXk0uZIuXhjz31+nEMblKsfTb21n5VhJ7+prz+jbzVBqZ
gNq09SVgNbumMXqTbXcJ4G1FSQ8qRKEymfC/apbEoz48a8SgP/Yl9/zfRHrdakor
RR24zGwWkurHcsON9swHRQ==
//pragma protect end_data_block
//pragma protect digest_block
GdvntudoqLoZXxWyy0q8cFL5rbU=
//pragma protect end_digest_block
//pragma protect end_protected

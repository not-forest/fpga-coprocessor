// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
VnxuCr+L9ga8mFusGbw2lT50ewsuS2y1WJt9hdr5hhsw+CrJLTLywbzsc2a5mBC0oNNuV9tordJb
5RlK3T+lE648d+cAZ3Dcp8gthkUUsLkSc2iNl76l9IDSoPcAmZzt6rUBGMkvUmKwg9PT4M1EbfI1
YnWAExOnVhmSqiD4aAbxwm0zcLRFkKmCo34vGKI/i0omlHgFlQltecXhZpuEiFhnbgU5xEbh/5TS
0cBXSJZhWt1Vdb4zMlyjNwjodk5xD5kkYgyflormCTzhyK13Qv9O8YW6afjSV63L3wBr21FcOlw4
32dOJ1FQMgLQ7MeeANs/sqbzJPNxgEjtdBIS9g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 15168)
nkf6+vkhyEt0D++C/7U6gSalCxbVF7tXwlfeNt1UQV3cmuW8h/x4ERtt1EiTffApzrsIhfVD9QKI
wSI3ISejyRF+HcaER8U7/D5mYglb2rnchXEXIO82Q8RaSooxGCVGlnC9YsrwV/P2avugIsbZYlRm
j/g7ON2HGWurtA4DRFZGRaTqvm1TmDLUMSJeY4q7u1lT0Hw4QIhteJWWdvOFefIySZw2qOxFe+jR
oseQv9FWsHxyIJoA3OFVN+Sb5lgp4v/O3XWG5hD4ShRP1oYGlGT5mG9ypYyp5+/qQwuu4k1ePB4u
BHDpvEahyeZkN0mKE0ZKSE6f3O/nInxC3BlZBNEfBUr+24SOFDFo6ZIqW4wV4mUcnRHs4eTOAUOL
e/2aEXv6dBc/izB3m4s2N/qP6VCqL/HK5yeVRKACie0+rr31RTGdFxjRuZvvuOI9Ee9/D5FV4fYt
35Neeu2c7+PI+avJ6/8IS6fIp33YdrJOzT7HOeJk2Yb6D61gcwFF+tfzT0ME4hbWWtAMZJlpRmDD
KdrTHOiYN1wPQjgSTx5S6JxA7X1iXql9w1xdRcrtZ38KkQeKYOCDDJgr3O2W4uYpBSTOiIsIanQS
NtVCOeF7qcNCUMFcZ1bzAGao+19pbCDSqqL2EP2LSopSEZdLJPoLEMpksE4n3m1wVY5z+G4GcOPG
Pa9dBTs22TlNTes8c9MDONZVFdPI67xzgy9Wr7uvgutS0pvji/I5qJIO0yvUROQQu/3iyLGKZV6j
GPRAVT50StinMJl9s5rmCgXL/8qH+dS0bjSplIFTzKdCgfMp/CDy37KfNOGfJvgvGCibqmXiwshm
76WA/khLEhqbtAWhq7nUdc2tQeLO8eUmpz5OHaILNRfpQc3W9ToEEXK0wZhminfxGRlP7L6w71g3
F5f2EfyXHEB69o/FASh3urYitp7+9DnGSHfpHuKIfK8hxuzR8ocpteHhM3LmgWURXOQitzBhD6Nh
YZNmtkoTmlsCPOQXKx6dj2r+VLZ+r3ITQCgIkIvIcYrizMD15waDMGsa+lRz0N3l0apxkh0hZLK6
X3ESQUh2W3u8uT74qGNFuhLpCirTLbThQo3wirIwo9TMMtxGVXTQHfxyOUphXj8F0jlTxbajKNt1
726y6VkArQd2cKYH39fwKTacLe62T4lI6muloaV9GzZmTc28lMqdeE/JX07zotQreBXQ89BHXbb7
hfdGVbzLBlLzW3dWIyIfk6XKcX2LfTeE4HH/5yZu1WaycMaM3kxxkDm6M+dIc6v8UszqcrOX+uyd
Jz+G3iT7Th3sdpswIAmfG6tOFP1XIPSojrRxf2kEQ8ZexGf11X2jeJSgyDXfSQhcPZQXbql/IVli
gmufFPWXeo+x3wy6MRjTn2tMWk2n3f1EBYGragN5xXkXG2Ac0Skz8QngdipL8rAYw2Zw8/6Givlw
Gu/2TXbQj1RAH0t8PiCs4hjeGDdsgejgjaVKt/K3h1vSB/o8UP2LP0AW5hm9Pfb3buqDgTGz6Ex7
91yRuesb5i+FOtSbdv4RgM58EYxWTWVoniWQMc+dyjZHDSn1XFKLYX52ja1CjTLCBShztNyFA7bu
5Ef462SqJ0WkahKKUInGU5GYq9yPxFLpelg1Ssczi0Oly8pIG4RonzE4n/L5s++G0BYHUEZZu8aL
pPVDQw3TpR08B4BFqourq4uJZZe88tir6OTsO09s4Xr3f7mFIx+ko7kUHPwcHYhDE/yNPSPY3ztT
qZLoQSKAPHgHy1uoU1iyB4xofDrnSmhiQDycC0B39oTMKDRi0V4tXWaWNxilKGcT/iQNRp9heCSJ
C5c1fDWBgS3Bo/LUGqo31hgfn/IaViPg8fq6IT2WsLDU+CH7mDXkVcQWByUGOAhuM93BtUc6Cl0O
qPvQN9vF0P1lny/xXiJz1yX5R34vt/AC9v4Q+kv04EEHXvD1pmYFxleYll0BWwvVHZ96NwZCuNvu
AtDvsbK7a0j/atIdFg2HzsvwrMqjq4WXudZcCqoBTQ25BiIHSXp9Zqq+YEeTgW9HmoMVimfMxhS9
wx3cgXsEJLqUq6PI5vCkUxERZzCZIaZj7n35NShWNNhwcalzR3b/6Vjz3uqVqxcXELhiZirigN2N
amsrmvN/97A7vl4GwPFDdnpY/aoeY+wpw6LVUHqn256l6s5OoDU2E1T17QSweeUB++8Z5znQSpeE
dwEPIW6XuFprfXqb3YFJCFfauLMrYLnDLUgrpm94dN3nrrj1siy5UeP8slbJ2PwTtH4854c2NGxj
PnBrkGgM/mbnIx5lV3BEQcpGCJNXD1IQTy7EX1/9vdZIWQHTAw6eb4jqVRMbeHvHSXHRHrgOqRn8
7lKoNvzmk8skxUUSmiN+jE2C+c97UJebiGov+W9mFtfCniTvaApvRiWnzqpzTbZ14mc81A16n1xR
TGEgjue1PuX1RIJRGLTH/maZ7EiWaLL80HlY0QFbmgHNup5xjsM/yfnlk/MCXLAHRXWqq3QFmpXu
0N6dZ9VtowopXvHVCHMpObKSGPv4obnu9xHMU8+41MVy+I+6qLCjDmJvL8MMDSW3qYSxmGLWzCuJ
SPUDYT1fZGqGyU3WVlYe5OeNGW367iTwAmLvw19BhgAlxnggMyipSOS4cnPZUt1WGLO7vPv2W2/o
5DjQqMEDz10ZKqaqHWR2ALB0QfhG5Vi7xi3xec0Q13UOPDk4POStpGIyVUvYbS9z2x+rKLIY3lOB
sGhD8IcV4DI3N98TUBZb5ZL4/l/cm/hYc5Ku2cLKU2vKggrogkxyO0R9I7N6VyMFi5DlGFmV4w7W
PGBJhhT4GvpsvnNlmKilZrdM0Lv157eHTN5RdHtGlxk0kipKnCR7USd0X8Rj7LaqIbZmdu6TPnbe
ep52+2WFvkFw1k+7EL/ZEH2u0dGGQBhQke/foBaS8cdH6MdxWjm9MvtUJgUqwuHaBjjO+WDshbiX
1f/+AueITqAoFJ2+We9kQNt7tegyzlQaCml09DBNlSL61bVtxHL23e0Y/NRRLLGwXK5JliB++FpA
jty9qBXgwZqICzoZOYG/XT0RLnVtY1Tka7Oc1YzIX2T2+HApTdORzE3FlFAD25IfNseRxxPcY3bu
kKV3vHTSVJ5GA9pYY4G8jU5i1yUpiRUwgDMdVUiy+D/7sVIZ+9s1gFShKK/r8VMtNT2jP9M3rWXd
8CnM7f4n9wu0fqIeBdQnnttglqd4AASKxROxZqRQnYwhXpRSaIxTGvAhWj9DzijsbPpmHC53oWCA
7XgFpRcL9ZLGk6mlDvTTtjp/J4IGmMTzR6CN/E8IsB43UFT41JojTJPuKO6wVIfxBldUj0kRUzBT
ud2uJFNsn8PuUWolsXTjwE+k+zOTF0h+BeKVuJQjQYAsMd7qqsHFzo4vOJkaXTUpH++C6negLELU
OOcbf80jEtFdpUMOxSCD7iC2VO2ddm4/7Lv1UvqCTjCIe2AhIl5L4pgaNfVsHNo6VHGXlytuMWIu
6BrLYeKn0D9w3llJJkVB/uk3DVSsBHmYBZWWec+ORoVAnXjoxgSAROY8IREpCn4cF9DzYJf8sXgh
GKVApb+IbeL+0AY2tkQbwhOBtqqD/JOx+2t/IFKpAMhCpCxSlMCs+/8e+EhL2ZUlVo12q14/ab0N
mbit4TuVJEHnh69qTfhk9PvDjknk6olQkJX+hWie26sFKhaYMSLG0PCzT+0vch/J5av3UGku7NRe
0ioT1uNbeouDxdzsLDpz7Quxz7fT4/4tUPUWzdvHnQC6RyIim6pkJClTaXzbq30GodXizl+gY3bZ
N6cnrZd473nBeW54kzBd6DSNGt0wk4ti6KOAWncAy3v342quYQfF4gzW4aLGTaiDIDUPSQNOGDJs
pOLnao3Fm8gJBLSDbwkzS/H4E9YIkC3Y3FcS51GnGWcG2/Vh1KqSu574ysOOhpCuGR4oOctTD9gx
/YYGskY+KGTNlOnyiDpypWcUwZAAEhM+AxoITuAanM5r2BQpzGJE+Ds6UNPYbmAcvcNU+Cyp8gb+
J6fVCtqD9DSG3131+G5Y3EzvwHLlpgjny/3Mg9nMm5iA0SuI675iGzfxzl+0PBa6ok3Mra8CKsG8
J1ef0FdO+pn56oo7Wn5YA++MaOVbmivsrMhxQl5FWsf8u0FIsvcYIO81V2tk0PLSsgTJQzTHV+FC
cI2XinzM7dydLwnIOW+yo/7xkUvDz7G0YQ3Xx3xZIAzk0eKvu+xTG/zmonvoAZaRwVIN5Fd1m9fq
+SAAplOS+QdXlkan1X5oyPxnNpSOYTz+CF8S5I+CCPaLISaYVw7/OnXyfc7gOKt3KUDB2ilRe1/u
gyNX0E1su1K+ucqFQaXfM5rIn1vQ1fhP9fHZQYv7x6e2h3xnZU/hBzSZe7TAQu7zWMOZKWInVdef
F9bAE12drPGhMSNa75ViZ2nWC+Gauf4HtsxreTSSV3eT675csZ4cGu/IvKlz5zMJkm0pJ8kmR6lQ
yZQNnf4HUGDREd8qTTSyuqAPaeqbWDtVOF6wBaGAEtPYR0rml9cg8Lm+1gKvpilidjvbhJ9vWnvv
mhXFvvOrtjs+rzWCeKmKBtoO06Fa+XeGyjYV2bUdD2hMSLAn0QGzeNqdQhQz9gN5rfbUM+3JlpZZ
cHAzEnYMMWkpIKYIsTgur9ntNOA6/CzRQGaKG2UPCtgQmAcRCB1RgVAAWa1t8MRnFAtWCH3lm4nB
TvcbUDti170v8Uk+ZMQDxXetA/DikARaPYCm9gPJs1dJ1Co+ZydFX5w2gJFM5+Asp60+ibwsmzan
fQ47amszeUfpyNiaN2etti+FhNDzKVvqBKAmtKgZrKs+D1Ha/1Gihw+/sO90kLJmkP9ERpIGEqHq
CWb0QCRx+OfuUY3d5MuXpUkY3s7sZKlFbki6XqpNLqc76pnr5m2+/ef2H7XdN0Dxaet+Tc63lT0C
GDLmFrOypOX/oKtjBuMOoIVkQlor1g8XxZR4nPVYux4XlsYeGPAcGi9YFBnADrmG+81NM703GZE0
D+Dj1uEqewY3Pa0I459gO060rE3m/zR8KfdwextCaDFDDobd2SJZ/h3H+hIJ87n4mY0YDmNvuiDS
J6a4Uj9BoIMdvz2/DOevJ6z/uub0bLw3ITKGtpdq/GMu4U4KPKBBcz9MOZFMBBJTjuhWNWZu1d2K
AeL4dg55aKBRX6vTIikRnIDlGLYSyUPBdT3YdoWpn1kqjjCoVU4YXgvgnsqMFk7J8GKUOwPtEpf+
UY5O8KfKRqRCloa+TCUPBioy7xAurnCA/u/RA0zulQGzauurenb4Ro6GAnIr61K7W7k6MliKreNU
wrzXdfotDcgolTrZA0/CrApTqgFNlMhDUzVtQw67a7cyt/UnG4jRYUqzIMrjBa6ye89LZR4c0d5V
+Eg6lU+uUrlyWoUc+idnOpLGAeAW4VK5smuiGbQu16jDIWd5m/5rNWYb8j8lcCGXcqw1WEwKmK/t
LwEqNLiy77aym5PlmyCLiDX5b5DSGUWbiGpxAuo35LPLmB3kl2dShEG/eQil0964e3tBB41U0Jz2
Z8T4HGgNelR3m3E+OXMf/FUabsZ1MrwwuuGBurV/ERpKcepAVP1jrplNOadLBjkyAJdMuy6uYcEW
POjPtqfAgqNKioQkd3XbY+gRG42gRBO3p2hTi/Qtl5gfb4KNedE1Ssnmw8r2EuX8ynosuePPsm7M
zi+PaE3cOejtibZxK44Buni4wnvTTX/BU0qUU9ualavgF5+1TZYNqkN0I65+/d/Guh1ddZsMnQBz
o5kxo3hiJPU5qp1Lox2tuE1XDVhkGmPX88glcAgxikyn/FN8yW2Gfd2RjO26JqV2dsL7RtAdJdMn
BLZd5pACe+ozYIE7wkKS1rKWth4tQDcx8DHO7IOVxedhn7S6xLuiHhhcOcELwvMbyYdXa0mboZ0m
sgg9TNgJ//2RkmaIoOr24mZ1F1v7sEkgHXQDXUh75Oihud5A/pRS/We5p5ZmX6q1777HHkmfZmQi
WpfvHY4i+4w+cB1uvo2yqcEe4jBV5Jp+WGscaxI2oB6gnfAuXIkNyeZ/wOMcS8MO8HKLLWiCzsa+
2sFhijN4qas3UjoizAna9Mbrul5reazrpZFsk0hlb70h6L1tU0s+/rICNzPZ7mwSEff9Gkdnao9O
2aIHA6t8E6APMPPPwRsxmf6E/R7Jd09aoClmKtTy1rvSaXptBbRJyL87QBI1KRmWUN9eUa1J9MqO
kQ+AX1tjf2Ob9A6KJypAik1OhUr8SbC/5Qx/4NYqtWYpxCMKZtReaqMNQ4vQ0SxzjONmhJfNCzuq
KWtmWRO7hdyOiAk2GBGsg6hFICGuJD/mbv8lEDiOZ7fz2vcJYyMaICsYlISy/FIO34QPWuvkAPzL
bmEhlj+EQiMF5m4uUHOqz1THmnHlGlFii8PX3+W/ZoxREEATYrNDwAZJjmwbDSfWMUXMaN7mb5XU
fFII0eML/bhe97SFCXGTBHMTSCT/KMLCT1nO5v6pqRt9htnrSygLCn4qgszNvFp/aoLuJ0uCEz9J
qnuNkm/sKQTJA1kd9CMVnFJc3g+rnXp1RuwkU9s3sreUGQN/nSeTJo5MyF9u54i1tuWzdtPP9XP2
O3FsyVDJqS2zRZSrLDbJp1I+EAX0VBaD1r/KS9SREJYpbdpQ52c8tj/wPMxlpWOGP0n7FqXDI2Ht
DHiz0T4uH7Z6IObRoQMrik8Lz6I9/a4nopsQopC9E3exUwdogI2Veh/RFdnvJ6dNRMI1IzH3OsO1
tkdURAy9Ph60gTIhi8FpzeHg3pJuUrxXx/758WhcrbUozTIPA0mrhQI+F4pdgjC119iMbb9gELWI
1z2jsYoOKsqdyRwtqG3mW3E6VEDibKwuOGkUGQF/HRq5RFbpq9T7yAUYce7+fmMjq610Vjp39y5D
00ZIwQbXXg2UsP76a7p6AK4O55MGnGXxXJ6AwIK1ZJ1JjuckOi6dPGWYYaXjFpOQbcZ9Raqy0Swv
LoEmKTyvR19ItA3skBHIhgtDYsgt3jNLtLxmhAErJslnnegBOJjBjkDuhGHm6NbrR0dipaPQCRD0
i47Fr4BQ9XomURoIhg8HBroGJPxeZITq6K6GJCPyRINADz0bXczSO1wyTRbRd1Q1Pcpio7ctFBKH
mKhQELMQagVpSzEIWsrRKLvhtZpqH1q88s2KGUlNqfhqmyHnjiFFfy/xqVyl+QgBAid2XLVNZ1sl
zBxzvuuVQ9sumF+8CN65CrEF+AD+o1wmk2w4Qk6S1SZ4mcJ/ZQWlsR+ieBRwK6tSDsFyrREshLgu
VraAqOg6xfrBppdvmTuN2KdOAxLqevfAsPdqxUVoPwhuk3SyJtyJuTvkwEO+21MXMBP9cgzI/On6
rK/akM2CyCpWm5DDi6/I9MsJOjPivDFk0o8jwdjB4LoftT4xyrTcrb2hVztcUNJVK2WEqVIYGNsC
fEMgmR85N5bhfKYKpLbTwOc+y7Kf0q4MoYAKnPlVK/OlFHPJv6Ar6D7FTKFt0ZUO52TVzNUwyqgd
OrKfRvYzkOYNNakAqbsioQ6uGii5wl0P5/PfBHtI1i3xcFZlGWyYdMwpJo+EXKtxExVfrke3rVBt
KEHlRjydigoXRLRpw2dDPq1pOnt/RLBPXw+kVRo22Bfl21/hDlE3m7DDgRWdT6HkVTM5hi+r7EvX
ZEUDVgOJDCb3LHkiMBFYDj+PkQb4jC3FkUvfw97VsscoZMOkQ7VFPRGyj4XIFaj2o7alXcfaIOGQ
W7EBR6GlS9W9WmnCS/TYL7tLjw2kjd9ogAoZNfI8kLfl8bO85Ot+SKQoAo/tD5vnrmFFGPLdF+N6
LkI9HkQPk1qU2a+1emlz7Ui7JABNITx/qVXvEj4e2r+G9ifRX3K5WQ+NL7V+cATc6PmN3MFgQCCY
4Va8u4SOig9C/K+5qNuvvRTpwPCqjrgFdchO9YEKSeSvpLLqDVO9uzeh6UxFPms/aIo1U3mqjI06
wesyKL1vL3WkwRUrW4lmBH3Zo7Kg2SiHPBUaVx2GdvlGi3eRJ+5LnsqS/Af8eqy9INtywCs6jW7I
39dktKMmVbJyxy8fnRMLoD7NQC/bQRPI038mPRJrYGqOjhOPcYkJfQ0ZlSE37ziSCU4sjf7IQgLS
aA6msI+SsOfjU2myi0G8NKY+Uup3RQT/gmnz5v0YsRfX4H0C2wcU7huznfj+yUxsOS5nkGA+PAEN
u3Kde9xDnpPPf9DvF1c+1qsfiHasaBB1thAxdDUFa7SdmCeI1dClXPJFMBdoEHMSnYXA1ThD5Ss8
iXsnyPdlKsxh+kAtVrehyCPftN8mrGdu2hFRp4HtU37xdh6+hfRD3d72urpbVX4raCHyH8y3M6f+
urpxzSnvXb2W0e7Gdf4dZWsRneNrSqEKGwWyhAmd5f1GeleJNw2rzNb21+4fNiuuJqfIfMWO7HMo
d2fPjYYCGDBTIuWolvu+KKdXUBrp/UEiuBw4kOL/+YDucpwzR8tWGs/xlcBYcDmpmzkHdlKJ+LmZ
p6mGWcGVxHtj5oMXF9YK2xZsTAewiPbzwMbRgxHRB3rWiV4jNsXYw1I5OfgAY34QG+ZHk+hP1jud
RuFkhR/yju/epaxON8DQmCl39kIK79QlSOT5rmSC1Ru3B6hMf5Bw3oZ0LMZInJGC2pnEzqQSasPC
aA0Hu3jUr2vtbIV/bG8Cmtd26k/dMv9uvEaY3OR9wQ8cu+kLtmTd/XiofNuxbnjMIEOho0c5hdqo
IcHjZO6GDq1F+JXJLWs5UcD2pPaSKICOQqQrWb7dSKV6hrxBl9E772lwuM7FFxp2+P8ZCYcYxd2o
gsKr6L1gdN+vpByeFvKhE73u9QkuOEeL22kNegmTjLgrIxBIUrq58tDSZbH18PScHbSsj6mfKdBy
8w8Ua7KQKs1DvoqnEv/CnAgUUphRkJsSFooiTt36rjgc5TItsqpNUqMLYWMhi0PE1CVxaqmOnTKr
viv6aftWAn0ifnz2hITvgtiObZc0xQkX26mXXdHZ6O72CnkoBrPJSyUQbf3pDWg/1YMSuFYwmCFF
dTdB39uOHAixpc1xQqbIryrYd0725pHjI2/my1LWq18/EbNiH1x0S+I7+0GiTxnRIaGLrQGGV/xY
QESDk6EtyaKS83U1C3POnu+mG9zcciBMROIShOPu5J3YVzw4IKkGP66ElToRIBqW7EbHoQd2u075
GMBrDA0oc2x7LGVDWQ29loUtnPH+nQE8iZElfssn0S0zihc2lA99Av567e4bMaEcTFz9K7/V0Nx6
ZfAfEp2lHlZITRrW11F5VCHgUO8fU1v5XuHUlrIinzONzTfZcOpudoLpPzSCl2tmsJvmEe931n6d
1fWx5HxihsFNpfW3eUza4PY7iPfl7nDOe2Lgpr+D8+jzH0uGcz2TA4rM2r7aFssdoMn14F/X8abF
7dncYmuTdov67aJlc4LjaK3U8821BGD97Co+6irIVozTnPHUfh59o9Y2YBpqg9rhq14cpzgnqREt
HrgQcLAfiiTOIj4BpcszSJzx540K8YxRA405rA2bkeDS8jJIEonB2WxQdFMib7ZEj4S1OpljRzOH
/05uvGS0K2dUggMfGob6cILRfhnfyMOAm2G4dTHvFhh2FBgPjegN5mKVzCwGF/g/tI7DkqDa0j2D
3cXTXCQGLGDrHarZWCTz6jqN4uM0yDJK7OiuKyPRicCxeQWE/uNCVuJYfTSdqrFtRbFJJzguN9fk
fvYa/8b8+FGgg8UWm8zfCFTRGR9QJRx3qY5o+6BzBBgargR90DSHOHMLdVD0AnsFQ4huojGpv9cq
R+ZpYg66/H30i6kSbb9ojmSJz1gVlYtOiVOp83fYxMQ/8uQhX7pYdRdP5cO3C7+Gl418XercE8Bm
/Lwq8JI35wXnzHSgUiBmZVGVKQs0nSuvxfOcHsGTQsSErd9U0X5FUqU7w8mEzptQzg1l2ImKAVvL
xRCkX/tly+DWhpF8+Fn2xt8P2wDA70GBdKqN4BEaU09WivmYVqDFe7FCiyHxW92bWd94/FroVj+n
74ko90SUcbZjwyUjNYi12Cx50am3W9PHN9uTXxwzZrMz3XyfMRkcxkEZf+MNkwnA2sU9cAwToQkh
o3gXOhTJ42f4OvvXx2xNX84r4lqNoN9SzBmSOlz5yz/BKC6YALcVT5v0nPUyboHkA9BFAJ0NxUIG
tHg6cvGgEw67E+RUddqiIxF/D23NZ5bBYS8LCB2qsp6tO7gfzKN1gINYgqIJjmZB/eE9dg4Blw1I
5PY4q1o4jKC6YLJRIKbi4wMNaoYNzKXCQq4IREhQviAF5+eMJTyUvQbVnTZXdV++x1HE9AHd9dN/
fYefTWsrDUt8UV/yN2me7VSwKJl/+KoA1DyGr9qjsjEZdZn9QDt8Lk5ST02Sn46J970M7SZkIibT
gL73GtZudMIQpLjPn9Omr+5qyVtU3OSb3PDXMwTX565Dy94DfbiZR/9uJ9J6pD6YUz4R3IxQCWZ6
/1x2y+6qq7ConkhoIklCM8/3vDwUoqKhD2PMpIZPivymxh89B1M2r1blSv5Zad3FKdxQ9jOu+Z5W
VLdN9YJtvTaHf1af28GLrW81gAQZ7Zvf6r7ozOyGvtwfVKX/sdPSH4+1bC3RGZL1e4E+pBWkpr14
yhJqVb6y0VB/Xq43KnfHcLbsIoZVq+WS3dSJG/xa6TCrGG2byrjTon0mgYdEme8HXf2zoeCU2eP2
oMF1vUL5tGwCuZR90JzepG1+LNhffyrhL3YKLyipPpfhCQvx1BmOqxPlyYZZqPxQDns7LDevxBjG
Tf+8B9lkBG9PgIFco53TOnUTrkw2TAhF3rDt0XcJUAmNI8dviH9eVXVpM0AfZVZH2Z+WWOIdbKzM
hHkHj+ehN01EBdrzMjko3u3YYwvbt/UXXq+4yUWOTU5FeSkU0vFnR4R5aRaTNclfRlnomMy9YG5M
gODheGs37Llrss5uJV1QPFCLL1026V6wMWRUgUTjMNCRAFNFYLG+FYJa0WbgJSyEu/l9izKP8KQv
fBy2G/lkq0jkmlgAWwiwKKWP31nH/82fxxry/UY4YepAAj/0p9XsJRvs0vjXOQZmXu8FgLb7ahEW
+JR8FyrEL7XGKSkdUjON0i8DvjG1Wk5VM6cwN1a69eyvzAlaSeuLJHdp5nv8ZAm5WeFKxcYYQOH7
HW0wULr26qVNMlX29bj4i460781I2rUhe1mlOGwPL5RiSZaVvjgUh/W0q7zL3AU8d2vqpjyw47Aw
fbcFc6Pwi9fneuJdXUeKL93dSLEZ2Y7m41Am7W8v+SQMKvVUz1m4Eq0X2+ApE/H0NaN7vNg8O+7K
9EuEZiSv3nBkIUCH1WYuSuQYK2NZhtJM+GVBiEegZdr20+7TBwymqD8scKRM6n9WrQuchMC40fSi
mbpy2unVVpGjPB9TQSxlfXDS5EAVkuroNAquPzLABvLyJxJDI/e0FOJQE89lTh91x5H8YJS/ui7/
8SoACbgCn17bw3U0th6CiVnSDg8eAOSShMyY107TCKWBT8J+6sYEVOYhMmofi2DjBVUYyI72OTso
d2K48cms1RfJNacSX9YfUqLTCmnGcJIRFDZ2DNW/VErETUl026xVeyT7gdfwY4N+kLwq8qKtOY0r
cxYOZosxRSJ5700ZXdnThKXxael8WhB/FjemDvPEzmzvcNROGuTxX/s5r51V+yizEc4m5ec5ZdMt
PHIiKV139dOX/XHzr6eINSyVrOahNR7XlQLobpgFxnZnDonz5zHXRRKn86pvlOPsEaS4mcBhDxA8
dtKmN2PbDMzs5LGioGBTGESY7bW3rui1OteuXexzJKiid+K2smLNq02gfVWXHGiZaAHmFmReU3ff
seVs3nyHvbIz3N8UT8ly/gtfa6QQLGv7r3J7l17nOA3+kDiyPE8ffbKhxRwwTdJ79ZgRUEIOyDvN
5KOP4LSvdGMMxn3JMH7dDoizUKmXvD6S2+3aF5TBw+X99GwylH+7GAEKWnHlj3cU2bx6mvs8YjeO
U+DiLVwt+WL5oe4mde/hVL9BzyGMS51qgo3C0z+9OFZ495eN2WJUyerqB1jPECzjm7KZL8a3ao5i
FwZC2OQjO4heboJmmn9blhyK2YGUv42eo0EOxag6lFkrzoaYJkYpualCl90r9Dtngb+iZenruL5A
RiIO40dUTNY9BKPqaWQnQptwFluc0SFqlKrzaHjWieucSpPl7apoEf9Lb1dcsChiZMfX1LMfnzG+
vV+mO+QsL0f94rDHSy30BkYxBIlA4o02Q7vRiKGcxMoWzRy95YIOHWvZXZ+UuHLVQQNEdmM1ea2S
+HGdPVHMdbEaMFXAxwUJHJM32efYmAAOpjAIzol0MLTMRf6tJP2UDYX3hB7ik043WyLGr8sqJ5XS
AGTqBF0lm55ahM6YVIo9eSm72B1Q31HndB2hDKr7mzGxbCQ4yAawqshFmts983B6lV0/jNjAYWk4
cSXKVnG3sNrUlauCH97eT9M9L+wo7grxE3sOZUDZdihCJjmCumpZioExC1W9BMedwmzZhcN/Cuto
pwoIgll04a7n9FZTl76u0dAfsxXBnxetoLqlTY16bwsdV0Bb6i8CCsMoSerQjW7PmTRbs9zbtYHa
ZUTQNyhvpk6iM7wziSDl16c22jnJDhblX0/BuOHW8i3t+DsiWA1OdRfxWwEpUJ9gmU95eupE1O2R
2kResOCYlHGCTrHSeLOB8voIbmXRs0wL48ZGNHeJxCg0gUGHbMTObL52tRVvbpZM3JXBqUazq6B0
ei1dTvSEugNmU11lSI4emjhC+88fNBrlG+1vzNRAhbXOvhOwJMnp9p+lyJll2qNwoqA/4Qiuqbes
O0leeTGz6/ZP7c2CBEQF37v1AJMybnOxeiOiCTuhCactUfEEX7vtfkC22tLNGcx+8Pmaff81JKQd
De/OOyh/iH+KY/zsk+cAbGntqdED6lwX2WniYNOoN2pbK9Y9VELK9omP7Tzy/veA+csa0v39YVMj
+oSEJoXKsmiJWDEGpPfF1RfYxbIUlOtjcpCAlnm3HEnsanUXshyUCzR2KtavJzc+WYToJDuFeKOA
Lpzqw8Ij5hK2wfV+3snCcdqMo9zithzQRmKVDp1RuDtcMmZKT4jCg5DoDVMb2x573HwgpDVKf7G5
2d2JBMEYVMv3p7P5arKkPycWCkphsAPTGxA7oz38zSfRyQHWsMawZO95n1a4c0lgwKMhmZI/MCvF
MgYMANgIvEYGqitx1nL1Bdo2m+5NFVnQvcAcePZ7RduK8qIHhgl3mAKfq+IiSqN0seFpAH4WZkvr
Eahf38C11xaCyeKY9ka8v1qcokPkgi3Bg5LLmXZzM71bJwum3MNnjki4gltii0zmtWnVc59pEaJh
JNDb7l1yXB4OhKN9grazWC8FL180tAfiUlNvjY+I3E8z/GW3P5OcEY147/sIIgi8rSxYEgKJVfly
5qiRV3nDGlimjlobKbY1goP1SLYhldlBD56cqsx8COuyFgpEqK+pLzhUo+0zozQUYtYLxTvpxMQT
ThOiLmd2OTEKV7bkb0jNwQnDhnOCMa+Lw3Vy51pBAUDegy0kaHcPgOmASYS8f26NQZ0GVSD4ybts
SYZ+dXUwZQw4uFj9LDhd5ZwX1cqTvSVdsm6weoE8FgFcpeL7hFVRSXIFZFwtSJGmBeyIy1p7EOBL
jVxo1PKki1Ndm5nK32tFd0qW8fc3sFuk/ZDcmMTHrmmElE45gBWZ2Q0ck6MktpTNg8cJns9r6+MX
UJW/d+4DH4xSj/3v/e1MaAGtGab59KFD/d1nyJKmsDLi5cIB+ngqHGVppg+iRs8J68eGQ4/tPHKA
YjgUoshle6I46shv8XF/iIPKAFpVsJHCCiViBCxxZfA2scjrMnWFkDs3VuSCjhO/XSjSUJTxGkRQ
c7UlYWQvRNw6ni4aHBrtK6BrAQGzBF/eZ003tbXqdGWnUmOpDhOhY/81rH1OSOzzKCv+foQ5ncgZ
XZCPAfWnENCKTQlgvggyGb0NYOwG/OLxwpoqr9wo1csPE39S7e8ATtMCd1y4O8SWFmdJd6gahjwp
5jAgCNZf62K1Wfta/481R/EufwZwRyDu2QkrZzIm3QFEwEkOy052ifZWjrwtD28mshO/g5MLC4Yv
tV3yE8V7KfYdRPspH0wjOw6X64e0l/feVZf40SzACjaPUmeBlFbnkCxiJ7wuFh11ohqT6fSI5B4S
UsaBojHDq5yaQrFMPp4WZvigxpk9yg2tlN3DPF5RIQiri00mJ9yXR/EzG7Ny2cb36OM34rjJ3MNq
dt9V1AdCvn9NcbZZLWn9fHDhjxoTGQ3xdcwL1k3pelLaedpblYWhYHItGxNXiNUUyOgc5P2PeXB8
4y/5JS6czay/sq43on4Hh5CMsBbhgJgrySQDtRXw+/NC04nEjBhmDcVN/8WXdgiTVDuKPAWAmn+m
1D6JQh0RxzjcGN49Yt9LLxHsdTOg27QwidlhJIScVrVDlO7/5I/o+q+b4qx0eZxZztYeScPuy92R
JcjXTOAWiCw1B67pzTLz40YGfqF2ybBgQQQX7fFt1oQuL+CRoHhttDCT62QRnpgNtLEG9fp9XIOJ
dMJCp5p9Dusjoe4Kt0Xk8A8LdsbQDgyiYr4+Z8RRh0Tc+PpEeryGsXMIvlSg8img/Ak4aDgMZFHM
TBO83RG0nITcZc6LS84mktEQl+swMzg0mUWtrEoSbid67i0kGx4HQIFSh2fIRYYz6vodYQVLj8+T
C6yUg6cXbN2kP2eFMehP/AgjOfhQYqdzynmHBrV0bj7/QP7xy6kiTvUo0XKGCuoYGec8TTaA07vs
r2XCQHjTbJhD3a9v214kNBTjPRYUiiYeikGRH+rUTLeWg7QZ/r2GABIt3oxc+AytF/lgc+EVomWR
67gxoLt+MyiZmRkcSnDr6zC5BFPHR2Dx4PUYBDFcB4bp5Zuek+vGfOmeCGvBNXNW9fWnYSvA0DEn
INP6O928jgbTGpZNL3bQJdxQsMklAL77iDZgjVZWIB1dSzl+SDTeykUlBpa8IMGEtzh4K8qMguL8
Da0WE4SlUtTad9fX1BbfZPREs78HVhwTKD8OTslYvWQHDm31WCI34oWPZQLhxNh93NZL1sjsVNli
zg/XNTR/QTF+oYYfuZzXJGa4stAvFWwekyFcJRW9fFmESB08kKC0NhQWpRLbUW7YQkMF4GeUUYT1
Xda5fw2eghOUnggtS6Y+UrD5YzzzEwi5DgnFzffZB1EwFovW2EJ5v4qD/GftMLGnsxvyPtMLcU20
IzNE21opBn2D4Ni+dMUFqRsSBj5y0bRC/svYudJDlS0FsndzT82ghBc1JdDzdWU/fLNFJQPaLSP+
xX8xK6oz/u0ZrlbGRHisVmCLiT8VTxHuXTQrbqnZlrym4nQtCKbGXsVcT1wNI/jufEJTSgX4QyI9
yXwbbTumioCyjXwUzqTiPUJKSPGn5jVxgmZih3E0iT02a1GLGiB5eZyMW3XIXeTT64RSioHH/Fh8
iS8fybeAEmMpy5px7efRDULQmBMDwJ1w4JQe7KnCnPqigEjGDa3YzWtI3je2A0VQKJvI32IiRkjN
zzsq8ONQhr2xQ7Po1jYD3P0WFiDRqH/CVLYU+j1gabE1taYDLsMTp6G/08rMnar72uF+e9DO573M
JwujDErDHcr8JZhbZbS3VUMqbAZDAY67sT3ZkvhiaUbkehCYZB9jC647bdDUt64OsLWJxroTWNT1
VwhjIwopmskGN8hQBFZUwsQQmS55Q+AAVAJwQaAi455YkqV3m7y4c1lEQtHdcxq9Bk66DTpy15f3
WpuBesbg4GJYkmJ8iJiUIeytRWFrbxC2yHMysRhnv41fV83/RN8vdWEii4OmpquTarhgbS2FxvHX
mLeWg3c25eyW3Z6/WUID+EyRgFyfSmScNYYNqik+amA3OtVEB/Bch28rUmWD3BwrcwIp2CjFeuHz
lBl/qPDen/5k/QHjS+NAscMIGATp57ozB4q/2asHFacrsIUCZXINNwSuyRqhhlm91V5mu1IxmcRH
WswtJGqG4N04/1Cy7lonvf+dQT95cvfkGO8M2ILjR5jhdsH8uNk6qr5jifZuIPDwnIiKa0K2jEg3
lga+arOXtyNAG+3S7SrJ4BHFh7kY7g96RKBDISiO6uVE3FwLO8RiuERz3zoIEJN+IweLgJrJLS2/
3iRFzvZmeWfQOjC9iiJF87gA6ysG97x4SCNruSza6ryirGzdQZXqFcLjsWPQCdBbrjQNVbELcnUr
/dTBJFaYZDAYEhgJL+lixLrHbxGktWfYF3AGBrxpsMrgq47v2klZk/aUhqg5wAWxppZfKr16AOjq
fLdyrx4AMa2eavcZRAExJWLbejkXxUFYItuNzfFG/l4+gt9ASyAO/yVxlvxtEs2+tWD4hImyFjuY
3kalTPZwGg4OxGs/nmQWzu5Avaq5on4BTiH2EEY04g46b0refacrlD/tHil2b7OwcRPgS0pPOjgE
KcQKJ5o88nHmGGkYAAjMkW11FiBUVayqmT6DTh82+f+ax7ngusX8L0TlHmytPWIKv04iufgRv2cK
oDPT15cWcG1WKnWpoce1NtLqQzaQXueAY9XwApa4ayfOXqA/R9s5CTHlKLxZvXmRSArINxmXGp1B
4aZUmLSyPZIGwZl2IZ0pIfeA3bk/+F1VosyJh8swbodWrxjpMalBLG9W+RkNL03zcZq6iQHOJGQj
tTdXDtbwTKsaiIThJEBwrvVyJOtQSfDp7/5hTGLxPvJ011s8jDjHIUYNkCX7435r01Tb290GtbgL
ilACLYf6NFka4SZsG0la2QAdv7fCvlKt0kuYhe6fJROobbJkdsknrnNbbzk2LjWqK/TiSB3h/Kbs
PqsXLjXvlLI7L8E9Vsq9hc592bHdPHGbN0npQOwbGii6LcUfc1Oy6zfGMJEjFpNoVGJhBLnTo4UJ
2Pn1YRtTBcQpeXviy9fJCEasE3WOFAqyv9rcTE/IhGjiWIiHh4GrTbggbgUj9FcGK94IAO3klOdR
yiVnbv4AaZpqWsf7js9bKLz27X08tzOyxZfnWFCU1jYi3Sg7e3HOBRjSJJCQ/lodwf7PH6WioHgG
rxObCE0d1EFNDt+9BkN6k0BP8g4QFrIE574ZeJGDMP0x/7YXAxsvuRObQS+RGeHrjoHpXsLLD6kA
/y7whNBMXe8g3Ownmw013ixUn2tTbu/Wic5OmoOXElruK3YKV4briwrNT7Qny5OdZEnTKv9hxNm0
rW3BJd2/0wz026s7WfblBWDZTBg5XfX4EnBtoAJL+ssJnot/uIBx9pJSanW16f1J/ljLREsDgBOu
0vnHb5TDbocIf86d3BZwKypOUWjFPtX/iOno3yJmbIHJb0yK+mnRaqsehUcBf6PhGlmgCNAZkWaF
im3xQIYDI3oFJFj+DebMDw0OfSG30Lqm/rqpcqZnLNO0IT8bvAPGZaHiueeinekptwCgtO6BspJ3
9o52Y3S0z8FHN8TNfFEmxcHZuNmkqOOOgEUz5vAp1hOiXrYXx0J6l1MksDCAeBzLrOLofB6NsyJy
JSRU3MQLLv0v2xQ2n+uR8nZHroGmq4sxis6em1uJDMkN5lGfg3BlKJ6PhmVBuH7rsVe7DMsxuvax
YDM+7LULAypNTzzVFFE44BRtITxl5hQf4NZtJtSzoWf7ZvoCS1gkuWi26OC48clIVrLubFTx7B/W
8KRB+3Gmx6sDUSLrQpovsiSHv7Cr+HwRMTpk8MNYVgjEzQXfiykR5fmWKwa0di7gU7S0I/Eq7tjv
FB+1ziqkArZbkQaoNe2jitc/FZeO59L5FPltaFjt5Mj5RHLy0nEBzc4nzt493rcBdzXU/1mqRbxO
9sGM1TD2PKqdFR4Rv482An1dn4tCaS7BVW5krXj1tIihFQa5ngE6xtegDceze6xPuStPowop6jmp
JBqfvRyuY/8e/ZV2SJm4KqV6AwOzWcubeNJyvqy4eNQNJiINf8dH8abBDc6ns1ZJCoBixGKteasi
wCfdMzkUYVU0ArNSB2ZRrfyJfBkE8vi2mp3ApL5w0gYuE4Z8vItLIXmgEbYe/RPwH4dpT6UZBIWy
5X30CptjTJak9VeHQxPH5e805gfAtToXVFN4elM0iEN9EYRiXVzU436J+OEHGSTOsBgrCNBC4AeM
MQolUeDNIosbzg090p+awO+fpL26AjClvK6jiOXAzZ57v9kmGMuT/e8nbZfazRIogMosw+bREjmM
oOZ83iPCHg0E7PbUxMaIOlkwqKnpvFxi24U2OmCfMRU352k0CfCngUIK+3b4Y4f//eBTL1MtgT0G
kuqcyZoWlAwcsIlyibwTpXSYZSIcqKWwx+FJbLq20UfDMg6dtnYQx7SriLdVD0NxkFcq9E9kDRAH
4xMas9Qjp/696V+c3ayvOfGM8n1Q0rKwgp7RcBlqqtiORDZ5uXC6TDlchubZQ4cIBxjskAlEsxhG
G7vKQjaI2CutjSfRHUckmWVmyYsRXGDfl7T0lU5Vs+luJvndXOCTaBe4An7zdURsOVrkAuHN9UZl
Zyp5lo8+dhxuZY7+iYxjMvhKv67y9Eqvv8xwC4/pzXBElnG4jhBQjkEUXR+fNcQAQCAsxKK2vd4L
zbkbj4UQkQaWnvP5flb1RFMzO5obU5nUWu4s089aFogoZr2UQP0xwlnMYPFk+z2pnNF8qHxnsWTJ
fdR++5Sf8zWqdsfmq18Q40VuO7zm+Q7iIUDBg17l64SdXcciRZfkwks22d2PHPTmXDxXWW8vlBAn
o0LhI04SJi010FYzl2X78CZlJ17Yzq8cgsGJXgg/LPI1FxLqHddItKyizwRsC8FNlOO6OnKgr01J
yMKDExJdRFW1tvMlb08+Dj+dIMHwWWiKtIap1OoY9lHgwSjqAogqR6TpvISeBRWDXtDWhK7W4HlK
ElGU4cakhjt/J9l58CEm6I5/tNtxANTLatKE2QUfglUL+Eexl5zwFmQf7x2o5c52GLSvxclRFUjQ
Y08iw0eGtamNPLm0kt7EFYvkltvDfi71R/RtTALuqNtwnH0TIYpvkVZ6juZs4DUgwpInSGcduD5r
KJ/sp3l6ovtb8BPYRCEAnHdQUB1qALU/cTibFNdVn5SjOnAOWXVsNevxX+f66zkI2R8l6e2UDmtF
ie0pQ30Ij6/JZAjwOM8v/FApT+YqT0Lu9gEf9oMgvDSaZDai9BhD47txVj+9Bogtiq8O+2SXATt+
gLs1yNhmuwq6zRI7G03rt3Ayp7++KFr1CsPkxPvN17KsK+iQGz4K2B83nKYaX7lP1TVwknYiYFuY
kX9stq/Bij5qQYy7/N5T/JVdA8W6187KhqmOKxOmeinO0b1XCpDYLO8ahkWOlSKfSzk50Mx/smFc
4ue833DK/rNYzR8nSMVkgL/yjWX8F1s0vaBH4ZPMx7z6cCIZy+yztHhmcFfB9bbYxL9qYOGPA0pG
nJIVuQS5eVf6Qm8OlG97i3CJc3INBFtIg7lISK4JqILcoJ93IbWNSY/+XVzmtrOttPYh5q1p6HGi
ybY9rTy+lPTZUUgnPyd6A9TstUPpUv3d/hUWRQiZkE4//lL0gGy2pQysJXpVyw7EU0X+hJvgZ52Y
DvMoHpAGTBmfl0sYqtY52mEdlthFz2uUwy9Lr+v7rXx8OrFtA/FEqd8y4T/+LXnxyvwFUhCk3cZo
o/3aOTr8U8BR3CYyCsTEHI49UxEb5X1NXtA7Qqimifu+FOEEQdwKQA5KeuBmw2Rdzcx6qJ7i9TDK
bR7xf01bScD3YITQ6o6+nnU7b8QneL7AVERW7IxmvElk8Zmx2v18nll/DOnfzD7eWMk/Z4hUmLXt
wa+RClwlvwqx7h1DoLPk+fBvHkOqNqeKDE8UUxOJd87EDHmApBBMw2j7RshH/ax8lOPOYy6EJB2D
CsVRi+4UnSmc8kw9PkeUNez1549Ysk+xMfEmCMxld/1pmb9W88wFZrpEqKAEac8B1psEYcl9dQpj
S2Ru9N/c080OsyX7Lx8F88sXu1vkTXWh3c5quPQyXI7WWcjr9t0Bqk+7ZogZPM2GfvV5rU1eEuZc
3u+L09klQd7SNM3759AwkN6lPjOo4dTPPjqNNKK73/04/0E3EZgUo2k9v2fFlPU4yPSTsv9hXGaZ
3fqDesj1owvXyy4bqxMEUsA5ttX6Szl8JhN5ErB+c6F6fXThgEnhJCfS7HoAf1vmocZ3BtR0vPtZ
cYOffs1N
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
qslF7KNd775G4ECz7UEuihip4jK7tstNRRxzU7s0yccvhYAXDrmOYRvykUMrsxFV/jYwae457Q0v
eT7AT1PqIO/r2UZGEg8uvyDbk5lveFkq3HJEKyAL1fC1FnBVaXQPolewryqEy0pEH0qRhJwiwTlT
cPrfgGmNmlbc9DA4LFGDoQrWve7Ci03Uj4Z0fs1zAGX1A6q8LME4/HHbvO3k1Pq3mR/ipjtDu2jF
PCMXztvvYbRTWMowM8zFeG416PuTAHUaNXvCV9gucGZS8PBfRaU/DwRpLk23YXVJYv+FtXyJ+XzB
K3v54tEwaSMnQ2JAFZRR5EONbCWQBftU/LBd9w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 9712)
IOdmMDLpSo7jezKseQr62SW99Pw9jSwrFTW3lSoaYa59AuxKU44X+nonW5eHA8KmQJPkxJlZ751r
k8ucjEiyrENDgUrpaust6ZeJ4HmxOg8ezehMdD50I6+WStir6fSJdxPR4OewgLgtwiuiwiJ/5Pm5
shufgY6du7oNNhhTz2ylzgf2XV5rEOObkdjKKTDV8VmCi3dCdgfivJp0tUHeaW6LzWXEMSwH68mk
TNEAuW/D9VZLzGvHSk6lAk4oQR4Hh3t07JJSawiZDIiaPqG6vAZ9KYRwXO3PkYIkJAnvJSlJWbuW
z62JDUb3YpaYIQWZCsa4Rqc8uwAZvdjXYZJl3izdyFNbupGYA4kM0HVLTPOeP1q8oMeQAhtavEXt
uZKto0R8AjaOKMDk8+taoQ9bOGkFRdCG/9JoaAwpXcW4lEqLv1i2Mtsi3cOtE8RoJJjkhMsFH9b5
2ISrVPPkLXhGvUB3Y/2EqBMB3QwY923FL+5unEJ16fNWuYBdICpwwdsJMsMw8OPma5tPdv94/cd7
10WGSiwrplw0kN0ObXVVPwgLQJ3sdi2nyChi2Xl8V1O9zVR3tkSsi/pgCX8t3Bc91bA+bplz4IFq
0lsoXdyq2IaJlyb/y0x66UZJOHXIPKwED/ncLUeTwihj6gA56IgJVcVw6lvNttvrIC2DnDxVeh2t
J4dTS2Q4LfeCGYL1AenhP5DNpdqurBK/jUJqbYJcvbn7jx44P33fGfcokvXhwOBT0fvmsOtOOCcy
wx4mQMwgcgur6RwICpiME7IsRIMIIiehl1v8PeO1oYTm2/hXdjNMVBDYM7GOcujnUj19JQswwsbz
Lwjq/N2Bw1SCVZSGSPh2qJcpYgbR72V6/qcMGj3I+8HrYLPNc9PnecEBWYRh6O1+KucsGjp2VtIS
Zqm+0ICiULg6S891Qn9P2fK9THJenyUk++KintIech8y6GBT261YNiOx9O6//nAQo0NWuGJGe/0q
y/ZBgscuQEYjb2RCffbYF9yfPIlt2sFf/s1M37mFF0+FN7DqH/Kw4+xBJZjY7jAzYUidIkkuTOyd
e5cPUZHHrccuwZl0Vik/exT8d7hkNqUzfGWWWcK0PHIzaqAGvetwZpxs11bRA50V87dRCcX2Dmk6
WscvDBh6Wfv6yeAOjhzzzxfIA4//rpyoN51YOBHN2MpStJtwzyguImkKj5NtXfaPgR5/RWUbpO9d
qo7gcJAjETiBjp43fxhwaI5ZcYG6Lm1du2MNgwQMZBzwh4ccMDvtSxkrhAv7TlTkHPgnqgQxGosm
Y8pybT+mBrh+2bAiKdt5IHXzO8HjztsWAw/A5zsH3tQXJJ61NiWj8HvKrDMHQf69kBtiTajUkowo
xK5yP4FXl03fGUbX4Z4DoAkmmsbqNjkoH3bsaBkEJ20V604cqpZiLHGHS6JfTBEx1WQU8Ninjqpg
nAUdAP4LhWhm+FTyeEZQmTqVrkmgyRRfgjf+086qmBKoJXX7am7RzKNxRGLdLecuuObxjMoVwOYG
r9rXntAdjVP90oxHLlDZep5Z6O5jvQ/uUwsdC7U9fVRpf1PVdwI2Sl9xBdrfXH82+T2esoMJOCAa
LED+yioEY8xM2rk3Boap4PPlqGW1fMNMO2kpphKkXdR/ASvYFFasTXpJgBodQsqZboICemwtd7nW
Yu0fG9ihN/23IdpG+05XlJn/eSkiQcyVYKbx+lmcPjYt+pq4Pt6lXtqDuXTk6dWa/gElzJ00Y0eq
HrDQoT9YZoEIXDxurvFRelNUaDoLrT6PKxoXl+b52M2IYeL1op5OgZQi2ZsCfLH1uugUd+uE5mbs
K5v7jGr4N9J/QDC7VAum1hqq+XiLMts1Ptq+n0WUrOzASkybVXE9p1UTHLson94xfoWkrrRfhu2a
kLVEBgALTRQaLuvjGduYlL/DD4I0h+1mL22HspqqIPzv3301gPhVZxBU9ok9QxVPw6Rehx9KxOdx
1WFOtmBlBhl8LCShlZOwjjRxoMLFVHgbX4CTOwXO8LOZccrz3QbQOvGoY/SHM8o7WaofwCAeM5lk
xpNktpLsN/xFWUxOc+EmfG/rPadvnWISmWoRBkmXJdhfOqgzjuiIVXqMLkn74D69hvkl25d6bvjI
1Z+kkBMzzYXyN3PCrKCfju6u9tv2Zu/xNZgcVwLLBfJofe3YwCBgHKmym70/0xkAl+f/5PKIJJ2V
mHnFskkjEpB+6STDxpN0EgGbntVCbb8sjdB7nchwm4SAreCTf3+WaX3xhyUvn557+c/O3D2GBPGU
1byrDl+TiAHj1dU6Yu7gq1IPTONDTEs36GNGxsKCF5vhwvefEX3U44cE5yaUA0LvJLJ0Wrgt8DoY
dP7axvIzLrxxgjNxwqyk6QOEHwMF+BEhqSQwsOp9QZCzIQdjZhMX7NV6lLaZ489uZMehC4OkmQAO
d/NsMjErA33SqZ06MZqQlN9Qva+6qpNvK1tFerkyPb7/PmE9RSPhDNMGZpl+w4O6jGfxBR30F07G
al6G4xMfvhjGaQn++NBSGdxNT8D1phf9O2j5MtMZQwqde+dXJHXltD0Uul7i2Jl+aiBS3LjaokK1
TfdyZvlneOvJjkbyjHgRvWlFlkjQBoLg/WBagsai1hvvI1p5J73MpakfIjBamNM4S/3z0zs7geu4
sK60NoBYheVIazpmEzRW2BuYNDtF+lCYC+bnAglRyfgaZ+9W6oxKb7yyNMhyKuyVRu0MiV8NNYF8
01hxp3Hl2l/9fpNqpYK3HNt/J+me3yM5LT8nnZQ2gpBZYJphvrptS9witSf4TJly85eKgME53rsy
zQUNc/hf+E/HOyoZPL63CDFogZeE9JpIGhf4zTdya0Pa+zzl9Itf7B9jTumhk1Cs5ebV6+hV5FQz
g3RaYxzCXxU/HUb6PqlVVV4CS9IJj+eNp2RgOqZTSzAfG1oVLmuX4MoUTzoCYaCWcczmsys2ZhDL
5qHGsLHC0qw4mQVCjlL0OAIu8XNkgHajD3BYAUDXUDlifDrfobl5nob2jyQiEa0H4HXyAEikZnQQ
t3aHiydhn77YoqvEszRE5/0h2iNvrU3WFhEPY3LWYTmkEdKitQbQxbF2O2aQYjy+69SNAcOiRndd
iMLo7Spj3dr1WLFEOzQwyc1eqOMNVsKQknsOKPKmsKWKHHMqnmZu0pBZnJjs34rIIh+UhSdLA4XD
yeg4Gsl0L/Inc7fC6S52sQkW6OzwqOHWuv0iepvKP9b2Gj5fnWwQiM9bSj25eNkUfGpZtHkcXLuD
V0CvfV+njLneB85j8ZcmfM9w+9e0zKG/FLb7I3u+tgVBIXquGU0LQ1YvqIkI7L4hMcBAvcZEa2Qv
pHY8o7bh8Asurv2m3pwrXAB0vxmos4mlbPj+rJUFjtS4tCGTiAg0vjG3/5+V4jsdhZ97DSteyzlb
5OBL1KUIvBVV7bOASR2bD08dvNJcJcwgnH3iUDr6f03Ln1UkJezm6/6nrYsZ5bOUQ8PYsXN/YXgG
pm6Uz/SzvK1aaKANFuOlETZr2EO7J8ZUfSwWSXaNK8tDKButZ/DYzy4mxT+s46a8fHE1KpZkZQND
tJ9hHnRyqijziB5ZOk2kbBBRpUhJcZ6KPsRdSJhU69tA4xyCaYNYDygMdtlcBjDsri5b+QNnvXf8
omvpGC7HdGVwD/19rEonviZTBnQaNXTJDVQgH7V9OpnlMvV5diHyBC0XtkBrfGeBf03cKCBibVMf
eDKWbJo1hL7n2HGhIuFoJAuS2bDU/yJF5qxtBi6Gw4vXaDggMNqrrhAcgnm07m53o2SkPS8zt6Iz
b/eJv6w6/StVQnYZ/aomkM1aQrPBq4N7ujutVhf4+rJqVe14A5F6EGxkjTiKyYbKpih53vlhQq27
vXhz9KqvRjxkdg3gZ65Os6NJWCUEbV44UHbCyYec0ZJ9JRumyQl23iLj6IN71XWfABEq00fysUar
T7lNChGv9RGV2ebsAjFb97eMuDaLftGGOkpFyZWtfql9oUH3CGqMR0AAU0lgzG/pwn/POh35ISkw
0wP2BilKfijxiRDxArb26BkqY9+lpAyZvdPWxNojPD/sP6qddkOaZvDwmAEr5pPnBscjajDUjPVY
RJrRdUmifmrpURDBZh2NQNm9fVEH33mwv2jgIRLBgCT1Qi0b7qXUpEgtxCsFh+fQ+OBSrWgtP150
M5uTY2csCnPI7vFdqNczNNJrhPlgdOcE7Mvuu1UHQPdJ9MBihh6eKLCz1Tm15dGOYABijl22dQhL
uJKtq6tbVYKqCJ6zdnv1MF5FYgLM4x1Z3h3PCkKsJ63Y/xEXt8jKNXSHpvyqHnQAgO0KOy9goo/E
0JZXhbFlYYcwO8K0WihJpbw3VUZd+DAH4bBekC+bw5IwSZ88Y60/fOBLWS7XzIW1C9sA3kYm42ho
uYtsiZ8HaDyoWnvbLq06zLZ3sQnc2Q49EVnqleqH5RIctWi7GV5WSTOyeh1CmvS23nux6Rg30jmi
mGjl81toMkt333uVU3spPjTYnun8JNXQygdNDrnxyxiqRsKsuV/RkoGUuJuyE8qJAwi6XByAUu21
Xsm6pG4zViaI2z/AhUtLPgYd3dAliyAOTsqVJA/bbQheiU0A6muSb5ciuEZmwsR/G6O4c1nKI4QX
I+DUNE7rt1KBzb1HHzjBzKmnt2ER9gqwz5L8QjaQ7OE18gP3ld/VItL3U69Yt8Vm80DRJoNSPGBE
1wlFE4IzVa7nWF5oDa0+9APFsAtOmDLFS35PAFCjmt40V3Uq8wUWTyriioRaAJ8t5YjSaD8UFpUm
Kd0SoAePvjd7LpYstcZvP8CVaUjOpYInQhNFVcNFz/jF5EY7F5wfvqtUvvJcd0CwN7qLrnA+vzjM
LuM1GdmsrEpj0qHv+94kW9c+C/tB/RxQ/XFx5gu4Urypp6O2zxWBIYq/9BKiLjABu+8/meDzNNFM
RfDerY3QV5a+a3kuPT+bdIsbAxooGzjd8yjz0TzRgWdvxivFGFrLFPVdOgwN/IC7mkWnC/krmXP6
6XQko8vbgdhhpypyac3VLfILaJi9FCtK/uowGSyoBaSKJ/S5eFVTuuVQS8QLdU2FUQ19plkGY4DE
LN4HUlbkEFBwLngTUS6Md3odjv0NTZy+1EClCWjK4P5pYW3qUpxUCIQ0O9ISEsdI/rXhNvMVkMC2
+AlndRhF0qjlNN3j6FAy+AciUXGrZR9s6+T4VhxyAQFuOQ0HQQYWWCy6vEpUfaSsvzEAWJei9hEV
qt2Qp0qtCn75C4aJHk+Jfrbc83Tmd1uZrmOskwiynJBJs4xBI/ZgwKuGlswhf57L+uiCSNKphxAe
/T1S3P8ffvKc417toRreUkmFuuTc919iSj7xd6eKg3f3LeeZ/WhHdFKtNuHzp3QU7Ugt+P9Yei46
NS568/Ie0Tl2vTZca258IKLZwmJfpOS42uY7SWjRzilv6Y24NUSLprVVW2SS6P4vXPAjLUf7ZREV
Fm5vDjr7fM6CUgjghphFvlR4TEHkDnbKH2b5q0cCvUTVU0aA2Kta30k7hg8MwRMuplVbn2eHJQ8g
179a7+E5wb7we3pK7AcHy0tX2wf4eWKJcRpk0gCQtTG5SdlyoivKHtDQS6VeeSsapyJalxkJSUvT
iLTm+NmwlsCbglX4jfMITPI4uOagFhmHwAL3nzcI0bziPakPScOvjw+Tgo4psIA54Smcvj5UcL9N
nrjZrqzAT396OSELSz++g69xjrGdrignhGstqRWzowag3Bizsj7HNpg0F7LNxSHSyekdF80XJ9Sc
9atk7vNaQNCx4QFhLl9ZCiAl1uGxTOl6GJVkz19UGiZRIdZnG0zZvK8WFYHdw9QPMLkx9Xlo+5Lf
GaG+G244eEJ3xi2EJ9mop5ZXb+ZjOIfdKWDBsVFLt6/kCerpL+lRh/zGP5F99rkk8g4lO9Q2ZXQJ
uSlb7axvWUkxh1jFTLACUf8J3x1geYDqdIMMj1Y0zKRxhNLvuf6PkSQ5areQToPwzqLUvD5yZqYh
jt98Vq6jd6HMNF1ZbZ7dNayQoC3p5BR0ZJJTvk1iufhgKuOiO2wFZKUcVovsOYo1WGNJFYwdz8w3
86/St0MHoqc/JCFwx+4MPtWqMrxYZIBZS3XjRCVEcqgGwkq36onR9J8shJx2Caqk2o0Tdh19ntMh
mR6XvsmvItp4OkQMyLc8CaHeqKe3k45yx0F652gk1sSVHGanX7QVsbkip44HkpcfewUXt0u2wup5
mEKVu9GGnY1WzuX7KOU5wCwiWRdPUCuvIuCZom+kLdpEsgt+k/q8EaTocGxc0IgheuQ9z3LGc/oV
hzdWHgYXd1DlDWoPsSz/Hm4q7/GTo2MxnebY5wQyM7uZXw7AeZI8iEBYHUT+fCsBZP6eZJ4scUdl
MOno1vBs6lB+kT95N8ihftPcrpJGaDu9cNBahqiwgIGR0pZ56CSAKm31/njuO862QaLgTb84xcI/
zXWsvvXfryq1cQRMVQeoR/9vS9AZ7Ppf9tNmT38Wqv8TlqqsMpNep4v+h6jwaXuLi6qH966x2UUk
BKIFySp/3p0Kz7eoPjw1XIga+CjA9/tIij+NgacVfpNZlagaij5wzKch5r/OWA7guMkOTBtPgV5h
4zSwDdpJzZq92ZutgpgdiMJhWA14gpV13ynBwcjG68zfOMhyNTMONU8bI852MFVKgU9Pso1Y9wcl
YfXAdl04C52zaE0yd1s5DAFexAdZVeZma/ShrqObTCf7zIyhWTM2PYy0Wv8p2gFgEsvrWK9wYrqI
JbGtpMHv805sWlWlOIrmMZPTlOD7Ik8JoL+luqK1UWl2lgzKXlrApi+PoIMGga+J3kv/ATFhVNrb
HsCzNiwWq4V70d/x+8FUOKUNHAioFthkNEaTNTcnndpkVB1ovctvSJtBCS7HOPx+TgDLpdkaGofu
XpBJlTW03voK3lXwmHCAMPhvVLVSwQNAeNHPincdTMkb2BVcnhJy9/R+xbCEkImIyjUhnhgVxJpV
h3b8CbzJe2BkoilDgvdb5w1oFQjEa8yOlJIa73UYXcejamShYihdBsIRJOjwikWBgYbj67LhvmCl
lXja7QE38dSAN+Prx5qDy54m825jrbEJ9ZQTYykTLukX4oltS1j2ChV2EsVrpXDbdYOWOMzpZwvV
68F7/ZLqO5zFSwZE5wZ/eGqiBdG0djzpNh3z7dOPm0l4UEEGrg7+q95Yt/NpkfzWhuHLl1gTw4uH
JFZrw+DbZ7X9htyjLGVYNFZZxY/l3ZD4bC0E21jSO12M6VqETZMSKHP700Jxc3HRzgQONrc07Emj
aiFgZ9vNCBGREkN3RJ5o6LJBI5SEzSoUQoiEmEVwvUPjXt1WHyDxyylsM/GXkTfeEv5OhXdEiV4/
gWBcu/nYgmGQf+BiEI9k0VOW5zQtMB6SY4hEE7ikZ/Vz6H/C/Nx5IgvkRFiRcHXEuYKayN+2L01Y
21/Jaxx8l4C6Jg+FJ7PjqM4oXqP+1NWYbVWJUdFKRMLVfJ/E4E6sIucfj/SdxiREssR1HRoRnShh
YI6Q1pJQ9/mDzwuOWJg/yOVs8qAHfzVB46zAMECv++yyj/rt6azCVqj5E8WJF8BMMQBC6Q4y5qFa
9lDKx5nEoSu8QjEsOHjLG895l8GPFpwKZYSblvCzFC0i8R05rCKbSHa3NU017vYaXvOSXPXq6iku
v8GlM9GedxA+6jAVHd9oo+ut8RlTiBMmR6C6tzXOVHKU1oFggvK3tIoR3GsDVHzoU/+FS4ABT+Df
GB2K3mJUN9RI6CeACxF2mW8PCa7cfPjQP4j+JptMKtPkJcViekAhqyuzDAXxo41TbvIYslTZU7UJ
ig8VmINn7u1ueM9Ke8zvM4UdIqCRgYT0XbHEI8c3f2FOBgIknCrpjlBk08slsFbUmOji0n5ZnAUP
CqSuQSGicLJDdTCsy8excat3M7oosPysX2qriaLQSoMxyhQJOFsKUBKxiKC204H9f16z1cwQ+tdV
coEf6YGkm7Wfeplxjc18jD+I4tYxTdLGSzVXT9teG0apUseJSWB4FUAvfIX0+JqlQY8H+QOxQKMm
KEEaghROM1w5mwNvB0ii8OaseaOynC7CxTwq42sifSkHOsrWiyqOcoGPvm+rwAs6NfCFlxdULBl6
NywkrxW/DrXfXPaR4SndtXMiVWVcVQwMNMgU3LPLKLGlL5gb12K9NMrMLfZrZ3xX/SUY2lse582j
41CnDZWa2mPaGMIHBa4ZzELpRRAamlZDGdTBDilgJ904TXDpaDfEayoSgHeJawNF+oCPBH0hPOw+
rfMniT4EAs9tR10w0Km9mIzpOfC6gGM4xnZKvsio18GC7TQYmbbQmGX1e5H8eVYjh9aFhhjgI5mX
3qNT+soihdcu1kMN80irT5cMV+pcBxmHUIQFmiTp68iTyuGdBEgvk4u70D19PCA00fKLCDORkGIU
6ZIY15OEIKkQcqM+zzea4pKO4IsAwKPC11o1oHqWoNDredv3UGIHdWFzM46GVosFJXoV7s40txWO
eYYSP+5B31Idy5lVnCppwASz6faq8vL/X1dwmI+2J4N0G706nfzFlRofhBKMliAKWeT3uAfUJnJu
dotYxptl3rc9r8QACAIoXvtvgwAp8SbwKKOh0g4UTWtpE0olL5WKNQ6p/sX6HqgjzaMpfC25iL8P
aXpVXm8x8F/kB0unR4zqDFnXKgP1gIfzZzgRaD5j4eTxqpm8zV8C66fyexLWm76YKFqsFcT31vCk
chCnO1Ci6thklE8YGXC6b/y7UmszIvQAmft2vC+hK7ScJgO68u0ePVMzph5SL7CGBrwF6gyFG5Rh
OA3sVGUUore73QgSsHu+gUKnkPYa5J/owXDbwJpO0sr1NutCcOSM2CmPPqkqGUAUnIOOYu9huzi9
GWDNPiWeH2J1IoegtHDx7VblPcRE9MVFQPqFpqKoX6AhVRfS72UQJX1/54zL4pulU/2QenVPZueM
Vw2cqkk84zk+x2gBcYA136WJgEgdpmvewX/1AnglyGg6Y4X7CEbV9h9gEAM8e4L82/LC6MTeL+Sm
KxMVMa2HD5kfgyJj3uvZtD3Qo1/2fwtzyQ+gS8DloUh2w/PkzCby/jOkwGUx05CzvrcK/BilG+6M
ApO9ub3Q9WEQae+/1eTJUUjG0xru3s4mVKkGtFiWHzIy9zfASBkUzMI2MtRiVWglYrXwF8vbRatA
C9R91brX8NaqwLZXNj7ClztzA3wFKDH0vyQdVNFHcvp9q5G7eLMw8ab0SbWfkqqeyWnk/7AZ73I9
YzTPc5uj4z4+YWNQE2vkmzYrTrajDqqmrsSYvF6FoFoseGV94elXK9hRVR1VTkB03VdjLk9/BLFy
fcgBrI1SFgzNOeNjxKcHggH2UQ0kvWU2L0pvVwY4IoaRvahzxcMmh64bOV6tnZuI28jFN6UYPspp
WDGjUbg+D4QXCNT1g0A/TnmlojTlhY70pZnGlxoR6Njs/V6l/tWp0aAzTH8pd79xHHScBbpiWaZ4
w6gWMns57dKpH02ejervwAb/i4b08yOSnTkOK+W71ji3MTgZRo9PPbWRMZx6X3rshy24HCSFMTJv
/7+ercR8MUh6ltpSt81/c0H0zV4SY+NWD8gfg9a4hAedju2DCuIPv+W4CTssux6ygPucV+oW4AkW
CzEMEHwj/pyhVzUr87sN7swrlcnTmCKJ2Z1iWo2Ilpjxv5kw3Pw/v25/sskTP576CNThfsB8lZal
obyKatxYAaDoPo7lMgpaffBp+w7mqo7U7E/C1EzB8yjhgWOexASPR+lkVl6ppF4oejz7NBJ7bb02
uExBu8cVOo6cP/jVFSfD7I+qMsLK1IxO/M/YCQnkTwSiL9xz4DszTh41SxvdwOZyv/KLkemNubCk
BkY6SALRNLDKdjAk/4+Kw0RJg67owgcR5AvmVd84wkG3ymHbn92fgLJCysCCIyhAK0WRVeFCxQj4
M60wEBtyNyYO+HcXelymDckxqsYiwUBV2hVkBN8cLQDS2oUdlS7tZm2vRlvXeDJ1Cy8lDQR4kVHY
aXeoU8zuUVisQQ8chdEBVSMuDOV43wn4BI2u/YVbw6CfNMHRjBhN+bSXOnsZ2c/oV+cNKqCFHpwq
/mdElaIoXsOQfD/bwPNq/CfSuORAjVXjke+aG+RbekmrlW6v4ZaZosTNN63dLO6guPHIbkMwx8VM
iBfrrOkCSTDT8y5zY7vjwheHkv6bp+Z/mcKJrrv0iL4Colqqr13n0rPYxXV0D4Vuct2qfAqpxfER
uDXoK7seVsCBh6rAczPtHSNOTwc7R9WgehcI5Ot0iQ9j1vjy6L3cP0bSxYGwuDN4Vkq1tKlODgmj
WC4EsLVNTXBAzksA1MkvKq7ZosIG5m0fUWcaq5x2GR3JGQ6eYM5e/RWpTJiPRkXhmVS+pPPiHsKq
M+d8nuPioclLARubBteaJB1VbkjqfcgsiKgoH8hMThOMuSwxx2w2bp+4r0swrW6ORzq0rLN1/nSA
Lcn6c7hZF5ffGCTh5UxVU6K0kRbXXd6uKxFoZHGk5iLlKhu3tdcU/6iP6z5pP5fRsfRWmPw51smI
n7pnPVVCZtlt230DkCJs5edhGCOsBxRXJpBJSgl49V6vX5KWbYMu1nsoB8j71HvcNFZ9xluTVOyF
hYMfhkC/qdgmHdpw+DH6Uy7ZBLLwsk4d6OFkN7We5yQZMAKNfksLrvR+ftl7YcgiwULs1tsISi71
tw2byKtlQnb7WR1YdqvynTINJKwnsDYX6Hqug5sFdcGekyq/fd0+1oyt1VuOpUmIJQHeO2gWdVZU
Gzb+bb8mDkxRcLjtoECAKcpHZz7fjNEYab2vz/sTBIzYXPDxmjSJJRqaDyyKEFhnd70baFz7EUCH
u8TiptdG3FZfC+Kxw9tJWYpHunl72hIS97VRHYYcbVUUGLAnB2/9EsYKDy+uYBnMr+BKBBN51ij0
sQPzGkEWJt/ChDQy637u8Tc84F1upS92/UhKmtzmgADOgOEp3hMCXtPnDzs9ElAGluG58VzcQeOb
1vo0WAJn9cjrA5G6C+xDkhrhjBR4XuZhFmOuLmFm9Hpfdtw9txcJSNOlHzIoVFje2rS3D8Kgz2ny
tSa6FJE/+SYNM8/3FB54qJ4IS4MxzJscE3f5iuIqZ1GDF22nx1wpAjmg/oAghQZgKG8DXoMNZM25
WfcdRK9ZgQUpvzfj8AXUzRqzqbovHCCAsejTtEm/XPeyk6fdBpUfoJPuxA7WeSEQ1UHNxdm9p/qX
uon7xUNUXGw0CUFNJ2Cpgzl27omKsTA2IwMzSq69OxA5ynXwTYH7obyTsTgeub5dFRs0KaC4gnRw
xbMwVndM3qiHZL2jb+JopctClEl47W2JrAp9J9AjBtdO/4QNyGlQNHAYBInKlvQ1Cnwjm1YTk0om
bZivAIV5hiwgNAOpxcoSznF5BWVlimFeuf1iudzpZDGekcU8fy92PqEw5VxuamKcqmtHdLytRuf7
JKliajXBDRhF7oq4U1Zbn+Y4Vd73qe+vAG8DlruK18HoE8upZp43f3WzzXnth9PHonS/CwngoKc8
tXD1i7DWb7gHWXwepbHrY7G33fp0uHuchesEyN8f6jRZ2rh7omFYaVfEeY5QpSTBqzDsdDiquOKE
7xWHqatswAkmhXMclq1cmPd8si6X4szgH/ThF3VxEDKa0OJLAtGI7rnTJXJBDe1pkxwvXzOCLk4Y
LOlXnisQBEHbwxYsYPIXD2VXpLMhcajGbjG998+/qqXIx7V95pt95eiatl0X0OZ6ta2NJURL70dt
iQdxaOtRDChL3c4iceBumtd9TvMOzwy5WEhK4a8tui2v7KJ/zT1Yc8ioPROshzNZdzI8EzQXLqJ9
sU/v79f5bE423hrWrnH5c7qaFjhMvgsb4UC9fiY7DTksC4wFuUoHgXw9f03Hg+k8ug92VZTqaO0r
9GCQjwwyegaVNaeP3smuSVNnorG34YyXoiPBYa6/dI3s9MpPpu+B8F2jhyr+HSQrQF9NPUUzyBNT
i3eHij2O3WZxkLkt4mE2Ns4cs+fN2sT24s2EIlkW9Dk+umDPPOlHyHkiTRaEBDsKtKwmufhzXsTO
z1MTLSBIQgsjKZVEwsl7amQ20TZjQPokvexslgJBS0kqxbjdNUq0e76/y2q/2jvH+XfqQVyVqv7d
4EM+/iMHPHuEBpA8U/qQwIVdXWQW7pPeNa+jTyXMSJCPUzb57GONnBjYNdcqh1tK7+6xaoMLGYZx
zALc6EV4h9oFa8b0Vb0NVUhsP1JfgBPXWszq21n/GSW7UtLyXQHocKQrFEx2iIRRHbYBYx8MXgIb
tztx92zFv4kWos5aAbysHhl/Xok7pcwBVpQ8GAubHr+fTxve+5E0vkI++4ag0AVWceZghlByPt03
d2uPxnk/CRpEBLFj4nWooNqvEgLTGOtyF7LpRMgYrtP/X5nN4jT8RXOZoyAeLCs9B3ejVllWvSL9
mgMpiKyBh3BAHVOyNlTY6wKOrE+xC30S71lL9/LVjp4JYSYikus3UETvJK8lFzoUdF7mRbZF7bAU
E1W5X7kgphKjWgf16LtJUU7kPdeiqnZaHULKfYDtQoOa3dgYGtP5rq9tMpNs5vLhZVZkNW33JbFk
rYdH86dMc+xfz8x38XLjdawq27rDhGXheGHMriM6d1FXZS8fNUyNI0jwKBmJDL5ytJX3hFk6beXW
S6LwVJdaNsSdX8TCpDZAJR1iRvTVtCC/Fgyd5xqEsea4ghzjjWILK4jobXKdMId70gt2GHho90Q5
nv80DMsV7x2MGBZkrRSiJO04VP0t9DZYBZklgxGeB4EWFP2R5M2mbVmu5e/NDUBiQLCKktSf4slu
DbrOWqYsuTsNfQQJOhMIcQai7U1c6sakLR9YfgQcVRq6Xvfy83Prwe3+ms54NHICGjC7kEhJsgBX
60FcH9PfnTUu56yjjhqhjgzimjyi8w==
`pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
bcQ18muyOi1YdHX9kR4fi4Y9hpbeNnJj9Dk1vn8ggb1g5py7HXgMECR2vUHzPeJT
I2BaCXKIZVnbn6bWseOyvyaRdi92qacqmhGt9YhtfEe5V9XqGKCZ9g/NS/A272Qj
lc0Nxu3eSbL084Sxba7hUHJ8zlR6ogkMWNPEM7032pk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 9296)
DzcBijOpRYdztaczVXhoxAXOa4LW8kc/9VfSpUPCs+aye0DHq6Bq1RieCBXvznu0
wiNrKNx0j4Y8fX2MVf8sUx5Vv4tJc1Ah3H1ZMSiZmpdOVFl3IjAsOys4UzgpR2D/
NI+yPqiO+4QZywwlAiDOHjMsib0xWzzo6PBx2KWwbyzZi1R3Hj/4hAoDWWk+DnL6
AOHnTj6QO/UC8XQqBc0q5PhocMSHJ6tbFOx1OowxuypMyCezulQJOZIhzXYBBYAt
CBB4+Db0JGo1wGxrADEwUutF8VRzkH83Hw5TbeaVb7Hk3wfgOd2ZgfTo4E1BSuze
Sszu8Iv8dS/mMZcKHNrpa8dYC7swttMruHdqoAYARruroL/8t0hhBfTIyIm/4Jhj
yEdAk+1KRyYWN75gsWjo6ohuiiDwqA0v4g0lvTiTh01Ar1Sg7m5ft0JgfIr4CcZ6
zm5jYEo32JOa+d/+nPDR7ONBo4d9bzoHYTalbGrzYRb016Z95Ozl3/s1T9/L5foW
qmZ4FJKvL3hNtUzWDiQQIZ/7DbZh7T9IrfakvEN9mtx90YR4zEhuKULqNxSssVjk
6hq7yYCsq3FVZbsETnBjhScIZA5o5oVCOYJy3wWt9QIVJ+MFfPV1iXUNcRR3JuTY
6UtbKKhzXbISAhmoV0YQCQeK680FFbGzlNhk4GarcVCrlhhZihXLfz+ExAlMZdnt
Q8nor15OGHSGexWOb7pMc8Ek3bW1z5pW7wFQ98M4VgDSMGjoRHDMc65xuT71vOvp
3zDtdWxqg1s1TIFHPvDfxuo3aJQB78ZwsqYKmmo2R7CPQhgZzG1nHerYTrpPsDnB
SQA16lvAAQgxJAX7aLnkyW7dyErXsimowoF6ofEmnsqRzhYuvMCNSWtm90jo6Zxq
HYn7t8/bcQfjML0Zh/6g9N1AqjLCAA5ixHEq/IMKHnRoY0Px1I1/SwO4QN8Xw8nF
RLfObTeOKPbJRzic7IKFL8Ta1ZNuac7G9OlotgY0t9SB393IXY3+d3tWFvqH1mW/
/WW7tc0Qly90tFGcPlA7kKCdTiQ9Hx0972zW7cCn5UhOtOLEgACXHsAQx6M2bpJI
RCiy0kn58JFUEe5VRLfsHCaUfkVw3ZkjjqtfwZqvtkOl3g7MzKxBTFwkCxbhaIG3
dRYLaHGPPuBeS+tXHWMlA3r2jxjDKj5nw875Z/a/hW8lMUEnHQhYReefo0VUkInT
+ay8mjksA1Chh1LH0wqVHB3nHgyBqwiT1sZ4hIOTVjkGlw21m4aqlifvTvvCNdnD
rDiU5F9tuGSsLoStuiqT1pNon/unBVU1OBzZNix8UEosd21diAJxcDXJE12Qk+tq
QYIpB7LnBa39FM5eeMvhSVsNlr2+I8bn3veLc9Tkw7FiceB/ZqbJTHDR/euHvOfl
1t7B7qno2hH+ouuPOkGv/8Ee3cn62edW0qH+1QBrwuCGjv0tzEaulUqd9gVqfxzk
AZWqccfPfeH+DTbBo3SqqsP1rk0F1j+3au4WIwx5NGg9gWvMYko9FFBsgx7nii4R
4Wb/kZ0t/t77v3YHQWU4Id29PheonlJXcKIQxlpSy13jzDVxpAVfguwLbo0Eh2fC
X6AUqHvnXz3jyFAgBbnq+OlCxzjGPahPNZYSbO8vNBHSUdXL1ApB2Qi1t+pbiXTZ
m9+tdm5qoPqNmZswLCdzIuDjfa3L8Q+c+cBgzNdjAUAAjGC74An/0B9+cZ8QGlAj
oqA1zMt0zFpVJg4HxsiOyByxqEbSYWUDSHmhWY4eIc4/U6AjskF+mqBpDLweqMLz
P55ivis36yC02qK4i1BvaM5aVNouQ1i72+zGleQQrd9+bFCaWkV02JOiuVBR+s0e
AckzzoBjEEg6moRZDWjy01HrQmd071wJUOrzE8T6BCGtRpby8WBKifJtZ8cA39C6
f93PV/BsJJW5Qk4cBojWIkbFrucdVkMZc9RhXfsOtrlQt1jztweckiRzOpF5OSDa
Uduu+i1Ae0ysBmxvyXFfkhbWrgUkqBl1mc4mmjcmuQW4WDtJi1x9k0yqNlUH4H9N
TtJM8MpTE02TZwlDcoK4VovsH8yMl8FmmMjUUSJTV8X2YYdW+Ps9nc0Kr2e1Mlhx
l7s6FzYq5oK8dUQlLVFSYpYR2K7Pzc+qzhWjHUb0vIRMeqgRsnK44VEuVi4Vjs0k
SDHaX95IG3aA8pdVQh47dX26O9wre0JoJnihZkIlktoWQsc1jMxU3j7JuPXKUJ4J
j/keVpGju4EmOvmkK2EfUISDE351TfEKByNZAFedvKHjPtUykVUPqMS+BVxC8ySc
HDajscZ+iO+wl2b/DtmPi1tJf3+cn7cbiFx/BlIa0dpZlMo3s02zqngKo2sfyDkr
Z89pG8Z2ulwV/zmBPyWcT3Z76pCkPq/RhIleV6Lnltdu4GV+N5f8zyjcfbs4KDyi
sx3Y+eRNiTVC4uMyLJHpXVM6Oi1BX1wUPAuW/3nnxXbMFRNIsNAmMZNjtgODD976
MhjkYnus3/MuxJA1CVYDXPjvpNasYCM0DBYZvrtp6lRl6R3DcKYBjn2Y9QuzwgaQ
i6zsOYxLlhL3jnlLLuZEO4O+Zkh0PCLKibXpb9XYD0XyJXOeVW8xwF8T8CCEdzDI
VSAU/ACg5tnZ66fSt9Qu4VjDVRtCck8mNIRgXnyhGWoOqE4Vd5pUSrL5W2gWquw9
1IBe8Tn2zM/4ni2bTW6zTZ+pqdSwZPwyG50ZpF6OMa+kwzLuKXyynoJeq5G2nidt
s85bY3rW4gxjO4EIxsiSY7Rvjsv3Lcjm5BAbvIQJprbp2sqJQkWbRTVoVC0j5WhO
k+3pgEpIzG9FMOb3jyCmkaF8ZLDIHm6EeN2+YxOzlwfh0Y8VCW/HwfEjR6U7l6hy
74XlNS6FE0As+slnx2mataEN6FQSa8YYhuWapBWccmRENe5X0TDJrsJGQ0qzuK0O
ElNYexFoFUUz+2ZTvjggK+PND9GGqsXTJBUYU4gRuDDiea7vsn58Gx9UlkRb3jgX
1vhaJW4XtPaI3NrxPkqmkCQQGmRHNgI18BtP0ZjKdqkdVmGeI2E7frgVykL5Catj
wKc0p4M2PeBB/KeYW/aRvVAcZDFgbUEr2jRggEfjHxuDbLSReHmXuBEsv28GVFpx
9jYutkOz4iJ/lWR3Qu+w8IJWkhYEbJ9W2Ka+nstcmu2kEwrSLXMbIjEgko7Eta9U
NMCQ0sP2X7xd2jxKjmWK2KhUbakOpTFXXZl1/mqv+T9dQGpNVO35snFItmwvvm4T
VcWfRNsGign412qvz5cF6mlzmePvrM3ls3835l86Av116SoFboZ39R7/33BWIvvV
A8+t66rwTUlaaApUAa1lDIcMzqdmDy8DaVRVxSjyAofuQLzp3YyA30CoQCo1PS3L
WPZL80kzGQlPKKKzDG60OYLZcMOCyDoYxY7kEsfnw827Wp7e6MBlo85dX0tDRjDG
8uqVoL4w2tt+HT1bXypvKIKP3DFhKeStWf/G8THOuUoszmDidRAPWJBexPMQGLUC
e3j76r0dJ9AkktoTF9FrdFRDxtrWxgD0VkhaU2TjzNj/y7aBDbodjZXV5wVFF2zl
mth6w0t2FFdy+e3/B1L+aVZQ9UoMhHzjcE4RBIYXBSfrLq8U9hAIl0atRsbMuofC
G+JSmGcATC+9gprkLrJzVrhTWkDYdrT1ydsmQ+9hpMZKhSIPnbNFn/V1TdvVbL23
/x/7uVhA2rxzvVrvv0NxqEg1TrTJGfGC0+vJtyF30+ewp07OzRVLt3UZruyzTxay
VX00qGsi24qn+qnAcf0hIOJZOtl65Up9ZfgIRsHj87PmNeRREslnduHkMBvTUffJ
Jtbapwogz3xSE+3Rof8FPb89tg5Jm3tl581CNY7l2Y2xVh730eOD0aNuLjQ2HYFI
UOjCMTbCs3F6I/EYPx9LinyLwfMRF9UNHm26aU1Tp1QFfjrcqjzinkcbBsyW6A5Y
K0PmGzxJWeOAlkBeGEj6zGVpb89lX6C38gsweu3X2uztzFq6aJf2ag823OTBapkR
PDdD9wDGzrGEQQbogylGf+k2FioFdtPuuofUwaXSvPWSz4qD0xOoByAbC2tkXQJr
s5yiF/F+b1RMorvOL2uNZEN2feaZh3fIg8CWAPA4WkHgUJUDTTlywxC18enBUoyZ
ohMZ81VO9dsb0/FXP2ACSy6sZVccOrqY3jTvokzQ+fWLoCj5voF4FSwyg/3VIptM
f1FZ7YME2SZo3zcdV+78AlawBTuQ/YThoeSw4CJhYNtQpUFGnseipzZNbY+Lx2kR
gDXeywRGBp8/UnReIutcmzpEYb2DlNpSk5wLhYhfpx5TWWoUlvzAHcbyv2Xe2NmA
lVJYtpqZKA8afWUu2Db8tV95rGED/FyW3djuh5Xs2eennGt2Yf1iUaLp02kVLtHv
rgwXoriMT1UB+1v+ujzNuLIE6ThpJ6ZRtofQhXOWmKgTRzzhiHX8dNQk+fKlltJn
3g4obWno/q2NMlUbdCbR7Hu4vSkgdtoVyGje6pHTtxdkABBCpQ/YiPH0RfWXA2La
nzBT2GWpwIHkG5RmmBtp7zxfvvxBe9ptCmUFArD3HoU/mrtsL7K9UTEOIzmnzO2D
1FEc2ZF+XyC3p1/k3t3iJaIdb5Ezq4He3fik9U+NVZchm+HKiqQVMTDeiVYfAvGO
ukiQ6F1D4EAwTeVNW2jx6oEJt3vZSdRWyGQmRhxib4Sc5hSA4F+kzLdsQd1kgM+4
HDX3aexmBageZSy6E1PGLhd4G1kIjtBEt+odeppu610sSKp7XzaiG/6MBjkmTfUK
L/mMNdmjh9rWFGAhhFR8EzPVOxFYcHOhxCzraUPKm5Rfi/X6IAocYetAqcIsianK
sLPpHCcPsmk6uOQtPEZs7ujUnmEeAR1mY09OenUog4XHiD6xauoTi/hd0JlSeHYm
5vIYyvwQZigbfwHU/jUfIJ2jocICt4zlfI/jo5OSscZfpsEefMz2wLvPWPYC4/yF
r64q+C5AYp18SSfJ2Q1mGdzeL4FV6tXWKDRLlsIgWK9n3W0VOHIwMkwGwjBzpZCv
Dr5a9uc7GWqeWSUInM7hvx5o9iHumc6F9VJ//EJghE5X0afbZCqsHlLrwKCbcM0O
Swglb2+jtJwhBhgjLMP0vRppYwBRQrl4FcF7kBvx626CN8vbp6Kb5Y+8bPxAb6bn
wXuYlBXw1l/s7yGn4NS1MH7vognp8Ws8TFdHo74DpV96yO4d1lOMUxUMFd01UrMP
uksNz9fMCZTq5LKl1bx2A1W6uv1aVc0DRhr2YzyBggyIBqeOK/YZIxtAzMYn3iPU
JH2t+/Y1oA+9nU7Zc376s1qvx7yNJWl1prbXfzjEcmbiA9LNMOiRfoaUBeR5fwDo
5GaVPbu8oGQ7i43j5eQJCsYE8vRQT9AKsL7IzNKsmJqSfOatdRn94PLdkG11N0P2
AF1UNIJdFndHa50ZFiI3QwVJk1ywwwJeRBZEUbTzTCH15W2pxm39BUcB5deVKvx2
pT0tFBcd17Bjrjc6H5Ac5MZFxC+Fy+1c/R9eG9GyQlAz3ucUj7/P93E3DSth1Yii
Xdl1rfNVUZc5wKxHyNGWx5oPGthoeloJWgrYEv9yE9XwHknmw3iEZPZcOAE1yX6n
7SgLKNWy2j+a6fO27K7RV+O74SDdNZAAJjHqzpiiEgV8UoMXDeM+j/cfu8Z4Q/LB
iddRW+hMKVcdLr+/dCz/Qn3oacAyQ90A3sNs8DfGXXwecN2XuvaCRQgVIWiKwumD
q2HdXMErNgVwlxE+7YK+BbYDsCPgHOh8dHEzn6Ij1Gl5X5+oMCLjgoWAQhPOhOKz
71mTS2LNcPfPmORgbsestXewCFZ4yWGgRTcgB/q+AxWLjulNohls28wV2GJnHyTq
6k2N+/h2cf+eoXn2LmdHzzy9yBBel4xgS2qPa6xCZu6vMEgb3qgxu5ed9GFNTTnU
P7DUWlY91d6fnzwsRtzTInX1vIsJ9HL8CZG833SjpdiCpN6bApMt0g0v33kS2Z9x
CO5RVHX09QB0Anh14YD6bhSOftH0kPJHye7/yBEe3hetYNruuz4JOiXJHIGKR0OX
nftfz4xLBkALQPrHJKrXb0X8wk4NHJxGDwfe8b2s3uZoCEIvL+9ADhSt//Wwxs4H
wA+art11P3EJlCvEixTrdOFvgo3jpNINGofXcmbkkSGfttPJp7YMXzH5nG6Ljdjp
LpEM1HH41853FHfMcUPOM/G29hBshLVIkXX2Id1NTepdZXMxpfrALwcrUP+s3fQL
5jP4f3mbMhdVLuNLbKOm/Jy4AmNS1R8P5pxYDisz8WIHymaRlJ21Tv5P1grXNAVi
SRyhnTOC61QSGsvQxF6ls2S/UmoDic9FCitYFHOvlSxGb1tg35RlzzyVsW7cMd5m
nhilBaS3kPxiDlq6BJwocY78roHlzTHQN0PNqNQM/knxXC1iMc73hYVe2h5lsRZx
TEkZDoVyMFsTtGZBWmNp9otV5jGYzCMFDQiDQAc1/+N2AkiPJiGw8mJnLYfcefnD
Ii01J8SujfbxU0nXPuN+aoeQt2xKhRPX4w6OvP76vuyzKsnLrGDujL8hDtCmLis8
bpEgBYwE/Pe5xNAfgmvQGdqcZaxZ+s1U4DLegc4JrwH0SsaoRRc0sHadRn25WmYr
KGVhO0mfQLzfFVu5WO72V4qIAVzb+XUTemrDdi/9D9/mUdCZ4T7zYdRD1pNyyznw
eOEgdBo44JyPNAN9Ilf09bztrkplbqrmMs7UtoDCOYt3enKu9FpGJkT2ZLJU1WBT
/ebWmNjCl9PxyOweq/LeT7ISGo7ciq+rfymPe0cEOIhASMyMN32hSp0ceDpysbv/
bkED8Ag4wPDAmUPvnHDbwLAsWmFZTVmWm68o0K2s4QuihHCK7/YNqiX/QgQL5L/h
iPCQimR2JgwungrIfCbYdGPbkKV2gR6h2pQp8Hd/qTVlAu+uPDCtIqCqMbs9hF8H
V2I5bfokWieS8f3aAD/JyQIGHZsOdrNb3sMRrp6UM32N/rg+orCC0QIDwzWE1I8B
CMSxbAk9k66AMuooifkf7QaALia+KuZlPoIG8LD/xxGcAGUVNxj88VOEFZ27UcX+
c6kTOtWfKZncIKJv+a4r57a6B2SxaWE3EanXJrXbuv2yTKIBu1W9hvm6opDGW2YD
0UJD8WEpz9D3qfDd8rWm4tqZoe9S6rPs6QA3tMkpSF8smOMg2HOw8Mu3IcrGo+T+
Ai+T4JLCN3qg1LBzI7SKd3iZkg8mvp7GV6XfaSIyGOs6d0+7XLnec2kAZmoxKU0E
SnoetEnDQC49+pePvYgl0J/R3CYcQ97h0f/9okDYjqfsv2e2SqZv3CvvXhZzuSrW
kxUBlMfe9+qQ0x4zYsnUxKvF5xvAwYUg2DUHGtVuLs7mHRiyMk3dgDBe4zwtzuBk
iXaG7y4yhnULig2q/QEqb3OJmmVqGmbn3hIRr9MK4KXvs1Z+n5eTFXYQjTvB+Y53
tMjBNZzXWNyiCfHE2CLHRsjDlLoVyroECguW7i/EfhsloHNQThnaviW7MiofDaRr
WWNtGv9pezxeMH9FSBHqMZ9aCEi2EYNE0p5WkVQWk5NFNqmkmry5JGaszzHJysOe
qw3Qu3FXglgkVU1zWCfyfwjlA73V0fPPOaArGNfOJd2GkTxV+3PsT0tWLOzDm6LX
5OSYFsrr/uNKAqRRV8w2E5OlmeUtUKRinb7kZ1dfiAw8lrZe7gJI7wmwdCa6GuTU
PXOePJ4w8mlbj7Voer/FfrtBfvXAzgb4tEhuMNe7qqmm9e5DrIuxiNoJbWa5gFk2
TY8Vke22QeScRQT5EMWR4ee8+39/3fgG81ainPp43TAtiouG3i5dQYv4ERYIYDq2
Zwz0+M3C06+Xxvtlc2Kgdvue1RkE2eE2ccjzwN+8tZ53nIRfG3L6qkzQsqEhqwBO
AnOfGWgL1E+a05vK3YjErPsGh0NVvliWPM0SEkQCvqSanoXwAgZfDXPweS9rGJxi
2/UX9ITyi8WgaygU558EPqLmtu+RTccqzajjuNE3eRpm3A53I2rTsGVlLJ8LO0vx
xCpfaPNkYBRKz4CDCOSeWOBkvlIRXVTYf3N4BvfjmLQ+PD8yVZQ7orDMAROPJ9na
GdWTnwoamquMNlMLC8bh2BWm96v8diW9mtCXYDmyYbmHKW++RHY8OhYeYZA5Smdb
08SV3bbr+54uvSEdmfWvmS43nRrEHqEx6GWiV7MyjOcVuzvfj++iU+4GyV6uDBYg
UHZef3IkdwhNmcaepaIcATk2x5MowKbc+exm4lDwawq/trsQN0Gq7vjRvDCiJ2ha
AYgARWInOMSwIBStVqgx7cvYIc/oK4zKO+10X/GKNAkQ6FSDsaSHubs6pM9cwHRj
K2KHDeBkjyC+HvrTtNrD0tEXx5LjK83axaosVMqAUX+n687Sd8DPmVFLKuzjgkQG
quv+ecTXUPm+J4l6AY7o49fI3D18aUnc1oesb7HJCV4NaobmA4BxLX74jcvDOxpl
fAFKWV2vfjunnk/q9HVvZ2ckeE7G0VOJpgloox1RPPcb79zwPw7ZEsbW7V1svQaW
xYtWQmNYggJqEOkV4f7ivIMN/D8nqJ/xFuHe+8VzQSurQEAzwadtjY27U+P41Q9+
9JQOu6gbhoVeWxlpeIEUo1aN8DY4fpZvaq2tmNvqeSmuU236JHgAzt5mcs4qzWUD
WhAtkH2OPclwVt0+GwX832VTCEljk3IsoVKLGKHl/x6ufqvner4DATHUF9Gc+iVK
X7yNW8a/i4RvgLYPnI3nloO1xTolp5aaCk2LMTSaAaeEF0vKaEbOoJuxNqkdtbZG
8IRqeXklfd/8Tb8KBjG0wSqC/NGZZi9by16D86JmVg9lJ/1W3cWExIdioHGFiy3u
BH8sQiz0+G6NAyPR+TXCrwEg0AtvTYVf2cCDTT36dkJUXFYwcWXLqpSvkH5lt71z
aVWdXSfhpnNuqVKVfa1GLArA2tufqK0a89LiKWNupDP5I0xTYi7of7Y3pljJPECH
uwtMgZeWrXXAm22vTUnX8ulinBOlGtWwmcvSFkUksvqrog5U31JFNlqh00ppYGYm
14JDectJl5/AFH9KSG50eRlxguWxNqva6ynLjxJ7nj6Ry9aEDp8hvhnaHf1ylfKS
mLMU/Q3Cw0vwn1PBclsdKRk6ffy4faT80GpFlmx72p6cnOOgUr818gKpNB8C5xkF
TF1xXV2IFFoPSA6qBMJIm7ADwgz+KK8u7Hsr06M95FRq4kWs/ea+Kvqky+Wx/CTn
pCkmZ2K62iBXaswkDseNEAL+ANBvPDjWCmReMqtRROSfNI1BmRh/KGGB4DI6aCiT
yRDGp4uJdFGu/vUeGAEIhccLMGfRg9g5Qr7l/Gf8Slb1gPKbq81Wx83vkBQKvnzB
AQ5xDJP9qS6AqSDsQPzVf84xiccS7Kp2IMxKSncaSFpt/4LWBU8ONXlcIYzhRl3h
kQqhZKdj/OSrEsPSyz2ucMFKfJon5s31PGlmj/5gzFVWAJe6YmZO1cXWs6L+hW+4
tioEGNrlw7JykN/QB0Ow7ZrlF/+J48DTEY7yoTTrCEomk2lX7vCj3FGdnvRh1wnZ
Fni0V/TbPFz5doU8X1FBD56H2JfZRtuEeKHek0ZaOU8ItE4T4b2dA5TlZ5CJPgDQ
obl3L0bPaZzbd3lRFbOTk5yuElUaiSIt2hQBRse3Hc4tAUNaw6oE6WMgvt48cotA
0Cwl6WerIC5OY2C+Qyzuk7IpYwA7KuoqHjRlBnl1DSD1LaV0VPNpPwjqjvcf3Bg3
dX4SJdzhg0hF2j3Afr9u4bZ+SLatHF+iEpg5QnJde6QEruIC5iYBIwYASBlIZdRd
3M8LiF7LQba53YHdsKoXKUMZHgEAIw4/E+n6ItUZhaWiieGr/6BS4LUCS34qtPVn
+0/n3oVNhfA4gydGFSA050/5kTVnFtQC2kNSnvo4vMbD0gUQi/TPBDhPmIhw0Tvo
k0f6wgt2J09ghd+vg3Z+zCtzTvVdVhnas0s2/FMt0cFsFz2iE1FZJQ54mNq6t+fT
MxP+uPrStU/aUPUJj+ugCt3DrPNq4if/C62hvR/kOzBhuwH2d0rn2zzxbe7CYUU6
lVZTMjckd62sqceABdLvh44Jz3SF0Nq/DJRE4vOgAAqw2qm3kVohOOj/TVLJaOPL
kYsA2SOY/EEkAgoTY9eVFYWuSafyA6Q9GnmZ1fnjJo8VhK0Erx12CSw+Fb6/J2H0
9960JUTsZ/Ko5wAH4bV8phuBrco7atoU7wGhzu9a2B4P9KZ0VQJZmoMpvUesUi36
UVzx5anNYhAqkCpw5SZkjP6/NiSwnTahbLW5ZliyoYiM56lcL6gd3yG3zGoNtwmp
BZBn99Cz+YhP5cIbvbjtRu3VAr+2inw5G5UtzNwHq7d42V1jmiuYehaSkpDcRQg3
KmANGM+rSviHR9PHxYP0ChlRDiaSFZUH0fRkg0ey3njbsVeC5yXLaXR+SPgcxpmx
YuzwQjt4YMdS9dZKE7YtLnUC6qoNDJd6MexqjwTAdHzvHU94aK92jKcyGlGPu+KM
y8W4eINWmW9Kw9K64RrdjlVXCfwgq0vju9mvjwozqvIT1dHfuZLb5L7cAKeHDDQX
xc9W2mYDrvWam+kXVVRi4ioJ+VQ7Kcr41NoItvSw9SKDzKyvHZ8QRL1iRbXNh702
8n7okKUeuaeBzKMrWze+PM/D/8nS7dnnO3MkOkIi+AjQvPFaDvpuZPVppCB1HnTO
Nz1tl/iBA3OApfloHz/w9yiCaQxOi/R1DAja5TNqIpzLFjMTzUzqjBz249KmPmOO
vAGibtS2gWNPDOQGV/of3X4MuEm+6JnebLxcDVpBlS78VfIzfJrHorHDpef1G7BX
aNmo9hV3Bk+377xTbINEAP21QF6Ddsi1k147EdUGtfw1pY17UobKIVy7Clax0+Ct
6QzctwXQ9lKLtJPWnHM6vW3I+LwDX3lOI7j3TO4uibpR/qC8Xh149aUL/hz97dMD
qM4C1lCfa32hGXDJyn9SH6rr2wXMVvCX+RwXXJciGrU3KpaZrHR9Cy/p+KKW3F2L
D4evVioMxO/NTBXVMQ1/LSpvbon/38Y899Fq4k9b0OKp5E5LdPLJLDZZXd/HlzmD
wfCFJA1Gyuu9gUApwNo2pdwojmeXrLWrRKSMAZYL/xqKy4UXFuNeY/iiUHPHUvdh
Bs6n94q/vYhOJcmEbIKILm2DY+ySBBNNtsZzbQ+msqu9ehN9YtRXQDQjbI9PYKLK
VgBWzJ8X+XnRb/YhaDPUN5O4u2v7tD2ZavMao7/1AUHpZZm79cF8mIRoFAMODaI3
i4TGTLe0EBjLexeb7g3cM+7XiiX9hEQ01mr37Z3xdTOJY2uasRgtDgfSW3BovskF
KaaQnTNNGcexxIuOPYTQXDCF9+HeRvI5/RIPLR5WXkOthJMZBqfp8NdS4fVW1J71
9ymFotzCD1ouOfxZVG8P4MTo9KtgoJ9g2pGuwgGVjQ0XARQdAExYb05lh7CxAWvC
uLWicjWcup2cTJ334+25UhYYTXBAv17KwCY3ZC8RVnMXazjLAVIF195Sb5jFi0Hg
u0P8t+KTp4WXgH7eO0vD/VtTK8/W7hwSKl7tQMEx+FiSNOavyqSjqrD1raynsF7G
OC1NnQ2MeFZASlPqjFVTzTiM8QNjTuVlTQk+AUrcrtQj1oMEccw20kQ/s7k1oQRN
Tgn1DpmIsQ9olaikubSk1ZQ53mFG0bBahxeahxGk7+P13VBYxNWukOoCo1eYkH4g
DbIc9dQQ8UfhaYkT37wZupD6JIEfVkw588ekejRrwCynlCgC2dbXPWUPUyIPJyDC
f4Ma9GCtwK6O+ISMTewTv8k/dS5OzC0R33SHhfVfotS91dBf9l5yBN5WlVrcOD43
S4XBUL7d56Nq8gb8Y1JTGuMTXX8fzRsHMsrenOO1AuCiJJVvy8Q75UgBry92TGI+
npEJi4fYYNG8G6xvkaX1m8OCuHSC6hF9GqwqYITsNUT4RQvnHuyYjawdLnNa71BM
gr2TgIOdWV5Tb8YF72XAxdrs5d0qKMDCm3jqZJQT18vRCUY6/Z4L5y0eOCf/iWXJ
gOUjyqk4CTBzEecznGkiq8ah1e1Cnbuii1HAQc3VVnhVNP92oKGFDoQzM3QcE3pq
1I99qOuSDGalkN4abYzRhcogTn3p6o5XF+2GfHlBf/McOwu4uFt7fwmL/+DxfTjd
5dzeLtugUgd9uOgGLZl0I9H37uxgsqfe+1adCLcfzQfcbrXbqHi98vVZie9w/TVk
mp2b9AFzrhMQ+NUw3lFj9pmu9/3qx8StHzRs829ZQ+FiCQEQpXOkyR0b+FeWCjUv
b2hRUqOypasTHIsTGyq3Zz6BBpQADybqFaHk8p2Mnws=
`pragma protect end_protected

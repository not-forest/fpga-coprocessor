// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
BIa/Odzy7Cn/vvPvkasy1MnAyUKsKN6AGYY6g2a7CPWRSS43BtegoQOJ2JiNq/IcAhzq9/gDooS0
jZIvJW0bB4r3BKgRNhaV2OvJNUzihwrmxHEKDg18GCXtUiKQk0YHqwmaS0Qae2+c5q5NmQJ5v4sU
K4m2o12yBvpQXtlaTWp5jceKU4QTB7bma2l8BwJaMK2lSl4bE1aA5cSKhPtC7P9xVwRSZ6mzDcnF
hVb6h2xvDmB6ZPH/igfl8NDT6atFiCMTK22WLh9FVJ82sgu6jJFjZnAodFVENHxci9NTzvQ46GfT
ohAUoWtDLmWvM7+LLpvcr7WMA1pUTQJCHHLEpg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 12048)
eErpuRWNU0WC0ouD30YDe0aJPEp3luhrVuCg7qVOrW5sYUuFVBGyRt4gRXFtvyKg8FVfhAqeifAP
GNn7rYoLpYUoRwcXhGz0dhzHZpHbNiEHrbRTO1/RQOnHtcS/z6joQZh4HtvwYQYA4WYLVRKx7uc1
cXXRhBT8Tiazbzcy8+D8++z91tfEbgDoZGSpiE5aInb9FMLHG7R+WHAMGhcVnmDveU4EkM3VwEnr
kK15C6Qxaw/D+MmNFcnKu9scXDO0rzypvp9BTTaANLR/Wp4CSg1dSvXdcYuGnxifGWZRQcSywj3z
8Ug7fJsod9hY814HQlL5oiY96qFx51h4S5rMhSkl3k9Towk4EmmnUC+WqsNm6Dw+wLCKYTfcThZB
R7roHygkkajHda4Lg2sJdUs1dY77E9SGyzRfSWcHVuXQ1V8Yfyt/g53RcYenh70yhZFMhq9SI8AZ
uNgcR3eDBTPz8vp8UniGPAoO5GutAzw8J+7kSl6eNI6bdf5YbqUjXNK607k26Pd6cTAGDAwdqLcK
8+iRXIJde8p6yUSFbeOU5nWSSG6K61UVsuHneb4zPUp8e2cnZTGfyRE+wrF8DLi21YG2M7bt6vNt
rs9le63xE8IP9VsOV+05wSf8kh7bF3yO71f2O+1O/Ol0C0wSyhBtV9XOJfQBrVNqgZksrt3/ZS0X
gdH7bJVKhii9FBND/m4/yYvxIusASoRHiyod3qnWQYDi4wFRWO615s/CunAEpY1aaGDZcqCyEF9t
FwyRnxMiQf38xO/gfPftW0IHN1lnjNZgy6+SEfNwH9sQbj+P1ZkR0yW4AR7y95RY3PvKzz9MenHK
xizDbk8SndaLEA3AbjRBifkG5MWvJbmtyc3zzFfrjKwc+gJvB9GGJTt9gd/A52wc6lZGjZIr633o
707BCvA7NTF5YWJ+gFwNO9xSTDxPI457e6iCmtTkKnZv2k+JXgJQ8C+DRo5Cy7mQrzHdtCG58Uw+
Mm1Xh+820JLLvXKaGsWTweTO7LBuowfeoS8PUl/jHY1EsAT0J/sWsb5qNNP5m2QECzeK3nOluP4s
QjrjIMUZ7Z5ZkUkk0D9SQgYt3GKeX0YQTEWuPBxEID3YV9PrMng0Xvgnrmd4871vuBNTIv/UePuI
UoTcc01MGUaHdiLENY2eCHckz39sW4+eOnhPnmC2FfQd54E0ilj/I+PazM/NGr9SCVDOoVnHA84E
Pl8xsxeuI8DYkayR95vfnckQDI0gYREZRFMRSQ9duNSSDG1LFHpGKe3s/AFyRIZvS3aADNzU4wXn
Q1rMWXYeFCibyh7ASoCnIqCVAbq+RxAqBJpldEQKcdnKSty6cfxRb3NCfdWWDBV8uhM5lye9frud
K3ZOHfiSfFSB7qNNb3onoIpwFzijxm3JYqOqDbMGXgq2oGNNram3Tz2EcTXtAcZEjpvkcP+nRT3K
vOhaPBh8P7dpNaBGXEj3nJpUIPQv63dxNHNOkizp82btFL5kI4PBlo/GHSB9OkbRDZ7fOP98Kd9k
6UX5KqJvhFTwee6pGCil4fSAVp6dMeWIkITImzslcKandDy8Xw0kEQ/M39HDQIyO+fCTO5mXLPqE
xMYPa67jRCeZ7VlC2oHzIzHRgwRjuIZ1rXgppjqeMr2wOFOfjc51KtCLIfX31FRu8GB4qW9bdpCa
+qCh3NPC1Oiohzn90R7gCkJyxFQyoqVfFYvTsorvRsy5z9V/9J/1zJgW3cdVctDLoB/Abd4bi8mT
iL6MFRR4+cHKoL52pHB3KQu9+4ubDkMLApqHUwQg9HfrTW2sQfVJdiIdhQuknbxIbRj6b1y2PmdX
DmbTBdD0De0Ih9QkGI80Aeqi60OnV0tRqJSeKYO0vtmYKw1/E5A6FMPjPMdLib5kWMzeBslFLwFw
V8Ck0eErS9b27LsQgOucDXQxs8o1fn2yxt+6J+ver1n6anWKeIrLfdjbfbEU2FSTZdtbITVpr1/t
AtvZXuM+AAVhwrgzrCbodjLoCDyEIJHuWQgfBQI0wVIp6155mPKk0tw8igiuNfvGVisJBdaXGUMv
p+H4+hUAnxjH08pNSbP2umb1BaiMQL5FuyoHXtf0Ou1U5mey3/T54qGeAK0mc7Hl1NcUNAOQjt0f
khA1MAXC8Kv508zcLqM5OaNWFkqxAgt3tBfNONyW2r9IsBBrTnbkUibUByMPnZOvyzEEF+LEtuDm
NZlOy4XoUSziMLlMuCqOwlJpIxYh6bydaOlamHXOlS8Of61TjizLRvT+u5mdUujQ5HLmfyNuCmht
WQ3MZ2lmakHUB5Ny8/zvyhTY8Ny2RgGX0WWTa7fYdB4hZbQ2VuzodJOrDm7ZHfoxUF+osEPIF0J1
dlTXi0Oj3otZe2r0O7Az2n6h7W6yF5Y/6cdBIVvq0BhigjwAdbETUzREtb/PAxM6QxU5lWA9vWFg
5WftR12JM+PgyP183JpuwOTgYIISlSs2P7nDi/puerImCwFbvb7CY2BqsFNbFAWlCzkOxlxW/eat
fwvpsnISARE8EnDWOwKV1c6nt1kIB7H6ewG3ZhVeMMxh2TKdiTzEAV+MnQc60HSrQLIXqBU+7phJ
ZiI/JuUpD1vneITK4vvHDTyaQBswfgl0nGRus0KnhODlZHnxm+cp+obhzlhlFJNOpNMOP2+Lg4uA
XebfgSeMqvrkPduURDl9whDhPm4x90RLER9apWp3vAIKykZuw6cilIMbdzR9DDGUv8P/ZDNBm2QT
CR/1IuN/4fFevXNmDVJeo6kbd3yPlWILhDA8oBKosLLAMaeqoitKRU2lX+ydsrnJ16c6vx0ZlGvV
ficRRerWMAeoE6kZavy7SqqryflQq0EwjlxC8+Srd7fQ0QXGq5l3q5x22u+TogRjQTYJPTr3RwOn
VjbUk3YT+0R4SiI3Qq0Lnsuf960wIsvl7Cq1dalqmczkE3IPbj3aiT7u3oEULhljbg5F7RYHMGtb
dt69yUMgAZD8BUiiVu03LHJvjfRXaBsFAt98L4xyhlAj1gQ04CdwIBEMaPK/cloUoHgHwHa/Y3vT
F42nWWrujBRTNNJue7B/hWKUR6JTwjnyXzpX+Yx1iV1YPunV6SRakfWYXSQsr/2y5vfUZLBstAF7
n0xOnoieMoEQQQdQTXctg8dUbK3y514kWvpzdHe8GRE97xLibmPaoaSts+g5vCE9P6kDhQkkZuHd
MPZKZB9XyPHP6Muqn17gDIdOP9j/gYVTWzi//j6njUJeJViGxyKHerwLdnP49NvmsHe2MB774+ZV
E/4AvFCkF10OP1T5GtxsK9HcV77o/m5PAqhSeCPZ54QaJQjU0XIlkuPpnJ8n/eIrmooQWhYx0Vvl
JtiKtUxtpqcKllDzBdJ0e/7sLpNLsGH7iMWTLXAOy9J88gZuBu4bY0n5SfQrArjHZ2wTrU0WvT6k
rAsYxJeqKroKMAbnFs1sJ0LG+cZWk1zyoE3D+OXMxnKkXVbyhX0cPwkTNvKIOlGLHkY48kOuX7SS
KmUnXdT5MnYSWiKqbLDPKMkbxibjO292ZGURhpMrTR26c8zpxCjsfp4Vsf5DeO72jD88/z/Ea7Wg
LdQHTjHtjrfQh25MtTV0reTnr0d9J8og5iH2VWA53dhakd9ymjkJBpjobpjnELLsw8GUvqdNj0kB
c2wSJ8d70oYC/0ppBOrCdmTRCoDrx3YIb7DX9agndmvCLYJXQ7dv0S489Zd/RKi4a2sT/3zf+jHu
JonJxxUmQLCNfulC9MQ12nz3/uChXbNCWP+oOwVWpq9SnqpLoavhgqG7B29v00y/ZGk5AKoFcFYx
WqnK6b/BpULtTHEXnoZ/a3qDrP/sZoZ9cYOiXdxmZywAaQfhvj2KiC7t45lLjD3MfKUb7GwPss6O
w25J5y32jf+kOvp6Npxi9rpfdQtjXuzgnzT3X/JAl1hj4P+TiE3kPHydSt+hFL80Jq1B6iC8LV7K
2GkuZHObyWDvfYq8jlj8B6FXd7O26xJ72xdQ8Bmz17q0+7AmHHuG4lZMP/ekev7MbjWCE3Ur1i1T
q+OfEbN1DsD3/l/KGCiptCteXjSn+qm71KjTtmaEutocjw55f0xV4R9VCiBJ/mw4xxo2mqjBVLN9
f+M5BlfQd8OiwQ2Ha8TPliFlXpEDBtL+XiiAWEZIUd8olADwFT69o0QyPJ5901occmOUNlbgt3N/
magFdVP/CPH+ozfR1tp4joLUbzWe+S/cdEsLi6jpH7dFAL+QG0Bf4+RaK9y3QGyg1M/0phlnjaGa
ZgWaGCZe7l9ZxQgTktoI4/f4W9r8c1bh4po5ZU1mSd7MPZqS42N4KfFnv5Bfkzx6pc1BAEw7Zw1u
+bAMBVEILz3/sGhiwVGc85Nz69u80GJkw4w1nIxNxvYG01ZlKMvxYo2lbv3zaVkeEwfTtT9NWmcz
WR+CZfGYtwbUgzEjIx2xH2GrXkf5ID9gQ1HQiua0YPezkry02DOC9p6P20vDu9uam7QmAluGTNvh
d7+1aGW6k7nmFchGERFBgME3mgjJIdfoUCKKjzu5GkYkubeYhSQ/IOc242nm4fDDprDj/fPyHwMO
Kt2KqqtfN/P0eVSlUUuSayJC/4A0cD+lNj74w3VJaYVB8T7nasHdhL4EjgtnxtCkPzn6ZnDS0HVu
kILQfEstoWNuGaDrO4TpDYgA5peh6knBGv2KdhqJSE3aC3jISvVG7u/Rh/ZcS1qELc6aHjNldxiz
VOUd0iwGtPXJSf1xDTUMlGSps+FRjR4k6swo9pOcdwSDXHU/uyE4Wku90P+KocY3fv0NyzFXwxdv
ffX3lpMqB96V+JssPYHweoPFbB6rinkP30f6+UCsM0Bykw/W3uxgYugjD65WeGHCf4HZM3kCIx7H
NMwvBQ1fbvXCkQ+smmVwzgYB6kz0iI3SfsUgLhTbqwNG/mZgAOeRmyauUIXgXmYaiY7uEDRTUKdY
pfJ3deAvvsB9NM+CIO/VF9Z9LYQCpnIqOO9aUkJ6DLdbez5eq/uPJ6N9dCWGNhhGuDAdhgxyc6w0
O9TGndkz3hUaSomz7I12EYf4rSqt7ofB8f/WQM/1ib+Pasd1gNwlUW/yXmOEdaEyZvFxjys006CU
r8IfBO5zZ+NfSlHZ3QfmHSGobFEKDTCJtUWSFMJhWykxA3fcgV4Zo36absqqXaKSIk2f4GmQa8EM
a0c1HrV7m4Pju1ZI1QoMP8a0osgIpZM84liBE+c/d4oFZmlTF5nEc5I4Grxa3rrNBnk1K6mLX/p/
j3UF9Eq+PrTIeXgB+ZK/Z0Q7Y3B6PQZoVT0D6s/St3JmZCXkV0X5LnLgjGpwevDV+jTq7uwtSX5C
xLeLBHFu53VKMQJH1uHNg19H8pWHC5w1ug3hOhMZ81M9ek3fM/Xu+3+ZKFzCXOrKkcStPZbtgG6P
97ibOgKY751svNXBwAFINHrZcecMUOybzUxumiP6J+sFaH9fD8UbdGrQIBtoH6exAjGEn0afYpMz
S30kWo8+N0T6ap1NyKWyrOd0Rz8xrN2fBYL7oH3ISFrHX+kBb9OweQEgjkUooQRYfdEnmnpWazl2
rkJa4Jlfv8g6s8ScAh10cV/9fhiULSAgx7EYZlAvujQ6gvWkSGmicZBk+DgKOcDNxwyWpIxolZTO
Q95Ynr/cJHnp8CMdHhhEpKUpP97q8kvztDCtLMKmAUiqA17Z6wOrWAT3O/ST2rlnccZprpQ30TPz
kxwnmYmMUu1k8xz9mfKt+2MZeUCKGGMdvSZK4ljJRcd1aCMu7z1nr0NQnsdQagSMobHc9pSAysek
fHQWgVGPnqRTAxDiZcbXxqXIvuZXwyIa/l5UZj1Im7zuDE4qlvcIXOpzky0VpFCKhxWZ0dO7JAQR
TVEKvmKRF/vJ0uGqgPagdmP9xf4ki16aVjR4YNdp4CGOZIkwTds556BV26Z8JhJub4HX9iRn/JaH
tzqeyQwbGOsWBjw9MAUgltt/PIRMAfFkmcJTEV3oBH3swqqGdiX6dUhrrS0U6trS8dsD+VU9Kwjw
l7Bmwv3b+EQuXEYEKlMlDyOyGoKwkn2FnZFuu5vO3E+jHNJONf2z4V1y70qzTTb1vZtC1gymO657
9li4KBRSMmwciOJeQ04BEa2Fp5LMpr9A5f8CaYditn+VsLRG/D2okh1VK1JKNOoT9ODNiQ6i/3He
coZA7ST84NOO40sscXbfsGDlrwbnDT5e3s9jcXy1wBO6U0dCPWgO6SeSrQn22Evumu2/6IY6rKwx
Uniu7efxCjbIqxmR7ncjZrTCBDESdZo5kanYaJWbZVhm6f/WPjtfKndQkMFeG4Xd3B/YUyGcrvxI
41HBrqLquSoDT9zHnyLcTm6zA7UNrxR0Utexw36sPpKtvuDDGUPWRMbTbHhGJN5l0aENdKr2klsd
HuU97yGn1iIsCytrOtCYDzZKMGvfRBpEIeoV5KS3p7V7lpoh/9Qu7qfRV+1eqmaq97IFu3I43V5H
JsxpvhP1pEepg9EP3iLbK21jPA8wwOxHWguy/SGzqGDukUpLrX4l/kLOtjrTVQJbeGrdW0YPVruE
ifFpkR3wwAHpTZpstAb9sRAblL5OU+XbSN4EVetoW2kAsetp51xc/RXz0nvVSrQIxr3XgBT1ahU8
Tb8Q7eVnvwpK5XFW3+GVX2G3N5WEihgiRy4ZYTS4ZMmxUqBTRuPUfMaZ2BIJXCWHqa8casRd7TAY
T77CztWCrPqKTJwepWvs7g9zopy3c8kes5AVsW9qd09SF5GuNcQEBxum9uPMcvXbOPgexS5PiFsD
vYn3DEq79gBXkoFBRzEt2I7rYyAIZ7RrSZAD6W/BfT7VrwGf5JpJWbV8rvox2l8xNoeAFDTEB6I+
0B736cMOm4GvuU+d2ipLA1chQV3dpaOiQI0eQVXlwvmGuHNjsX+I8+23cWkha4DoLlC3uGFZOjdY
0BVtANIHuqXv6t9m+jFllhUzFH4uF6B28e1suVCjpNPf6ftQMQb9SEhGDOIB5CdE20UJjGOMmsE1
rYKQuq3bE6p08+akrkIGbV4109Ur3+RBQpP/VrzUxFwQiF29MQjJ6CDr7FBHBy/3FF08mikI4RO1
DXY3D9uyGOFdfOr4YB29DKy7e3VGTxd2iO1x75vaVBzrGV/qqiYBgU8j9CfBg24K+6ihcNeZxqWL
DO+Gbm7XTcFAL6wVpvtiLRllP27zqI3dE261qXo+lZg0tusrKuBHitaIl/G3fyILxSG+VmQeSoDM
HPkg9sbHXzqp1h+vmI5YJofhkq3GPKVLBHPK94zW2EpNJCdP+2htE++IdyMxCj06VSAyQQhtKwPG
0GD9HwLr1NLliMzaFXE8EGg41UOLc7syan3jepQ6cO7VOAFDOXxB8znvByACUxj9L0JgXAnBANHm
m4aZ0UQnT87GMGZ6JVTEJo2DztRgH1TEhogJDvEgmlx/sbfp5pwls+0s9/vWM/U38IiLkpXmDvmM
ZZWc/ZIv0vHy/N+tWN6EVTzM/IQkRQ0MsfccNd4oOLLxKvUMFStkz8OkaZL8wc/UPLEncHuhqnwF
gNm0AOi7K5t4FxrXODr1+ISNc4wzkm4oS6iEcXzf3cwx/KK1u3pZZUjwbvyihrFMWw3CyUC7nIqd
9wQSrE7uDUZo5hg102GpVjzw7vHQMOQ92o4NDVqY6xKm+hgYFt/AOkLX8XR9eUKU2egET1PuznQx
BMuQYWgnfZfgPLFAgV8YYBN2Lq3gUusH9uGuBMku1QUgw2J9CiLxtYpRDImic+PiMGSPnV4bGzhS
pLmnsqBn9oqMWUZqd8DgevsHJRKN7qqtkQKwXbpxx4KewrTUxc1HrwihVDW67TaUSgy61veyRr2s
hUuYpzpVVjwFFoni6inUHrHjS7zkrv0h75OyeJk+IytV4kwUWX0nyto/i+QIQ6grJMZzMBbTweKD
0mdIPM5+VsLdf/LW8iATKv7CwS6DrwDlEnQhaFcJoxKhUQe9XhFxc58hu3Urf5EJ0inu9UVSK4MF
LBYAdomk1D+tpLroHm53qqKeFrWzcCaM8unTY4uSWrqMbb0BYRrolBNBZJe3y0hB39tJUpdvgreo
h8IRXIBqh3EcgHUf6+xLp6Pt4GDrF8IdWAWX9QcXup0mnqS+Le6WcGYhhFmPUUiyTaFNf+xVcUl7
OivmWzQA6Kqekb/kfVUoZbtF3rRTXuW3qv83AZSqTShB7cvi0up+qg3DhHtjY+iBXZHAGy9Ws3QU
acvk9/0dczFTWmc3uZQwkeZI2DobxLDjpDrmI10YSVuWh4QiI539mQyW1Jl0tj4UFWkUEeFOgg4p
S9/EfmoVf1fsB+9NxJf5HxXYtCWrMPaVKtKFFLWN/2zl1OYfbUXxQFEM/qZumAX2ZpYtl2LSK0oE
5rGDxMnCKLQqrwJ7XA7TfyTJefyP/8IFbNPVVQSiPhuSTjDMK3mqMiTURa7OdEVCV/XOdrPqwnaw
3pCsyqwMlgv2/DIhh+iFhHuZT7Z52I4F2o4YBFwhagBiMRcnYNcSEG/OIeNmN+O9zxnnSioubAfl
iiyJw06TEx9Rug6yseQkoTX0NM6wRr6yCCo3eOuEG+MfGMzkOJ8Kb3eeVSjo1hbRVMC+XOqvvxLX
LZhxxE5/RNE7XNmmdnXXpPyHqKmqWD0/X0gChio47rzHPuJ3hf7qyh+OSAeJaA18ehyNytE7AspR
Qdya5vxu6Eq9JWj3hpMEh/UxDra6+G4K1B1ZBqlujeL19KqXEVTiYIvrv0/6XjTJ2lQd6UsORdFL
0+vTcz4wLl9avoSD6E/GRJm7iIuAd9mQz83tzUnbAk7Z0m1ZfwFBiFxI9XW3bSQEqBIBFtt5geC3
cFOfRz9mh3dr2epbnz9b26vAR+dTEEdd5TUbHUuEG1fj6j5g0Rba2Ij8kg8U1gp8Lo7G7XZ63S1+
rPWLOv3sxV89M9o43o+71f7cjq60DqbYNaAR8c58c0xVLn5cBdQb5qy2JrEGcUT35c023/4zW3MY
qVp22DH9oZkx1jhReOGyetTzdU6gQsBMot67DohgR9uRGtO/l9BlOJmcFuq4ixh+OKVavHPsXShk
sMZoeUCCKJy3oK/i5ovnPLLe1XhRVoqGdR1hzbtupmU0RWZubzg5O1QoInW98KVneABPlWoMih5E
Xl3Fb+n4C7sfj+38p1fgjZOPfS3DXHHK0PnH34qHlK6QBbneIQHtuG/4/61Aei4CiHhQkd6iFuuI
gJAmIs5NNZmR5Ywkpy5dXjqRDYV6v3GJ7R7Jv4bIHZ8pabNpvVlkuqlXAha7AkYaRU1up3a/vmCc
Ja82ymIa0M+IUcJ686IQFNcavoQO2OrNKq4VGe9dPNZzuUj1IPOBxTlD7HAx2U+7Sdmrojcy2wU2
qZO0+vSC1fP5bSOP9REixCs++zh74Csz1kqEzQaX/RQQDFdVwQO5P7RHZWfidHM96WBvP5hr6mKV
m7LohSYNWtCUGY0HIyCjzOCVOWWL06N/ifrJmoW5f0wdSA0qc+GX6yMK0RebEvnus6otyXMqC/Kg
GPGxxtXF7UTsMsxQVS/X9KjeFVjYy502BBbEffWfcmjCUyvm1xsbSFc/gHStG9R56qGHn4Za3sUr
WDEqq38poVCK4vOT2fYBBbLOTLYoMZg8Eur55Kwt2vKfTy7AiSET8hIyThd+9G393H6gEek0NJGX
H8tlxmBliLE9iXBfsbU8ypdCL01xdZwLyYJv3qcATaClFW0sR8ZZPGElAPcgJqx6jm9kD3Ywwo41
v4tkqW5cLJRkUk4SOMTf2nRHNkFwUpHrqs8al02Y2SdhKFGRI2DF6kyD9jQElX933PuNG/SLg/c4
P8pdV7nslfLlCoq5hY+ZXsdWJfy+QHMbDqXWCKgKq0zMLbc7OacvAqT1E98H2e2vdMR/EnoaW3yW
fNhxMrvuhr83lrlxSjHHhffWO5rRrArACT7SCgwi5kt40lsnZQvnL0ZBk+3B1SEV3++PVAJBl8n4
PYh6ReWjei+QXgQx4Xhdw5nthfrw6cGBP4LT9SK1CKgJhUEDDTz/oBNHMWBjyUdw8NzLei0+6uKM
QND6ms3kTdgJL/DuVrpLVZVysyxPSa5vEovOIuOjsiREnbbbn53adnqFQM6yiwrqPYpa7jTgqMAj
16LcPhiM5nFipbHWtddGeSH3Zsvgl4RjlsL5QO2t52i5+6Hqq3ERDN0uaYpb1JG08t2B+/+hTWIy
fJKyL4nXmcVXZYZWDVA3b8v1JEHO3T9DZkyfqdbwjMaKRXrcsO5jfis/Hyq/lQaTzuQZaUKdxPvf
tmD0CrB1WnMQPfqBibIkJFtemXTwrt4/FRVrTBL+j2KYaZOW3cEha4J7s55gYXtO3YoXY2wMzGmJ
NPLp81l7bsc+O12qcVVk5EWTkL7yL8mm+OPaiOrXAOfnvwuDTNSgWhDtQwcpU7grDOBMxpJxuF/Z
3GjAXs/YcMeWdwUUx7iF4XdspIeWgYmYVnvSVx2W1MP5hiSIg6dhwJJJzfFfnldEyCgi1SbrzLl6
qu5LVRrSZD+/j1XVvg4LjhiVcgIvWrf6dv99gf1EqxOJqfea1YZXPnlOjb5mtnRU+1cF9N0jFZOF
i56nUykQgurt62jtRq3Ehhd4mMguY20uJ3RER2Zp7BD7XBD3wegoBHVt9k0pBEkeGV3VCHcHyt2R
FKYXOnJ48mEgXCUXpIP4eW42oo454tLn5v1Q/LISTp1iPqU4Pb9jGUw0LfNi/yg2cOL7Dz2RLgEn
CQrWCeGXbN6mTbRLZLjWIcVVKcK3mL44nKM9pAiZyXB9TS1Rpglr037f9EBLyMaTVCli1cejY6p5
9gGWj8EhvGCODdekqyQQDcF+qd5H6101jEo1+9isotnGDSWfHahk+0w9QNA4MSDVHWzSiNFwG6wi
FJSFfsuAaH58eMnSB9mTS3IBTiIreKGJOTErhVcfWegBdwcclwRAtrpJ/4bBJlH9cFrewLuQGoUh
EnUXcSBByC+dLkLhA0Id0iRpN+M0lIMJBs4DztE9dDOyDKZxSORvcLby02JmrcGrCRpM1DHfM2d8
GYsJ82YZ3+2s5JrTrmX7MFUG0P68XjgFvysvESviT0fqYYhyEINAooGTvJa+CyRA57HedR5YfFqD
kPnAxo1IumQjCHrHsKQ/ald2LzA4pcldtRCLEpROpdUkUoetYlBe2u1NqiO0mtx2F0TCdsOGgBCW
RNWQTrrqxqiR/w46lOYj5FfZo1blKDNSfq6NQ8N9C6VqjjWv6pF4a7ejLNvy4LwHrEkMKJ6uDjbb
jOXpcyMTEJLKvYT6Kmk2JxVvSN3YdLTgkbez/2mly/aA3O9OkzlR73feGpxlWaFBYAJQiaAfNCrC
lDEuJSmzl37JfAaWoJeL87XKa4FuxuBW++EE9RiGQHRiAvRf198Pth4JwL7gZwwlp7OEcAeyaiO4
HzfLzC0UyOADXgH1pEoX3/rZcQyxLjnN0JDIjvB3BRtpH4PgR2GLYUK6z9GZNXlPaAYgP46pGsT6
PAgwQBWleIKnVKitxx3fNY84pZUrEcqxUkeeZnfKdO32wKLD1zTFIcEe1DvqidCAhSGOQAEsFsyT
GFUftjdOC5+3ypeinLnJavA4qV2t/O63DHjhXkqIK8oeVp4pnXVP2p+FOSXdRr2EhdxTlKpqXI76
8Vd+ZUV0YDNzpHkDOD5gMgt1s0xHVWnmpA4NRCuRsTR1qBI+E06pSA19vEE5SnypaQZWzn+E2s9p
wZwVmCjWq0Zmui98VFEksPGGdmsGlBad30ZP7R8/joCO8zCHoATbpXV229aovFZK4jxOZg1rAMs9
YRDp5efMU+ZG1Vvm0DJf9909j2H6feRT6HrHCN/QThGtAhORm9yrgn/AdhLukdbBwmSN+8Cnu3+y
Sk0qIpmTlZ7xUCUI4+yVlkuJS1rzQz11NhHYxC2QR0EO7OtZC+qkywaESOEuFh1H6Lg6VSpRUaIK
PNIEMdMq/QfoD3pngZ59XCBBGMH0F7MxETrN+0Qz6xk/9E2BC1n5joA5KKKVQemNkzGil/+teE/t
zXuVcAcy4PN21FD0djcSz0UD/Lpm4sGs2KNKA9qfP2qp2nG2l8QjSmKiFewcU5YxSNobxFTPmfEM
ox3tflxnxTBQTCa3FrhKgfGqu5KU/nm7FfZstkRdgdzjDh6qx3Vte6/oLWvLLDDXfMjANR/gFMvO
Jta7Uq3dl2RiaJKGGjxeDu7YBf7ee42J+AnPtGyvEFz4ez2LC9WG0MjATJb5WUnN7XfSjcd7uswp
xpxJZ9Ocbiwg0uyJhJ3/zgpGCLGP6Vxji2zOwhtIkHmipnr7JcXbrVHlxrmOaPtCHcVYRzL9ViC2
kZi74vHTX1Qjn4A2KgZC3HY+CVBnHPreXZKfHSp7kNAZC7cIhselUtIpwHwEsesOqX8Ysq8fvet9
+nwcCbgVtwKIWhsBaPpb+4HJs5XMyyME5pu4R2Kza2snTTOpa2JWsPPhhtvZYOnJ1iAzfV7X6WYy
vRchWNH/yl3wZ+pSSiF6RXZf2Pf6p4Isq7nPYGsL5Wgyvn/DThap9uiUQmCrt/yKNRamiV624FtE
5z807tfluHAcJ6HvxQNgEj/bgs03pCTa4LCSFmfEBWFwBYERyqnqNr3RjmovFa3EbSk/8uK9li2A
aJNESDCl+p4qCUYMUwHYwnNxqMRnI6QlY4WORXD76jRZHd7ksrjOCBD5qnPCadgyvqTazLcjANCA
+/LVfCs8bT+qog/xJ/WhMYvslDZVhP3TiQa7P22E0mF5bb/JTzW90a4Uf+SZ4aGoFsr+gwofB+Pi
78RX+tdSjAxFqlummKeXEFRNg5bBEtUGPfqQNCljxFtkGnZEMwjnQKPi63sBILZ4xblYEvEjWnbx
Y+ohcyCHsdKFHSjWL25o2Uo8sIU+XtwrYFcYkmPjS2kSKQJVJonZd0pET+R3IghpkhI/2z31Bm0/
1NdEE+rtqGdDZbeY0DX6usDhh+ut8CYj+UYjnljhWZQiQPksY/UPi6Rzn+v1TQeS1ZGGOLJTbvAY
dUYS2X8ZV9NwcVjQCbs5Rf+7qppLYE2TJMwLzAMp7abdIYMQln4aYE/nUzoOyIc/PAHG045QDLAg
T6e9Iu6F42DjCwX+UPblheTGXRGybaXkQrdSmCW8aSwOw1FIQYs7px0k0Oe2bNPjSZY6cVLhBOnT
uYiNLPVwWKX+K3vxqDkSi36IWQpMvIXavSKL/evM0JqwyCE6OccqyvhKY+4XtRthkn17MseUAMXp
pGmmRS1+pA1oqTBpFhc4eK8nB1s7RccMpYkV84hwx0nQehe7XSkGWpFJSHCOy9Ky3EN+H6gSkMJq
d1klE801Oo/nH0BAW3hYVZpIzBpr8PmQiYc396NNWtjnIBXVSKIV2b5SLvhanlHaBQJwEh7Mt90e
eDyMMgoL0ouPUyxOgwocsxQplQp4pufszn4v8faUr1CX1vzz+YdEellrKzqQEZFObOdgQzFcbRXm
kUoFJBQ54ypkyw9WdP2DeZBgYFknU3Yu6EFsIbEyU2BQoZ2WGPAZsUfZ4fkFBXTpfjp98WFyoFt6
ABlROGRfXR0O2mQdYTBtrQG9cjiyZ/2D3aMLOBLP2gX9UsctlUdrleCwbs4KzYEj+zexOL615bHE
whB9Qwt1iq+Er3j+Hiv7RNE34dK3eeC6xhdq+SUZb8ZH09rfEdlzyj2hy9YtlhGGE4E+J3XIEpb1
n4sYfkbZGuN4kNs7qxPItLi5Yy6fxkvvPnVQS+duRYkBrkgToMdoBmFsym+3l9lbbZOa04rOGZTd
HaODDKgzF/CX1czYLau2GMqFRNALPAL7ZpMTr/IkTXfxuJAGSd0sdBRX1vQxvKzKa3fQABN8bs9D
xKRrfBJM+G62bUXkxNYlZeCoWY+/6PmYeZiG7WK1M8/2r4VHGF3gLvgT/cP8gRj1R7XK/72jphf8
K85shWKzLWIx05g6xUA5GhxqPMS/yR12NSt5gKI6fpgEYb1VsqjEUrGCqg3MZla0lC9tkihis9Ji
xFG4BnA0ncL3F06IKR444CR4+j2iKkuS2z/HGRHtSOaBXdy1LWlNFJ7IPgz42K4LbD0pHRLweb8R
HG4H6+buyZXN9/51W1EaPlj+1wGGRcCwS1OLX531nUynGDv0etlnTSx9t/u9US32BRuJQcnZgmhk
e6Ma827XRJNcHmToez7ZNsTIFHxC+pffrjstQkE4Fe4VX6UIfO122HVUli1PJJHMcWCFrkv44UPl
AKNbMIQXdFG9bHZiWZDW6khzBYgesq+7rYsEjsoiFCi1h/LIkAqv5D/phCIwRKuIQMPBwqWMyJFf
YMO+O+4eilor0eN/2PY0UDzOem0AE3xlcogMeAoF069IDXn4hzsFg40tq0tK/whV1tYzhKF0QJs9
GRRvL4l/bsE2QmQJ3uxaNxkblFT/QLnYyZ96ecZ59v248mS/Glcn4xCAmO8cNnv4ygzpSahs1jfu
gnbOu0RcZtp/DRu9btBDmZ37k8JqtS5x+yrU5tDeMwpB/gikJcE22xZYORdPzjjOb79wZIrYAYE+
V7PpMi1sBeGUFH/cdbK/TqvPrteRhpZ73m1AAYRyqcYMLZV0rhBFiiaZfI7AvgtDmx7fMC6XdxL5
jmlYMB4yH5BEGJ9envLgcA5onzUV3drCc8rC1oszQ3N4ssnQWeIE1sUqePI0pvIlTw0bKdapOHa3
SnZ8Ht/lzUFs3Nr5nTPLHSM0hdO3Aph6y1rJTPyQ4ZzycfGMbuGyOZskx+yi3Z+LJAONS3oKvu7K
RhmQh2eNibVTjhYY5VjY5k2DvN3CTSZ7JRr+W4rrBVnS/h3OpW92SYLgnjITgXdpPYwsA79qMe5O
AYjXPpcw8yjHyNWGAXgbttVmUyu/XvmazO7HGWi2FiicEZhG1AiHZKjhpXXxpfM3AVNclwVAteQw
JH36BHIA2+sIKxzT8pZGG6P96E++ZfMfjed36D4Ir/rtC3CnuvbcuMFpBcLmaBo8SKQhCGtSbJwA
9IcJN0Tm3UD4tpZxMK11Jap7kE5KsKnoOhEXq4po1g/X0FUQdr4Nz5XpYK8NFm4yqx1/qORpPape
jUqlaNGDDslqEMru5gwAON3AUIAMwmeDwVLh2QTODUkq2HkfrO2C8v6RKjyFAqys6/nDsA1TSBv/
p157Ms/+ZUW4WP9jpAvAv3Nw9bks9c1uZL1awOnKRtfNYt3JPPq72kuQttzvMeFpQ8HOYaK7mysP
3enuxOTq7PqJ25rXtHr0Q6zuv60hqt+IjiPf0NYrfSnC3EL5WmY5+rChkAADMCH+ds+GOBFOfwvT
IebCxD9UEjsL35eiOUibvKEgEkA+59RvBwU+yLbFZG0Ysg+GenDvjzthhBctl/lUBBJO5RlTKB1D
tXIyeUzjlEBWoCi4fMcMWCPRdwBTxuAGP2kPzSJddMWywACzt2SUOvcCUADIsRC3lamRwDI0Qwoi
ivmxDxyFAw5obwAvVuaCF+0E8R2RVP2OL0MkkA5PG86vXhUOFkBLJq4nAJ7/AE9RCkPvIBHlVGxb
KZvTokfFQqgW3XDkWrfnSRyLthIyLV1yiaRG8w7lgGhoZbYmG1+woKYoufjvGdqKvTLAGLQQBt6N
JbWet/+48s7FGUvgZBEW+sBPyHfQv4kxU9XqH01YuBM0SEZwzBVtS5qa3swQCNFK7T9TV+P71sM3
9voWagKvyQDS03ReVB20YqhpsQatkLGpc5wXc+b1TsSs04EWrjz8IMtml98Ty3jf3r3R7IYjEqUL
ITIoCqrfHyHWnrAVzTWk7kAfaDUh9ducrjDROK7FuDsbO+KJsL7Mah6PWAHSjfx64pVc1RuHd1BL
WKVgGhq5EqpFji1PtTTF2C81Jdr/goSe/km72pjO6qFbMqCL9sLpMmlxp6XeFeQd+GLTI8ZW6hGC
bq1jC9ajHmVFRfAfVyiVBRZ/fdlv1I1R9YZpDsu826kRomumY9jJ5uDweCsLgAyEE6pq0/UJ38vk
VDw9TnaITZcgF48WHHP0dO6xMuPDgLdjO4XxRju00cmp8g33UVFg+i95EYXUxNzmlIikasnyJ/hE
mVI1B8wff1pD075VoyXPHXBLOCla
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
Lxig0oNpB3AIlaC1elINsSsErR9JGjREnrfKhZfiG7UW8dFBBMBMraegtd1lyUI8
DqMZgJdWJk2vuKkmD7XCu0A07TQq6IdoupMDmL7h9uABLqjOeb3dSl+V371yn8tF
K6b4gm4DBTDkFpkMdM7b9i/WjrvAD0tZ5ysfpSXZeE4=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 48640 )
`pragma protect data_block
JeHYop5afdptIZH+47W0t7BrLGcuF4cjTtYrZqm3Ky6W0P97KGeY4v4zvoWaPRNx
zB2bCdkLg7qu1mt7/egm+FKAE28rEJQkPBJTgm/1p8DLX49yd3w4QHmnJtQHDyr2
p/ALPU+/b05gTcIAAzazGjpCr7F1hKPnbM110sbw7N6iygxx1YYC4l5HmNIvQimg
8Gb+Er/0Y7hV43s/A92PiuYRPC/rx9+/S1idfllvQxp9+9GbChbi3AtCU70/9IT6
pSd4i8/gqv9QbQ6kkFAfJ8vmfg/XNNSAMoOvXiLtbTRsWs2AX9b88HerPFqTOn5v
XKpWwv5LauT6QJwjXHUqmd0owisR18OrIsP/EmWHZncrv0T+klz6Fx+hKHs7av0V
Eo2cHHLGwbZDw19j5+ZwyHpv3kqhab4EZhPPk8isi8nHnC+mw5r68kWcbZ8ocUqG
lqBykOQslOmBw5wko2xLIPNosBXvQ4ERFZ3nZ3uVwednif50c4LUAL9bRQnpEOHE
ENrwhMZ6Ql9kBS6ciuIhYX0cWsipJCpKzK6b1n3BY/wPJFAfrXDdwuLrxUSm7juz
68phYx4b5GZd4kcwX3UNbmUqzn4cL0FnTCOPIwaix79RfEg5l8WIEy7g+moSQqJP
R2PwfSiaF/eoeANTIVSRzeafDau/WojVHJzWwbZK3pEb2w9bbgNYaOU8L0pNMqyk
tLUAiN4UN/omdA4GsnHv8N7m/rYVvub9zq35805qo6HCSxfBUXXvgar1xC5pOAlc
OwquQC7nusUJVtubW8uC04tDPks/H1rcxsxeYSR8pkEnKqWCh70lkX+MgrqGGqo/
av3soHFsrvAulw7a5sTuXmZeYOAhPYd7jrRaXOrkSOqjPNKfeaJnd2q9YiCZ6u3o
jytmY3gHDoPSlrZd3CCYNDWDJQ594bifAqkNyimKV/4CNcN8DHoCmzyv0gZJn9yz
1bD9/6JRjaHW8ihNfvTDYoZJBtG+iNuL7IMOy+OXmNqh9TP6lQTx2G9L+gT/bvq0
H9g6wG9ga6w88hzj3E5ahsSP+ck2WI4gLt0VKBGpnhFMvuz/+CxVKuFkhPhPua6x
iWnEzeRgUIe2Xh7KTeyHTdrehAqipFM2p92mYlR/N76Og0czpOn3hdLUEkmr3YZJ
ZAuqPthUxp+7uelFm4BrqD7yblIZW/4agx2Xo6+D8wFos3HQFYzxYYMbBbDAPRdB
pLN8pcgUCx1T4G8VTSV0w7zKkG99CWLZFEA8H8LhcnaKaHNgVXGCwnWEbk2J2wIA
T4dWaKrd+L0bDxSeclABBwOAVOpd7N8QOALm6ej9StCkvf/eW/UB8/Ib5IQAtPOJ
0aBfSOG/eSLX5CT5Yxyj4mNi2fzUV5ajqWPG/H50ARqck6xWRgY66tSrwLphkGDy
tNS/fWJJht5CkmSYSzIdYSTmacmGEQ3vA8H1CqVaDN3I9JIYFXSvGyfneujObNj4
FfzoLi+h5HNV9d5LY8app8T93UaLWfQi+dCTeYA3T0fPG3ZQVY3WbITSv3sDNI3+
79hvJICZOVh6j2oqhklMfGqFgpBRklV1/1W3boxqOwOqqdFm+8M/RzEVUdx0O7Y8
QXmlPGElEMZueAnTzhPYzP8Efwy1ioXCwDqQ7RvxlSkiYtilsN7TB9GbcZKMA5m+
rPH9Vyul111J8TBzfU0Hd+jE5eAY9/OjXqQCzAv9osOMfxiLA8oyjtdpeIVc9jGj
R7gTK42OKCF21JDpOsfrnczxrGI/4AKixpkYswh2hYCEcL10bq74M1donUmcbdQX
8bnFgPIiH70KwbjozXcbIbVOFlP4ymHilVVlXk7QpqcigouJ0p4gG/mRPAEQ0nB5
WrRALxwb/q6GHMtAIIM3DR5Ls4iIktXqjsUzfh5yVKwSSF/nw/wWc5DQms5Xl0u0
4t02a994mtaCSfgTEpvbpn3DkSVpoQ2XaRwz8zfk47vGN35DujhaLQ44jyjWEWBQ
WsX97XFLirmZf6JSUIelyvcpgq3OQamXGO5t4nDuvg3HUxrjH/eM+m4wOeimi3kP
77FGWUid6pCinn5n9L9qCyU+jege60cPbYJvhUUMG5gX4V4+ylKicZflryC+wnef
kMD5NZ2yU4S6QyHfr0G/nOEeYv56kb3iKtB5AhiHYMXZaSoYbORnf5t94tLS95V2
KzMZqrCioOlfwV4D/zYJ3CYFnKZMKQTWbd7VACGwXwvro6WMQ96L0W4XI6l0vbhc
ddHKZxBg/ThMQ9Tt1TvhKiZyH1Hb5nJA1b0qfedQcUq6zemnMwyGGTBlmh+4lRRl
QFOuLi8A1Bp7JKaWJcbCiUOaXrK6O8xLtb7Qm+Kfc977TqQOW2M+yRXw50TAVU2j
VauzELNuQTHQH0nHKJk7EJs29IAR3fT70v9zQexp/moSy6B3n1mTkNsl5dTLSKMF
uBLrLLPeF/8XHPXhC5y+HklMvothQhVyzfZPjOXlhP2nNbi6/gt7gTmxKMCbzgJK
940VmSx19KGV/l2ICF8fV9BE2wPDWkNJgKmFx4QvxdtahBRZE65god2iNCUJ/tsV
8Nuu/jHvnUl7V43REj0IL/zlc/Cm99+V1NkpmrOwlgZVzoZ7tblajvfXuWPpD+pv
2dA9xbBmbYcblyrzwDd5NzretttCdtGQUSLdwlvWJKled3SAt/n2+if2/WdQbhiX
vdO+zhIbzlYIcWv0afxEQ1AksrcEVoCuFquxPqMQ/3Re3xYePfwEIiNAF1XWd1fs
J1fDwB8nqVpDLj0p8I5LkIQA3yGVQO+V/DRGnI6Q69RteXvfdDY0InsIowbOuYO5
mCoAFFdeqqRTRdnj+XvzFIpzssk9h2eBlJD1rQMNL2WNQUS0oJniJRoKrr58/VEe
Q0IE3/twYPCWwu21NSTH8IN8+Hc600JJSoPLtaMz1K4ycj8TwfJyGyPSJgQ2ndcB
yrojpgZhjRvI5SbvDsSxHwvELg0L/+8CvD3TFUeuVS0VT0MEDVi/Ify8YLreLuBi
AqawLuIN6NzeiS/lnKQzLcpfzWwi7nx5cNZlh+9KqzZgM+VNbHDBG1uWyOfh1SUR
ZjUziWye96Bnr9zqb6ni4YNd3q4BQWtRS0isfazwUy9rQZ76qnrGYmZ5IWjiypbX
EH+D+jLBvyx+YYV4S+JpEQjTvUaAZieeQX4hPG9VV4R5VZvU+gXw+rDZf5nYZrvu
xgPueQQDdDf2Xops6Ktayatio3TLMuTS8+QnMOz3wARt1iOyWLSezrIO9iW4cWYb
TBPnX8Y6vpN1EOfDX7KDAt1FH9vTfAXeOdxM4Za9JAvjacv1rf5JaVFrZbhLAUpj
SOIfIPHptJuPcI57peDYLo5JyGkUDfdqm2nnKCgQv5Xk3cSHz8Oj8RNcrqtsnBpj
vbJ8fIulDsQOGYy8TAGoeTqS1PxWDDwkLzI0uvl0nux1lMTBhB+TnRGSgyT6Zm/o
x2yYbIA/67uAjYuGvgG9NDmDl37M2BUXsBj+6WnwK7z2k2EtA6dqWpdawDIeU5d1
wMN9l8QVLLtjwG0ItBmM4aiWcBn6YotpmfFVuHQfxGX25pm3on4/OAB/KaM6TU1Z
1kPeBdHFV9rM98M1kCXGt1y2+mTE7SmMywb9Su39D1lVZRWurrgrcJjDiw3ddfFG
s7NDe2hxyLHCjSlF3N27V2VFxYmtZ/oYUlYjApuu7KL3JMws90fifZhzZkfmRRyD
dqNMTE3JlPhsCGd1TOJxh3MvUpc4C2IAIlXFCUnDUmUtvIZUT2wMBwvdCZbslfm1
am5japO7xtNduvdbl62Q66oAHRowT5y39SNqtHhx0ybk6ZWroVYI0ybfGR9FD3KV
veRMt3eff+8OahFy8lAsFCYKh8efLNq9YNIhvbVQPyCRH8qrEfz/y5M8d8TRqJtx
3FdZN7jBl3tlKtxTb7/c3H0a784ws2kk/9PL1JxXgiwKzAB0YhI9mHIJ9IhqIQof
Rf5xa1nr0N+UmvVSSJ6QO1X72oDxvS19GC+3QB+WwBpxX8Ahn2swTZGKuTPOdf3/
0ZmGTmrxxC24X1mANDdJJsKzIUjkMhzBt2J/1HDnbg0XBmif0Nzlq/rQfeA1s1ei
0iMHQnEF5BysD9SILLvbCnZCj4DyoZ+Zzgrh4bFUoEb9DtIls8DdmCdngjXcWXM3
jI3l9xAggIijbIYFsE6Bg6kTwXzs6Fc1C0TjNlq6g373WL8i/s3nwg87TuIMLjax
OPjd1txBSJacabbM1SaCTm/I+ipDaiJlhkSiaLO6I79+QoqgJnl/GBeiElhA+TrC
bXc3GBRosPakHE0uPAuwBo389NVeGKxNIkBnhr9ZPpMV5K58m2d6Os0xclaGOyJd
dYk2dDDT+01db42l9t0JhLgiRRAlnzFgwgaRU8Y6TL8xnkT6jVCdKg//oNjKkbCf
vzgg+cy7XzS4EUElk0krxsLetMQMtxq+BxTIjSTfIcqyoq5WqgF+s6IR/yvVzSxI
O7NIJpSyTAYXD1TBX3MppjXYBOtv6aZpqdYtTY549X0CtYi3crxoz390ghq6ZXRU
w2Jci5qqxreg8NM1W+y65OHoIjpS7u4Rcw3eHGRfgkBnfoQQRr4GL7j3PH4jnJKY
aA/yYbpeR46wbYrbA1XrESSNcAHexYYWY6h7VYfyME/UncKx49ntHVpBdRLxyLr2
DOXecA5vhRKOZnNhtMQrg3c41Adn19CmtfUrnE44WzaUi0yzY0S0hpMOeH+RJ6zc
CfE3OBTAIPSKY/PQYUdHqQvkWg377/77T7ArECf4pLSPrvKu40QkwoxQBkN8HfAO
K7j/jhmQqOb3GmbGvWWNdCpoE6ML6mYIhzy0EaRiXK7DR+zf15p50XiI5/pk4j0+
9tY5a+lZdrrBckOpVECF1B7q4Yv9yCIKRjCGa3nTCXFebp69wuKPQxg1kBKuuCKT
InrCoJo+Jjxth3P3hV+M7CbY0Dkoo9b4L0dDq2+6pRyysP+XQLDbQ1ReO4yR82cd
TnOu2Xmo3nxGz5y2Xzu2u5EQsjEt1ZvZF+rdR5831mxED4fjuB2IXqodZzCxJmcR
8UkQvL84Q/TWYKyqkWeLo3YuUa/v71zoarmOJWNakXTV2ZpfNxE5o0uynGzSCipD
aOzFvoRJDq2p6wcK3GupxBYAVPlC+NJdYVFSE2H8MsPCxiehc2FAp7046nozi/kC
OuROe7qHmJtQjZ2e6enMI95UMVC7Eyn5JZ2Ja/JkHIhxIdgCN2DhRavBInj35k5i
pzQ64qn0/9Ken/pv2vMwSTYmwiFepz4UR+AhacLlEk47h9Vngv+DGSq9HLWWy2Ue
NOKc+ELKJPzhmWEZ7i0K0pzJabLtEWvtj/e7mS6jAmWeQ8B4/8dW3gcLqMxIRKhP
cks+zYeoE3UWLVmHtyoWClksqjO45dJInjyMviG7yk+ikOP2lr8/t9CxMboHtqib
eHmUiUCdIEviRQ3q3Yn9hDZxMmXLKhsngVcwRRNDh9EjidFMy6Twm5sg92x2T79d
k8dt8tTg0UR8DsoYaFe+ovGMy5geZoCY0/6JHr2ENcp+SswZtMwl12l2giE94OKc
epMWq3av49AR8UvTFdzJ69fV6LeclFVs1bxlaoP8WbyJsvSB1jbxzjrZ9gD1fT9s
oe/KCWEvij1p6Sf5mIAVfWjVVKXMRHfu8Jb38xqiWwslQK1C5fLpr4QZ0hbQS+ZM
olouNQlYp6dwsJ8+jKVEa5bMTMYtw/XNzVNyMOqxXyJWVCeyN2jzxT7Y2dvOGqSn
lqPDNE8Pjqwro52ViedB5rFqfsVGyCFg6oRA4Lv6nvv1oAeCYD+DdJhve8MLAj0Q
EiYwZpUV0xLVocfdrVPxJSEpjl7lRcc9gaz+PD3ZxVmPDspGtcNzO7qYXHDSTIVI
pwGd17+2mok+s9xFWU0mFU11d8ai5hz4PrrY+ReoTKqdRLvTwogqqDnQmTEEKwVw
NkXmDbXtpL2V2qgHAveF60f3w2UXJ1RwZxT7SGPeS9HEwkS3HTrzLYDN/XO+4/Yg
r2atv68a5w0V2BgyDkCiEZ+aIa14enYVyg4nB1M6wM4iYpoDO2rLOh3DRDIif7cn
+tOhdPJuFXIhvHcOLQHhqGUs+Ik688RgzTc2F/dx7IC1LEH6i3g0w5SQFH+EC/2+
0xO/ANh/tWCwcvOfMlSnJgIpQ3s+zI0PxIiXhj35scQHnyTGjoSmrMasf2wPLCCP
T7VWASYBArknf1N2dFE7Iq2FTzBNsDeWm64/+zniyhwc8gGrI7xpOa9caou5fWW0
PJ6nNUDIyhC0ppNaXP7Z0w30U9NbE7ghfxhaxhRqiKm1dypVA5++efvMn8vw2SWd
/KyoP/MBkNMZsmJDXYLDBZmoiUmUhy0Y6Kzv0ZkWn+i6yuIB7NmVss63xZdw/enN
wDzhcO/P6Psv/qfFjpRtoBSjfVPcM8nFK7myY6eSyV8jy/1eoP7uQhVAMXjckwFq
3TpWGYvR9u7aPAaRi3ot36fZxCf/dt+FZlvac+yGqFvtAeA47gnPLVnuXDzMMr7q
1CEYI6mL1ckg6FLbeMcyph6aR4WwptdqXFEnIfNMSswmA81IPbSy2TpE6lkGF4zW
hXE9MtG2HfaCN/4ZwZtYRosDy3tLD0grPzZABIJRpImmCRrzgnrqsjfAwHkemj7c
voOxGXH82Jqu0pKxKtqvuSy7NF2JtRL57Qik/amAySJVwzN6Y914+Pl1JtH7fiHJ
BM7RVCXM3+86JT+53FFkTb/+2usGs1hAQ0ZrTzoPKbS0hwY3vEh9UEolKnxPeqTO
KaSoTauFTirk4yUeF2majqS1BkFj9IUNrkvvOWb6WXDClYFoaRj6D3m5D9Y76XY8
RACwfznFDB66x+zOgdZM51yFFvaSjE37idXQN3gopkXXfdpBlZiHQweyvFoMc6oi
DY+HS4dUTfzGK6FgkOtrlXXCb5HuL/sHUXTtArvjdr2k2h+ZBPY2o7EJ4sos52va
OFUK70FpdYcu1JERKGeJRZYM3GQoe3uYr9zyLAmZcl6ww2XWJQONW/v/cp90yqKf
OkVoZx02Jqfwx19oU1FTFzyrp20mjxrlcevPht+20/fM9ozeNUj1O1xsUILF0GNS
WZ4bMQ6Xg/bdkUs+PnzzL9v2xqsnk8NBB9DILl3Vx+lQnR8CyTSDwOJ399UY0im6
yd99Sb36QcQgKX4RghMd+2+QKqPj4w0WsoQAc2aWXHCUPcoE1Q4LJ6iX6B2m+QgI
FrzSLDEW0D11vEtKre0G+mUWjaf3WPcPZT/dZtsGgbvlEdJ9bQHSS5O/CMS+CWKu
P3ZSfnQTLvchV2tg3J6oyRueuvOpaSZqxUrsdeLfx6t8CeXYO1S4JIqssQQM5PtI
O++SdYq8ov3UJb7YlgegyWlrX4Kspeg7ofT9t5bO3FFqtgm/QNVwqUtq3X5H+FUW
M7Q3bWuT+6in7lTwFoSrIK/xyuPk6Z7RgO3PPmvVAUrc/T/lS8bhsDxwqCXq5T6B
dkwmUGn3qy6KLag7qzvUjhZcud9SEkXg1Uqn1IQUt+wRpXA5Y5YBTZVdepAO6x0Z
dbVWOmisDq95xzF48ok7JLlUEUViTofeBq1eftE7wf5WInMYcSrM7XIrDKX4waLf
YlUXWHuZaDEk5874wTNYGobb/2/gWvW76q4IGju0EDlu1pFJFMP51wx18kU9q79F
eXUIrUXgi+YtRh3EzudPbBfCF+0HJ7S1dfwrLqIBadDxxHFL/b44qkkuuRtHVo5+
77ACDbJw0BEx4ro8MTCGeHfxJ+t6PsTPpv5DFXBxfBK4JDWxsbUHblzeSRgh6jjz
7oJSvEwQ8hJVBtiYVFuaQZD2oXxI6Xq/Atwek6SXrvZHrp3HoBJU3we/VgsS7fjQ
COk/F6D8u/3WSGNzCWspVX1czBLl1yjoVYu6kFsSXRu020dJr12/NqtjrQASMzVz
/JBxHhAP4l9t63ZELc73dXNd192g6c7nuhApnFwV5X/JTuspqio+4PG1sRIkexHZ
rRmIA7oRyQE2QF88k005gRZkRd7Kin+NSOFh/uDKFPKs0HEAMJIjQH52t5rnfVKY
1Se+PK0Vaqy20Vx7j3wi6gfqVIid/fQ7PMJXMGpn7mWOiPtDZDxRV3ioXSPpTFcR
3jQKAydcHyH4kaaxKxCJZBeK/jp581wmnkxbrV0wHavllEBVERsqtk1U232wsnhJ
EMqb7TajFbDntVNI1qDbDzCYwdGtJbr1EB3OY8kzX3iUMaHDBcLMEXg80phJoWi6
ypsnDnkJNXcI01Zr5cZWdmU0MLDrhL9tPsqSpHY5csKJ9sKsyZp3bhnLTGvUFWku
iyiyOuRRGdZ0ahi6aLYtFLRtubjeD4ZGNuR19gFHr2pkr0rqKOXATpWKrIlCnzy7
6t5JeZ/xltaQgfkmQv5XI1vvc1stOsrb6tkZXl7lJqzyLsD9mfG5UfrFmzoysYI1
2TMtdRLhHtkb1ucsOKQCelHsHFhvHVOwdmZctLhg/RgLbBMmnDFYsYfRUS3ScNij
9rAqYsU0yxnnyzS7lxJ5koIfMVJEFT7mix/PXF02/+rOZfaWssEiYmTDgDfMaSA2
YOfNPKHvrcHpZLqT7YmAs3lJ8QgsygmYLke8kKhnpefTJPayNECHetaquUbTOqJj
3t+ez/UUtH14CSckmX1gEO9VMrIIOsXAouGlYYgnSYvt1n3yqOScYaZEZp/EqCSC
ZxzYTyi8+rAVWW2EPBV+2Q9eY4/6RUl2X9QxIN9aj4SmAJJpTN2RMYqPqH1X5raY
GPAnrGxQxhJL66cuaHybC0Wa+ymhZV5KkjDXOKBX+5fGD4p6m23QULOeJu30Cw0e
gcWVbwyWj5pAKL9yFlQF9l9i7IUsUHeShMyeOtlPAe+NIym56rbaF5AmCrm6iFc4
y0pGmtGK6CUKCv989muuV8P3wtibk+QleN/8kK/jB1bq85n6uKJ+X13ON1m11Xh9
qQKYyf/Tufg7p30BnmQWOaqu/T1FbfqP3BTu/DQj70tgzpmWzu00+SM4VgOLEREI
/JoeS2ci2Xw+zHOBPv14bJSr1RDkcsoGhKzPCgOoxy159C8XkutMIhNcHTtpQX4W
6/3Gs17D+FSRYrreI+S7Ih/41e1YPY9on2RFnKNyiI0VA1W0v1UlAGx0r+QK3g6e
N0rkG/qXrrY9IrpGbotMnJq104BUhXVYTAzQsk02NcaWmRu07pBveIBplmK8en81
mWps42RSDrtg8pqa5S8RBqbTNS05MmF/YUVHOljxozGbJ0LM+VRB0c0+SEHribAP
BhpHl4c5yLSXrzQGrwQ1uVDkXua8GC3bP55h3VofYPa72q81G5CNsiH0+WvZ7LEU
nlHJvATo9ExyTGGaAleHnLkY31kz6dlle2hy67aZWUqHDZgE+obXp16TzDfe5g4O
j8f6y8/VDRb17ss2Lru6CMy9VZ1bx9NlxsoXXuOOFh0BpGWWiiM/OpKrXOVXn7n7
YdiWpEekrt1bkc6u+7JGJCtYTXgj3FArupmrcpQopdU2BdxFRRNeYytjkJd3B58x
9ASErjvZgADP2SMN/5kY2GwAyb5SyEFg9UxDZ7lpUCH+Tmy8ULurB6yAXfpfJSXf
YXPvOqq08xdN8vqvDWIDPBwIOZ+ussc2tAc3xleKnwR9PoEjm541kiFwTvcEUwv3
9j6AaQnuackkC2GV0Jcyt8v8FQ+4sPqyuOw6AZmDfWblyPQZvwEHjAttdBGy3Ysd
hV1AJT9AAxXij9GKnNU0zkuEMXWOARmF/7NfrwBRu0GKkG+skM0D+alT/FB1Cyws
/yqHgu21DQ0NhqsvlgdA/zP6OZfq/CHEzYSdZloPF4YbPvo1V3UAT8+tc9ZVSaLM
f30vTjiS8p2iVkDjwH8TTGM8nG5b782TjHc2+F6Ttz8jW8IbZN1MWrKjDtWebP7e
bsixpd3wQjGzguEkQIPlQX1gAUQ9BladPE0aX/I9pvc5XiO/+t6mHEOO0zTvpvF6
BHp7W/y/DBo0FcJftDVW8Qmep80smWfMTxl58b80WpDi+pa5YLKqKV1ML1nt9ftl
JFVG/l2XUx/fymETAzCMt47E4wKsbOz92IrIUPr8JNPCLeP7dY+JxKKoHv73Gke/
4CnkIyalA1l+xrvssmR6tN0MbyJmHLJHLMja3oyRsBGC1J3e3poY6CfbjuaIgBup
TpsZ25Km6OHZpWmbepyXVOVuXodPqBPzN6XpaArOB7NArPOckGF513xEASCSDHVl
viQGcrTDhlq+burGokeb1ZzcOqJwIih1qaPlVft4cuTk0oFcMUjA9vawZaizJCuu
GthFhTttE5aLaZRWQqpeLK9cg4NqfBpDIBcWBqmYZwxfhNh4WF1it5wXfY9XXwPr
zkH+hWUW9IWcc9YcAfmOXQXB0YdX0AOOoGzvwLKwc2XabKYsKZDHt5nCWbf/AlHm
6OXflnt4ug3tIkkmqZGeo2WztIclwsvRAd70T4eKY7+LSeNnd/V3esrEC2adpXRz
TMjsPfwgEKGSrWUPc0SCJe8AqU86F+nl4GCuzzxJH1Uh9QmPULWgck4IPk7CWtJf
cTQ+Fu/jkhPAmvesggmZIAyQYDYXakHY7CXDjkUOKscPgUNdDMBCdDZkR1dZM0wD
nPZL+bYDAUpyXitALItzVK7UiKIXlYm/pwUSqTIqohOnVZM+mX4C3kqYqnZgxsRb
+7pMx6sZpiWrj2GcLXb+Hgh8vOhH8mtcdAaPtA82B7lNScGzefW2hJij6oClsSyN
2wNyCmBUaAsHdUWg0WC1F34f6ypq4F9zPz7qZR8YNZUaZywsh9q60DOMwRMyszvN
3XbstvsQQg/AIt4BumO5T5EEonXniCwFsZtoz22WVZkCczzkx8lWCL+kzUYh0w9E
OMtHZ7rvAK1WANEHTthMSb7XEzCW/ySj64YT/abBygH5p+QHTzFlOWnhngg+g8ka
wPGkGAGqsUrZcvEHO6REiWi50QudN30rbCOanHFNPBRBePH5ZaQSL4ivKFem89/r
duBLU7hmQ/prCg1LVtGA6wr6gTgL3s7U2lQexB6EWcpMJsEnLeG+iNG0rOD2JLOM
acCBvvic0ORtCPH4ekkvR7PbXKLz/gUrQCF4JwQqYn6qCtUibLsHfghOFpue6FH9
z2GdFalAYeMc3SOlbPGG6Htr1k0Kr828a1fewCPrwRyIdpj5zDayQNjCJZJqjg/Q
ANiydDwoSKR/XQiQNBp9aUMJek/0CL5R9D7Aebgt0b7I6r6LPJHegHO9LthZmYIV
Dwo3ry15LuPlTO4dSwkiGTj1SHXFf50pqwxJWkU4hKxvRmDFJdtgaffCdA2fUnKb
PIV6kRd1fRZFBpUQNcLOuwr7qYf7BLe5sp7seQ+3bLDk3bqXWwec1h3N6SIZjXBY
NyUWs/lG5KcGyJkD2lfzg/MGkHJ4RwUGQaJRHKO44Q6n/8omN4ZfsPc8fni0ih/j
iaEtaptWvlZKJ7jL25bFxyXpICQdu9XTAwHm/XowNSdBofgj+8nY00W7tx/9BKrf
q/kc+sAwCJgkOU0xK49A7W7nNirKjL/Phb0kjHqO8volcOQNF3VuNKIYFxWwnB92
8NROjfB4xlYKUhbTG3py+w5fasZqk38eSdAyMDUxJdvtmKMAIMe2aPa2Nahek5Od
2+wN10vbN+00o59tL+V+R0+yIxmV4yvfnOkJDoy4z5Zt8LnK5AqfDO4GeV/g950s
VtOHCJt1R0seldhDMA2mMuWMjOvBxjZRebeD1GaWcojeoDJ0v6XOFux97jgF0Xp2
QTX/qTcTW2E7grkKyO04zNrlZZ8x1WwWR0fRa8byAyN4QB1UdEncuzaoDPRq4CZy
rJMBk63yRYql3jO7bPx9VDOW6AAHoLvY5rfy4Mae6yyFhCHX2gndcLi/SHvpBF70
Z2zd6qEtOH2LCvUfEAl1eH56ONQp3YfWBc07IAUokuDf0gP+W55Cz+tslfYYeJJQ
MfBSaWj9Qtw1YA6mggOniikTCYRjL2wne5LmUCdcwiFSApS+/9WwrfHy0C2V7IB3
1ghYH8Um+t6p1/ZMiDBwz2G2H9nA3/2fR1f7tRzhnVLrbqk0q36q8aEVAxkBFINf
0fzjFiD8LMDB1sdSgiOnVXLkYu83oFDdaogzDH8BheNoi4HiqA7+gAVwKwe3Xz9V
7X7EUqQK0kp+3isCTrp2j5PWpsJVB4LtxxKGEOcbA6jGy75vHy9l7edGkJ5BqpZg
lBKCsCFcv+0+7To9AtTZXhptuhl9UEZLppFPQ5XKcR95yEEXRZPmudnbqJ744+I3
uflUN+zTWuYzmJ2rWBsvnDkOGVHs6jMHrnua8dm+Q1g8rjvlBJFDke/acW+gySAS
OFzP+hivtx9NdQUF7HhzdYIbL1hfwrHTokE2rpNjqPsdDI3w8pJ5TdFPuZ6jCG2x
XoFVN68LJjSjSu8Gu9OVVjFYlieL9wJkmpXQe9QbhRMQJ1aN/R0hvh6qi+LZtpp6
HIkc2R1a70fRIvzu/WafjvZ3+H2xmnWeYmjLW0d0taEe/b2LEimzutQhRH7t8REF
cDqfAGpBVwD6D08MLUiBJzZYsysiLx22cEksWX6bgHoG7nBdMzoaIPrVY5OffjgC
SXuV4CG1Ls+iE8hwRhpbhcMzcpiJGXYkEsAg3xz1A2J+4cPgZrPV8ea5x8TiDAtg
+xPjpMyyrYa0oYz7MCisgYTLv2fIrsHkKgNCm0I7qRtT9CJynTSo/+tpAIjptQLJ
2IWH8r/Hnat73jkHf0T2kf7mO6XFTiLfP/VNaTea0X8+YYlW19g5OTDNaVGEmFEG
8Qy4dYRISXRtQ5K/FxPC4rwdu4DIF/iWq5jSSPVYRS662YNU0sgm1TL/WUR1gjl9
/SrG5zEVp/6Z0KtfKy+3+gsstSIK3KqEMBsC8rolxGMDrrkXsvx5GCTuipcZoU53
d4HTSGLTpkVakS7vcpwtHJj6wldZ6gsO5LgYg8Mag+0GuOmadP0BP9OCR/VA0yeZ
b3n4Z0F31wVEtSr36ZguWr37TFzGj/7Rze+IyVnj2fUIaCT5bkmFPsnKuk6cWhd2
Qbd1RhwLyALPoiHgDNVS2yQrYKCW6I2xxFzTe+qCkmCbE71LMaw9R4y3DjKyH9Xl
QngMVEgMB45LHN8n9ITyjH4WQPg4xZDalrsIG/3ECIcbtpWA1qQmgdAHap8CiaVk
BxEzRfBZC242FZJ0uqEP8sE4GqsKtjErlBkxi3Fo/UXaUDUjq3zc6cC/sBxRZmRw
CKKVcqVLetBzZYMNuMNaNTNReU8cG9hpMGj7QGahdkUQ+d3IYns2iZNmYeXXTppc
av/GCoH0HfzQCDX2mjr1npVYh5djbsuycZzH2Ml9psCyEr+5cXCu34MCbh3W7Qq9
Sq5IIDED7/VfTFoP6Wf4B12vhILS4lXkXRHMMCnrTs/+FLN57nAWVGiWr3sIWxFY
C89pBwri1Vqjqja6i2T2mMaDHjcf6d8bTEnR+bSccXFuKXwKp9vqgRa7sPNeo7d3
1S+JIyBPbTJl4gmoEpEH2GP/ZEbN3a58leDT9g3BStUUF+IRj7iKE/y+JKN+omxc
7UqRQ9t3H0dgNvIDwrqf8iVQhkNUEJmvB3q6CQKQXFcRitQDUVxwgNnhvOra1uYz
8NuWV+0WK7uiqbP05k57Q5XKbQgrOxm+Zu6cOb6c881EcvyxpUD8rHL4RYEFU9wv
FJsfGxwzR5z2qdV3Jg5RaSe620KNjv8bblVO7d1UIbjg+vNlWcIn/DPmjqvyz2wM
rZ5+P1PTkjmUaEZeYO7ebUE+k9i0mqbd+la10xzS/Z41mpFM/FolBtYvHMm/5DUz
A8/otyOwPctMEsoI6zzjtcgL7W0IsrrpHAbxHaLovLDlzTB8N4FFis4CjXge5OfE
L0NO6LUW76szaPkXCOZgaaEZ2j89X6WU1TICDg+Ie27yZnmqx+4j31AyqpVTQSZC
sTN3e0Ch86GnvqxxEavWf8jl/grFsUY9xaN+/uzFxitA/CwYquzdrHE72BG1ggJh
OVupdbeI4C1vTuXFH7X22CQpPJAMeOJ9cFHVIpjVLn+25l1+00InOe6qo+732zAM
Z26jgxa7D5G1vOKBdTO/iC1iOzcBSE67V8n6noDngsa6k++JT4dK7CVOqp8JZTGH
CTwcI0h/49vL2s/VfHfljJ8sPtKz9lKgbRTG9NY4h+nvg6Q8aeJjG6A3+ae56gs6
/Y/3oteO0K++bliDoWfed8cMYkUpKoGCSG4drAE5ntf9wHHBIPMT3V6OhktnfNBJ
EVYaczlGBAu+EbdGCQxmnN9SU/jRzWfL972mPzqRzLdSFAQsrg+vNpXUyCaoKTPQ
qhmwBUj8NWujnE4aINKazhvthAs8S2JzNy5CNFKNjO5gV2yNqh46jfggJzX+WLSo
rrK+Dy1v1F10cvk4EXIV3fpSxJa3bAifzIvebX5Z1VxREWfJTA0Ivh2S3fd3dHi7
BFsg19ss5Dm/WuzmnwNYnxGv5LCGwLh7oR6YANML2kWUDTalxu3KiB4YclNH5H8L
VVZuZ+0N/4L+b+KFsz/TgYkoqDx/sYRriyNj6DoUZE7HJPrelJIQ/e6CpOqSPjJG
fqhZGhbNOQX2ayT9WFAybvpMQfD4B4vVxBlG7S8+jIPjXh49E4zdEC3Z2C3303U0
E2kNwX8jx5genNdWyo5Fn8cvkShw1uSqexxM9LzUZ4zbrONCPp0oO1q8W81Mb98f
/HkCLHcMTYW6zAXZdekeC0KJ4q6OuuCTKsXkfTWHqPuYp8o7n1zdhU4mQVPUNaTd
ZOWegsjxx1ZK6stJc3tupmEm/PRRadE4/ZqMM34QKjbr0felIAHwcbSaYToqFGJi
p3HaQvEyCrqYj3QMviuy/7WJY0u4v1akUUawel5K0BBnh1pZgJGLdqHXTp508j46
EkuslzgM+W3TQ4So9lSlgCdTXdRfBLWYmlJA2jvxH7GboE03SYWUSloRn4MSAm0y
tfd41jY+JstTG6ec6Pvs3DwfKPtMCbQeLdnqiaob9teI21udEj4J7alenBdstM5V
isXuzn2OYhyEVYS1S1SWogQ+0JNTM65yvHeV/yB/JVN+oWY/7v5Z+0cip3hogrbO
Ewn2/LBnuiIHYHNvkpR08RVUU9aY9km4ZXpIa5xAU1+CzokJwq8GU+vpA++Y0jwf
0605pvSMNYJpL5TOQ5ZhKAt4aUpt8HRkIdURYQGRR07dc/Eb6K5HHxzgNzzjk5So
Jozk1GDdzA15/m6oRidcS4VRAQUjL2eb2CpVXzs6Ue9xrlaa/x+YFX6EQwR8y1JQ
OzTdoU1e8Ca/UDBMuHu00758b8kjsmZm3JSdAAGyl1+yABjpu5QFYw44PrjYnGP0
feJWH1Z2qRZO4vX5D038Fh8SbOBD76sHMtjbxI/MMheDPOhALHNuis3F8lCSPkwe
zEtWCh24yO7IQ5I1Dr6zMIVVxoCKW+I91blxLzxAxSD3U8ThJwh8xDbECTJ4aY15
PGtLTRLefPN3YfaHpbAz/lm+31O7bxWgx25Mrrixn2qk7BZI5RRVTEi5oRVzUBDu
ifidN1z0gZe6hdbe2Kt78mKUZIBkxwpUB8F5HSTCyTObX2PfXIgv9xkq5BImzK03
2EjHlJuc0+j9aFvK2q20nUSpdnrG364wBwYLHHtw80mKx7Xe6FQ5nxzZpr9Iq6p2
F17n5N1kDBlkj76sgNfZoJS22rklDC20OZd09wjQpbHdfCzPJv9Q4D0pbDq7Ttsz
vVwNenNbi3SWcwosq4KcJDg1rBzkGHSPd0YQkFSzruhbN0P9vMcsgYWQ38ySuFKu
HNF5pRTsJGvAwDaUTA66OSicRahMXgaHuIpXJESCK5AYqOBN9h0bRUIG4T5467pW
QyXmyCZz5e4ZW8uwhuOrtur1ftfvVsieSS804x6FMn9FaB2+lYzJytfg1nCgkfAa
IYKvSnOd4XZXR6LZRD+uNbMbIZzCGhacNrqA+RFviIRbude84aqtZwZzF6fsye5d
4Fze18EMxMGGE0ZQwsQ6OIbCdWCFF4+Jz8tTHuMPai9oznVSnhfdy7PG+DGgQkqU
ZRLjn5v/ZZbmBtVz3eiMPx159kqeevoU9akZEQx7iPDAv+6WWOfYs1rJ+ZLlK0bl
WLz+oruwr2CbNreBmrfddeJhLuvmYmDb7MVw/voklgGT4vPjMvV380EUgB69nBks
g2rgyI6q/5xsT3tYP/A3KUoPAvzZKWxJR4Eu4xADXc4CNEcZ2x/ojTp/5d6kb7AT
PPhzwfRCLjsq7I6/aOYTFwZ1S/jp6/aSWkS/N+O9DVyzIaRkSwlTP2oRt+zN3WqG
mXAJNSA08UO8+vfQr0CnRKrqehfl3mhAjkbCAjkIotG7xDuE+0+j2m5yAsXWX0aJ
5B7eblWt7YJns3zqPQK8Kn0wQ9kthdwNOfAPHKwUTE5xyZDDBomppyMLDAFpiAXW
ObcietCcu2ETVqqeqBz/PzqS4M2lM9q02bV8brClUfllpinLuIT2i+YXQsyjhKgE
29ew2md987xMemgjzoBwqgvY2dWTG6oIC2yblfns9ugEYPsDB5LdrSqH4qHZhbDh
aU/vyzVmg940LuMvPH0TAeoAsuNpvVOOdElhi3yYNj+oB3Crkdn1+5oOyiKelh61
ZpDvUZv+X4KR9vbbV+rQUFPRxOSGuPc1aHkiGaJi/n0GQjNFt6Ho2Y7NtuHTh7CT
w7OicjSvNa4uE7liB9wOTJ53cdWEl6rfmOW7w4kH+wbYya9zLrLq4zo+sYYddARa
zrQCy2WbGb1cruWRXu2sIS2hg4tGvDSM4NvYQs/rb1BxEjCBDYb2Kyi8CLcZ77iK
P8KG/kc85F1F5j+nrFSuM9xB9JM/Be0c1x0q+8UURLl6i1GDMQyjpJe3lLrdW3zM
BCfhP8OIE733LFOZAsScSBuRC9EsQZMdlh2mynR/3x55V5AGTwHNfnS0IumMuzX2
jqyAkF2Fppj8wrjjgNM4A+o0XxA0o7IQ6CiLvK1wWJ4YTQbU4II+PfrVt3j6xZ2F
JdyPO7wGuC9z/qL+GdoTTR+3R1jMICWiiDs/fxAczXUrGtG+zHWwH7sTCndbjZ0P
Kwzz+NuityPtGII6MIOrBlhHoWpTUXpHEtKk/5066ECSqSVPnopAQuxt0PSe8veg
NXzGjvikmlFyJJuDvcq7rhMqOBCl+yvXVdEs34sWxAO/sAuMZK1X6sVmMPpnz3go
ZS3GN49Bh0nC9g5gnnx4VmlUaCamMtxoJocJxK6Nz46mKY5Fa8ob2Yvejkku0bDJ
qyuqBi4ZpKoinl4vH1lgDFl0peL82Z7LtaA5TceptS+1v4fzj5RX4+4QRq7YvAgo
UASuf19fk9IRFZZ+hvMil/KKsc2s1nWg8jxguEMoFoY+WV5rStSpWlsoXOdrfO61
rDkFYuhB0UEEsPIFPwrOI0tE2E10MLG9phrUVZMaUiddYRvf4wAlhHzptzXr/Klz
VzVIvvbT5cDCpS9fUuYjxTQuBQZ9l2x3UB1+M/EsGdQG9Hv62YYun7qQNIfWDGeL
FxrVQXle9Wc7Ttp9TGduHjre23+t3vX9ZMal3/+dnHf7Td+EFpOaQBU1jC30PwOy
49ojqdGUxVuxu4ZZ+3AbYuSWZJzHmikJxLU9HhER4R3nrxoE7kh3Qcu8VQDs5BoW
Rk8k+GLz1Ke1lxJvdu6IFti5lSQ/x1xtZORSCYQNNKDy6im+od36EP6IFvcGRTLB
Zq5m+lI6dVP6J0tRxDDTwve8XrwbLpTpcJoEsuhaqVrE7TLNlEjjVmmMemvs5t04
L5i+9g2djosY89H4SA+H8PbeRXonU2nXKQjeTdmxL6RmA2hiU6CLGFwF989hzcI1
7W2YkEWol4+9ZjEB/q+0YnnhV1kl819DWFTLpp5nKXmmV62G5Rpkyd9DzVlHsYGO
kIYVZEPCn7nrWRmg4YYAfSTmY6PVWaZEugdxT2pWoN8QAkMea8rp+5d9G34GJ/ji
UtO2qodKqUv2RyaJFECIOXFapiQGLaj4RgI6znLIJ7BrPEQ6ahxS7lCZbCcXBWN0
J8A/REvUrtluyJHQEpPjSfKZP6UOtiXzeiLeauNZ1VCFFVWgmTCVp4N/BkuKGwpC
VLhVHxK7jzrz7zi+r6z/VBoAzcbQdq/PUr4smI/ltRrCFZD0+0qd5BUzjlTMDE/9
41H0ciisyqF0/ZCN//6Sah+IRduA6g5kcia2VI8zAUV1XVTbcmUK33X5nKLAwB70
4OyYM6SEZrRAAp+2hWKEOhF6PUyY+gf1Zqt+d+KK1lBq3uhXqG2a0iGa1SEk/PgJ
aUn4/RKiPnv/slAAirTDrgFICZhWydzxl6Z2wcrvbnihgfnsGbViwcYdKmu9s96l
9hMMWC4PcuX5p96TUaSnb/FPz9mYVFpcdrL0Aljq3g9Dgewh2vAWPrbgmnmG4q2S
SYgc2PnFsnx7whwDT1si2MSgWqr3HGs49dfNN+XPElwOPs8jkepkrEl1BV3GUABU
z3f8ecZqTGZUiu5vLvlj0Q1nTIB1ImESh8XB7/t16fbEflAaby2gq7fQRa55bYd+
CkTNykEvr8JW/hy/3FS/kNrlFHVVf7vqim6xqdx2YSWyw9p9fY1Bb6TO4fam3LcE
8Swfd+ExFWvhmlLfgASL7hrBvf358gBIhy23rxtxrzDxOhc5hUpYAsxfUu5lTaX1
4ogkimgU4bbkVkjHX9isavquMfjfHG4viZLlKdQi85Wdse+vHRLiYyqQ1QhtlYvq
NHnjq0gRq4wxizhy6uPjXN5N97830aUrrAuMF7ZQMqvUP2Sx+iGox6AafAOWI1Rn
5fUELuSLFllm0BT8Pmhzv/0MhX/4LsEwyJCeqw7aOVA2ZEK3aipkblJLrMhYqwx/
+kzR9OIe0KIoc+58dyiBtE4Udq/E2PwMnYaFaIpleRVqzuVtrkUZT5ENCcDp306v
a/fmpmTZXqHVr7AT8166Hnv2iL82GmTKwUuqbICIQWuP7H9fUJ0OT2XJZCoR5GKV
byaphGWY2izcAoeIvPLd6ZofsWXV+fPRES+Xk/71oMX7RjJVszb4Lb9hGSSuI/FL
VZTS+cqYyMIC8V6xeuBkCpVRAQIQTKUhlAKd0u+3ZPqdzIsRaHrZPX3qOlCxHzzN
PbNdTqY1/jexP75aSil51jbpAcpH8o+wi+gJ0kCoHm+pEddWL3Rrrp8E0AWNAEcO
rqyu9MgaxiWx4aLaaAtuqomJHD/DBzW1Ehj9gQvPgAEg997wvKFEAkdGN3efi8nU
RBqjuSm3Fj2btwefp713umPmFi8IEt+B3YfF3GV3qt3kBf8vcVKgMeH5DJujbso2
zp3Zk49B6SzRO/Nw3EdsGWP/KqGTgNN7QhIOp9613uvVTqXYCQUg2sAjAFar29/r
FtrP6E4jkcLgyVAae0LqaMM/XVHjwyiMfnn16XyQOPCcvz2JzmxwvNLBH1GLgS/R
kaZRy8ONEcH7WKWEpDyufozQAyxeBR4nWqqvx9qKIqH4krbFbv3O+9yCK3FiY6TH
LDu8n/vdSy/lCOfrKv4MZyWLYK6tGMCzx74Ai28cooTP07IqAkWyX+qV8Sbiv9Ta
FdgtjZXHPpHPjG3gFXsJGXaTU6s1ouSFdYyEVCzcQ4Pp92SuCoCPbKp2mmTMn54V
qZgsLu+oq5CSj3OidcdWa+xY2nTuJOiFx4+XhT1njrpK6q3+qyS43zEcq8WU9TOe
kZf9NsW6Iqb2Jw6/m7V36Of9QM0vcV9k+vZO5KQIJkCULP39Wj3qdg4+FQ6OjkyN
9C7Al4bA3XuF2SovYt2jO6+1+XFSb597m59W1WRKWx1htZqgD+dm9tqwf+76U/BI
hRnM8oOJtmOcxCrbNp62mohbdsnuWDZ04Mbcf+alAIobJt7soMDWh0ObDCNwjRoS
7YTiAgUm9XkGlCGIrlatm5wpYHdoF5EmOhDW3S2IaNvo0R+65aXuPDO53dHxMRu/
QoYSKFpZqfA9FUMgHv5LnQ+WNWZiAAHzSZj2yRFXqJxz6mOP0r5ZvZcrmHlR/qx1
wZmlZiwI6pk6ND0at0MOR02Q7XK05t89NvGGwRdxdezIMTDGEDXehNmFJbyeMmOR
OkK2jT1UQ3DccPDUlxtbpwaUVfiK8hzckEjBTFFqosrFkGcZZqwG2XOM1OCCjuXo
k5w2IwVa5A8lP2vzAKm1rh3VTZHlXgwQj/PSRhc/6cHDM1VbYrghZCluBXZkdCEX
siOWU6iEoC3jHikJkacNkKnrk5HD7tonnM6h4/et2Y0tBcHVfc1TGQC8Hv8liens
VP98TFJVVdvyIF3AwGD8x82uM+qH2Bl9qiYy7LbkytI5zaNVfMNVrQbashpfIYQ5
MCtWBHfvy4FMv5NXEnSA2q86Rk9DtQgnpiCUicRHCbWALEldHcClwXCyFs8n9yIr
xc+lc+P4K1O8D2qVAZnYdcDc8zIguK1hr9r7it3sOUM9ODhw8gJDMA/E8VJToQWz
nWGJDn4LTmNwxcFnXUoF6470xZfU/rkoRXDb1z72nIB2Q7vTXTPCaPWEH76VOF+v
kNsYwimt8aFmsk25bQJxveqdjmK23ShoYVZPjCgmSFAr/IphX2/M8qR+KuKHD42Z
0N4X9CL9GeD8TjZbCPC6Ihm5GNdNo7TaDAa4O/Bo/FdCl33Mu/tEOsEvB12NI1bf
69xPFI47XtAn4EplkfSGrp7DAcIvjz3Osp67Szs8YBDgO2cXg1Rj1cRUPmst4IVr
SZJgwc6vNeYHXkkzyu4CWUfDX8/GTptDuNcRJK8HznibseSmjFpLz2l22gebFym8
4UFfXAkvqTDQQs4c1YRzBgYvFlZQ4TjVgYUrRZwR99ALquZSpAhmSqCGYvfX/CmW
egWqpR7lIdII4wDTNgLTVW4vKq02eAKp8wBeLjvo2o+5HbZmcYXdHplJItzWPZ8b
tAC6l7lsnJ586w+tj+5nfbThixIVVuHN7PROqsUnUUlezj9GVuEUWIxJ0ll8IBi2
33AbFJa/HZpFSODnOnewouMErpmU57K2iA/ZPIIy4eL3I2acC5jR03NyClIzOTEA
ilhCUp/RO1RtiRIOBU1x2mG0NETOnsUGvIkFbj/81mE2YGs+rBWIe6xzHlvajLjM
hmJ3ANBulfQrxjF0xHJ0IsEZnDsxhYLlYeYFASv9drGsBhJGYucEW7Htox5jU1M5
HOqF6GrOf4KJ40BftYwMc7SyZITindZyDFdu7xjdzRtj8Tgj521ETuyvRJLvZMEt
I9d+XtkuExX735Cp2TZsh9r436PTh44zTEkqKG1SwLtzhAZwBq4om+kXECi33ygb
+qAreMZFVi/siqvP4JAg3nsjEfC7kkjjgUdET26SO34lxgh42V9Mv7hiP2kAV5+N
03D0wNckGSZUmJrlhT5qrLE9keIqT5RcXyA/ofXiJhdWBd3PhTw40A+yfWZSRr4G
4hcwfRm2yT//XXMj45u14hIn1HolrzWu0qOq4CUvVDQCEnCp4RsCypDzCYrZLqnP
xhAwz1hfuZyMgdYcZiPIfT55q4Rdq0qQxs3hLbmcjeu61IkUwLyQ614f4o0wkd8B
eAgrZbM+xRJDt/oNCnWpWom/NxVajHw+ShznKZG3ocz8ZrBtZx2g+Z9VABMdX7S3
HoioaljoO8+O28CwZLM/49wV1LQmSASnKsueYOLAskH9QRr+a1u2Xl3s1pY+zkUb
Sv45TrADO0mQfhgK4kwrZwDNcmmcSzJvZSiQ4zT0MYyW9XJFpK1eAEuCWwdgt4W2
EiPVWyNJZpIAMeqy6BB0pgc/bNK5q8yWE2aP+RD0ttUwJSn/cGretsPJt03tAQMz
uklx7xr8jdzotk85Un0qtd19tU2Wg523YPzvBK0m8IGPZOzmMQ16Hj1gtqdF5+oF
swtyeDHjVMARuPqgtDIzqRInYZ1Enq7z9Bb1tJJZ+OduOoVaDDdoM2sKIeOFFDdp
yu62fcel7miLSzqbOpqDrHSgD3xItSoMc28QRo1xmgGQtB51d4n53sj5CaIfVXcn
t2VvQea+Eibv9egBD+9eOo9P6ujKdfcQDgjEC0syUGQ6u63Tuo56hSM03NQ+7Ynh
r556EkUpol3xs4Zc7IoN5MoJBBuAa8ji9+OFj8FDYLC7uHCbneuU2BEcVRiEj/sR
s/unoQGs3bCsBCd0fEimghqkLM+f9Eqq1gz8a9xXJw1j1+K+F6Vmjw5b91+fa9Wb
xj/IJGQSSldlvNEDbCYxlZ70wGrh0Fh/8Ea5xh8TT45IXDPjyFqekdiBaoQLGwlo
te5WYeNEUsOC/OFdr4t8gePuGJHC55Hi9g2wnqV88XnLuVllPT5SYunTPcDjNAOn
jWFknPdMXtWuirZVc9czmh45uOnvWYWW+nW1fweMoulEXKgMWVudMK88OTlqddo1
4uUgx3iHFPMQJVKVIT1PdnrqX6m2khG7kJcx9r3yQRJGHszn0KD6pmZKd74h1h7E
BZPiMrOE5C98F21wPamOP76reEckmcPc6nzqqq12RRjiU8UiyIKdQ6pYkH7xH/9z
78vo20BVDtQF/OKM27RhYIFWKxcdN2Fbcw4JGvNcPKinPle6Ylv6seEesdcNpVPY
BaLouTx2E2RFiZJjDeDvQl0ozy8nK2b5AYG5/Bzao6UnK05+lnSck3m66bdqpFAH
E8CAvH1kIR75f14A8I+rmdq+nm/rm7T0ReMy/xaqzXBrkNZ4RLpqBItmIAzITftO
84hAq6MssUZf05YJQHZNLCgwtu2MfJLXieZ5quVsGukvZTu78+zzC1CTu2NZQLhO
lEDPVtnkgeqVN3Ri0aUsrvfHhewbCjGkCwM/LhCv6T8UGYFt2flSlRWm1C+LJDib
EJPLeOppWtAOurf+rAvxq6VnJYfzGtoEYOMIP9Ng/CWJ0mwjgrfstdUvooiuPkoW
QyRFGS/uYSMZWFrwg9Bx0Wf526fx/86K3LMHmgi74eYW3BIJJn1aAywOZXMBKyvJ
w2oGLoqP/LLhiyLHDel/DKShWFKOiKH4erlDi6GL1bG9/p3s+aSU5nJBMy52H05v
s46VG/7p3p/qCR+muR2BL2P9fNs7NvAAjKKxHiOPL+Oz8ZK3tOvnJd+9Jk+IDrx7
ACF11taCSW/i+STYuAhDXImyxAd+Udnx739miadqcv0S7yqM9PWaF2lTqaPKqEdM
QxxF1hNO1Hy/yrmMsj9wQSFcRYyk6mpb+QdeOvoM0z602asDooGML76tRtO8wpgG
Wqet4rgKdyI54HoNC3p+7lbibb2gs0CHgOCO4HQODzLJprrRaJdWFYLbtifp8Wce
dQ8lzZJU7sKLhpcCizeJXYLIiU3LbTV74+fa9R2oVTZ/w7/PJjwJxi2G2ctXgI8L
j9+MmLqdeCkhGAwdSf7P65GLOoS3/04oLtIcryt3BSXvkFdBg2YhuvCE+lZEVfQ5
OqEzftSZLA0uYwWVj1HlYRJrHmG7iXet6AfQvTt2TV6ja1sRZEODlF0y9nRXV90R
5EuOUO7fs8S27QlIf4T518XDLb6m2NggXPsCCFPHLaPiLZUpWVn0yUgIrXNQN1M8
BcNS7ZnB/4Od1Me/WG2TJ1WRVq3AeSauxLX2Y/KgyWcEj4HEoy/vuCLN8hoLvAJF
yVG1kiKoxsrpC/viRVUiLJcSjYiDKdyIV7NhSmKNn+b3famtaT0e+Ou6UzXVgEN4
NElNLWS/vSnvKvUrRvFcRL48O1tHzHw4RsLmWrZqFNfZkkPz4UpES6Y2MD29a2PP
FYwdCtdkzs1IejGrNWkZAUszwmW+u853P+p7zcd/ctNmmBDnCjYVKSpVhFrjL0Ti
eg7Py/PgGdVTzRAUA4szCKncT7QvYh4P2VsLORnXqK3X4gmxvCCY1jfN8QFtvKFS
llYbpHZzsFL9irsPp/8+uljL1HFHcOkoBCSsVWiKjNMDK1AQVN3k0GxF96xIC3zv
BfFHhEmApOsUd54lK54WY8RGtRrvIx6JLcmkn2JaqmOlAge1YDrAnEZAUCzOKE6T
DMd1JMDKtv0WoMewsDyZL/lW2nYQ2jLle3Cj36kchdoMu1i3y3BsaZV+fqZvuzMT
4ZDWsDxtK8z0sUsSI2pOY+42+WtXre2PLIS3T+1PHbIJ/Y+KwlY8+xLPHIrta7t3
sohi7d291S1gYPYd0jjvE8SXcHwdmvpgXjqxsn4MYhc5IyY68p5I5Cfz8fZoLITj
hw2yEt1kon+F8mWGTi9QaqeqhlFevRB/MzzPvrdk0/y5EwMEagSzIgswcffIaOsS
H1MxA8Fy9gx7KvHaGAD/FFgLAe7qgEzMRgn9OQIgk1dcV9BCXPK3AVYt/nW6mftG
vUL6T3bJ8oSYCl0uTy14VAj2/pwydxBrzxWwaHpy9392M/3B+7QCqNQ5GrKIew+R
RZewlvI+BEevbmFZYncsenlEaROC0Q79tOLYpNatyiDVhFQbGcmw7Ro8aVMe9W9K
aoqlrvV/gBW8XkqztZs/Pgy19TJjhRJjNXtvhDxM71F+SsmLSVFKEHp6lUfdC0da
ef1DqgQQI2kLIZXgf2XJdBq2UYl/n/Izzk5HHFhXiv9L61NskXt5nGi83OPhQThR
vU+h9XN/Qjv62pJPcvchMonpmxGk7cRpY35Wfjc25MfJ+87Y0pETfptLeH1lR4sH
it51RmICfVgPlX2gLFpSUG/qS2bmuSCntttn08FfpvRhkOkNzyp7fdpmpnqp4mXG
WZk2PiVj7yoha1JL6x9fk8AAp/BqGgEaw0H47gofsWGdXP71qhzoVgxKT2M3wi+x
2PX1RjdAVRJzd9FSIEUSxguBrDYkCwTpGRKxIPSJJUPPd3ZmNOzIFSM6ZsQc6x5D
G/t24/sVe5BWRvSIzAJoXZpBi8Vx9qNG8FoGTnj8ukjRXgc7ihda86wOg1VM3dnk
P7b1TZLDVQzvQze9AyGr9JLmmoWfTjguDi98GWiPHY+DNb5JE3BcC6lJ04Yb7O04
wqeuIsWBgTyW46isa1Hz3S0RZhbbMLJFjBeYaBkbGAely9i1A6O0szO5kelusewe
9YCBgD4R1PLVpF+bbh20lxOsW/VyR9VuLwC7M/VWQkK4RfqL3KQ5d73l95R3yYWf
L1Cs++eya5PQJyqmedKwD2mxoWs5F4ZKKoACn5CmbEVKBRnS5lADDCB9v9lMQXCn
rOjd3fg6sycLGT/Z9nkNj5d0SDq9HKF+fekie38o1KsdzmiL0REOtSllXQZChdS7
DidLaJwD5kqxRa25BfETGxv2xGX570kE9mnLDDQBOPMsG2wQs9BduoDwzvIAcxeV
WwHunKhSkgDGKlzW/rQgj+s+wfDC5JW7RGkaeIFSbSj2e/VK9yhuPtqm/V5h5j1y
BEIQzv+yiSD7uICAxrOaidx0IyiVcpMdkiyaGdn+R9hMZ9Ntf8SfThbKYqCfAH6c
Rlr9iziB/qW09/o+D2ptdYbGPJO30NrFJW02QzMlA5051VRO9RohffBDYYJJu6Ze
TdSxK0LyTCWXj3YottZaA++XdC2slP2FPfd+V+TmGhu7x5vcRCc3VrKiIvVaB8Ur
HNqg8HlQHwglpfX75VW4yUkAKRgwhpjbAWtjQsc15hbMyycWo6B82GKBSGoImxoB
5ylXewcBHF2UQWIz8vSMAqTTh0ICv6GDADeUEtEpZQn9ShtSiQ/9cfqESPISJkqP
cdl/C5zawoxIIXCEazs5LjHmDHeJ+AWzJUTOFjKvZQk7Pgx5Cpe6rMxD9BAasxaQ
duj5M58IpHMX9m2Z6jc1VuHKNDkKPUNiTR5XKPRpqd5Ft+F34SN8RDUmtiWNABge
gyVqGND6MBR8ulELJTbKemxZ50WICJhw1vO2USUsYUDNluBKklufKH9oMF5du4q5
znKP1GNO0/j1CdPoHFZlX5/6dcEkmZ2Zz+69lTp9L+n+OiX6vxn+5rDXOcHY64CA
bnoOO5u2DhdygZ4n+NRq02y1bVw+cSF6hza5aE+5SROLauAXO0oQAGJtgX7g8tvm
Svod1Di7N0v7fPvkwWWyVrGcPFFxMzgCuSLorO721HOFH6ym103E+MbDQpoNxjEA
xDThmsTj2pHmdeJ21rPHkmIAiNQK2soVz0uhPQwtJaINZ8IhrK4nWmVkkm9Jbb2h
WMsE/sbfP+lrO8mKWftlgDUPyBPYjHFj2W2p+dlIuGnuEnLN0Ww6Wlcrkg/eyOR/
06t1FGE9jNozINUnwp4vYFEmtwM7gwVtCHZLaC7IBzUbW2BNTBRrCyhEqMot3LUc
OP0YzLuPEWhXmy1Bg8WRQ1Mof+Rv0RyfEVjA/lZjR0lJqTeInGX6tuFhX3LHHHgQ
QzTsZiNwylNLfvoTD8hxoBrnnKHR48c+VPRMscDICEsL4QfQoMWrM0ZgQCKP7jWI
iq2uzMWdEtmrYtMHYlJZk5eJMJWHYEwtWYiWoZ9L9jTGgNysJgf4OFTcGrwwWI9r
JvaUOtVxQjceQRdsDQpBMx/jUuIZn2u+0UN69gvxKCdaetH+4Ana52Re89Suo80p
ktrS4CEjnOb7vCGAh/BsJX3vzTsGZkl7D3HpejjPgY2IB7yaKTeiErIE+V5wUq1d
gVTOETRumDsz9OfFBY+p3hgN3/hNE6YGxXZa7aeN2LJ1ckCsi/UU97N0iPMR7snD
g6laavmk7exTcTyiiiTpOhEgNVRf81mff/KAhU+M1nELm3vEnuO7yCmdz9AA1D50
t11FGbsGXqo9hlKodTgr3XFGM5mXgGVdwEOhu+xdHLov6GnVkhGIv/jXf4LSBSl9
O4fq6e1VaEr7sxEjnzc7udi/l3rKsCxROabNiXp+7wxtzMltSTIxKmcLQYYP/rcY
G8sdq1YjsVE1erP05hom6eN0jKRW3RwSiVvKYtVdGcHI/MCrB9naQWguoDt39MMk
pvpcYV0tij3049C0csL0S0cJ25rwaPqm1Zy4CcdD9JffTIo4GF2po0JiOeDzYvNs
BLhoO8e0T/BocTs+QsJPUIVLt2KuT8JcHBVyuLObgulZKsIchY8oj0llzrcGD5h5
bXz/6gAwiR35FZmm/7I/MM9g8Wzyaz+tj8vw4hSI66/v3oFkqPjfhiRJruQfjSk2
M287h2y6Dokc4rJCs0zY8ntufrk5+U0XRQva1SeCZoIKi+lw+kL8JWLprUZA5Bna
YVMuIyetIaVSAWygn65fLtCMpHmitggCWb1ZVVOmXxo8hYGmm2T/T+BJ+jLBe/zx
v6pLIvAMTc9qAT1gYhIBYpaWr7j9PoJCjOAq4PB9pC8kANlSepkaHK/TzMhbc+wC
sOThLjHU8W6XsbwsHupVlEl9qlOLYNNJDkDBdPWiq3V9t54+OzWzctCMnUE+Ylvq
ddUp7YHL7ucMiAWOW0Blsi13Pw+CrYTrnk97ekAAF/V2PVrM2NNpmzkHXNLgDfmb
DkADX/STHVNI4kFpkqGq3/rsbO0vsl1u6RbAAKyeyWIn2xBvvQ2sbEC+QywHdu4i
iUGzYxLaGwGxnz5UQmMigZqoSruOZ58T/OiieXOJ6rJze67ITI/yqDNITLazQecI
AbHDv31CHFZJxio4VNdx6zREjg7jJctE39f3qiK4aVLwO/389gqyMQOaRs+SpQC0
hz9yuT7FjBqfKRdWau4wl+Z5ToQRvpOTxsxdb3gWsHX85VYOhoHmquZds78MRQvq
fIcgYm8KxP84O2U0sWiZNtrr9PhZ0LVGq3vzroe3FTltt8TJA5tmmlMOuUNmxaxk
F/rrKJtFnLn9d0vZG3XfrnH5sk/rb1XUDgpvBcZYkqUpLjh6NguxZPkQkQHYyVoU
uOk0h5w3HN923J+2t+4ZrR2Xfw3JTQhgLQcc8wvmIAksjxpx2H8kIEE2CJBBh0Ju
C8ip/FEXmyZ1IsMNMQRYeNagwaPEwKNZ37xAo3HRl1+2UpNnFjf/GCnF8EvfMNc6
jdaq4N0guFHjVnEpc3mXnJ1Pj9s80GQvy8KnS4QsdqxaWbVQwwoTGGyuaJeAnvfT
yHnaZ9xDyNSXTI/0uXBNwxvKCmGd2Ci0MGmVnryKY4za0tvzWMRBYuM0RT9C940C
eaqA5poPq1evdaVcqRWII7xenBNEO41o75rNZcEoOvtBbJmnu0lofqCTcAs6Loyt
NMcPAMBOzjtziXJ7G6hfWIDm7R0H2ZR1taXRI831yjTLaE739IYpQdtGgIcv3vpO
khpPYPJzXQIBGr+EzkBDhdjfc3XyRYHdiiAcw7kAR8AQkFN08DIjikxxZGWrN3c5
7ddjkMlJMAK/jnyNEigbyzJnQCi8GivIYeGMIfZI5HkcxOWeG5RiSn8vrtp3LWN+
yR7yXB0DviCBD26gRWDLV8rPMraLusqJc7i5OSgQxoU3wUD4fpEzumqm2gcVK95Z
Mv53s4Ol3Duc3bYWfcPmfYvq7aGwdDCDF+4b7WRsAsXnorpcDrMo6VK58TbaIrhz
svQxrwkl2io16WzbQt1Gb36MuGjUa1lN44kvA8MRCDZrFLpDvsIEIWM8zuFzKXzo
3YBQ2XXM+rYxo4lTcQdqbxSx6JQErI8zMEjg2f+GDPkoxjjXNvlJVjQuzZWdKIRl
qeTjRsbXN3m+UkQ9lU04Wr8B6PoiuCWACjzzQJ36/o6c3KaCnOzu+Y4lDr2t8WDL
XeaosQ8OZe181xjq9onp3dOBJJ3KC5UZw4biIOD8dZeSCcutS/eBzEc8NA8j9FSO
YRsih9skh86vxqUiZkOJRSndUYbxZdCulFz+NruV4KsBxn9HEA6HhrP/ZWtw0n3P
nTDZ/QfNQANzd5tNosNAwt++RaPkznrD+ACiadA8LoQYsfTsD3BZgrB97e7uMZpK
tMMYYGeTOyzLPicXant7ChQZ0gcPeaD0YaoIZ60eA7D2IZU/6tsRR2/buaXo2DzN
ZmuzrD5ZDFagFxWCSDU65tGMz+oawCJ5IBGEyY8kE+wRXNpm8B3KYH8Ir6B7kKGx
VsltPP1WTUgKywW8UpJft/7nwgtxd88ky2tfu1AV9xvO2/R8gZ/HtS8qDnhD3Bcn
tkg9td798ww0qKB9Xn7ZG1NFhkxQ7Aen8ZcnPsXZM9QjeTXgCmH0sR6bYJ7/n7gU
mXLOD6E2kJgrEzMEZ4a3y5OX+K7evNFuuPsbxem+n/lDYhkKsLNacX0WajgF/7zz
zBjpTOiZG9FvQBmmqSOa9Cx6TyrndoyqQ9fN1qDzv0Yzu3oRHaIFhlixMHz7hs21
4TSeckSBN2MVsGQXgo7Mz/03fQMGSJin7B1uZRiXDhK074kANeyspveLCBfmqF6v
4c+ZK23igSUdEenavYyVH2eQ53PUqNj8I4MqXxHn8bb/fgRaNJDOJMgg5y0LHgvW
YvevniqvACgiiP0l/ag9py8khaIriXNTOfcRruwMmL9vT0Naa8SD209v5SeKp60v
lvYcVvc+ARmKYcARTiLWIHyWvrEm6Mr5NbuuQ9SbI4688n994qwMlzGqllSNkNCr
BSkz8wHH6+g+efFYJyMP7AapTZuYkSMTWfu0uiQ8zl18hoXk0PDxHi1Nbq0KEHaA
rqojakrsxKUQ2NQDIgBN3jDm0StiRzR9JevTA7zHqygi4W9Yf5ve0yPWj5l/sfpM
T/bk0l6kqynCVL8S7lbwJKpoY0vuCQKl0g2ILRVYEa8YwHqZZIo7opN/CFszdSGA
aajqlAw4A0Uta0/pg1D3ofILtzBanrdUf6lh2BptA6zZwLxZwMjk9aB5KaCqyu7V
cBa6ucyRwnI/UQV0tOO1o6hKIxKJnef7zW+pnd6/zbI3zN1HTM7PA88w/21bIUJS
xqRwgyKlqgkq2hxy1VPXh2P0tyZ1XzU+nXYb0VDz0NMSTyoe8DMa3guAhoIexiqH
p5IFp4ruSjIZO+Mmqtg/onnpfMs36URPFHSNSP5JhIR8TloXTYFfExxqZU3WEyv4
FTxhheXkZ7ZCmhHSuR15HuYQIxW8ZwOQARKPAzvshoNgo74u5sbPHlFrBCzO1OpA
pPlCFY6ArW9ijLcTiV6DuI7ilNfVKXsKU0kze7QusFVUKmwJMUfAVhxsuixZ78Ic
6rYpNoiEeqHhU8TTpIjN68KPOIDzB5QN7Lhlu/e8Oc1SPFs+1atXWgqs4guUaIP9
vYdyUI6Aezi7sodVmyd9mhBU+YLlQjxorAz02yRQo65U90QQu7db3Vsxflzlswz7
kRIsztBTHiPWqZ3Cvm3+T+t3fVbhh7whkz9QzwXaihYEgU+umxjWy1XI1snmZXGL
2bej6c09P8GETTQ9Dj7lfnr5/asB0wBcBAKXL/1VydzyDACL1Cio0f/ibEFTmJRa
3dRPu22jzwht9XuRSmoO6JHTwdcDWd7v6Nt1IBwOb++wQcMTZUaXd8aWLRscmSaI
MD8T0a0O+8i+REZ32E69XsSvWLzcsohkozwy5wcpGAUZATP7wZVqzGCCiyObacTT
3OFlrRwGZq+vXKBz7FZLJ2tWjaIWJsCC5CCV8mgIojKMILkpiS63ZooxZouuJtxp
te0Azjes3sYrbshXjZirb6OmVdYOUrmSfCTYwtFGws8Y2WulE0yBeOfccnoKE/Mp
u3VLd9h4VhHF6j9ByiyElK7vmGhxpjhM+4g+coKtQLFSmVOUMmScpRjACSllicXD
22QW058sXD6aK+HZvkEmSwXDQDNjicDVl3UEdnbQ0XoUhyYCWyp3ko3MdCuK5VLG
+hxV2aw36SBWg9rpJcTpdlVMpyABhaLMAAsj7+G2qR63Y8LvvpBt9YYIUFCA02H0
iWlsB2n/Ivc+k33R22D7OOjUXE9/AaQrWB/zvW58j86Vzacs/oTye8iMTNtJbPeD
H1TMSmhOQ81KdCRzBxiEa0Or4VaISRvNIQx+ek/hEWDqiJAXepid0R0tEllbfQWb
fdhzJBl2mJv3rerIhXqfqFg6o0OisZdbgGXIKYBfaDHVpFGKVAkoB1RgL38T2V0a
RRmOAExGWvxvDhK3+u/f+ucV2/s1EceQOKk1xzX/UAPeUN4fCx3qmZjJpH/gohMp
ssZ5Wi7OaJCoflk7FJut7cGG5kE7/CCJH68cP1eyoRtIHD2aBjoFLoMs4XH0i6D/
JBIxcKtXg/wWDvZ221A68w4kTjfx7s6mXF5XfyWb657qgT1GZYfULHonyOUCFm8z
Xr9cLPYtlef4ccbOKwVUEAZSzeMTNEJoZwKhNi3E1C7Lthuwd1a2uW97YYUTyP2B
zVITSQZZISqEA5+uZ8V1dA/Hxu3UBjhnmxicKopTXR1ap/GTOLefIVS4FM2qyeqd
58DFpg2mCBXiTTDEjUejioQaDjYQwt++o0OFmAX31mTImg5hg7wV7fYlCso4rxrC
2KvRCmEcAZLkaUO7+rg5gopSPKsGiy4BfSpYFP475KTz8ufff36WDlndC2SdeOF9
n1Ow4kKXpXwotoca5nPJK0OTylJDP45h/57qBQMLOMD9GBVPAI4F00JWmAzPHljJ
xM0g3x/LszYFHn6tnp4YkH1BakIoIfdQ/iw09l1Pl8kzQzn523oXyfaXTJy7wtu1
ANwSVcaLxJk3Go5IxUvKl3qnjVDO1pY0535kpEgb1TNZGmh1SxByDjwMNoF7OEUM
VDDLdXQ4f386on4GRXEiDF5uUXzT8t27YwpwuVpkwY/F80etqOsnfx1aQx8kE4Tq
lMHXyOiPmovZq4AxZ1dvrQyGHBfXOWEWyobDrvjreIoIcMVroH6rqYDInk8siVbF
WSDHfxiByG1jf9m5DNF/Q43m6Yd5/EJmHr1Ik0zPDy3H9gW8AL+bgtRmYztss4VT
6sQF71cuAPZpR5xFAxJbU7NwQbpsiqn4vRq7+jYn4PZZzYBDZbZcqg48J+sdC7b/
aLhoPo2fjatxtERp0lItJz7xHmlM8eZTq/8ZJp+nym+qf2NUqA++8Mx0+/7JvUD0
l4GS33KcTvvOBE8N8Doc03B/8YJxRI6/WASOvyrj2S7qE15547JjqMqpT0KmjCP1
ZAoBzaNUidgK8Gbb/jfb3aGOT/q4SD95rd0Dp8nK/TWDDDstBazz+PcnJdC3pAnA
fc8uW7CcC/pMUrRjQEfAPtFQPmOIoQUtNHDMoMqXJLLQmR7R9OE1XofceXO154/E
e7vAq6o3nqQmqEmpkleR/rRkLm2NDfrXpdWfx4FQ9q3zxffk6oz9+1Shpsh5zWxq
L/VeoFKmJYxFI5XyYucuJ90z+6FYNmD6FUxoDV5m/3Z9s9cmt/wiD2LlTE1sZoUE
gZFxMOx+os2io+LijAOo4YII5WupBh2PqMiFP6hRNSTLGzq4RQxTGf7qoqjF4PJs
bjpK2nTKpvNv0H5uXFBV4WWjZs85RNxHerubPGTIm/piWHmUDZWd4PbLU65TdP2q
avVa4yRcrA1R2s0g5x4FL2kjASYzdqVW4/Dt5lPxRiRtQDctUtI29Q67DCk5aVEQ
zuN/oCOF+dr+xkhjjynHQw7ugGpw4EdwYlkpconzjJNkeCAVw/m7FeYyImnp3FIz
B1wovaxUhcZi6O42SFpAqfsnWVbSRvtK+dxojusxFVmC9aITiPPkW2RM7G4XhD6i
tcqsbsCYH0u71JHrMXt1OvziUnGQMVl8ETvwZyQS+PqrS7G0+Tg8Drqv0spl8z+U
zdEBNajxBGXNKuwrIo836ix1W66UgifyJr8TB/jivZhx310SxG9myE2hKMoPUFc7
httnHr94rPQfVSZGsW3aMjNxlSPnWME8zh5TY62AFrzcA63jXtBd8BOmdx3puwUg
a+rOAIQv7R7v8GKDQ1UFiI/a4w+VTiZQoA+oLvod6yUV6hDujwdNXg7X8JYP7OOD
PapmFZArwpCGJhCywMVoVZ83I4B2MyEQUjjDnhLP9FXF4PPYQo5RLgZadI7d8L9u
6aB+CIXmOQPVPAS82V8t8zCfsGvOpiXmvUuXDng3m0+GzhboQ0LwTQ15QpgfH9Eh
c8z/Y8WrdxcsoJrpikBCRNeUSOxVHVryrSQpgiefgSUz3oTfILjNfy8vi8JXzRbi
5AvBoi8XsaTOl0EQxMSjHk7cgOaOdvRO6sNcxAgQr01xprzE8LfzHf+/merpdmdD
H/AkbCE16GsFB+V5CNLme7kOPZK8sBTKD+JkjcEnu9qSQxiRe9d1uxVxz9a7nwc5
K88lEoZyQII8tfkxzO016eQ6vyb6ApCnDWfCSHHCugizy2Jn3B/vUu++D3wgbyPb
NIMBivskN+ldi3geVwV7DN1OapuW84QPE3C6OUcdvVa2rBeCL5ku+susOVrgdzGE
ZmNUJqDW1NUmwDFLjLIqk2pxDG/mp8fm8kGejmwatgwvJtkykBw51bzhVjUw+gaJ
+NpQ+dU5NOiYP33KuL8pS+yca0Bx2yG9UaJfSApcXWcMl6VGhMvN+W60bH3WsWK+
Lb/6zV/QgOyRgrNjvOECC2EGscf8Rv4A5mrxUJnLCaEEz1lnGFfzHDUdaYMghHsM
mD3lRIDZToRlx/9e7/eK2cAGLuZjdOM9AeF7rHGKL/NU9W0yRUFtDOq6KpcSUpzd
9Y2bJuu4aR7O5sM3rD0PZ8vGiqvpMU2SV5KscPd0SEI6wHDnmi88slKNmiDBVhfM
lXWBFxdtyRZ1iKgHX9u4k2Kw93dIXrrZd99eLkfdP3yX/oZXLn9N6UjyXoLlFgaY
mk0ElaFxfb4VNIbPi/pHU6TC+rMM0qTwICK/kvGPxNu007+02moW+Pjmrtgaj1EX
/2KoYs7KV+8TCjcOw4Dm49fkUjAQUYSCN+L+Sg6duNtDoIMx10d54oSk9v8v8gBA
qblTdG5/jWs2O3EQZ44N2iQkc1i+sm17IBD9yEG6QJBbfaP3RV1KK4JQktx8j6Uv
IPZO3UFvr4ofHqsEt/xIjgIz7aaj7aJRwr7JBV2WIjqTkJisik/mmwFJyRne3G5h
6f5vHuwVTfJtQ7rxInwRGCY9xuwfWx9yHmwEpBQbcPg8fKncwwUkpqFk4YRuk1+9
sIkyJYKDvwM8g+cPCXjnCtxhm7q8tV0T+qlnvGz95l5HsLWxp8WNhXKK+C49H9rX
rKICD0/BxD8M6tj5j4HtpyE5y2TTwS9BjW+mMkh5qla9LzPF+YYi9cK9V9Khyifl
uXen/9Myzsi2nzdmuZX80clbaNyh7bET8N5YhhKMTp2ZXINsn77eJwKbf3ZRHgcm
sxt+GJ/rkpx2YNxOvbkMpm29p8sOn6TFS0D9LdB2ePI8pSlGBTzEQWaSap57C5Mi
b3vQPUsoHYV1THcdeAcCubzfFuMP8igvKdqxYd7arzWv3HcKtYeLoWHeT411rzVN
ZjHWbuhB31QTTNDU9S/3oFPV57NXfo12b9VTIkDaF/LU9+k63k8i0pV+qIKoc20Y
AstT++cxrCMb1c6CGLrF9NRJ3gfmIkyc0aGuPmlzdo9HU1Pz7L/6uNGY2dhwcE/t
wvNT8LnjvgV/MbG8Vkat8cInAA5winlxC47FFHqX/dtzsPQcUGbThMiUHN3rrnVl
d51swu2MvBcPpUaKp54dg8ZEyySoByZn9fUDIlxUuJ76CnsQAhR1SqHRG+UwnFMW
sCz7KqYi1JWWNa53Iey5Yqv2qw2a6NSNkFb0Dd3WTKkvc7i1ihwTDzocxVNawahC
7cc1OlquBDDSDmp9/Fv+o4TzipfG9CQl/t/YPcUUhzNXBN0dyEVuIc40svno+vm1
aMVggwXp7AHcDvXrrDD3VTJ9dphucP2ZxZfWglAX3UqCSY80SMlCzucOKgnK/SUv
1lh/ExSwarTDAgNO/BZJ1Cz24iOK0h0xMJZY4vkJNAH2bPy96oWmZKBMiNrYTilb
4t19CW1ZeU+BvDV6dXhsXrPl4O7cQJYctd584uSWrUe5ekXz4/JJfRBm7pjMDce6
M4T4VfgimohqVEQHTDICea7vG4qhx4Tagxzb4uwZBdvg51NCMEN4z234xGjPllyn
6sSIwKc1DKoLhf+J+Zw5dSzg8iifhAwQTYvsAPJRsmg4dxBQjHvi8803UI5aBjF5
5yaskXTzft8M8FkION8HIEN0P838SSK1Q14VA4/71RY02GFrwvZp01SComCXNvy+
8UUscWltctPQC33Ap+kQ+yBlMfMplOoRMHGng89UuoceF7GFIHt51eyzP2/0zjrg
JkamxQ/C8hzRljdkqOHGC+Z8njARVhCmvzop61/EagisdvJ5KtDZ+9m7LsToVZJC
pcUQhBDnA9dpHYKycoNuyEuTuZfrgb/aCquW6GU9lRlI2Uy1mLsBMWWCrYeQH006
dqInqbxUrULkNi4wNh5kljYRr5o0KDcKvseQFKwLM8hs+SgPEnXzfX4Gtkv+FtPZ
Pvj+LibDNCtPdiDDUlOfu7ZYOKLno692t9n38tJ4V9wiV67jNBe9lU9x/8mnZPKZ
U9GPEy7B/Y9WUp7h58zt1tivs/UY954Mct8ylfStviV9jPhEN0rK48K5ufAoRzY1
05dJb7SzG+brJc/24Y3EzK0IEFNN8kby2WGcMhDgsBhudvz5psIvBHJ6NK9yorHz
Ho6My+TBZh3cOyvFErfx+7oxp+vKYoKzyC5+Bm5rQDQuVHd7PFOe1o3uJXbCNspD
YTa8Jgg/JC31b4ycnRIDVMmSN20iJU7/Q6K50ntcYnF7XwKc/6UvVX4Oy9vUXDJJ
Fa5sBxXIsu0ykpS9EQCugW2R9I1S9NN00t/W8b/jXaa05baxNagSqZMf30M+wehY
oLB4c4sFWUfw3tNDReLYB5tp5u7vbZjWQrLXT7nTziopkEdIc4lseyHCWICYdMNH
w5y8CL4gZVRnLnCERNV1G5rz5RYuiWL1ZxPNeLijaeMssI0BMqdOxc2t36OFsG0b
DuWUaOR78ExGtCXh+Fo+C7lNeTIFSXdK3oiQI3gFY+BXsEQoqZZ8fnuHDoc1HMgh
D7RMVrTP9bmxgKj6alpcj1L2cfhMIYJQXUXsx1sXydhVK6Jzwl49nVCW8qZ4lrOo
guIjTFj9cVZlmHChHK6x2+Lxp9Z0XTvHdBGFfRjuUdW7YDkp9wbe0Jz79eByNVc8
Sn/LCXENnlySRFpIuiqWD/9sy4Iq3Q5USYRx/IQBvImndgAeMUIuF1yhsdnGxOe3
f46xxDCtbSstbZDDq1RJ4c0l7UgvW22MVv6Wttz7ZqL2GnVFpLTqVajWHwaFsDv4
FqW6b4Y2a8Hj5Kz5vy7o8ysADWmSd4gZxHLzT/JtV/1WQGGyuth/VAZ8he/KXvc3
wEhzxiKjsRH8DssZ8GQfdfWA4B7vgqDEV7BPc8sXF26EsmxStnfOgKqz/7S111wV
1B18OZNxFvOgIqRTTl5DDuXnAqs4eCAVPsg7EhT5+frSTgq//lvme3n3o8MwepxW
v9PTtMhzT/VItx+pCC6dxXFvPtAEfffJgLKqUag2uz808D8MqKZOKNTuJc8WQOYH
fpHT7GU/7SbHsbfnmlOTfXPYPEGhicN/sAVpIFhDFLJnKL37mgpw9z5DNlNcNVK9
orC+9HWnQ2BI9x08WqJ2F3YlUqZWLkERncA/iq9z1oiNJ9ktqs50gFQKKtPwy5n7
tN/dg70Y3e/BhSWbaCasLXNH7clqbWgnkiK9Z+9NLiDumr0XNjciCi6dZjeIt+Mf
4BsYCSSEFx1VVggPxs+Ynj+9PTo5RLaK29EGykDycd/KH0G3nV4ZJ72WzspI6jDS
/Hd7U281dd19gdVdpy5LEZ9xha9xDlggLpUyRF2/FX/2Rg5yfP9cJTQMLE1CGqT5
1Z7Ilsnwe19erO8g9CZkBr3ulQU1Dfcm9Bj9s5jzg2wYpd1rtfiyQ8DrP+LAxib8
z/eWfmygdHgJ3HFIlRIGnp+BUTUsbnnbfAdCsIr2cBscL/ZE5yhxri91RySXJquj
bVlO6skEQ2cMnE4yMjZz2TseDsFou/azePgZp8dr4X6GlK5YrTGWC95dm+byyKAz
GIUAXoYmWF96ryy/H2m5O9UvChmpxmBBQqICEo84zl5uYSl6TsktPvRo+4GumoXO
4FbG3EPOb2QhWD3qRlIwR7PH+Zsj+42jvNhZKYY5vLhEHTZ9bhzElPj8Nj0dhdFH
Vhed5QPCrzfa3QlasQBB3sLgQJPsxiZnA7rC74JqSjLUwmsFZfzWIYQ5o4nIBGxW
3N1qLMTzErTqtGDgW6Haqe/8B7hQE0f93NIKlqF8CMsvqiMcKb+Va4hpYR+21Sfm
LdQiVezgfT6k43ONfCWmf7CGolL2d2cDsG+cTHVT/lyOQ2T2miTvnTb/JHM76xEe
VskoirW5WyCaSbHD+YW0tP6Pj8XAuslFVJHfgbyf0nDk4sGruS7f8seqPwkE9/a2
gBoEZWzDjINYYn0KQoQFtaRv+IKarlqBDeLK/pMFss9sr197TFGL4w+sU4zYM+sY
yTxR+HyhscVdab+pl1sx012l1lhEjrU28lJo8Lqp6bF0/x+lejC5TFOVnq2Hgk9u
y3tGYm+GYTxFHqAKlS+ClCe0Iw7SKaI87zBUX8TDb4EQN2kyKjcThqmdJbdpu1B+
lN7QtXw9lrKZLnxfyXFZIzocOilohep+cnVS8uCfzJ0+Oj9BtBLUF6TVlH0le3dk
n707wEyZ9Vz/QNBikxlqwtOJRkIyYLuoUiCvnKMlnmuG+SU/zPUsA+VSfYoQcN8V
an70u5xl2FVWgAussf3ZvdPn1IFbYOD2jObYCXq0r3JSGw+FMDK/aBIwT+fITJpg
WbBkNv5ARRlJeE3VLZsyCu+8s82eFIZJ1SYM2dgyV0Gbqbp4ke0fvHd3mY/B61gi
B2+C6YKQPnsZ9GCAH6vUYcIrTOBs+NCK4STPkCTBLSH0vbtN9xaETUq9FnVXnY2Y
5Mkgc/v9R+CU83XFgPHXTiF2owF3jNGbzjfWcr39Y6tYuRUsCs2XUmewelR/dahO
ndGsYDNp8E9iDqm/ibS+5NsB3zXEu7HbT4os9X69qyyM7un7+q5zhh7eiLoX4TyZ
vZSVgMgz1FtF8S5BagUsIq/gY5BgcAqvGa/+g08kiNA+HyquJVkbMa+uaPwKFmyf
bshysVDHtt0GtG8/cTHkW7MgOJ8jRZBEGFM7Cb+kp9ZR3D6Ms2F9xhF7cChO4bh3
xJdstboVbQh+s00SJOQTVQPQA9bjyTLTzT3swp1qKihyx+ioAWXLlfQky58iKSGd
0Cgz5J200+9m1gQ7vPafdW+b0C6+g5mnb5vGZn9yE+1VJlSQAcILos9/7qOr1TZY
V78QVRqoNaDqFUm/76X5uTAgIi6v7itHxCaVxzA+aN13bTgVCPPwZjVMBqiIzRro
KWLXCncNe0PEU/+VXROJA5OFuH+/uFLLxX/B679fHeYB22g5W9P3E/xnoG1807K5
bokEomhrZnfluR80w3cmPFl/ygmx+p7RCbNNVLwJHXR4OMjs6IyWXsOe9h00+e9X
OHDi9I2K1zvD2t0mtZZMHmtaNank0TD9PIHRyT+ryp/W5GYA8dK+0fZ+wVw+929J
v4/DV+TFxa83wkjq0zaNXqXPwi8llOdoelDSlp2HtKDOeMAPZbWK5HvYNudOp8/+
fgeNRZ3r2geOtAx3xGI3CPNdwicri1Ps9nLzS6QYRDgBL1r7nIGXZYWp6LF4GAzs
ulz76Pv68szhk4CQ7iNU9HKQhRNnLxTZ64c1X4R0HwS2zfCABC6hXFdLUcBGUMoP
CLYzUu3mXKtbOUEWNJFLaon8govgSYuTRoIVnlynVHNgcZ42z32ovTWroCUspqr3
wjGVpxogNtGv1QtV56PC6/r74fx/aM2ESDUOIMobm+KKmibNunQBfZ9R+4PiT3nW
TlXjtfNz1pjH0eNubQPHz9/9owiuXVhjBs2sBk6xwxQAb0mN3eEkSESNZZ9KTRAx
NMzvrc3DUt4zlqW76PEbQz3OPlblFjImD/sHXRg6VR84qul3zuUzGr3mwgtqWaAL
IaiRSXJjJu5uBQ7QvXXbo4JOdDcWEFxVJQyCAMCx5FAiTtvfvf+QvCekOPyFdUb5
DELihBB+7SdmpcfKcCJg8KfdCBkEnwGfMp7c++1vpTfKcxeQ2YJe17Zp0OZr+o9T
kKSpNq5mLhWDD0HIVQw5NkMhqwfFtN6mVwgO2Aq7czvx3VH5s99Afw65h4RYL/Fj
Dq3xhLUpUtgFFZYSAhBFWRNvzBx7dNtwaV+5Dd8nMcOxBXduecE9b/ZtgeWcJyO4
6DDJPcpFKBXE8GLl3sezStV2cJcmbULbFWZcFrxzNAwgJQZX8i2JeGPk8sJIMARx
uNVwSPkqs5Z87QVmNB76ENVJh3JKbfqk7Pqrt6vXUGYdXG0RztKvnX57NocrIKO7
HXI6PobkDQMFwjT+8qwW0LxmYKeHeaMEVlA47NCxFKHd5go1jYHwi2q5jV8HUyP2
cLMC95NmHmvjpvzdF4v5pTvJDBaIU0u5E5lcjDfgLJrvVleyDYgVTCRy3u6sWhbf
vVfmjVT0BfF/ZLM2p7WGdaqcnRgD9xz+PW6/NizxD/Oj+GUk4sACqxyUuTHmItut
GxCM5j0u0jEobn1yn9w69pYQDMfFLg5QSRo2QO4eaIg3xKitmdXe+MF1XHevqms9
mvF3whJWVUSDNicZISc9pmOOAor+Bort2X90Di/G4r6MqoA8PUjRTIlowBJNd8LT
SwkeVKxnljfBujLKMipRvQ2OAYmPrWviND1HhszhbENIkoAIHouCg2VsMb6VKqMP
UJaZBTCUS7bhDgrV2BXECN4C+upXNv039xLbb8hqSHPbrW2vduwUY4glqMn47kxs
3B2TY70yT70O+j2s9aDkWxwh+00sHNU4744qs3DoAr1RyFM+1COztD5j+y2jpTbt
u+VJ3aEjLLrZF3koUA8OT9u4Jy/zbPuh96FZeTIsX2WnL3qi/q4mXE3q4RBqOHxN
K1XTo54rIhAjZSBf/PdzCO5Q+yODy3CeybUSQJM+IQm+IulXWNaxM9zWnmI8Q4/Y
mTCl+4gxxKzhwprjaWLS911vH0EuinrrIlCMS8HRXuoYFLlzyiXe1kLkrm4C9JW1
261JjDHZVUDHGRnVh4a6JRbkoxdJiiEpbI0mSB2eSLt081qAzesbeSN+Pqh3waww
JYVsr6JQ0/p4qOlwXLwtkXobNRRF00ktCko5xshyz+eh8oCpVYK0Mk10Aymq424d
Bd4q/JH3w3rEbCQ3iaH/C0armCnLuPmvZxSx3PKhi/ZPFYKv5VThJk2wVp/+e3u4
V+UJ4XnFoQYVP00zNfCedpi9t75qsc1OB9Tcbi5FP9AdCSMKAVsCj1S2ZykIB8GW
vaLaYEqqg+y6LQb0ECbkRRxQru2bU4+QRscbEbvolXscZfSdbLtudb9Xj1kqECxg
6eIjfZcqaSRBrgBLZ623ry2hWXwUPCN4tR2B7QhCgDnpXmBdtGEiyicWjC2AcQ9g
a0UxuO13TbVi/U+SHPcFntyKB59VbIaLS1QDSIYNzpm/Z5Tqx8Vb/UgKuR8K5lYL
gG284u8f5bFC6sNHEfTivPqVUx6vYXW+LR6QuXXMgzHyH7Jvdev0srEH+GcBI1wQ
aaM9S4fi+WqbyP22jccXyxGSDS4qZOC4uwQTvahnCIuAwxmML0WkFdrcL4KXYtYn
4fRtIlrWHKA7CfNpwHcK1L+YnpvI4Bd+E+Mr0VE3MegZlQJ3jVSW+6Ybcx+HeYr4
7+Qw4NVftWwRkRGKGjKm650Liz+xqhCZolxiElBxsVCBd636IFaiyB2Hye1hX5bo
Bd+SVzyD7wexlPYxn2b/5H+T6mLztNwA4zdvqxxhEPz0CKooCVkMdHGOyQKK8Cy5
HD1BuRkhP2ZmWZJr+dWxYJImEboK/nMQrqOeN99CHhsFOtGJc3tlXsjNVeGbvk+e
NhFcLX8FrLQRRNW4gpYkth6FBEozPmQaF1mrYBFixt+je+zOfzGJNsYFDRphsRwL
eRlZoVNgucuSfhE+NpR4lPAly2MKFOiWwl2Q9708HTFy6lTzuTGDpKiImdym/gdq
oqPgWXfFCIhyw6bXcx7PXThluE+aIpT5OcSkD4ioGt4WGELDAnMpC0f15kd2mVFp
6YJOptiNu9/OET5BvbuRQogtXC08FqWE5EYwXwT10kMCHkm3AWmr4rEKjf7hGF6L
w+x34ColNB7Djigp0l/ROue7qvBqIDfQbb5wrg1V8DSdYqYfstf9gz44EOTcKRT6
hJFUqzl25SRA+4NNdIeQUGCwMRe0JGHSr+BLRKxVOy1O4vNbCByBHkrhanBufW6w
ryJK1bkxbkwIcUBmMtqLK4dsaGzHjuZgcdvYiimbjyBHFvot9/uSuUezI8Rlvigy
Ia6rUOvSBY96+iMU1DGITBmGid2sDeL1dzLPFqZryMe+KGaEhZ7ycz/zK1UBKUXF
r2DyqrAKn0GJmMXUknC35j63/WqInuTPFNjyKeq5/E/qP5tPFkXJTS6vCgCPSfKg
M2wXwr438m1z3va0TJW6nKrn8gYY+MVotfgFZ4eqyJO1ZPWxI2atIJdx11570Wh5
/haQNd+gV+t4I1nTJ1KkvQ2IxUXDV1pqAz5IOGieAO5AiA9B3KVQtPsJunmKG8Xx
kMLZRJsoUTi/Kv8yC185iY0jTHtKOA2zYBmz58p/N/RdCzbhK7PniXsW2IJKTlnh
48y01IkFMxpHH3pt2QU4ZeLDa2+o0rNRIuJaf0rpknoJa2LQkvJeoeEmTwMe3+Yq
UoyfG5OAmia/sQpmxzGBAd3CxGb+NGKczpVLSNpQIsTRW+P/YqHCimZE6wKS7vrz
6EblCdde/xBLjVMNl8BZ4Z825QrDTVGPcku7E85AJAu9Y5DgV65QpDJClofhGltB
7UzttozovPrd7K9L3Si0HZs+y2qabpApbIfPkjkuaKQKQFglxvfAtQ6uBsAskck3
5jVsUwVi5rb+C00JnphcdetI5WUTZ9aUgJDMFKaktrs0VjqkKlCw3oRgkDm3IGKc
Gna2PxbwAsN+9nIhneAF/gEnuSnh+s47ktD10fRtFmXHZO3foSxOMhB7wmDbsiy5
81FF7CmVDE8SA3hZIhJOFG1Aosxgc2Csd/Mop9z2nfbC382/cdlxgJ/F1EBrA2KG
wXs3G5CtEsznpRDj7RQ1NwfsI6om/PyROjhG9gPpgvfFTytQUkfMQvPJd7+XNmlj
5VZpYaE8qFZ8zjk4/BqAi4BQzd0n4CCUXk8UsbFllqEhINko/99SmTwvGfs6eYWH
qcFVcdcYHKVruwJ5wMN+KI9Ws4zVFrJDZewhRZPe1S1NdLn7nOJzR1giDg9buLDj
3Xh29djQYx2Pcoo2IhCY3uJDwxFGCUlJItTXHBBX4OHaW48Zfm7Gm9XzmpwWmrEU
2VGWKhlL9tnDlLhJwL4YizpC7rqHHGAQNKOnDnhjfRl0cMtDuYQwLXtekQB2ceyL
zaHAOE24vVXISu6J6xuGMtZ6K3YYfl+W7BOuVkWXnnS2BUZbutXs6moMHaimg5zj
gnBMVY44IyFAoiW8OI/R71z+iAwTjNXRAoIp6t/zyVgVS2Oc5I6lfzMiYHNXThEI
X3+SB2IVrb2EO2yzk0i26PiSPVQNmFvtKLO+2Yfjnv1zgaVtBIqWkbAoUvNDvYr0
sQGxQWi+minD1OyZnHWkIcX+rrdL9RmSH9rDEvSPMNkxqpBD3JqmXc5SIYH6FK3c
agFqVxm7YzAT/3tnihXzulIrgxNl/glxMzT9wsJV7TGCLZNn1ZuueN0wqtdPDRfT
gzdSpKfEuUS79V4Lt17szyW0n/ip9vRhYQ3r+J2b7Lq5mR8WBHsUDgw6TuHnjT5u
KRAK0mX4MFruurnZR1HTEhfzBMsXiEnk0OpU2uBpZMMp5pvcmcTBNefB3pEqWwCk
XxzHriCLN1G/8LH3TwsMI+J6Eo97VR/9eevyFMV9hMJHRLBS/aysbnIDNPyQ9NWY
F+LXdrpl8TBw+UGRJEsrGmJWJuFaLrNRe6slkh6eCcIqtRHnXWidWj6b0pLv5QEj
L+7MTre/Ifeh+X360wBHLSw/ZQBSYs+cx9oeKYQ1R9F91zFr68ugTf0qI6RYeMhP
N5J/MyG/dt4RE9PdegCokIYVxlhZR625xfGRXg0G1TfIVKD7vl5TUNDUvZcnUJvO
BNI4TnbTWKXEBlDXHUHjSFUWcHZ8X537JdFApUocngzrmki8xCPQvY0Ss4C4Jg+G
i8bjOt7lyb7ssrlwYCulq0relAodgeoxdAAxEWeNZFCod9zHK9595DABJ7FLylwU
E0GkqrDGHMC6n+KKbBb4pQa/36bjYAf1PUia1PLh0ViKhZxOCW869wEzA5FSejv9
I6Jwy7PprE872wJaHx3c3BpKBFo3WJdRz2P9sW3GBWfayJX+vlmCNS0in83kiWxD
7dB9f0/OXJJY/ceq4jV1j0h7ZZV98xL2UishmYNKnYQdkL9jJ0zlWZxz7sbsQOqI
Fq/Wo6jFRw/z7AiTFf+aAx7hY0vh8FElR6+HC189Zpvg+uTxCQnR6zDUJH0iC5IJ
P7Yh7WRn/r2S/D90BdgyNAXsQb2WvNhK4p0ZmWuB3Y/r6E8UVNSetwuYvFJi0Yqq
DmkEjvuL1CkdC7BBGAFESmUJZ81WivFLBazpU4id8A6tGvJs0KeIlIr4bT3Z5p1j
XoP0lMcRs5WeurjzCG150Tv4J1hzi8M4hV/H37J8n9zki6t0w6FbWM4kIwg2woWc
Jwsik2we2i1KC/7sINRLc75nFZRWZL5qqfOP5ktGJoeoQDJwgZl+PHRE7K/Hb1iX
/OeCT8F9DETzHfMTnCvGuzVo5Xytf191fPP3LcnCRs2o8zapyOzl0/YFrnxoRKau
Orqnb44VMuEYtcZl9c8Bt9oaoKXAvBMN6v8wtoQfNkcjnYBnK+8A6Vlg3GRFGk6M
HFJvCGO1wak5Br0oLcHA5uT5NuI1HcIMtDQTAv2IHHw//F6bZcbVcif9MdaSOrhm
zqUMHd8hTLYXCRHzbklRUtltbF11TvqqZInVaPYEkK2TT2BsErYs7qTsyp2/Tm32
L8RpmIDv/jyNgfW+g64AfCISgzctHbw+s6a4peN1xq/vnK5PeuBfi++r2loSRFOR
Jkw/fwKGGIIFgZvr22LMpdUXFZtV/BhhG7yrSSAZP5tdgagNgzFea4vQPTUkhfoI
Q0h1jG3Jckhmevyq0+VjWWymvx/30RMgtQqJrAsu5IUlTxbuTb1SDRdHar9MYyrK
UXxohf+AWHN3VcvIBDqBVqdwHa+mHbdgPxDTqL64L5ZIfZluEFGXLmZw9h4MGJBM
pdc5wyneOaJSODN9XqAYx4+QuSW8hPcaPp3kkPzLKU9/e9syl2ZHn4G72a+R4Hal
xIU9v+Z8lfGeVqWXOAKi5biwHZSrQq2RuWdNKhOlXP/lImTM/rTwQnJ0PwETYTqk
vK1jg6Mc9nUakTMKVpXl+Hts2zsxIzsPJa+MAkBJKDqUJtER3z63sEIDr/F+3NLd
eX6PW5aGuBZqUvgS2YbaUnEp4X93pRA7i34zFwBklo7yKLI7a3zkWyUeJeFR2lp5
p4i7sHbbzEHXr3rS6qw0a2x5mMWFEXXiDr83KAQF0AdRuM9OEzdqkdw/EgLnfmAA
ZNhUagbXSqGN1qwS+jCKLHz1sD3j/ayMMNJlGW5p87I77+JuszHxh56024n/JcFg
U9l86JujDWOKp7oDlohOMe1mf0MyqOreLk0Eo6/6Qwy+gIHsQlxbx7AWVOqVR/E/
DV96wqW6yuwpFml6yY7BW6z8/KNmLfEgsL01hc7Ht6PjR0wSit7pzP/887ZD/pKY
agaEqDrm/yvuD2QTVBUy6GPc0FowqePEVdoi6tPCf4MM/7lLV3SFXdJRoRPFruas
iRVWmx4pknZzYkSwDdCDeJ+EihW6EHSa0UhTIj+381nYhT/Dh5yx2O2C/ctbx9aO
pi/rZFEnB6ad2mwPY7d5Qb3k5/bPqMw/9rlpcYtL9IVTu6yOY6YTy+BBzjbroO4O
rpX456aOSa4uoDTfl9nXXVPFXT4Ye/u8d8D2xJ1SUq2ig1kh31nQCaFUNt3uxdx3
Xu9KZP/xjXt+MEu81MTknPV46l5ufjwdA7StKJXKVpIufYrCuCN6EuvDF1PZuTkj
KaTFQxem2usHipFAY5Kidx6NASFlR6YtLlC/juZZ4WX0vbQiK7PnoKSQWAf87wf/
gIhxEN78V7DbN0SruvYnUuk5bNMBpoqjM4b6bHfTE+e6FkWGaAB8DY1H617EAiwx
DvklrrqTqYvVixio8jECrXMmS16L6+YpIJWIHruek3Q+603ac4b//pn51CiJFs+J
8ygPcShM+R2ZZMY1v+mNMuw6f9S8CDYggILWdd2NJP9bheQfM3AcCr9k0OBaLGAM
F6hDW4s3f5CB9U3h1NE9dn5zmyLq4sghgulVBQIU9f5ge5COOOzTWx1FvRpYPFcm
YqwC6cIHVLwYa+buGa/SXhMEhOlbaIRoiTBUO63t7NRPwah95VEgd1zYp37lKThz
2p8DlRRvknAPHf/wAG4Onl+6wQKaIRt0kIoerFU4ojajMyS+AQuUtAglrLsG7kpb
tPtj45neqvaZGG4M3RFgGbDIZ+Z5aGbltsb81wm1XhFq2TDYleCc+3mSgZpF/7lc
HMgLNlOo5uqBsBrNoY6RLY2WZEBYmWmrSJu486tHKKKI83r4DtgM6TLsnHaTNP0L
uk+Wm6IoXvcZ84724p/NyBMbGxo68T6zcNFfwZ+8nEkyIkwVJh92He2d37c33yvE
KFQk7n0faEEa8VhT8bmuBOYaT3to6sw8oltk0tWEkU2nITnNF0GTxKrop1fvUbvM
vKqfCKppUOvM8aftUXuNDFlOS68Hm9fQl8oTHigq5HR7ku9gYNzXZw8+7kPsqmTQ
0e9rKd+uf+Le1YqzaUfIAqZsntCDh7Xr+HNgOAXhd5bRtpaZisMqdY/8Nmy7yf9D
Tl3ZyKrWPNwFk/MZXiSsExk8gbP1yJ0Iu3vlCHOEe8+iE7t9zVe+nmQAXlFtElW8
gQhtixgu+TOPHIsgPBGZo5l44kEpSCnhHanf8vExxQRjdNJbU/InjnnBP60jymDY
myaow9RtzwIMTKHWFelhn5aAZxNQAJbRtVzrxLRC6pL6k8TAfzP93C4NJbMkIo/x
KI+tEkuFDNM4e82/Fy+/9nP00E5Cka8fLSAEvXU2zixpNXZLtaLzy6rxF44Qzo3S
2rnhVTzwyvNHEwjZi3xEEpI+FW0nzOyq9Vs7U3Fod8c1ule2J4qnt2+gu/zbNOHI
Txa5hNgNYFLx9zMwjuxYWLFys3Jfg0DI9ql2RxFdj8JQaz/S+QMPPhwp96vTU0Jq
R5IlaNJ+1FHIwG4P2o+FpQ0L8cZyUFazdfoAPO4nfTtF1WI73hfsT9TuhS9R7CK6
P/cCzkzhZQrPyBaD3BHHUiVXR202ey3aTeFLr1EPt8C1sIKy28B+4bstJ/AUelRO
uZ1LAzLfGS7GTU2EEpuJq8TTWUxb+pXk2LGNvqNoCn3JlBnDXHUaebfjga/IEK6M
YzWVVmN1lyP+XzQfsFj8akucQWTcpaBUQfWMURBv5Uod8wsE46DeF3Gul2RjYehj
8hCqWil+g9nKyBrbThpdTJifXsr7qr4yW4QB9Akhqdp5P8kBFr8DlmB1QMlAvLfD
Drat5u4vr5KaY/OA8h4oMEJWrMbdqoq2yTI0OrCOMCJlyQ5D6nnl7RiQbSQqD0J7
yTgFgcFOMkp44EMeLWPuxNLUdSauwJ/Js++GP4M1kN9RmvI4Vd1xQ/XHnLqx7K/p
9oEhuaFeZHA/gW8w7qGmrLPAsuyjn8dxoBEagSaRcQHgxSl1ky7bYjA7X6U8mHCo
/n4I1OiaYd0qeQWnD+N9b5H9yqIztMOw9DQTS8JFNAafTR75aSlA0Lb69GnQ76gI
NTSF3mh6kUy5lu0q96iUnpitf+XOvfpyg90NapMokQaAwrJM6UaeoJzGVliNU5sl
3A6aYuWmyZYMXSvqCcbmulK6t8+/5GWEtyH98rGw/wV0u8ij8esM6IvcQ2BXmrqt
XkSGIw2gCssO2Hh1ASgQtjsbJg5iBYrayxhQBBbT46mG0bojc9rieRHqOIw+Qel8
n4m4gy73ztLBKB/+qTqiC3UubSIXacS9Ckzdu6hH/QXWM0dADxO+vE8eM0G90tb+
13/xTjBXawCTOMP7U5wMKsudPB5kuoCPwenuXuUttwPjEUjljssVCJdycC53PlOV
gYT5EBn18cssBOmXE4r8qgJo2pgbFeGgv4aMHERloACyO5gIgiItAMuBhWE1tWjf
0wkVvimB9ZOvsetCce57NlEJwiNzry6s8SY+lO/fTn5C2MHvHSJLVj11Pi9DQhxm
PQYzWGUudqdm//CIsJBwykSnn4bagtukoMZFUDT8u5uzLDzYrvwwnedUpPm5AMlH
kNF9lYuKCfB/t6LM2JD4rTvAN62hRQ/3CwwZ1c2kkTXC+oG+l8CRnl1qbGCx2SgI
14doCfWB4aUh4pjArNOOktGZhnWsiiwMAURnQw8vtWNHm8DVkX8RVOjhdbBFmK/d
ysygv3X9sjhV+4jGG1nEtSrEhty4Fmt6xa4GwcChXwI0lNLDgV3Ypoi5/ZkDN4ba
jobMcq0cRKoR67/zs6MhBRfoAfyFHv5tozt0EZO8L5ZKoSOex1sag/arGK+KInKr
zrvHEz56gieCplsvGV46G8K2glxeUcb/O9kkGfWu3woJtWp52r7SfTP1kFRNv8nG
uU5ZhvaFo6fG8wIdK8Ov/kC6goGTkMOz4ppPiMU8PH08pUdlnIk/6MevXBAe6i1E
KFvS61YwxmE063JFhQnbpuLtNX85mY5SnUiF+618N2LyLUpO/Q9AiOmGg3VYBI4X
g+tVJJZIHUZ3Tz2VYiXw1HkjqMrWeA5cYrWQKj6ofQn5baz8oxckcUk4FyhahwUd
CdG1ezEw0SMasK9DqiRlEHtqVzFts40Ygl1zUE/aArfEwRm6cbaJJXnLkhz9A4dl
WDzLwYRa+gYTBgLZ2mrTdL6oeK4ogL9xdIaGgiPzQ0w64IzTWy2so9rCkqgoCvDz
DgVj5qSKDUlcVqEqwRZuGWtahL4oCDh26iB/g9uNixZRKkR8d3MYbz/7NfqMOZSS
Ea3poJcI7QNT5aVgDkWFmBMXS2Ze7qHsunssCxOAnRNF9z+Rv2Bci/JEzZ1ULOo0
o3IlRf4UOXdH4iWhmcff4gjNARK2USJEmMBK4VJt/ugXLu/VCFa9bTkrSx4ksYsy
f3KZ6Bgqcc6p19xbRHQFvlIQxkWw9vBFEbisljpZYkhiMCxJT7xVsTxoG+6aPGQP
uJq5drXNZL1mTQ8qYovMzOGmDc224DcaE+ehxFiKn5NIf0f9I2pQFwkdJ39+gHTh
GpB2CI+6N/yX+lOf3uBZOcN77mCUnJ0GQ3w7RpD9fMGw5mYXmF8Y/jicZXunFaTU
ZaItkHIc3e90XyCeYnWYKajdBdgTeugFEbVeETh9QW1h6TEuIzyyAgePfVPazeEV
VGNQEQA3J0igpf08hATRxfWjdC4md8xdwKrAGKYWkjwW5+E+l3Iq+WFJ9jH6kLKg
rPKfk/N+Kphkl1oHFu7U/S3iHldFpuOXh7Hz29sl8wJTPvd8plwKgSZ6GXrgser5
0udZJkPzGKKY9znFZoWvkR4pYAJdanDPBGOT+HwGzTn+g6jWpuEZogWmL8kDHh1m
+zLO1TC07sRtkAquIcUYv3YChiAKj4kbTUsgOaEFJKobQ8SSkymqdDm0YEXCm3vi
l8u94RLNHdZGiAJppB7k6E+Py7iBGUyEcB4PKa+rvmDWkTqc/Sd6DZEQCjpI+wRC
Rg/yEw1xAahIsN4DImNL5+9mxl514SSpADEtCK5fz0e3Tt3hixx7eZuHMhkdqrE4
mjjgSlICgKk5W9WczpTjrl4WIOHbtJG1UGa4+ktJx8+M5OlQzRJ1cX/fhjOlawZV
Q4r4kWaToU/Oev6Xlc/JihN02hnRHveYRpQgTZxqaTyK/hg+mMqUcngcp67jeAse
mAbCdCkMCVap28YgR78Nvsqlm5l9DlTVNL/LPphpdcFWQqYwDizEUMEiLcWFJG21
z8kd0SXLWTyeegLmV4/AovOBjnJhnKa2hB0d4qgOofhB/8C5REq49SliIksaPRzY
SteZrgmlbXMOCGFaG/1b/ZDHB5UrX0D0Vqef6gpUpsIx3duS69IhoSxrOpfVLefd
5PBOhk/U1QGUxRIfE1KBkjLyVnt2twCfZxYWP4HOFSkTDK8C7TxzlpreFRsaEnkw
3THUgUBqTWTo39Ax7BnRkYz9csNEyvHYqkaQK3W2nm3EmeCadxZBlXsDrn2M/fIP
ViycRFwxcBGYfopzCRa6VtKV4mJQdyECWWkI3Eu/G1qtLsswZgDCXWFl9FaE2xr9
+b/2JdkwdKsUlx4MjBWKj+hwJ7B3A/lh8Qs1yx88sq1SI93bDXKz7TSs/qymzbiP
x/TW9/wLvCM/IvOuOX79wSKg2dGOr6isO3d1SVD2Z8YYEla6eEmYWX/ha1MYctum
ah4ew0UUrlYrhqbbCj9uccuEovbz4pj7HXjRWuc1qMMSQbhWZFdRg/udE0XgzBJd
OLBlHUHrmYLPWVK4t91L9x9R3/k42HpaZVWwv6JUI6t85hDcWKSUmNMBge0LORh4
131pqd+0Utlii9hgpKDp79Eh7N6IiLpJg52rdMmblRaBosD5R8Uldo5ssAcb32ci
g3Eqtfx561x3/DhOJbl6tEwrGZjkzOtgmRPrkgVzR9yNtT2x5+7S3JwqPGMSnaKO
yIVY3ISK05VvBuRGXNTVAcmU5aAbp6aaFyruNA59Yn+q6ebAIfiasoW2bF2B+2oU
enDnAQYFdfP6agLMBVVcSJSlXNx0aioEMqS5PKyNQL5J9wMRXOSQsZlZsu8+y6Q1
JdngX8a3U3f6Be6GfPy3IbtjgQvcXvHJtiptPsZx6L65jgAoOglwK1iT/X429dJl
Z34WvhF+ATY8NMmRb+T2KELk55FWAZMcRRcSh7U7c+oy3K7qIFHtRWFCjYwI5nGS
obKRLspu88QTUyuqUoFM8ZMQ88TGOje6U15Hgd6VPm3GUZpawY4t9XlDFCjSx9+h
KXy62nRfBia/XwFO1VsU1dMvrZTcEfl7u0Pf9OVm06k2xRKqvPKJgXTv4CKRJ+R2
aoNDb9/MDaMmbMN7PP0uaWpk5YW8Pg5Ia4PurcwOYUtT1HRsoHEJzcpcLDLwosD8
Rpplnq2O5Zg/AtVahzYcLX4MO2KLIYdE61bUm4DqjpR2seAryfd1FcmEUeG2OVtg
yokFzRZI7uleln1aTnfm7Wdj8Xt3hghBHxjbEiIJa39lUXSMiFJS4APemyu0azGj
+k5zPeFOhdjZozoIeOQLaFYADX1KXDnEI/qaNHot7im3nPQ6BN+gjuLSOmPdSMQx
BNoa7DTl7M3apCT4fYah7H22lbjKZ9uVncvTD77R/xPGlIp9TDtQMrMDaqJtXp3P
WMXQVY8SgCo5kgF1hFWnllEY5clLbM5CxrmrkO6rGCMuY5zGlc/E7L8eRut1rLGD
QdpU9xxkcF7jy5fy4LVc1xP72OYbCiM5KheTUwYpiyRhLi0LDoVakHn3cxA878La
kY7+4pJoVD4d18Dgm0w3oz5UHtIqCvhkSR0fUuUfJirhtawI38jgYJB7jSOHarmS
4K5ZgVp9FUW1V4BlTDHPAyPoG1O+2MyURGFmTVLzK6dljC9ivBsasKQxZwLHy/hd
u85ygsJe7AyNraCxup59Cxjgy82Eb5OnaDAKnNiyPKfYgmf5LQPBi2oWF0pL3Vr3
+vagaeWc53+H2BMIR0LAas8jV/z65nLDnd9WMv2FLTaMHMmi0hfZ19xjVr6YYMpc
aeWmThnbyWG/19PSMpKIBn2m8OrSUq4x2CJHex/qTzUZk9BDEBYuTtSrC7mB+Kkz
TcjjpeooZ9cDw7lZfgU23aau6X3D+P7r+eBDeyMvvZcL35/FXGo1NIr4eEaKfCY3
KA9uqegOy5/Ju0MAVLWaSsDM7KypPZe9Vtnt5USj7k1bFdzlNGNptuMbwDoyqbCa
ULZUcuL5ge6Vm05UFi7bFL38S/Ylhys6mP7LwD8tJDqGc8NnDnghgTlGMKfXMyAH
l8WSvMzg0+NLaKfXfk8wnTO4TIwiCiMZBpn+Ycj/fpiyQ6xG/n+ZvS9a3bz5WQF3
UyuH72BLiAummnK1NEYeAGBM9g400z+5KteMNsUzbUGog917SKoUvI/7UuMilGMT
+NhyYhPBVUVGg0e+47XbTGDlcM7yFOGvOP5RkxH7t8otH+0NfTFNaRnWzkzWKBI4
ypvsqbPMtOMLFL8xSwal2rPDujhhAL6aqD+1KKHJnxlZwkiefMe3WItda48lo7UU
hjr+6wI583gbhGUtBO90K0v2eKSENRqNxQ8L35Lyma7X5R3lHpYlzH27u/4xmfcH
ZiGo+tUNLw1IEpQa8HGzbv6YpnIjnCfhpLvGEc9ddHH1isXDFeUrQJTbovoatVxo
IbY+jfe00UG7EpCF/1wPG+Z6jDA9HLQ9ZbVTUCb5ExCBZJ+8BIDBuyp8WnO8DXrW
VjLcdgZcTHXMPIb6uQcyekhCDiZmkPDnhbf9v8dHvzYDZ3JE2EjwFR8oJy6E9D2H
fN3675DD07LAn+u6/IeTxL73BbGm39oTIBIFDz8o2vjnFS7J/lQck/o9FYvHg+4D
gc9vWaPyPnG0QPFr0AguLM17/kyu/CIE8Gq0GfDxnr35+rQr/WyarmurRrcaPUOP
O+vXiZEtiiqc/cUJoTvs5LZACyokOLD4JMNMRXV/643vUzes1jsyFJrTPwba1B8L
X/xCxxcBs7TqoK3Ukm+lve89NMCDJ1cg9UaiHDXSS0Gya+OInUsXbfcGikm+MHsQ
b0s8LXNybpAEBK/kJR8trerSmeif5GSQbaNVrHPn9vaXliEKLWToLA18dTob6LxD
GA/az7Kix5wX8osi+6arfcEOr/i5VbL4b2xuyML0JS7U0GP6JtDbifhUF0Hr6AZq
uwnMVSJNjinrFsWVoGL2864Gpvj/47UfDr/IQXRaGhl233Cp5x0L7urrhScDKkIV
W6Bwt6tUXxQ6pTjR+7QjZ3TvixyJS07f3QGLLSYJ946i6GiuzWnhF3xykdQaGLrK
zjo44XJWJDx/Oy1EMS25qNf/h60tQfc3VEhLHsXaF3COp2qhFx5ur5LGX5ZWIPqE
+FR/N5ie/RT7cejlxNDSedC7Ggj9xi9T0VpNJlZaZWY5lCxL2o7KIqGQ/0hCJlAw
cH31mrBZDODp8jygWw089bPei7An/7grl6LymS8/O8O5Nt6G+ooLUzwA7JHVPpky
CgrlRvpQRnwZ446bO5cQOB7Y8es3GLBkWzagRAb8c9S4atNQmUzwdeB5+xrduOmK
LVEOMdLhiFTfdVYQFuTsMMsWRG74c6Dz33zvpnmPg9FOyXfESdrbs3xNHmScvugh
PgIY5hkj0Bhevdx+llJ6lueSU5IpYsvM0n0E8wAju8yhkeUKB/vuRo22v9CkJ/t9
/7NolhxE5qjvPYjxt4yd92aqSFCWTbfU53IXFJ1kzCbx0tG1D+c70PE8S9zEE/vv
JHE55LKtMvYF99fXMGavLgN5Bp1BHarfF8E9BRK84UdEJza4c4F4ZjgbALIyyHyG
YSG4Re4ImbM4QlZHUgJofjrZwTNj7k8Qc+CkMF8H8OR+XVPIchPMlMpZSbp6Zrfl
0jhzSK0kEEQzbAXukUrxtRWNpwNEbVtPpsDR1mzBSfxlLeWuLHCZ4NmcMuEwf6zE
iXSyadL+5llE2k1lmrkBfDj+jvzu2MSYXdUvX4qeKPXoirY0vF3W4lkdOmkcuuB3
UFcSxIN4zFeYkChNBxZ0fB8yWWNktd6VodkuywyLnSYRJJNNzvhpz9meZtOPrH25
ep37gGwMKRZX6kCzKNFzp6Pg7pMLRIARffhTni9etLpfyOYR91BEM3G32CdVX9Wa
sKWJT91m3C4uuIFYa/xCg7lHfVgYDrjq8gCSi0lQwsdSXviOwpyS7dQlPxwykpYF
GeSmFMXELJO/RlxX4CKupofJ3I2J00P+eMbInBei/XbMPk+mJcU0VAsC07JcizhG
kwz9axLDVghMopOSl1yPO4frUZnJFSiHbjwNRy7zvQbzwDzbXUSpp6rCBv5ZY2cQ
QrvHlfOoeFTn3w1NL57dp/VNpCQafEcw3Mm5fda/1u8cnVXGDOM+cooJPICF6fQV
YDXLE947OW74Wz4h+f82Grci6Dd/xkbZZ/v7RSnwK5m3kk8cXKf3ezbRioS22jP/
cFuKhp26MoP1XbBCNZk2NX/GkWoiwqq7D7n1nxkW/CG9cC6Cshl2BNOASCWqe2xq
fXstQuRGdi+lcxLeHU61xDfXdblJudUr6XFUQVT/rAUUkTh/+gUkBbme+yJ9145z
FpDZJXnydqDUePdTb4e9LBhn3srWGay/AY/7J4X21imJyW6uc8S4FsHC2LM6M9g/
6h7ZHV5lCCGUWU575VLqsbU1RG6XjjrI1pnGE2N6Otb09QEzYi0+Z+j85YSfIt1h
0cBvNj/GHhwUp9HqweZmGlLeh6Oc6HlbZbyrh3mjineIN6lFvputf63xCUPBjDxg
G7L67zBwTT1/rwffkqtKVhlFSXucA6Gf4uCVcxWi7Pt4aCRZWwjX4SNDoUbb52VC
GVT3tg/EX3TlgBzFp9uNpQjYrCtfLd5ZNRvM0rwyFOnhXOZ7cpPh+lVE73cuWlND
0pZOY1KLBAwNGTvB7+X4xPWUa4zkHVkJ2+jlQMpKKKTTIkiWqHZmrdghBr5JBHww
OtBsKoqcA0QBRh521Qd34XAp/n+6RCRSYu5jRQ9jHzjsEaeaQuTK8a7NjqN5wTSs
OyzOhuX/zMbftiPM06ENYVV7SH/B7nmPckghCl7Ty0Nu6SI7HsMrsVsp27qN4Lds
Q7BE+gfnzVYIUWcriiUxN4w7d3BeSDms0scL/u1Iv7FwTP8j9RF7fScG2ARAgnOl
gLuwQe1/gLl/bqhNPna/3O5A/0fkoeOTZHS7NUfXr7r/LvOui/VKdsxijzlIPlD0
yuP3ZNLgc+BYCd2s0nSWuX9H1XjogdQ3zoSMkjM4oVZTAeSgCPYh1JC7Tpeph7fH
uoaDESaKgd14RrRANSmXHNOudYOj1SSUSbSOLmekIF1NPKagza5KxQV7/lBJirDJ
7pnibrkDI6Qkh50Im1sczMJVL3u3X+KEPjX7B4qMweVkURJCSIr8HdWKdcuwYSGJ
taVfkPyDJUa51aZBvC3iLt/V8UBj4kv1tHhTh7PJarJuR1MX2MvY0JSeiARtm1z9
s8FWqKBNuF2LmrQBh5CIyKp7F17FV8NvYSghf1BSpf44f/IJhmV8GLH9FH18ziiL
w14jMd6QTXgmRBlpOr3BTQ2eOUH8IWKvlS9RZYV5Go+KfmvFDqGHZVf7x6lWsNRU
5Z2bUS++yGTDfzCvJyQ66aEVSDNExbjvp7rX2BrVAJwZSXDuVjaV3XVWYgdRJ9zF
r3if6Zn+CvgS3hspWQ4RB12F7zs2ExFWwgvH3u+i6c5oe6GDRMMWNG4udsV0nO6Y
HUp3ur7SLEPLX9r/tRvfhdSTm1eMKT37XdloAtpSZf1+v6SdirmVtNAmMOm0jiZ9
COEmOZsuHfVlLdgqtUKZ7egnep88EYL2ni8Bbxkl6ZbXA0pqJ/eNLuK6OHz98gIc
+e9/xU3IzGxPnhnOOCQnnQhQmBjnINr2pX3+C7GoY/ZLJW4b5skXlGXq2iHJVXIV
iW+J5+f9VtNHf4BBdpeyYilif6mo9nYrRYmyrhV3JM32Rl5hyriGqsj57jj0Z2Cn
8Tfyedu56SPT0RuHgh+UPrP6bOJlMYQssNwOY3xD/X2bxa6n/zYfF3P+BjGDgg8i
fY4XFS92xXgxLzOQH2KJGtETi5vfoRgkkt2ekAmsRSp2n/mSJ+os6gNhXH6OFGcg
fgOJBnIfck1eoCjRa8wXNHubsY21c3XNZmrVigoulxx5/3NN9iZFoyyuzhrJN5Mp
Tu24RxCgFu6SNlce1wSFCs7wuQFlyCUBZA4IvZvsd3E2GC9NwBs1Nw//x3rN/KDU
CNd/0LE2hC3y8Yp1QpGMGRvt/v4JaZoCfSO+FKXH+zJWcxvjmCLGjS/BUie/HyEj
vORjxVyC8i3H5EOxl3PlrVLk5jWyhLQ77F8aPRSLxQLTxb9KSgwrFXO/DmnKCmNu
LE6DFM2PfOnDnSaObzLfkJf2YvMSLhkqHwkofBskz5vK2ZUY+fHG0ruhZdCHxoM1
tMKkHBqfohn2W85gWtdlZJcgHxH1aZqqpCaxmk7oNI138pLSnyOji2H4fKs5WS5t
dNlv1e/qQF0AvqPhvfNdBNSYQN/aK/KZ3xuqkjYCyaaYNnAoWSZyY5vQWy1pJIx6
lp9Uzk1qkH5yh5Ilg7R/JPi3d8/l4emeGQ1JnTrYE7i+BNXAVyiXJLRS883ou7Hd
3xGhE9UIjgjSJFuKa029GF5BTWhBfmpf3+P6WgsgMdv2AywozCJBcaMkPwx518Ls
DhI8AHU7M7kX58GMWfTDqQal9mb2TigenKOJLTh7P699pZzz2vZsl1Lx/bySb4ai
ECtvZ09qWLtY8RLaM+sM2pu2cGOVoyk68fpxcNHNf93aQhsUGhmDoz0ecc+vo15+
eqUA8uqvRv5F2EHIxYFF2siypnZcUcYXfbcWKr4rcQtdvCUet0JJfLmqcnnrDMXe
NOlVtSWsSYkvfltTr1Rj/AgHP7ViskHCjRG3i5IXVNMEkGpBADjEo48mgBSXpDXH
eruM24GARrLp7q5pH+Buhq3T63zThJd5TE/wlG4upsgn0Ycjuz88uLqXjW9lIAh/
7Fw6CkhvBMp5HjxMX2KKpkMGnlBrNJSNZVLwhXc14j2VmCiWPD1duuoCs9Xof3XI
V7dN71lAbFQj42ZLxabSIXCmNwcHrQ7ugB5kzzJVoorpJ3npM4xfoMAZ+wNKLfYI
gG+sXLjXwbo4/IKXdU2uWrI8bs+xrnU6UGb0IdS8EUJL/UJnhW2l0m4eXd3TGqk+
rcghs8YS5CWDod7pw7QO5y3op11A3VWsT02zwbLYzUnXCK5cHvw1GA5+XPGGXcP6
cwmyigW2CnQIHTo0/iO0FmR7y89nyehzm7ADiNDXrtXQ2ZGD423xY2grS5W6f8gZ
UGiEwTzxmfUSJGckJh7SdJzIAGgGM9fls5zOrn9iWxcPv2Zh1eta8qsstQl5b3MX
lEzhvtRf0q+Z5ZvE1dTOiNHLg7nZ/OQoW1CXjhjMFULevi70n8y4KcC1jHLvrkS7
NwrYr3AgGGIVf+/HkhgYEMpJLPF3IBZfbjRmObjrjcWfO3QhBXL1lEMEAwg1NrSD
yIZfPklYJcN9JX+WqXn+w3JHS57tNSUk/K6743QnBiaCRbOHnJ++y7eYIEOuNgsG
kwMCHAOlX37tB2j0S3Gb0Q2njTKfjndb8/BPevdZjtf6MpHpsG1HZNfDcAjwgmSx
eCIF2XdtJE3X6mMW9LI9K+DCMFHVIFvuBs3mANlPL4a2Pf85C6w0Ruuwp0QP/VKB
Vgfyi8dd/9pBetgndelBTMfH/Nu2gy17Og2kMz5ySutbryxZBfKzSBbJWUw7JEkM
xWzJyng6Ed3V9sJHK6tJ1fREau1MVKjgAgVD7gEcXaR2D+8yNBhx0jqoaEbbSuX5
Qu+RzjPxgUjPVIMBN+f0aeB8Olmi1Yeq66l870+BepJRjuAOWb72dmkySDJROgAB
QDGcWWFYsW5b1O43JgzJ1p5Qqjs0hN+6yybfZDVV75XHjY86qDeUfjxIik8iypEE
cLUnwV1tw1a6wFXBoHomME3g0RWTndvHu0cRSCZInAKrONFpG7QLn3wgnZbB5KnM
UlRPqHxBzUHtZI1O5iv5pByDjAjH9/gUeZh6sFPa8/urZAW6xIN6ksun0R3uHXBP
QIfOKY7/A6RUKFC53ASddXIrN2dbocDcDUxh6GvHhJ4aE3YxUzmHRnTzClGGAAG+
w8O7SwP3Zh1L+S8aOrkHwyN2He+GXBTRl2ChgHDSvbXHQIaxb9/8kvrXn089txQ+
Z6prWTL5++rv0zTnwLsmdER462L6EVx/Jd7Tgf0Z2TlGYmzcJmvCXyWqHJADr+lh
0+SKxc31UVYFJN7jlEPdBSVr6rBsP6Y/m5hOmo4zmXoQXnikFdKlLmcnTZsj5JKd
AFwnoS0JFi9+K14N/qpm0B8xuEE24cUa62Rymhux8zhBw3azk0cSuuSGwcUIPQzz
1bljxcGj3YGaMEyeaX3aj8j0a/bt3JHr0LLDFrVkEyJvZsoDoqhn7PNjrHx+EogZ
Q0d1CMuWmrT4TeWFvCekwNyO62mCWk+wNy90yJWd16cXYA3TBHozmodq2Tk9s0gH
tMKJ90zTwuQSYXgCrKIclzkg0YO5bophwD/RZIhgIspLV+LX8D0KUKmbol/Um1Fa
l3EBxgt4GEQsA13Pd0FBYPmXBUCMTDQsg29XHdnXDFpnAMhpO3veanAsUHcqV2Ey
U1sQscmiI2vDkIIyxM74pWWQ2tWmCzxmK3OPcregt/B1EqRrWnuIt42NlY87oMY5
kiYmyFk7ExpXm7ixJges0+3j5x7AI8IBCR9/Y8Nxhyhj9ZDILvwlKYntvieLQliO
ENDypC8UJpVRrxCCwnJWsAgMPng0HdwrWDsndQpzLPFPdaEBYMpYWLmQfJhHSG+s
+bzRyIVQcYyAJZJAf6RpubViKW+0CogruIqZ4mOgYS2AiQgXMiD/vWTBwIAwQBqE
sefhJH3AJrLVxPbVAlCRf7kZKzfP86KJ85R45AnonjhQrH35TAqz8Y/yDdl5e9WK
wxodvsLVYTc62vkLTIwwWHMN78vBEc3YaZXBxT7ZI0Z3FUt9tyrRYoyvRBFVp6SU
bfvvqxurUDG9/ONCsdsI+g2njX2ELfgNGQwkpmzM0kMprka6rOliDbgOSgIkNZYK
XmwS4vzMmLNmGTaj3parI+kB4KcajPuKL846y4ayUPMypeVu5gEAU0y6Ob6C0aBw
DxZUYpp9d1dl5VeVGZPUa1FFmT8AQelO6bTPYP6ClqX2taIsjfiiX4D8sMVutQaQ
TsA8Q5U/QrukpHkm4jAqrqPzgaP83tOVxP6YkvjFcmd9klWwiy/0EOOy87LfgIzm
Wg31Z/yMegOMI9iiNTDS2rFLMi7jVZe/5ibflxa0uClbpQ3nHBkea9J7kjatrw7s
YntKwZe/P2nZBn4bhjunhHsKymgCrwitlOlIls5KZfNcJm2as2RwWN+Q9D5e4FZ+
d638mw/4h/xEqlKD+tzz7YZCgrDaeXBbBMFi5of39RL2qDxi4qDQsS+yDppJG9QK
EIrS7jrvYuN+ZkY/rNZXzugbNK80r5Ul58BHGNDwSRXpGt8XEjZWT881OVeOcYHR
mma4CHhvx1sqFcjMRQJZ6xnQAJgZEWcDhE0GdDVQAgnPD3MRiLwm+O1ku/jLQl0f
Hp8fvUOKnkFhiukv+cDTr3qxFBdFjeETYj0scZ0SuloHFuV8LF79nad5hKEtWQNe
EbfsuHQ00nnBOSYcbfK3bcWaGDVsk9W9gbqrzfXSxRprv/LEY2An7sUUBcnhFQ8n
gxRY3fK9j6t7upjo5De9BJvpLEFSkZxG0lk0J9w/N9LYsLZnAf7HSNDz5dBMVuNd
0ZQHO68mcjQRsT3SpGpW3d2UlQDJ/TqqG/cKLot4EDmhIPTx+36q/YyvDb7Zy+kR
GbSN/L+vMmXeMc9LYyZXMhUgQp4JR0JPAHa/w315t+XsLG2rBqykO0Q9+fzuTEYP
bhg/N8WxKTEYpncn9IXIXQyK9jho8pgACNBnB5X+9w2mJno1fbDhDY+TZ/vlvIDX
Z8bH0Cs1a0KUWDaYsRqFlZ+8FF20mhCeyyCmOs7Ql2R2ReBV43zWMghYAobKRxc6
yHfXRULLmPSdQcBhiWnAeoH/2NlshuMXCp4zIUZG9I/vyefvmgMAxLcjzpneyDfw
Zssv9GL9ZseAnx9tW3xeKpo/UxPa/J8fPqaFaVslN0xFg/NTEV5Y7aF4S7uCpxhg
uI1vfQI/SxUUTIRpyWgArmepJey8k4DizI4OJ2VyR5QGB+8d6JZWnKmkGHdR0jUB
Xyl4lv1t7gvC6QCLGSOOPMhVVxvVQONk3RL0lSx75X578auvhqY1gLiexbGXChao
1dQiaDsA4sw3ZIp1tH8uSsJUVTTck0s8tBqtv8lso1BQVcemSpiAoxYVVO+O/7Ag
QIkMLpvWoN9YKG3cv2XvN70zv8Ig7WBDsZE7O0LVGHqGOSuJ99D8Slj+oLyytWMT
CnwYuApd768qggD5mV1+pUBWezVIgItiyNtwV6C/2AHwfgl/qQuiBof3Vj+ccpcw
e3rXIGgobo7DHGD1LZPOYl9A/BTRoYXZjnqugE6r5t+fO4fHda6AeAsTwbgZXLkU
pUGt9QVdkl9rln3W4JuQUIB1UQMYMyZR1Cet6hOB1yJfdbDYu8w5WLI2/cwHIzai
sU6ikjHZp38ESD9p+HRWf2yzWgsRn7Djk3utGWxVYCk1ylRESgxNbijhxQ49uKtT
Gbn7svkt+VHsywAKjb3zJQ4KZxmVTZ+yFlr539XaPZk5CFKoGwnGxjUqYZ7zPcz4
Y5WBfGgXkS30et6skJuJcsWwV+YlXinhuRIrXfC+cOCXAoiU0JbHWmWd+XXk8iOn
QrxOwAkevWpam4cSjVpI3xnQDSuKXh+wVdrZ67+lIkauODyZhzA6i6jNldbFfCBr
nIJG6Bk0W412Y8zcEiPrVTRlkVm1hDmj5+sTCm7qvghBbNWPhMszY7cVkjqFuphu
qOy7DiumaU0peirJzyyMPviPMHqagqs3nzVZLPnoV4MDjrJxo9KAI6Dx/6IVqpHI
XMKCTht4r1JR+9CWAXo78gmDsBaB4R2dFYCeb4aLObw5yP0hA8spOa5CnBySY0kF
KRELyvB9v86ggkY0hLlJpvRyMjk2f/LDcK1y83AlAEdLqIBNah2xbI0OIowX1cP5
1D46yQ+EWBoqSD3hGIfx9fjaItsVsjBEqsPSnnVPzLCQfin/GwlPbNogSL0xEgzE
3Q5szoR7NRk8Yh5dOy8WOxx/Pa+KNwogyROYvUAhwyfb6SHP1EIVYnVUpnp8SPR0
BeitIEd3+j/1jMdMPr+R/60jf60QxHmjqZXqDXxm6qCaDO1e7oJIOdCyVxQzefWY
vB8E7Ayxp3ewIGAsVoBZdX6Ujb1IOPqYltLI/ssmykZsHLkatr1URc5nr7LmpWIX
o7bhhexLCGwwt0svzp0KEBPnGOsrWgtserGznz6gIjVsPdPCqexw+ucOnPP1JXhN
uX1N2X8lrsgXCN2/NJMqVVbA59k/A7DqKl7aC9vn7Guy21ThsCvRJVlA1Nh19CM7
BJTaKojjw0zDrMlMNsgfm1Oupa6+BFyX332JhZSqQ6fALWMNOoIviub3+9hPTca4
V+H3Bc+NX4jQZ+jjFXt061Zk61C0wdtls/KZOdpmN/MHbEwuKHQXThf6V+RYJVWn
ILJcUSYMyeTMLwDEiC8kVEVLVGjHBxt67/TuyK7p6fFgTcL36w3AAY88ahBVWa8e
ul6aKlzrPb5KYDKku6ekoAJ2dq0OJAsRoHICyoZ7xexuXyifGt+hbRXhmc9d87v4
8rlfYDl+tpI+OKaMaiHJ0E6UUmi/eMdos1WAWoAatpiEOcvjS7l+OnJ7Gm2JhF9s
J8QGF8PxWViAQtPGZx6phQtzqJb/3gWOhGm/5MbaPjvpxXsqvbab0mZEmZlMCNkT
C87I+tharv0NZEi6JJrUy510Cm6mUXtjks91rjmSk29HlW014L6W0p46dtJrNWgx
bzhGESKPH4HhUJo8/2C6mY8407RhenhfkYdLGhHWxX4lQpzABnXIJaYbv49LwAuq
KvE7TW/IEFRIjAu4PS25UEGK/iuUllesDurmukIRhMF5VpR8fQB3rgF2wBJ0f1do
4pfs18k7O1n1slxotkLI3Y+vEjC3u2aWUALf5rMPC2m1OTdYQ3F7WpJZ+eUKKxwo
v+BjgG/JVanQ3sm7yI0kW5hzAjSPxOmQ8loVErclnlsUjI6ju4XjxafETeTCHYeL
Teum//7SZTX4QAb7Yp0uffKUtjXBG8I3dQmZ4PKmrECY6U4h9bMdhXja9ZjsleW4
AS3FNVb89fbZJRStnvegAKBMGwqAudRvSwAWEpgdRO49q8zgZQMyoEUlJdKOJ5yC
o562NxFoKFoTBkpwfVMq3MoAeSI+m/CsTHq3SRBC4FmhsjXyh5eRp2pqBxdRqNsv
luobVdLnf/JDpknJhtYc5dRoVNkHdQS3esjsnrhbABeO4N/R0xgSrkqGSgo3qfXS
cKwg9cMHgKoN35AHZN9VQbeFzhUbV3aI7GxeFEq9Bf/GfvA4tqPlu60lnG6nbhA4
TjCf7oTbA8hd91FvaIp05enTRjPDyzviFTuBwwH6e3MWoiPUebNIym8c2wsnNbGe
4nL/r2Ytd2BZb6SEXTLGOgYN8e4TZrWATOTdCuoxjs1kmE0S4kJdsIvmx+c9byIB
/f/LEqE+pE2ClO2xJUj2HB3BUIy0kOdGKbXJWKXHLyg0vTuu9PpAdwPOyr6QkCxb
LT1ODGEBjxCwwu09DQ0DqwqAm4Jnwjp8v89lirG80DIPw+yz9gR42FkOQH6MlMev
OZiJce1bMzJMB1wCqkHLEybZDJwqJlUV5kV+BflWHKpe+FBf8VRyJmfwIIFZt3Um
r9xaA9LoRS2zmRMA7YgkIkg58S9FYjzElB1CNIGF34dL3+v9xVSSZrJgpku7iezs
4FI9BI7i5YJDpjoA3nz0DZ8dP4FNy9wBMDxyJANX9BxWeW8gILVFDmf0lR4O8KD+
OjrK5nHj5QieAM2vcqwz7M2Y79ZdbDpMxNI2+Hb4mm7QNPP2BA4H89Zx/rglus89
eq0004fz34OkTHHvR/2WyYTKGXKZwMcDO7ApjrnBcHyYdBII4JtkuQ4NJDYHdHrJ
3gmjaRK01rTz/UaVFIUzXu1I3udHZXSVEqRzXT1o0NZHFrTICjamwnTgpb09rz8q
XmxFl8psBPpBP6vONxOL7WQKXlNW1hHJ7RwqaCRr9USd4mKxZ0ZRXmdBNsuWXAZ+
M6UqVnMTUs/FWegoORG3vr0kg7gBs6HifhZogyTfVqVPb43QiWBL0tqYOZPUKEsM
Zn+ggrG0YdRU/nelnwSFiQ27lie8dTZYiFGvXW3266kQ4yuYweHFg3QaMMtXbEmZ
3mxilK+MbOmIgTQzYXzK6fpUj36px1xNClp+PJa9/DAA5At+xSVYaRuvmNS/kIC3
a5ZSl/DDVJG+FoNPyQCpzh5UVPDkQcYa4xocqWqFAtk17N1UPk+nmZX3BJ/IDG2h
mQ1wSgdvgOLlS6r1fthJ4SyMKsiaMnDUGqZkP067ZT/ifNPNw+j/7vkU+YTtZWEJ
L4ZazZ9UF6ZMGa1xqAv2glJ3PFqLezesizrMmnWfYBqnGFfE2ClEAleu3VVxTb07
ifu87zJ2IciXi3kZe6tYkKYd/xyTHEN984V3lg7QdGFCBHmLKiWESjz+d1DQfE3a
ahWnwbEJiLgW1VJGwlq5HAQEDZkRAd4e4b2F+3tVHaq68mpXuYVBvYLdWFzHBSYj
0oYtC4vWdqsuP6kFsfUlX+expv9SXhA5/C/Vv9oplioa9vhg0MA0BD8pZQWqrN+p
XZLhbmYK9nl6ZoOk/XL8kNWx0Pl4y+dlbOS3EOxzOcSVv30mk5I/EeNGuofC5bUu
hfe2Fb8mw/l5BN8infGDe8RNilCSZT+02yw22s8jyWh7L38JBeJ+loqay/aCrrOk
DhyQ5y0QnFiT4BqD/ca23IQupWA+qNrw5yQnn5sgyes7zu1gGpdraj9HMKIAsDUi
X8eDyPe2Tfr3H6/W7Vw7xym0lQiAAYCGpLByHn/NyKSvL+WpzpQI2LKzI/+36aH1
MF49kOmHcWS/pjQv+H5/l/owtT+BihAkyqA/hit7J4RQVR96DQv4MGHbV7IH2y/g
bCEPcXq4ADfrVXxise6SV+WuXmrSb5fR31svinl8z5ZLRCD+zjzrl0C8kF/LEsok
9frSuHgsreSqfXCqabxce6uMW3+tu9obSdhPTkNMIPQrVqOqBzXVrIkbJw7/jfXz
L0wj4n2w9l+rutxdPB8UqgScAYsoU8deKcrlPZ00Z3VUYtelrwvNuBlxeOAUzx4j
LuchhR0kgaB94I+ypT/v/6cip5XUzeFbnWsLOkTrzeALKPMIJmBuSz1035pHK9vK
G+UHpxClUxD5G5REvr3qgr/HEmB5+NIASmnfVeElnnl84SuWTfKohYcyPYVrCc5c
U7xl54UXJoYSO2lNEbtG2OovfT46MCX/bhPpbSeZ4asCu7heVPVAGd6dX56UnXlQ
yDCG1q3ZlaS1kxAHGKcAroC+PfCl8/a24qj82b69aI2BGLHyG3zXAHAkVm9tXSy7
1t0IYvRfVMX7NkYaXNxnikobhKO+EYMfrYbNtKafAoRClYvSKXGjJn9pIQ8l7Gi8
o7hEdQZKUh9G6AkENlTWuWM10XjQEG0kog6xLrQ0pTxh8gyhqHANMPkHRlEI4ysZ
pGoziw/m+sPiLMwSxscvPPCBdPkNa9dTy1DAkYyukTUKKPAb/eg/AEmBgAaxktCR
eMEPu1YIldGJcfukQcdrs4gmsEN00yInf/LdzZ/s2x4pxGXal4D18U+7UZB2wHLu
8Py2ZPTIztx1Lq1ACEvt6ANRy2kSkb2PsBcwXFzyF+B/J1wO3URIDc0/JuGhZb92
LuGlA/MQNzCCrzlO8IawVw1PERIzgRVqpVg8mk6wfc06+z5XeOGHbvMUXguEJSez
8DM9QGoU1YxDkYpTgyanlUF2xq27lyDc1E0oaes97+wBXC4gy1RV1U6d2E4aN/CO
U+QaPXr3HiZVDgzqKMODmowvDiYGsVISQ0OxpC5g+XWYDSAFlukcAVP/RFJrJZXL
55Hecq+7FSORXYcGkC7MCIRNCqpdLtN2FbIikQNE3oh4dOuUWvvg59KMvjhrx9Qr
XoQWCf4lpnoTIef1hJUe4NQYR0hZpdIPrdKQdrgTIvjOwvveNG+goA27MlY0LJZy
CjRFyjIkOK82Q0e9amFpv9vqmyJWEa1RniIpbsdCeNM/qtFEcvZuNbwEEcJ01TnC
Emfq4Xw6RmfgepGgJPt8FYJM6JAoQrfrTTiB8sKqi1H5k/MATTHgI6Ug0FgODhIk
nokIGDs+CRMH29leIo375ls3Q8SSKHbSXKisExOqSLi64hEJDR0zptp9csMfWR98
AQqsPqoEnTBeFy25QCJx/vn1qeUL+h6nx7nkc+plmK0Q/l/DpZHyMf665SCrS79f
4urUZTyIByr06hkqEXqWMW2y+MJt2CyvgGSlUi/8PDQIaTRiz2dFiCc4RrVxbR+t
PYWbFwK4fFQKi1nKNcapQf/QlpiG5TGhacyyxKmYCgTnUCvsSlSS6UZlOwYU+ctY
L9OHySIzKIt8Whe8jb7+390CM4bO3DkziSPeKSS/1RAT+tIv310n3GRWWHTkbszz
skt4Vq8Z82qEXa/6uKP6JrMjfRpU41oaLuCiJKqPwx81EIPQbZ69hEXTRE0Y/j5S
orbxZgYTARUAJHjdWN7SUxNMSAXT0PwjVCYl9QpnMMOVR80T4USCICXWuVJuN2AZ
PYQ/sSDGGuwNcvRRGHuPWya+T6mKf+2/wtTmCc+aZeTaDAc/6waYl1MMddC7tzP5
nz+tdwn1S+NWn1yw2Oz9zWge2BrNwV665MhpB0dUw1LM3rQrsJWbuMhCRZeSsCZC
1li3MMahXm5KRjJv9dciFJkW7EhLTt6QFIP32u3HBpbGaH9Tef0EAEFaszdJgUqD
BgJ9JzaYSjPZXyvj9abryA47ZZq6VRtXVJQrVPJmagBur7+SoZrVHopMJwjPopxU
wJDjTO8P//uv/Q6MJxAPjQ==

`pragma protect end_protected

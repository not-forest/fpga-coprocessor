`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
T+Hiz0YeaRZEI8ZRNqFGX0tIYyvdccMfGwbMPsmKTxo3BbqeOgiqhW8/iyqar/lp
XZ5DxfY1DUMt8B3t6Tv/uFPTN+QJTl+F/4qPM7/gGtY6KAfyOjCqeSecjp+tFip5
3wGaScXnLgSCUktHYpsz3W/Cj5oxcNUSgJW4S6AeGqw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7120)
gSHOWA1c2ivHhTxgmViuftcgX0ozRmNVYN6QyIjHh0GI4Zp/GbNS0i9MgbpI1ApF
3AwWqeyHDUMpCEQEJeLasjrhSVTuemdGDoYPz6TLp0hDWWXukidmJWCS59OuPLv3
PI72bWGKhmhkYStqf1p3Bf0rkqtHZ4RgdrGSIH33MiRrRoC+OCRfOTHx7NBGU7z+
bR8/S0DwYnTvwboUJmuFhTFvI53bnYXimXv8dekDoB+0WaXHFBSU0mWokhsierL6
PO4x4SswRTeF6QWpRXeUItiGdEypBy90MdfZh6kuR1o0yaxJ0u8lp2dUNk6uQRMa
nyXdyPnXEmJQz5JaLrwxyACnenl7RXmoB1CTKLaEMsCUyho82DYKsT9Psqya6m88
LnzgbXKS/LBTEzt8oURW6OHNVwTrwtWClkLpccK5fPhInlOSerptQlTa6FTo/HhE
DnLv2pdRh9cqYMnDbQeSATNHMaW7ge40hQ8O/aJExE8fnsO7rgFlB92CnQA0SIid
heILy2cndyoqTsZVV0n0XGQtZFRRMazNHG0DmbS4Vze5djwqSOMLWpa9OAFnD2AZ
HdrP33eUBPAJUwstItilEC/g5JPCEf2a+eqPVSv6/WjbopBIQNSWOfsvafT4eTtu
d2qYVvbbHPPN6TYgvHTv6III+uSzBbdrAGO1B4y+G+vsrGBt5nZdb5c8Ecy6/KkB
2qyEB2urfH2zqWVehWhoOMbs08+empg7Sl0BcAdy1wJgTGiOgIe64FtJVl6IdE92
Xqw5XVYojfzBP/kaKjVC3xbpAAO7OWwQ+iCsfa+Nb/vxwMKaC6jyOGgZjF+UvGzu
M6ygZKJCy7DMWuXkCS6xPKTvYfNB0ucqKQN2GjC/KSuHBuAURe0ZRNjIlceSUu9M
1HAgJxsOdhifpQWsPVgN/I4IYK1NjBt4raDYuy8Y1PjdaWGvWnxWAVPfhrCJhZJY
hUZicbLKjoanGjpSghJ+Ctl9TNqXwXU34/dVw+Vr7hyRlPA/dA0i4dEua39km8pN
nPlg6EVvFMLPnVT3ZPHqdPSaM14s4xyLQHMvIJGeHFiaLmYolvqLnA1ndQAf5OcH
BTMyqlnjnzaAVhWTmMh/L0mTqWVRoGv8CVToDDNl5LjIb3SxCNtBEMNtnYZLEvPJ
lBeWJIecfgbLPUR04K3TCiF7XG1XemA2+xGfoW0/6wk0JP/UMSiwRY8D0juvN7nW
ICY54xGWqWoPK7eN0+FSTaamWmIlO7jGUj4qEunWYAXnD3Mik5g9bPhhTWyvIPjg
aKW1UWAqL3B0AhUiZQi6quNpknzzumwZ0HWEehs5jGxs9zaMtsOZFjM8q+ZiuIbv
LAFKMKoO/oG/h4gj/CQ6QWf+1kLwoIRM+Jvt4BZC/qavBU9lQmNROjXbJp4Sp36A
W0UiMINydyCEDndg9+yEiWboEu89lnT52SpZsQCXGW6FnuY4R4JTtjFvFURhavWg
MDKIMWV+Eaim+liLnQcZGj4/mEiy0S29YeXKmfXFkZnkQJqo2vilQCiRKz+cNarH
zqft+r0I0J0V29Mh6nd7kWW89uz1NhBNNktr8h9wQXRi2+rEBC0Fdhy3kkyKyD6b
b2rTRnHb/D97Xijq9fVxtkXRSpZIjgOMiPNwidmCHLBS75Nn/9QKBTRkbzoM/kJY
Aun7XbaWbzm0dTmftSNIRgXjF/6RR7GFUDhdNQO6uhQCDNcRbFNV36y5wM/qrYlc
FLLz3BhQv1hLLFG85xZNAXyS3XxScw1yTL5mTjzDj9le7QCNlcjo+RzTgDpHZCv1
QsBOHefvYpGcG6zq29AnalhuQpMP+Ig6Vz1CHRLVPtBldYNevkns10uftvf2iPZg
p8KYtsmf/73yycfTR9CbPmMrxO6lizEcEqi6wLAWymtaKqlqzpECikAUG15tS0B0
fCwoedx8wDnOS2p2yLGwITGXY4D5XcZprKmT9fUA283QxYVhp9B6GNEdKRsCYKYu
JoCrdIT9bonjgHh+oUUdk0OumYDlgf5xvhsUEEIFFDKODj4ryAmlzFHEelOJlrMT
9qiSAhK8aF66xN7yeQl9cMvPX+/b2pgXlTAxmFRxfpUR233EAFE7ZRPkv1z9teDq
OeaZ3dYYmS7IqtYvpV5O3ZpWV9+MniONtZr8hH5bx94UsBgd43azl7BLnPr0LMqk
ZQPHzRGqcxfvLGLTafJVExy+UuD0kTrq5DG11paQ5aYCdZHpl+sgJLxRnq5mkrLd
QJ/kn73o4Tb0tmwa6zHAWpy3tXZwOR/m1+mV8lGxScSP6rYMxc+xCKUQ56QAqG+b
ybCsqvDbPw/T4WXPHv3LW6XKTfM7gvfcPg/sa0QbObhaPTqmBPU7VZnyGKDgk16E
l4wsWtpcGgPj031UP34u92y08mAdHOdyxpZe7b2ArahYHZDcdzZZpmYkj+ACooO8
99fM/WZDEcgArEdzsM7J0xVGN9btj8MPY2J1oDAyv4bHOzY8E7cphd4p5VbW5enT
UWZ1jPVf6XkVQe1mid0wjw736FaD/oCUa+BVclayJA2DYq7jTYBmDJJVBIvtQN34
Q3/QPNxosWGo+GRFDBhbnYQTZj/ZwWL3KrlCCMB79bdDOq9P11c1lPYZSg9NfpkQ
IlWksb4B9N6LqkI26FvOb3/KNmHIDgEvq1YHH4mXD34Wqg8VWZrJ/2u90XS7MLUf
C1hFrsr+V2JaOUt/zZ61ULF7AJ6f+gxs3qMmLNfiYy9fXxv8LAW0D0ZofL21jzEg
0oaJ8tmPxeKOy+oiOwmkm9xuFvZDVEYZKsm+12JkDC2/LDFsfHdkMbmXiJWX5thv
ADndDGObRGWVHAkybaxcEYAYjA9EhlPogghkqg7WPo5VI70a391VBjHKcnF7qQdY
DARswFn+TDpuRkA7cb4sO8Jv110GcxIo8NQ1mj+G6hJL44Sl40NtrMNdm1D+Ii+9
g85kdXPwdWy4MK7njDWcgtiJB8LgL9B87ghWhMGyD9PESAG2crPYE9W5fsy3QzHk
WZ0GrOOC57snL9uGLoXbEixJd5Q7AoifeBZzs5CfSUqc8FDqgHqT/tWeFpvDQmTF
v2CJjJQuLqcguHd0ISY3HGVTPIkVxlnG7DfTXfbKLrSOu6AneL7QkbGpVzh+AdJS
1P1shYDBOA5svW7RuDMCsEDXJ6ioqfXjd9ywiMrbySy/MoElZHVqKFmA4jsIezGU
JVI7HYEp2G6oWKndfJqifQ3SHEoymXoRbFYQo4qfJC0j0e0gqeDdtYE19BkZqYHb
lF0rlVGHEWB2dDTYUpux9oCJfNxsfbQLzUTL3rf9WMo83yXO5kW/N2iQzkz5ZD8o
9ZOCuV1jiSYDLBl6teE3Ck2pSPLpte7gKhuyW+4Qs5fb0j0eRJJz04qBq96S9lR6
3pi6ltATugXmoRC3Ej/P0Fg2ddSBZW6RAi4qZ//8OT9dQjEZiWb/S8Dh8yhxzWwr
237/q71NYUb5taLj1ly8y7XpNe7UOovzDhXcr+qXhc4cUaAjbfaMlR2EgUBH6nGv
0ONW2h4xHiJFtqtqP6Z1jyRprlEJS/vr7zSB6wqERmTABo2Ihe1DdJSN1PsWaWnd
5T1/mli9YU1crcdOBJr9xQB+WjPdupkWw2I8dZSv906qNgI+VM/4Hquw/XiFxHsf
tY9BwBJfsKEHZaZhoqOkrc/nm5JOoHqn3ZJgARw6aGiEPclPv2EVT+w21J2no0uB
D9PrI/lV5lcLB8NWoCJlH7OAc34Fgbs2SdRuEBSCT0Y5vO/KzD+5Jp4J8TGPxbxY
WsGx5AVmWNw63MQgN8tZ+52snyEYpVzjEvTJeon52Zcm3adZHFsU4BjtmeMKQBvf
apQ0sSyqCGFOiPCfXVgL4AXCs3yX4k/nDV3hUQ1ANHLNUPlE3X0LrDVzvdt+UvNF
i/+JKvGvD6vSEEDtNTW9uxw8g/bchvZ2UabIObx8HAYnsS+GwgRA6etJ2lKK9eir
BF8R13RMg+fpqaKF/45wlXKpKW+vRkeWCIYDC0KVUrIWdQm2BOlX4GIbhO4B+tsN
rOS9wJDRg/0tOI/LjmKEyqOMKmDCw7Y1Zak8mllmwdtnrCfr9hCZf/qxBG5CZUf5
1u77aUwDQOBMRa6bngCt/krpKKo7LRXxZeizdp4qb2PXZX+F5xly5pDknUocFspf
5YERAvVCOVett12iFRWMFf0nyYB0LjaZ12UmEyLZ52TDWRoV1urr9qVwCe7AktLF
8TIqamhEVGdKMUPGVk5A1XuzxY1Doh0+oEQ6KRswT/NssTMGDGzT8G6itUbZ92vi
7vflNBBSipUha1oNbYy2hq46XWPsKY8fULPJ3jNSFkjHwG3LZnA0SDyYQhww1MG1
pR4A7WLYulJmoNwY93ijeueqU2Yqb4KJtogTgUAM7sv0tFjOcYCMq4x7tTw7Eq4p
HVxBD00wOShZoMeX1KSzMPWe2MZCRaEDmriPTEDfnMpWhlZcEDvQxbpleKEWtrsW
Bwe0zZMxh9Pj4g8r6y21w5vxtmo/uM9nzsTGqHd8ntYtdENmJqNYsLEpwa+HH6bZ
6Is3PUzty/odGPNE2v/DHTaDYcdCY7NYHtTlcNfNdTIaDIp9H3ncOxMhXh52cCNM
8xb3bN76Vtb2N/BJyUDRCi/9ij0mXlAtF/nyY37uMb1inoMQiTwMr2YZzoAyJlGQ
Dt57yv5FFiWTWLxzdRUN7wihCAcw0Ci7crazoRCx2Ius7XsQyd7sGK1chnbr2AN2
fRcjWiLZqLL8VZ6rmCNu9ujO6/riI3HDzhW9yzHntjvwMYP0C+9CAQphjdz/deWv
9NYT8gV2M+KIEzOwFf6VMUlsYq+KLpiTwsLBgVx/8Toza0LkJFfYXQj4yjUUAa/d
RGJ11Rbg16yvNVpXql4/yjFXqbrwLBvwMLd0KUjbtft1fXGZ7cSgvLxcfOgR8xbm
zeV5IOEUu3jc9cBY9op90Z1ZYKwZyFNkvyImA93CJVSW8CNX8BZxWQ7I3M6liPFe
UX+CH4Cb/Bnz1vztCfO/cg7Er9gSh1fiaoQXi+74UA3eEI4VEKwIIDfGQZ2U6lw7
dN/yz+aKgRxQYm5cfTaFzFQMeTO7oRySAJS7RE01bxCVZ8SFX4bsCKwhmb+ZCZI1
jJf/Dt/2lk/QtnsH2akWo5bby36C2xE+WTGsYWSgDt0cTYGGzv6/X09LP5I4CVoG
nLZfaX1Ys+yzaMd1f59nwZQMnJyJ7Uc1I5r3lvj04qC+I4hbysIv/rq+/j3IIQDJ
fIJR4MAtsRm0mZv5cY0vsE5TomqeoCqs+XCbCZwZharCgW/2o8yo3KEYBxQRM7U4
outP5koWGvHDqZjEy+NfhKrmC75yH/kAGT4GrCZ8OsMsq/h3KpUuzAnmSYfL8Qfa
D24vIusSybJ3TjuPegoSdDAejE0v7LCkKogH+6g7K7MB0ULjcTWfinXZTIIcV5lU
eJ6bjeFvU7eiupvzFvGqeowgu0otT1kNV2h/fIX7m3ebX4GXZLjO677wNoKrbtd2
E6JjBP4RPvvIuWDSkathe8Sl0i3exHAp6GzZs7SK9DNiqRHaMyPCR4nJLai1OlHU
4uh4ergPseCgV0tdbCtUBoFRXp0OHCiickTLaBCmBv1dsy4T+L4gnz8G0K2pBWAa
7HOMA7UieUNF8TfEGtjWMOR/qTNu7pe+26BQ3w/OMQVOlFVY+U3RnEHD+dZlqeCg
xzFW350Fpp1zGBWu2F6clKlDTxN/ta1h5+i/+XsKc9Bl5KSAbFHBGDv5rzfic2A5
s90a8NLNAta3oDDCG6oqlwE4ifLi4+deKFJr72Miohc6cMjZyO27RGMquyqHFo+8
LN9XVQlH0hXHAglUP6eCXgz+RrrA4gHfqqRee7Gf4CdcKwBuhJUXpyXRSIiH19Z5
LYrf3pe+Gnn3RHLB5iaGoYsCZn0LvyAR+JzuRzWf88Q4DMRm+EdD/GVmqkyJ6B7R
GzosE4Q/TaL0kjHY1++BcnZ/JABrY6JlE3mUQ/vQ4lsKbAUc/m6kBNC5P85/4Rgk
3wYBjKMHPtFMN5c6cl8q07USjt0qXTZdUScB54LEiVkYI+VjCGMlv3l8A8anRoA6
b5hw4mDXUGQJEUrrvpBQQWnNjQkFqT56EqxU9SBoU1gfkhxsqmsxp7e7RaARNU4p
KuNgS8iMTzsReEmSrns5CC4kgtanjcpcX+tYmao9+BGfiYKEIv87gMD3Zp/o2CQr
vN263blPrEuSCaH0DZiIKjDSjTFQrbQrANbVwYUW9jOScwrB3WryuELYu2I1YFWG
P+sb7d4NcyXJ7zsigcudGLfA2TKZ2tMkFlHixaSKSBDt6EoXTtec8hBx7xPu3M7C
SX9bvDSO33uT5lA2pjhgephWMHIBTOnbBbRMTlox0ud4aUjrotAu/HQr6IvrDsVl
Wq4VjB6+xTCY7FMoLSlz5w7WNySnWeUccv+Mkgls2IeYBTdvxd1Z3/i/N6LKpybe
9mrEoEa6tCzMQ8SC3bLniObGgYzSpyqTZfxgHhNxV2h+1ar6jsqvCmDD2gS8Hygl
VScml9mYEgXiwshtVuGhkDrUGYs5fFu9pdL/TdK4X8aGH3g3imws3BG6+4GeYvuq
3Yot2RXbQbWngJgH3jAdIs7ojFy3RzN1hA9hTLY1SWbM8LWTFwKc2O1whmW5CTmx
4Dw2ibWf77v4bwttc/pcQelTKWidiaJVWFViSM3bBQanmGn82TrCM3X64cr+UKlm
r6tEme4b5mYn5Q3AWYzVwdksLQKrTYmggCADnAp4QMReNLw7+Xmgjc8eVeloe4+9
0k5Wrnwv/tE8JM6Q5KurjVwbYkTJiiibBGU9pSlWOSg9O6rfdZoBom3SPyu97nEm
m8LQn0bDhe4jhetwKxg/4pS2k1TnEFnwt/xhB0eMLjY9TGNk6mA8E2zlG3whqGwr
6uOMWqKhN51MMMAvM98ikGJxZiX+SstUCnmvqxsvA+hcoUpF0mQZrwwYp98nmBaE
SbegCzJAJr8d2II+898XgM0jiYUgc7VtGrDxPvk7xZTR108YiA98vjQCnaBnN+V6
/v7MTfh5Pccy1fRCxPg8udNJQ6BhJs7SXrFzCVYpK1IvXTx9M7r92D4g9NVA2/hy
0iD66I2/pRkz0c1otcHoINQ4s1AGPxWpGDZLVmKaWwWzkyf/IQGMonrr8LUJBz6X
dgqRxmRxh5lr7J1MVCN+s2slWn171hVoIc7OI1Ga7PGAj6KiqaufT+MB1C7ycmNT
l/MKyfsDlCwcSffju7OP+BwxJMKrSa3hbIpN9phZQtyPYEXeEkRzQoYaqNzxRnqA
c7ZcWxoRHHoHPcckgO+my5O5RAEs0mOwPeLjXzRttpg+ASsVdOw0l/gXL61i3wKi
2W4aMzwtXv6yGTxNZk7vCh4LVuDT4he6h2wMAmUwlg8Q0Uvs2GL5ng/mBKm2yztm
X4Oy11v5W1FTkHjzRzaIB2B+FWOWuzQ6Lu3Fbsghvv3wXrbU1oQvsZY+lsrihHnV
7Am8MmG0239vRFH3iK7ko2/uax3jRsACZYC0xYeIaEPSBir7DOrIWlPSWfpet0ml
ZlATbtCKOMtEQnqF4C7unItBy5o7ioOXQQ08hAXYF7TVTpBWJq1hLM0Je1wCFwbr
U6Qr38gXOKt+K1ML4/oGzM/rkmj7j886iTo5AXqmuKJ+R1Bj6ACGObAt441zQicP
U1qw50AgKqJHCxfoM+HkVOO97SIeNtwqQMaXDSMtVfyna1LCL6yjFDg5olsEc3Ld
RR2HIOwyYCXhKjE4k1bhhC2t6Os+TL94yRQoC0hAT+a4QzeXNwyj2FxlgcMgOh56
frmURRlMRr4JPw9WPfT/zb8bfwUPyP1ROVrDAbqqjB50dPVsOSnyCtkIwtI3msZp
M47yajn6SyDb3wof4gPSSV/e72wCC0n7g9ElqE4orTyIg8lztxwKIZMR2K2Rvp7e
nYCqbtRrXdg0SOVHTJchx0Z5m3c6LhnXGUgTpaVjPOc7Ru7eHhmi34iAjoTABIAG
QhpjJmfZ0OK57n/hBouAEX/STEyVLa76jSQAckSIYh81n5cBuZgQpH4QGN3hBTd7
/vNoTQu1Ynu14EBl5O5H6zbGbCCFmptDx9wjVydJlQbB/GhireYT8N5jQJOBN7dj
fwVi/QMS8V1Q0i2+udtEukszb7mbTPOdykbf3MMbvMWiJaGxiljU1hKAkscaHgA1
azs33K24ncX1Xr1bBpTXgWol3THNP8zk6wWHXSoNUdNE1Dib/N9ys34EQDnQknX6
JmrYCjT4i8CT+BhFiGuPKRy55CJDiEZyvVE/tnOPrv16q1jMH1NTlrkwIfJwt80t
SZ0pKIUHsA68VRVjD5odSsptiaF18/F3IttqM1qLaRiZ1VH8l+ptYOFBn3iGuZXe
xh8Y3M9ivLVHz1OIgWw+h5dW32ubvqvvdJ/nQSIbR4eIUrzLem0Tqoi6Hs/fwirs
S52ptBOpikY478+92PCNUCTI7zQqEBU2hFiwzrgGtY935YauURmLfEP/Gocv3eb/
qJ6xWWXjKqgC/94C11AlEJ+qFcpo7D3bHICvXGxEuWUK8VpnRWLVIE1iOZF3hwjP
1gw+d5NJxWmMXqtW2qIfDqTEX73gWTXa8IFU1w/hqN9v0lNZLC9asOiRKnMszl8/
59Oo9+X0nO24kd1B/YNWxi3lLWhs7eVYkQXuJQVQNOg6gIdevD88ewfVN4GFZ6JM
8P3D4BxGGlclw1TUaX6tzLzjasKAO7vGRDaf/TxRnqnoWTkk0KrDL6jwlBrx8ek9
eAmtybVs5gF06tO0MkPndo2p73VFNu3tH6i0cL2OOVTY+PKsYkJdRz0oykfePmGz
ulz678bw1ABWyrQMR5r0xVN3w5gwc7hqn7RKACYpUKM5umi8+97Sa8LdCQYecooH
znihV4eoKJsPWqdDAIS9asm61NUcz7YaGS8mDMgA+qchQJrjxBuoYZ+VUAyn8Zqz
8nMfU/X40VhNVeI+hKNAjJnJ+8GTKiRMIt1i0DACqv0AqMSsf8uNzlfmm4B0wlQb
F10TYcB70a3Q63ikd5YsB8b64DrQ2ZW7ENzRQld5ZjqpYjJlLCZ6R5N2ZsGLA5Fq
0p0KuugKqlJG1fJPFxNSdHQUDtioMpnqzl5NxToiTEvWUzeeit+6FciV8gSFDrxe
3PtEnuzotyace9Zv2GTGENCrCY3uRFPN+3W3HzM44OXIyYmCB/5B78maAl22cXdb
52LGzR1dukiq0OSagxaKBcyGThaLH578/onjPo7yY/kOmf3IOoKBnVlpRECQwoR1
TBKr2eRr/6qc37+ugDalfW6G97ymipaWpfufWk1YrNgg/xeJqMqYq4fqMOXeTo3Z
hCKs0LMXFLE+Q2H19mDxR2K1anDhUecliQ0xbVxpnTVyMadT7ZL9knLnlTWE1+mx
8mdJzzMKOhlfw7pV7oS3ers9AdogjgBzIRCyjAM5fVXYlBh9GEsANO3T5nNhlUK7
e3UzrX8b5FbBPZ2zJ4mLOA==
`pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cWzKEZXVZ/I4nMMQq6QN5FzvI2M6NTt88JkaXfxvQrO0f9CZQ4gNlcldIyOSkI5X
ggxsBxNamP0VUXpsf+SkCDUmQFjj+6GATKq33z8p234VGsdOF/pWBAD5uXKUmisG
HlThusdBiK79QE1vLLAB/TeZXKdpib6+BE45QUxNx+E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10880)
OGYN3Jr3bibO1W4OPxgAIhQZS/+2qu6Tyh7fOb2T/33QqtSEx/7KqY0rvVeammvw
G5ThMzjfJBCQU/sigsfCOZOJvYuRZEG08L6JvjhmfY9h/ag/pdjlZObwm9P7Ayor
IpJyZ9Nc9xJfNTbpWaypAMGoLUgRSDGuX7SSlGfGbY58nQstmze7X0cJfUdAc5h2
wz/BcoUyrCJpGvbFsFXXEpQRPumGKxT1A6Xwya8tRzlYhLiqp2aV9+kGZkzmOaui
Pr272T0eDq/3N4KJcG5T0LtLew/yQSFsSAwk6QS2EoOlJBNWeyGxcBd5HzEb7hFO
50yKBrW8Zeuz7f9YX2Jue7G4JbxInDWcsfTaikHeh8aZvImftR+0L9fiMdPLK8S2
oJbspQ7FkVxPEGLB7fhy5E+KX5vGujEHjzYqWMt6b/mvZt/kRidZBFAhwBP0/G1S
XXL1Kvd++RugX0OUjX6K1CzS5vKxglsuo/Uso92f8dd9DfQGq5ITgMG84As0WJLa
LUqjZuoktuIy+rCJ8O82H5Q8lSTc16K2B2J7nIkA5xNg7vA5DcP9aHNPwFpd7iHT
qJMaXWL2vdju78MLC/MpGV//OBTzTyF2cO7lmjoVu7h2Ulz+ePGeCrTMp5sLvsBi
6b+/lQ3muJ/JQBEYrytu/EdTK0DmZrhr5kbspGsavdtJftVJjH/OJ1MxuhQzELUy
zKaWEd19HYpsm8BtCmEOBUYQYM19cExDTWXDRzf9tpIFWzOOmKFGOrxqyR4eD2X5
dUbJsqJfHuIj9JIePBIVE249fo8qshtO43PrEoUbjw8GScUx45FiXfPb5Ko5b+R9
3y4Fvd6BW9qd9hDpKTeYH7wfF3UQkPLdC07DzAvX/299T9kHrqKXQiWX3bLXrOLf
yygFm0yL5jeINeg1393YFdiPGUdrJhzEC4A7NfcX6kCk0JLcK1dkoi4tcVPHG+tr
6Zn8RHcGyKlXjkfQhGlMn3fa6KVTEe8RpdZ/AF288ZFop0uRwKCE+t88z4PxCxR6
Wgf+VkW1/6awV6wki7fFAIBZWxMyfxWwquXaCzovKNORneAO14xfTaQvgKuceWxY
H6jY+sX7RYR6SRUEJyVCa8STf0ApyvxzqaHJKNUMgPqBfMYOEdtm6zD0oYmpt0zP
nHhWci0Fbvm3kHSjmkP9J5omwNDt44B/HDOZtnXCyeC+vEUet5KfeberuPbiV7CK
32dSx5HkLlcUrmuZmP5KJ/b2C5/v8KK66k+pZDvrvNQMJIfnlDWH3JCT33moOlnw
KnW3W1FqAQ6vGtcZC8EAGIxs+K+Z8qA8ybp1cGxolfufj60m86iJNpm1ognUSqgm
sRGQvSoOSWwjEm0JQDhDC/Hyujb8Aaw1BkQF3sQJBAwh6KCq0mH0So4sDWO4hY04
0Zv9kktsrU1Z97kQ9qV3KX4XlcKHS0WxDsuPZIjKVqpCQdWGx/xdcj6nACF37nkv
+kPTtu1+bWICE8LlvUPINsnmn1cust0iY+LHSHAWUbFHE2EtjnLZXmz4/kyWark2
UxHLGD8I+3t78qfCJHikNPFMCjs9QKkkOZcgCk1qcU1CptBN+bIfyVxyYnNsoLCW
5/UQEvDEqkDZ/AlY4F5/6GU55xqj7CgH1Ez7ZAqLti0+xP3pygXv1wTQrCZNfNKj
Qatsg9Q9aHAavG2DAQB5cuE+W/0Mettrh7ow0Pm/2SGguN7t/8EcGn/dIeMl1vuB
5qsff7oTimFjGi5qYVai8TWkpj2x3sle8fsGEqUy6wJjpeOm2yjmixjhuCn9hBjR
H85OtaWJ7L/mN5KlygfBgp5miZwSAoLpuw7Fw8OObmV1Oj3YQLzrk7D/0JB4FphO
S65dS1+P1ZNeswKs/tJlCCFrZIhaxwrXlif6JsM2cuYlitYMnGDymDdCTX+xincY
RUxE/qS7dvKEQIsbcuPDgW+B2Rfhu1mpcY4jwYGfethdlI+2s+x6gv9mD256txti
IE0EjLayUaFgyK+6q+G+ZWkymKkMuVkRb3wctxsNBPEVtdbmnAn5obcEYzZu5FQ0
eKyG1g+epE7V3k5mfWGtjmHapFTWyk2XpcVYA76VtmsspPHQzR+m7lw5NyISSXxR
hsc0IksL6xbkOGMyG8slHt5u/6Vp+chNxwtZe9fNNcvvP9aR/mliULSeCYW+Ox3o
4z+2gYbgxZC6qxXQNcIvRgVVRsuI1SgqZSleaxhQ384fqhHwkdUqImJaDQF1TDr1
LDVfMnJLyKEMOme48thPQhP3I4C3NL9Iv38hIWy3uUN1gAjrAdHjnAFEdc74rwP/
mbzhebuYXHpDsFY9UY5qNvX+HOxoXtUyMMygi958BvcqajIHBwE12Kzi5wlmBRWW
qQXrgMgEPV1Hm2mlM7+D5IalgFWv1rybPjyPuLzH6ialT3zE9z1a6kb1KVhXgDIK
W2paDSvZ53/HwonQGa9EK69j4L+6slwJe0smaHJh8ReTlSdPnThBXtMOFuftU6j+
hAMGRejceXquEuCrgaWmnwa+67igedA+zZeHSHafp024AiRIXhNFGsssTL/VHZKz
RAMj8TPd7HthzadbMb5YhKmcBwXXYGJ1sCFlOzE6qS85pzE1nIB8SqnCbGo+Om0j
UjKBT5L2f8lHkjrxExrqTWXN40tFX1KHqBHwmeWxzNor3JJ+6kr88KPuNMhDJ+/a
o9ntnunj1CPbbyxKyRyYj/Y6+5E9wa4N2eQwaHT1cAI2dx2aaGkAy7PRMu5zRL1E
4acN8XfD1FPIUyb/6mGPpxeOHro2QKXVA8c808BS07xGYjzn66OiC3MzX5JYy/RV
guaM/yNdHvcYQmj4ZP54St3/9zlO7W8kmWPljpIKfNUcwzr/oy6vfh90b8ItMJHA
Lnl2271BJrSodVJsHMBxrm5QT0ynzmdumOQmHv0ErwJd4ZxD8U42qZxQGun+kgpv
XqDaiPwI40HFZ/zmSyRiZS61lxt/3GV+a17iSdxBXwkYyPJlIwyAaB9JH4radvCt
Mott19SsE4e0BIYHwkOXKHRO5dEPLv7Cg2IdGNU7BsTY74Wd11rhWaIv9vhT2vSm
hrNg1iDKw1vctvwnYQu+WHEQ+pS21Vo/kaPgYdedMl4ebpW1fNSpA6b42WQPzDVk
zwQpdXFe06BQt1ZIDumLCMyRhWrqihDm5IyXWiRj0PwQ7jwdePN7FGTrfbg5snLK
PvdD7eAcfXbm32c0ENZeMKK6vgQtyxCldH7Ot785dTXDg/4lKYBilx/oMaKXEcIb
B3emSnmXPt0gxogodLa8XbJykMXiIRHjX5sw+uD0nwWv5X2Y4AmaeUccdWNLXm1N
TlY6LBcSzeUQE4w8mrezm0Q5MEz5/YKzZPOqzmRMsMtXcppdpzSv7AdN5+c7kNYh
69WJ4I30hwWhd4N8G+ESqJFOrulqtp5NRGXzfUtxkdYcFrIe5wJmDc0y4uxgeJey
ERAbkBeVdnYsXhZI/vQSAw4WA47a2/XOkzKpw4F+vZHBPcE/4BWqzmpy6FXIMSUt
POfq+sbtVDP0PzA3v+5Hf58e73BUzxdSKoWLLSLhVmJv2Z51HaZ+InJ8HVcnD9bf
MVkQX6kzEx/v4m4N0ZhY5gsNxHWayfURYfDYtEd29PnKexVgEDrP4eEKCFtgAYyk
6l4QfP3sLPhgavFkMj9FlsBoFALFhmx08ir5twcRnte4MY1/zpzd84kWdCbkJhpU
xSiZWphb6PSKvm4N7RobGJ2B5j3TMoXWE0RNqr3SS3gwNNKG6yxRjpy2LcXBSS3u
voYPuw/pdhAHo2UAqSOdtys+WWKdf1Qm/a+7M5SVeNCjdt7ceZs/pTpAOfeRJhLX
1dIZTn9fMn2FaAk3pySXD8E9KmGVyjNtjN531Fhpr2XxhVkjM/ZQEPqRClfEY/3U
uJMdSY5v3y6zn9kWjpDuf44Jpx3iucNky+QYAbiqzke2K1IgasPyeU7M2EfF14nJ
Tjj4KeL5sM4YDSIFvY8w03MlRWCxVKVxTrkY1lQABYL70977CEIfrI9/ruRPNL8x
MZwFHDysk1dFZmJ2HwH0uRoXfV8utsxtRWLCtSSkiaC4zIjGVb0X//ZzfWTuF8AU
1ffNLoQZSr8PqmMfr7ZwXG4/II9+GgQgXN8k/7HcX6U+oNPEFAzQiausGX8F6kq+
kPbw6l4XFx4oA5BZzRlS/CEvo3NAjL3d4q1xV8doYWRQCaAh2AGCr9gpU3K6NmLW
5838P3kdVdutuSAC/NnO3hvgkNYboorPjDs5qFtjLrZX2T4AdyT9EBCt62rUbGT6
eNoVzFgkJnJ8XTFsCZFBTFszZUWRA4NvYe+aE+QkH/tQQqqcc0+RRQZt6EUIDtiZ
3LoM+tAzf3eqhLX3btrXDsvKZvr+mIBoKZqK1bMS+ciUXVu98Y0GXcG8J97aVcu4
w2P5uku/tDaz91wNgUPJvv3aqHDaZ/D1JQAmaAvTbu7o9O3ATkXwUuNTGnsvXJ1G
J4Osw3WX+yIhWoed0LejpbQVQen3uRTzNt8w/oR/7Wp3pzrY7FPB5xFOtU9WQwy4
rBpzDO0h5v+jbyWjo3SvJdeE5Y9X9zgy2qh/PryZShUBdLZtO++7Oi3+2hoctV0Z
V1uiGy2GWuMFfkymLUSEQfT+Xlxew4gPlYEgbwkvFYw+sokcs3DG8ao7F1o6aXeM
XYOkxxaCbA0ddg1UJyTUKSdG2NRYCouuWfGWNFqcBSOWzkSxHHvL7hIFqgOxlJpL
7iYj6rvB5icR9IiSvSUwI04SgL6Se+jxlx1qm/aWcqw02dlr8d/bc6gJ8qpf6GxC
Qj7SLIviXHCRg+xXZhpaM07nPkfURcN0sUiJ6pFsvdjKd/lTEs3cJszXsTKO3zZW
qAxy4qW5rLOmIZfAi3xGXrMJbfgRJEsuPsnu2Oj/zoz4KFenm9P49lgtohQbDVKB
6AaMZWM5iBjoZe48LtRfhMkZd7CaAsC78dcSJITwA5hYV/PF9fXiEU6bBPPDmpeG
gngNW7qhbkbjM+0if9I8TUSGQaypael2iNg1tFltG60z5r6VaxgTD8oN04p2clY3
bY98m5AiUYp7JW7oJ/ff+hFz5YKsO4f1Muy94g0OlIai/8sotU7hTqrLbIWYRKFd
anPben/9yFBmHT/tKjRMwm4jYzHT5gmZMgum6XsQsLNsvDie4MUni+pkGGBICpbI
/gOYYNT8GxQZ/aa50c0hGqI9Y22xu0EZSFhfsraZ4p5i4LfTMJnvngOScPL6HY0H
tlI2AVqJ4/xh4idHRMzsm8ppNKPxebVvEBimeVsFQYWeg1jyTu6FKGSML6blo8YF
RJ40RVU/7SPhRpeCMu/prnf/6vbXcw/VK3TtBo2b4XSYpiEb+UHMNvNUWoFKLHcp
7RpZVNBwGd83vwoqJD3AIv5ea6f36ELi8awjjwwYJ0G1vpnrAZg/foj7/Uy5aPpx
hHgibNSk7UjyxTvAst3sCIu0/3Z1/P7awr15PpokUhuY3EL/EAmNECyZ4o4otbR/
XzrJ41+jDU6hGBCRUzGyd9baA/GGNe0nJjDrnz6Ry3CyfqCDbNdPy0JmefUWkxgg
SKgaitOal/Xo4OFUJKNkaO4aXdO5LzRuK1QW1nVpdZTcaQi53Aat4xEoCov1ffsl
Czj+BkOnw0Tbdw0oeQawLKEtMZUdCWLYZpR3BrbK+JVuZs/vRmZeCA38rqBJkvyy
ceXJ8NF4TB3X0naEhMqmQ53eEboro5+J3pULoSgqNvqz4MFUtBQezpfg6MMhYL8E
TX17VZ24egXlWmoqb9dLpBSC5GF5DCAvKLU6CUvLLhBz9a57mfQlsMnQRDX63TPh
Y3hQZfycpaZVsFQpGq8x8HgGS6/17TqWcva8V+WrfZMkt5QXQyZSUFOhStLq/Hot
yog2ECQNGiyCCDjWkY0pEL2Vjpt+JUT2E4TDR+tDVL0UsLEFeb+1cEvwv8CHfsxl
T+JzTy8IAkJ85r/TGohJbuwE2DHu0q06J0H6bI8eggY1Zw25z/k/jDNxcXM0Pch+
VGpJylrvE6A7XEKKNGukEmkOa+16Ejzo8kQS1N8YlLl1HPJgcV/RfNxqZ8KeyB/R
sGslBUtJMYgz0HOGWJ3Wx9MgJ4oJeXCcKFMPqVYXSwQtKvJ6Co2o53k61Yg2bkGV
CPD6vTsX+4HVNunVUdJB4o1fz2TgaRmo2puGF/3MCZubLY24+M8l5VeNQbMiwWXy
bIhKuEg7/kvWMMypzP25kB+RdqNSOAq9ITcQbEIiraCz7zHEK0TshJKFlcRep4gi
HsLxG9B9CFYt5OZNmkBxJSyaaUuIZL7ds1OPsxSPUB6ET1UKkj6tuz2MC1mFmTTY
6/zCt9JXvqbE5/08WDcELJYadAhL5X7X5BI8j8AaMtLWpa8WSatuGwvFX2EMsH9u
vrs43HoowqcAxkbaXNB945uymHn2j86SKbQaBiJe4IRxdaA5TYNCt7SVXg5DOF8Z
WRYguZ0AeHJg//W36cPRETtCY7lNMKHsPvfm0tMcjn1d0YxpSyEFEgEcsW7WJgdQ
97dSwZnWtvhOOWsUVy8ok9Z57B78SG8YqDIj+mbanvmHysgUQNz9nBCL+kRN3os7
WgJFuBDBqh/PlJZHhsZxY0jvYa0++5/VF2f90PbWxN9jPGgIOxA3WBnlAHvFe8Xl
Zq+mFbO6j/bUNkqTdEMF8nRmdRkWqF92HPRF9nnQedpbKhu2eyMVeHqU1xCRvf3g
KuLarfJTLCHWtJpyzy1WLmJWwUYqaxkiZpVy4AddcvB63Dd6fa9+xfW0KkLYn6lf
MRIsARYgYrlyCXG/weMNaDhujFE51eWu5ZjHs4mHhnvuTaXPUpgjADnLtCkR+BCo
2w2WAYimJjAKA/inFOpVLBdUaYztBQF6crVDdysX0LaLZMKpzF+N+ejzLLX8wAOV
XPUQsnrdWBu7AncB5WWssJYh01ahUnv3COi/VF2OBp9wyenybQj+8Ptgi+vk1+gR
tP8LGgsmNKFVB3HKz3UEncqsrznP2g7lpxcCo7vJE6k3FrxAj9h4xdn7dVflrHKG
4PCh++4KhnRWS/aGDWfQ5ZpxtYMK7gNzAlPuf1wKqHT4cVUKKFHObniM3SBnib1Y
gh1qUBHoDcm+VZgVpPkmC0yHutP8wtvxWFu0KYKHdpzQkcXaCvQ7tQzKU15I6yZ3
fx4EYG8E7Ge6QE9cTwdZGdEcKRrnBYnuDfnqHR+nklu7ClaLHYjkIFEIpRCijBIk
5FmvDVhB1UVISBkKAaEce08XFOUTQbyfz4QTqG0tsExGctvNsyAAnLkid2GQGePH
HHgJGbTteBWaH20OY2I1VsEtAWBjPjhUzhbbpm4Q00faF8mqQpp7gD/Al03c9fdg
Cq7op/qh0WFOYffoNXnFxayef/y/4Kt8CsfE3gJ1TQY6nFc02pmrbjOjJjNQ6vdZ
0vvHJaXuNO92IlgbfXlqNbLUZe3lCyM4A8t+TNfJLYRAvXwlVpEz+oMMK3ICxQqF
L0H4/QA2nwYwdr7gUI342eHcqKVUapeBVWiXKnJiHDk+eY+TfayiZYzwMKy+XFAI
MHfj1i3ehOQ/LIdiKwV5kZugr8tHwZao6SA1Pemo4knBa2QYUltk7WBQ1mrzoskO
4mI+lszS5w1Up0nCmBesJzPObcoSOCyNnY6QGZSwtpzZeJDEEHlTcIZ57DMVV9RR
0zzBjtq5OjABEkipROaqq1hwnTtJ63clNeGN7IwzXVhEvNueYFDnthNP5ag6IsNA
97D2m3pStVm6ts+zBLj1ztMtPRrPjebEkumYZyBmyXHvBAqVaI1fn9MHF8+yfvnn
1jhhFeMC2cfE522vTS0mIQqWyKR+l5ZmKBzKgTMEy7X+gBHyR09qsBkMS3hP8XWi
DwLbiAX9RBkiv3BdSoOUufYd9n6VWzw8vW6eUe1eXcMl7Rzg9YjuCwH7BxfOZ0+m
T7G3IXh5W7Q7qHaSFEcv4kPgSoBgvHxZTouJli/bmIODrcidA9bVJTt54K84bCJh
xAyHQRQ96StyWFTsSz6egIPMRoAfSBR4nUIXhgptkxtWBwyNBlJ4nyGuyO7CZDfX
qcabg3mH0VNozvTBUNR2RjY+QUbUwrvuFhMUU14f8yQYARLEW5vSHF6T/qCkEoTg
Tze1YAocGeJvu4+OnSHCxS6SgAokEn3sdc+b6VysUQXtoU2DF8WMyjNCjYCGTNn2
x6W6DhKJT5x+K0fxNxW8joqA3tnvAW5Ux60gmi3QvTdXb4SfKNvGkENjGQd/VNl8
c2yWOR9yb/1SOoKmDqV1Dwu+v5nfS9cokPmxuMMs85a5qjpf9YcXekaqHsDWWrC4
C+TzsjHGwZtIQaJ9eRsDkJ1qJj7RXe7RJprZoTPsnC7Fb3EBZCdjtBMWhyGsjU7X
DBgAOxlsOgbJ2l80+/lj1qrMb7hIcynKjo1IXEX+rpJbT06nw6OjLGrVmWXCapI0
rYX22L73qBNj6ENj9zTebE2trjyOTNVI1nKPltA4x2bR1BoC0sWivVLlcGYzMsMr
IktteQW0wJ68emXPv/f5WtxLwZ3OQeC6NNwVTQkEsj5e1ijZVzM6cFcXWJXv7j29
syHiZsJ7XUVxI1D78u82Yj5oN/P+K2wtQh8e/O001ZTUcadLtfidPRhRR4pWPJuL
JPfwST9sGzyKv/hYN57CHIfD9Ut7I1WVMtK9Q9N3ufPEMywdCSRpOkRy4otUjGkE
Es3mKAq+/3sCYeSImveTeR3nij0/xNBddYJMdOVrxVK/tbDiJEYUi4gq1KGMuHlf
QZ3dLVM46nt6qZwNieGuar1PPPy44m/4xZHW33sWmhsoO+gJJBMIHa22kMHRrtNw
4co1HWsM6ZPEcA5giY5FtH1xRq7C/eqSr97vX379ejchlYySD5VW24SZDvsRuTwY
RWed0C4yXEs0vd+TBL6UbkmHzKEs0kXZVvNnjfWjnyw/yqbybd/Ks/YWdqojwN8Q
TxJpnEpZ7KPahPtVCRwPyRMrAktYyQ8Qa4Tq6/vfMXCPpgGiH91abPbL7HmLf9Zl
ATZHXokQzwoviZoLfaeTJ2bkAzlafPxadErnL9Eo+hYkjCHDY/oGPcEZQBQRehUM
hFLj4FhVrWTS200TYieZNHhbdmBNMhLjMdojBn5MebInCL+YrkmXiVPabeV5Dg9R
VupGLuJqJFC2pNaMH1AeC4bGkLtnpnNa2//VmydIpVfBcLeOKqrBcl9nASXPqSCb
y70qO5xoPbeiO+zMVwXwNzPvY0QRQ683f6UdpqlHxpuoDBJMFoPb064RvnmM0fEV
jKOPU9THzbcO+MOGXOvnmGItTUeFqUfxKYsRQKnus0HnRkxRRTFbu/SK2EEdSggb
Jl2HXIpHMahDMQx7fgP/+lXABhNO9blLuMm3YiqSpha+zUXXxmeQN99oGSK4z/Rq
IQWyrrGxlm/Smv8gAFcqe1zYpBLXXILiRXRE+H7lIRGXsEEqHXzTeqrkMIwsu2Qg
hvUBAPXnhjyXKos1mnUDjn1Ped98KpXmjetHyluBxKSkCHAo5lqnJcoAlcCyZK1f
GuUFBAfvxdjsDIIBs/S04hED3KR/KJIGsYzrYyDAilG9EXyNnStPPxf64jQnSbfx
X+j4yBu+Z385PdGSt1ffXnyjANBHIPBLPizM13QaiTYH8WQZA6L/C0CBp+VpvuHd
EeOwv7k7lYw5FJzLmZmPlQHapGZ5jplx+miSFLtq19a9zLnX5OdUbQOXEfA3oQKB
Dtrk5bCDPCbn+UbfRKCWJznX5EPxaOpXTTc8IOBEs/CYSiRAyGhOQkkpRIHd5WcR
G0V7Wl58q1WXqUaU7T+YBkr7rDlAMdDtqEsDi9VUmZAMJoPsqkAe7NsOZkNVeNXU
svhm5I945otAXUzLKdSTa58vtXGlEEYiE1QgrEfgh7uySIUPrj60lhNPhi44VTQb
+Pg012FJ5xz4q0hNJcOejsNx2BC/mWEOO/Z+DQs8VQjzKJGosh1Zl//q1BGOQlXj
r7pmdMnFWIAF62AZ3+amhqSZ50WI+Mp9GLNJAnC8XwwnX3nUHLCmhb4LcOZMUkQ1
56lSqbSexk4WnVIy8fbhMkODLrGCVWi2C/koAZ+K22h4WrcMHY1zaJDa+5ieVN6Z
4/pevmgcxnHgU/9uPwbNLlsMMZVbDN9ezrtzb2Ks/TlPiCHsyYZyl4KfYL18rP3s
BJJ4o5LlS6KORkMOvmqIO4wxXZ9HRKWj/MB9FzHIKkG02ORDxr7kA9eE32/TXlV6
iDJsvKMXTUYR98rrJjnrDWHGOZXq/ZUWO09Ktz+/22PtFO/2iRmyfMntShCYj5ZM
TJoM9gIF9NSmJJdJU4ANFtr2iwKyIRtsFIta6ZOawCr1Q9/w9XscrdSYJLf0Ggyq
LBIJLDhWDBOmlt7qrhnLXTqJDZA7CCRVCmxDvjw2dzs988naDhVfVIAqISynr0q3
jhsObmmDrvu/Tvr09Roqba65e1sVkdOFEX4WOmaZyRJn5A29hGhd2SKeqs16l9on
LZ8C0+w1aCdOJYv2lk5ir+0NMWMOAq8FJJvKiTmseGsEFeWYMLjK1lYGMcgo0yBV
UGY8WzcjR3e72rgIalY8PIDw7T84cTZLkJFmMgJHbiGBRzR3IGyy8xFIiLGGVkOS
MO8S8vt1T0VzDQ8KDOt8pEVLKLqwWQV7/eGG/Z26uJR2ZuegCE9j7dL8TG75JVJ9
jsM8DN2RGTd6ruZQyiLUgpCsBk0bWdEeda2ckeszmWK8V9i3v8YRDs6zVecB++Ot
C2bBiHo8oCDtIQOWuJUGNBuscJtTNxD0dYfh93QKIzBT9pIzbwNDcGq3Iw8S68B4
NUQPfMUOb8i3UDI0xRG/bY+8ubdYAh/qk+Fc+AfPrkF8cH18mio0N/QA2tAq5ers
ljcCgMSxItJU8kfw8KBp5UnxD/r6OkXKXqElS6fNnkqSGAFXtVW/wg8UJLnJuRw7
rMNZ5XtTWJ9iUFaEeb2MKqVzEp7+rwPPgok2e/+1M8KLTaC7kUU9vPAh4Rl4rCdL
bAo0v3/MQX2OcnS+cNoW5IMf9Qa4p0xl0gAp0rlC+II+t3UMFu2A5xWFHNIn3Icj
acw8EqAn7WQXhHV4u3IkUYJxfjbCfVD+V69xnOxck0aMBVYUxM++XDwcdNiMtB8b
327Qua4nAvW1TTTWNq/gEm8VReM02DbLLq02jdIt6sjA29twWehGfxqxW3UsRvTW
oSluKoBribQ1bBsgS83fHGbBVGGcKwl+BxDHiNjR0RrF895DdZrXKZOngREjSa3h
eYLE31je/tWvSnwvlgbgScxZ5y8GMhsnP0ubmcPLylFMkjxMKfPE/U+lStH2HYUK
JnoVd9O3vP7xtM6KvGxpMF0Gp434L+HCOOelG/P1p+t71K1uFgUsLHSEihhPODGF
jhynLQCNC1niaH+JWIR1cebJPlL4kqPNEDAoFKCqfo/85WH34qjLAxGVm0XqHihW
RX2VIiOM/jNw6IM4MZhiIhEMGVR9lHztkQj8LeHRRb1Ys1QV6nE5gTtyolhXJhyb
l5gGj4aVGCvO8qMfMAVMr9y4DSiZ+zXEdvgR+TM8iclDIb1shjWNKU731Bj2xirj
M2nwIqfxYfKCYK1aBjl6sGa7NkzsLe/17m+3HmG1kwTsJHArMYtdGhApSEM18Y9I
aewc5+Ef38ohyM2SkpCDRchMYDjnpkDLCQkTXLH6/krkQ/JtKuC0i5ADycVBUacP
+3DnAfIFfgm+38LK28Y+qod9i9fnaq6FpuFHbLWZ21Yh/XSzxujyW40Z6saSxEyG
trWwXFyx0S58cWmZLtVaply02UCLbxfM9vh7zxZ7gLjgdrzFdZk8DGKPaqg4wQpI
V5KE9HXg/CNb9BXXDF3UjO5b9G7GhcYJQTpLe7O+Q70IJ+4u4kILes1Zq60vRsrq
I/iZihaONTxEW5ZhE+gUDU7jHDePf8SYHWoU1Egm0633KHufvGtXcI7aRbppJdDu
oX77v5dtuFXkBQHNRX3C2HtZjEWXWUyJGiSrzyawf+4SNTkqYJFy1at+kIq6hvbe
6CewdU9EsxiIv6ywxS0m4IBPX2Z3uVkh8G38HN5F9f/y95l6w2WjbHQZlFFKl5i4
myjR/rg4j8oCPkNhjkMUF1oWr5ka0vWauAPEOtFlxfRDDLA84nNPj5BzVB6kG0YT
ao0bTfwk4jUIhf4Itsg2DHDSrwAhREAw1rl7H9o24CrQKL/wQEoiYflSZTt/ohvh
sWddmyMLMCwZWm9HIwlmunYHGA5qBsvbk/mAf86S07V/2pfDZ7l+pKjDfcrA8CGS
vVqBsK73gFOi5qL3ASIzvlmA7WwlenXnjECmK/tCmzMcYBCSROryLoj/b9C/8ojq
wV+6iBbEf8Qynbht2n90VE9luAvvanQEmPQjp2Gf5LXjE00tHZuiI3pm1PsNcJha
sLRiZNAfoeFcc2OJklYYkt7Gzju129k13ZUXH2a3KIjafFOagzW/elwzjfwAFWWN
ddZi0t34cxlVd8r5AT5HA5zcmnY2Ibgc8WeSm/MxixwXvQBnY5UqFqHNONLW1dLr
RJeZiGyYxPvQJasAAM7mQLEUanH3u3+jErCLCalPGJLAkx54yzLGzlKsyxCoR2MQ
mtXC6GogA2E5IT2Vf/lqPfQcIbpAg5fHh6+gJYhPi+egKQitL+DtUTFW4v8c0MBR
zih81WruvrncU65PfjBD70VNZThLy0DaPh+PA92D9dOCbYMsPpPC7D5EtBLXKo4o
4B0i6E6dui33xKRXpK9I6wwsxhlSz9d4yT8ltBPUrb9j6RoShLxZGWj4mC3vQFmX
UweqxhlA8Qzu4C4p1w6kYuWO5sp6ahFw40KYUxKT/3g+j719amnMZQAwPx8ESM4f
cAbs+InmZ5SjPk5VqND9BLsIfEf17iB8CiLzsm3O/f+7AwjHb38AycuJt9ZOLfrN
UmPPm+VOPivARkYtHlPZ7PWqZd0tvrFyko8QkvVPyRzScHZG+y2UQ6URKsLLzdGJ
fd7YTYRieWMcoh+9E2wPvhNVVEs7szgdnCF4O3ZYS8MpiGzosjTjcltEE6ocI0zS
epMyBhZURZ26vK4Qu0NL+hvj5oGTDaCIpeehm31ph4ihjV8aPM7syJxcQbsYRuvE
3Spu8d4hAu/4S4nYQfbI36nyO4y7BbZbkzCnuMj6gfsRYQtZaJ4Zk7DXVLkiuj3c
YwNeZbxgEV7Ux8W0JP5jeJdSDcCRSGCmuyRPLPgycgfR3NXnE5yYTIPItpkIexC7
2foy94njEQWK/K22P3H2CHThdKsWBFtb2aAenDWDz0tuO55hQvJIFmwVVCHH899k
X7W0SjuUFEj2j47oNtobbPsC/8oZPzR1sixV7p66ai9hp95h7kuRyQDqvfkp26ZL
/5BEZKTfmnyGln/Oo8HVWrAwDRojx5UnWC7X8OVVAs2d3exmUPk8mLHxdYSjlhVl
vsOfoAiD21LlwDOa2k7+q+UA5rfuC7Lo60tA5Y8FS89+pSxzjsqWKOTLP0Gt95QY
24szB9MtPo0RF7wjcB3eh8Re+9fwf/8VWDaASfWmGeMyL3wm7x9Liv7VCa4lFfm9
c5Zo4ySPPe6n0EP9hcDi1E4BbdJ49i45UfsP+vxTCUEDW1Vkq46dUM0rWXF++kLI
WowNbDXpHlSY5gp2buSzMopknYHadWqBMZap02Gtv54wcjmP59BEr8Y5B096+Pgh
mNFI35O3T/nzi5rAM0ovC4VCF4V5XT3Gd3eSKQH616qVviF7G+4xH1//otl8qA2x
whpaMGKJTBaB6EkaRx8W0KO4hsdTErjEcvKeZ04T6IMcnVMVdm/aDV7VHzgf8OiT
lLM5zx4OBNAiB5qvpHybtrP38ZILzk83DhPO885xqe9XQMbngNRv+PD3dAqjUq0q
U8+T4x4o4QTn0jkMgXMM02QPhKc1v2073xYKEYLPLqj+v41idWs19rGir53Z7Yvo
DG+QXQo8Xu8xPorVkJbwAHA/4INYC7p0sARJaCl9Jr4axXth3YXPEKLTKjU08pPY
sTVA0DKSSU1cxYUQ8waXsnmipjmojtOF00EkIAm4y+wLDODCb/pjQXTt08Mp3L3C
X4vMuejvVwjg2FDj9ifS5a/NefvsUXbO72YcZn1rZnakSDIepAQasvNUeTGpyOL+
5U7+ZLkBbTTttAnG8PZbUwGEVKtP70soHotaK+1ktfgIarH4+FvA+cw0kCkEt+S+
xvhf13vXhxc7/w8dh0oh4tVmkmPS1NPmD23N8+DFI81Bg2wT/5RTS9f0khe/nkJ/
XGeNbMSc3IBujTJ4/EQvbC5fUVJQv3Jlp4BLoqvuCJJWFwdcdkDOARQtQJdvR//E
lRRJXwacIL8L3YpTCbfaPpx5PiWPh8D3CRUgVjaqnvKRzmEvnxfsg0WP6ouH1d+7
bE2ZS304vy6ys4Axlb0amwqBhr2L9L+jWmknvrLbgZ7SyN1iLjyS1R66tFs8LOA4
dMzntDjSfdNEJzSgDuVIhCBV5687/okUfeXbqMVcTgc=
`pragma protect end_protected

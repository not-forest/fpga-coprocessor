// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
CHRx9WQBg0h28PTnm1Yk+FyNqUNwBc/m3JyLcctIe7XuPuDxJgMhjOkAqIs6QBKT
uoRrWa4P3CjmFg5oemPGw8SVZ5BsfpzD1XYzO6ZlVX8a3L9SgqrDW52lPQJUkSGH
3mZXBZ2KWTCi/c7yBtJ9tHlHjFYoVuN5EDs/XoyTnxykqh2FEx4C42E57zmrwuw2
4GZmnhmTNp7DAql5c+K+al0jpMnqg8mfgD0ENTH5o0cFgZrqx3jr81IyR2Hs7+yO
RTk26TphakFR2WVflU0ulxo7nG7V5z87A9/OYdvd6h1EmUDN0VDJNw/M8JntfQZV
kD/3fAQ8s2Ilofaxn0taBg==
//pragma protect end_key_block
//pragma protect digest_block
34nzy/o7qcDvDdLr/PtsZrTFPMA=
//pragma protect end_digest_block
//pragma protect data_block
xq2n/M+iNQEh2Q6fCIBbTVZmltpt8YYzENW2fR4Dbu7LXGOoIYI6H72b0XtMnxyz
euS8ItQs9zu2rOULKYL10tozdfdLz0HfOKR77rcPoE2Px0vS/R2jBV1vGUf7OVDb
7iPsDNBxM3PBt306Z9Zk9RPn8yrMdbVfyGbeoH19USWz7E1Fi6/FyPbaFrm248CV
hffjJJDNO1S++eJRHk4J/K5H5rOx4k8oF8oVUID/5UchvasejFoAzJ3GfkE7LSl/
iFXAtTR3HKCaCh3YVIxav/DsR3bOjPfhI34r8f6IVBYLFssI5hqcVOMh8wBkbouO
+KNJrkUpJezCPaD/1vu5WU4yuu+KO2BhUYDtWHsCy5TdojhLAWIoV7xLw16UlETg
peNkPlMFFG0uZn5+iCU+34vh8EhNBwoFGoRIwpwy5lYoBJQ8qLL5/kW1mYGnKF3C
1AWKQkNVbQeEUawSzWN0uNP1SG7UK7J+d3MW2j1IzHwCFd5pKHzvR8LraK9oRIvx
1DXVinvlGuC+2WhD0odcc8oytboImR5HgGNscvMzwDMgD5ZNAGjA8lGBaTkNe3HC
eacf5WT0K9cBdCTza4oBSJNp1PvxmYma9SaTQXJYzTEHeR8Y6RPA90iFpZcg3cGR
J+F9xcmBISCnXuNRJkxrjBmvPFZKtGgaN8iW435ii2Q/n+R8GSc/MUp99AZOhET4
SQVXzqJsgcfKSznHJPd0vf/0GeZY5vG2d/iG1LFIwdxwA3vbErsjPBu7zV1QEc1N
cjrZaB0yptT9nYSLbnNKzu6EmRC27PB+ZFwK0G2ctNgkE5a6PM0UMj/L85TgHCbu
dbPihERsIoWexdZ2I/daQLCfbKJHSgo6XoTjedd4ZW7N7OgsEbul8U7Mc6tg31Ru
PnskTT+Dn8sHj9OL5Tg8VtVqFW9dQR9q+5PTQVz1QbNqX35YmaPi6Iej2AByVUAk
j/ZE3ok8S5zolLrbZz/+44F6LvGE6b6957iNQ4xd40lzEC5giIWM3jdqPoQ+okAK
KrRvkUmbPP0OP8EkGEn+GtkrpG8BA0R1UZCNl5nsBHhwfS/fN1dOp2P5oarW75pq
Mq7BUCb1g27XeXyrPS4mU15QmIYyCaxsIoVECOn9UhL4vF41ywSYbckYKEH2cv4R
BaW1uWYuLoPtbkGg48fPSRZltHxY76cy8diws/ER+f+3gvRhPgoaneHXGkOqJPcJ
qIdWjYhAMBQByinzH9HcAobz63XIOVrK8Wmg5KujIs34MjFVvzOhmV2Rek4AiWEx
O3tDDG4WOPIY90FBdq1TNI3IPq9v4fNG1lHt5rbkZhXrbw8MsS+0izFU/LMSBVl+
XiwGaAmFNry/1hxIiTJaERpK2rKj4VG0cwSW+/ZkJXSanTqalUlD5cWs6XQdWqGK
1Aaj+6y0AJGS1Es7ykh2mNNYskW7mcZ4f7FNm/cxDUeMG1SqIAht8CMuyriKnprV
UQ0JslpD7ySH/eeqbF3w9UROVDtyvwIFh8CC9Ug9J5a76t5WTOd7tJTewsz2Duul
4haVJc4xmGFJvukd5myAWCCrPcACUbyFHZbGlDkbV9M+qbY7TEVWNZItDLUWC6P0
nXOwbo1cmBVPRr3n/cKVnXu0iIxbfv2lIG69Sn+Lb+PMRYUmhrol/7EKO3ES4RX5
LkScr33UxKn5Ul62di1Ek0RVSP4PWdUttpvjJLO4wtxWA+2B0GYx3P4IbyQZbege
mfhjHkBfBXdzGl/2BBEHE/PIJMPe/7LQ53+DDAr9Og8YAji6G3ejQjjVGtEg7ppX
kDH17DnTPW+qv7kp8symmTW2ginyseS3yWM91r/WT/ziR0PDgYF8AIfAB3Jzd5zt
Dp+u7vGRuAWNFLq18JZaUSoGfz58M9ZwA/+2rzU7CW3Ss8vcMXlYIRWbk7GNzfG3
YPlk4EkEIqBw9xWP9JPQR4MmBDS9zx8zdKUf5qtc6wwJsUs9rMSslTeAiOOLR+NA
sGCfqtOzFMlOvVgDY1q8O2bCi422dfchvFeUTlXyXksSZWKQ/qhOPj0XFthGHBCN
bsUqgZyYvrcBfEB29OirFQ24HtZkdALOJTXT+AmAkJlpKU98tPUlEdFxc+Fd7X5G
P/3Fkl9fFMq1X6OnjG5Oum8wSDRotwGDTdfAa55OtR9pQwNZzhT2R1RJ3R6lAI1o
SAfFE9gvkBkAJVX+ehP7eZNVegikBOmeFRcGDjIaDGcUfHmhNz60tnt6L72wP8sN
Lukyn53wRlWhzv/sUymo+K+jbjAoNV652uaqg74AO3LWpcV/O9leHZw7QDSKYdke
woRuY11f6VsaSarVV2ZbmWI+8ADx1n+Pv28F1riv32ALuN8wFb3bh4Y35DTXVCKx
8VC3ptT+DmnvFBTfoGkL/t8CPT4O+CYvSk4CNrZzuYY3aDobzEd75XCW94EGIrZl
5TqkbUuuPPqhgxbyEiXJzJLoBK74Z604IKEekeYPfl8kqvpxWwZJNMN/hhFwcOdU
CgI4cv1qR96vLyasyBbsxnhkXQdN23Qpe6UH9s5wL87St9lWO1ReCUX9+F7e93BL
YNz8WQfDHTF27l5Kz82DWViDO2+pXYjrawEsKQneW9STQaCU8niZc83AlYjv6vwz
le9aUCSAj/moOEV91F+cTQQicN944+WDOYKr5Y391yEhTrRNRukQITtr1kX0xg7W
9dyrXVHRWipruovu65AOX11ZToao4etuQRqRR8h5GaikZhqG1bTk+7FwL5jN+2oS
E4XlD5jMnFB1N1nZ60FIO60V5hJVH1mZPL2+QdAoVV9IwRgeidpkZVdRPEKtigYT
flSjczhAR3HW4PW4bt5xJxc63WKDtbJ5pG9HJxIEFyZ/Q+kTvKMv9/UbdgO7eQNk
u8wUxuDU9sWGqCCk/ZZBxoU8pD3Po44mDpnze9l7ycWbdr3DDqEnS4cXwga6vvkw
FT6m8o3sEdO6SyHlU1+oMv2nCXDNji3WCxjOG1vA7KbI38y0ZcFEjOJ9Lh8maNcw
4+GJNjDA6TTEft+Gz2YPM68jnsFCvPUOAl07Vz08uFnAgULZv0IBQYDZXM/Q7nsf
iuiMRpEOQ5HQ0FPlOAjpMzVMDEXAHmuMbrBCDlMvrnAkIiwu77BgnHuuWj5jzwkN
bDfrVNZDciTlUU6ffqboWjmo+ZXfIRklxE8LTOAas7CqJeQ5zYujzON7UjbSfnBo
Kst3knxkScefa8N6oALPs7DgiZTt4n1h/gWWZ9BSPQ61URl+7B/g7OdsOAyRgdTL
trF8EUDPb09aqR672eilAxUaCUoNRuzF9e7ssm7EPkxApk9xAVQkKXwohnljqFv4
XluCNN0Q77FW/ViHpBvjK3lePx6AoOVn9Hd/ncBeLu0pYJa7TtuZkdjF+1KAcY0A
wGLQGHAd61M4GVgUyLQmZLraFGJ69/U4Um4uhw80NAWxSaRNSg2Mv3cb8KGzWXln
Hphj9zHdrsIWxm1lu+iQ52sgWGP04chmJDIzP+AsAvoyGDSBu47FZxrRt8bpMucW
eCZtkNVkVys/SyExJb+iC0jM5LVTcE/EZnBC2ShMz0FAIMmESj2KxVZ/ISMj+BJp
s6sLJCpXTTBovZGwySv8PgnT5rHXLSVK5RSvcEIZkXClfJ8mYNZQLlSN5KI7J0NN
T5V8ua8+4zH3gBRiQ5ymvTsn9d0GcoYJhVfKGE8e63saER2kMcZBHrtE1Vq1prX2
QF8n/uKANrM/6BL2AkhsngJ/hurp4sk0yhTUuiUht61+GLu7FRTEnDdQrzrh0C9T
+Q2qk/mVlMJuJhFCM8KJtN5xKg7kvsng3KneK8pWBFSGWyu6NQjyRak5blRjcobT
0P48Vh6B9wXRvrIN/1Qqa4O72QMCnyEv3DciGNRLttL1m4MJSH26oAFA9+oVISK8
RqIZzbC4YWhijTEzShiLHkto+ew/TT+4+rgmizVQX7RAJ14vfDp9hEqkIPW4d2P5
YwpTSkow8UEHZlu579Z6G3NnQE/tWruK1ASVsRNtiJXN9wTSGmRXsf2ufdY3cxV6
AV5Kwzfpt3L4tEPoB1Z05QWWnim5YsitPqqREssgjF6m29ewWy3Pknj9DRNrJnMg
F2Ox38Qznv3nNNVTV/Qpv16EyKtXnclKSDON7TFF0RyihNvfujRCLM5e37/9BlzH
ZIqhHYbN6h9eT9EME5FmkziuXqFvL/qZHqJHoB6n/BZ2bNpXMpvDv0NkSJZHeBwk
BkpdTUIVsaypXx3PkL4fzl8AmDNW11tRiXQsPK+9JdjciBwHjYRGO2tf+C8oKlBQ
kOzee7TeuiLyF9Xut/AIXwxlxUOBNkVNoYHw49jVsuU98sr2TzsyqXdPKso6Cq1t
BbHGAqmZDoSGW6s9PK49Q0tjW9cMuYfV5fML6QThtqQO3SS1q4RExQQJS9zgIz/C
qEmOMv9yWyeg1H6WQSP1grZr1Mk1SXs/CxOA4Kt9yGLqLkPUv8Fgs5RnA2mU2Oq3
IyxUkt3Tfg7Tfa3wDuCJuES6iICQgel5Bt5wXbNhVvp7+pIr2NDVGrDOCnh+Mdrx
reQcHdqbcdrBxTe5aeR54zFs9uKAgTTjD9a4w6qF0yCnnk5KTq/Zu9qNhiHQiHs6
h9YIMMCdYzXetiiBI+YDWae2jxwN0v/Phc8z25rbYIcy5cBhvKvOAx3tloFoL9lf
lHik25DBaviyllH8aa9WfpxAOw7sVUCTxj6gx5zmbcI8IO0CRyJYOCXFzzEjhqx2
uxx0JkKwqCyPetptPVS+RSslknCUM5KrnN266PvqNNBOnSV7mCrVn/BB2JmZpICX
5sdpbUtiRRShlN2jKtTmyHGBpKi41xdH01wH+uGa3vrDnv1K1YKnNi58ePvFp5UI
xFnCEQ2g+5nHrA2RNvN5OEle4ly2GHNCL8lqD0FZkgnFp4tXUWJTplpjTyyGDI19
xf8dshR+etduY2KXC3Ux1b+EN6Q6VQA6ZQ18w08LzxgtB5km5zH96mviFxtMsD3V
gECb3Irq2IHK+yp39wdHWKU02vkSYvixN8+HoFUJdQzyS8xIwQkE14Mq1aeNJzav
GDW+ABhKNKay9hM6SChXC3pP9BnVDD5grh+NCx3dDI1PXAsRfbLMma4OdJWiKCBa
cGLvf8H1iVbLH8fB0LBB9V0TbrV4JLLNx3GrlARMgAu+wnr5nRlijno1DovdUkrx
vDAfEYHVaPAzmZqlkKfUzQhWSngBvQ7Qio4q07t3Ilkp1EtGU0bjYjfnHka74rZ8
6qHFwsJMFtWgI+RS+hUH5ExlXSmeon0g7G9Um5M0ChRLz+BLewKqcZPuU8n2Bhqz
QCaGowgAmofq2sFCz+Q3HSnFS+K0DaLyW4jzD6cV7DTuBj0Q1Ia0r7+Sf5Dcyr12
7qSPiVXNY31h950Yom1a3YeO/GVqVUPJB9zAJ2kfXC81M/L0QdWfhiVtsUe9HtKp
Dy1XhjUap6Nxd0GcClgU52BFEF23uRJeR8dlqzjDyN6qd6Jh3EKnwJmbEjivHRpL
ouCwvfMWiIDTI+d0CraIGDGACY52MGcxkm3LV9LWHh1hPGfba9dFfyupQPSAzp66
j3wQoMyaOIhSwh3BQrg4WEt18J3QXpmSpM00OXqDAdMK4C7tX2SBiZCNakP7fbxE
ejA73dpCuVRGaSFZyMAv7HJzwpk98D/rG2+hCL9Da8MFVYEqEN/3SkWmT4jOwBu5
LLekTn/rM10cFllen2x2NFdZqMtLVYKutW716xZAHQ2tmO+6rekUULZR1jeKS6ee
v3av4UiyrltYi0DssPDl+FVsOQZCWjD8/azq4hiocvRAkb6M1tRfYfQwssfQ8eeW
yzPC7TVVIzaE02lZ6ypI9NlUg8SBNBvMHFzfcl2NmTIQlnIPy9NR7V9CvQGaqGZr
sIcbSV/+4nGZrC4z+J4NGbrjX8NbOnUe/7ZljtbYorG/jbcwbepPtsqimcrkhMHP
Do3UGMYFIavGMoJZKwc0aA9Re3N0X3PwET9aKA654pD7hLxkwvZc60tjTkEssTP+
dRG989gMeOxFLljX1pVC8p5X79fgkBB26G6m7m9x2MEz4fXfnt4Kd+cuREh48zeW
0SS1s1nxb2r2KeIWDgkmWPlfXhl7ayoiBWqoVCHZ4RagwR+Ja+ZI6aZG+6zg6g7O
TBX2RiOd6FbfGNDb7DQK0sH7APkHSAkRFfT/yU6+fTZVbRAiW1pxGzxwQSjfh77r
P4ILUwZ/gtLy5SynPIgqnZPIFSJd+b5ksVkf0iW8twN3GymraX4vcaCCfbhxg/Ls
Be5Hk4oCWui2/jLs5jloiMAqjxb0sYzAGoZrZWLkK3OMLBzMQhs13+iEgjhmiDHb
9tGcMiowv7S9o2QXgpT3RAOiP2vbTYyvjwgCypAMe/mTkGqFUcKfHbA0/R0oGCey
5tn1IzfcVmhA3EkxrqxsSOXu1Rj4t4MIRVqpfx2r2zuRnLzNR0rNxS93w7eiGQ/K
G9hfbj++JZYFXlJhwIBNk0zot3QstW53ucKw+8EyC4AK7T4IICfwgWnqH2qBrlFo
VY2/HvB1tTqA/KmmG09GAusF/kuTuVs8wY+fmTo0QUOZX3uiqHhUIYMVA22lle1/
PM+DvPqLQWOkzQ+ESzUDNA+VdiJe/er4ROquqEwj+unP9LI2QJK+6m8mQB+uL+e2
WVsimQUyAHKwhwn9y7plN/tO6rNTS61ABVkBsUXtsMcj/cKffGDVzvZjfnBYs4FL
NlpYuAqMtSpZpPeh6p+nWYfhUQXqVC63wYClOeD/4AO0OWQRHOtA7ooucPjDfFNP
PmDTo1bwwScdp96eypL+fxVfmZb26VoZGwlu6is9jcnACsE0fXt9TV2nUAVlPyJ2
AWRVkRBK7LjNdnvTPs5amWrvujn7EtnzNH3vQJ/BiUKIUmp26qCLaZQ6PClZ8P4B
v/OnifQKZmJoazD2u9GUThfuQ3DGjyAnnOUfyqDW6tih/dWsbs6vLxtRrT/jpuZQ
0EnnlVIci6/c0a2DOoZPq7cibyBr67p6DAdybZ4nP4zrTxFYL1ExYav3k2icTbJf
gOvGo6gRy2cYcxYHWZiw+UutUE++fhCo2eTImI1o/zeIbMc2nGlezuyDAulAVxzN
asVLtJtYv6/ItRMmQAisg8gz626XXBymZev/MuOQtrlMFXt1iQq2t5h1HT9pxHIC
tleRESM/V2/f+joDrSiotm34UPfYdXhd7MLRp8TNPk6C5Y4PC1KOpBTuk4SCQEKC
6/oqlqSz8VGmaP1IHmGwfPauUrPN84YAjIVfDnA9MrtdokIXuNMymXEt2VUfj+LD
3D/4fSZIuBndHUmy++WGzSoW9mSMOi9JWPlxrqSWJ5MqdmnNrTnkeXyn5asE1z54
N3jAOgmdooeGxZYgCH4TjIKwqZ0hM5QmC034TTcqHdllA72uFk5SJ6M5vqRM9KE6
kJVySGDlYpRVZxR9A7pJL7Tgijv9MDJgakAMTa/BCfK0kWQ8yxu7sJx64hhKgCaq
J+XOI9hPBhMsH/TReRnJbEwmxdIstk9xmFJix714ah2CPCnnzk9vA63ucalGuZzY
f735xl0O9xBLP+XsM4pRmu5SYWTMvmwPqfIBgqfTt1L/4RYobyn3Bbl+qQBvB/It
T/e8CuZA4ki43N50ZCKup4MWNOFUlPb62uRAr4Eet+NeuQYX5JSwzPsCyfmD4iso
DbZUVrupxfXoWY3hVFDRfYcTdnfa0fI5w/Ap4h7SfRrcoBVOIBn3NJ1lDKTbe4Fo
Zi7JnSlTBYaMcvrOTZ4gG8BIauUvQMr4o+h/Z8QlpwOwyuf6rEQVc7TdD5nGAuyL
x38yl5SOs86js7omcspxqNOUua4ng6h/q2LXaejh7FUctnD4XkTPIHYWc4hjACM2
sza/y4nlwbrYidk0mAayf3t0TP6Pri+U4A70ePS56Gn9CqGF5HmDbNXMA/DlCQ6Q
ylFE4PkhdwJodhKQaUKwbW/fGLTftPtED2MwKmgu/3cgEcdPg+vnZE6qgsn1bscS
ZzlyaV/RcwyuiaCzbRUxS65i/0XECsihEK2ATYT6/AK4Rz9CUrgCcRcFzf4qiYVM
HjVptgtmMdNecvxIeDiujxqW5yxFbLycfFz/jF0yzT9fw17mNvY/lRQE5xUZGcPJ
eIPYwbKarKXyEUyY6tSISW348iuyTuM7v8mK550PHb29bJrSLvpCZJgZ+hg88Gx3
soQoMdfb+oxzdtPFjhF7tK9zrK9LnPDm/f3RcjGpDM+vHc9R2B/WU9OnZzeDJ8tS
P1ytfdJq46K8Onabq99eRFCCdgSkV+/gNoptyg7daLQ1mG935jHkoz2maLsv6Vt8
C3cGYniWIr67TqAKucuaUJczF+lplZAZVIiZfhtNbfysTV4tCq3OPvndIXGVGgck
73Zo7bLGEdkPdgcnvbUmH2Sdg+tXLACCoCnc2LrtL6+MulkZm9zTKVtm84hHzZYN
mnL5ut8no41fosNbzcG/4ZQGNWLxMZJjd1mCaFrSdi6OFH0DpfWD/sOrBavMv7tK
PYlGYWIYMqiIcE11OQwfngWZ6d6eETOqu+Nld48wx8WP8i8rNuYohHGncTGjv9QI
rhy5z54wUO2rNSPdZNMdzWa01b1gvBE5L+YprxUdDGJMFsS/E2ABMsa11Csap4B+
/YMYntMPXCYYFfXRM8HlvtIQ2QuOCur1EXVTev3IDsTnJnAosjpRld+tXbR1qtOw
MKymD+HGsAZqFRBjdhisG/ByQSaq/2CHFrQY/LSv+avcNd3SfcQCqQRyZnLngegE
Z7zC6OhKTcCnBXmM/WQeOpvYMPpRVQTziiTAVH50/mzyp0g/eN1qzpyQnc9geFQL
qupi4KLMY3s4R769lqJC6W4Gp2nW6x11v3CQk55dtssOsttboV+M1L1rihrDTI/R
ae9mnpMpTeU/sz4LDgo3NP07AUWRVX+48jZ0juCW28nFimfuq5P/TEghD+UECR9M
tk1JhmC5YGcanlQ6LhwM6CMxGRbil94oeaotZHZxv7m9M5SC14mk52XhEZw6JLcv
XNhorzIfXf6IVlavcEbPv+GQX8zCbNCSs1Rj5L2NFPMe9A8VL2EKtZmDhCIHUsbS
X8P1FgTeeg4nFHvEGfAvxfV+Q7uXMkyhbwH2pWuEH8+KPqhvPsPBfOQX8w9x5ceq
J3BJvUzuM+uIloypGnLgHqwskxBmn7SfoGCmEObLe1c7vBAX2ZBqcF7kQWzWelX1
/2peEpKrhf6KtAOC+wZ4TmQ3+1S71nn7HSNytPDMWZqfl/v+eMC7N4PtusOYFkiO
vf+jUw0OaKe9camZRmhfBeyVtSutBhoIaCNb2n0Rl6Q/RV/i4JhT9lhDSGs7MzBP
1LZ31nYGoouger2/xkkmDJi/eqf3In7Mn+kq5WXffHFEifixYqtQ6N5dS1kNDby+
HRI28hrTaSkJK6+DS/JxaapnqpZ3oCJNv5woB+/GUXX+OXvJFB29mGikue1dbdHW
fkPVe+y7gEn4pu5rmyNuqWjEd6PIIhr8+rsBpIvd6LR/OiUY2sKWxXkaFr4T4a+i
mSwJx16GMFBBi9OYdrik6C1sk5ighEcC7AbMvPWQeD6hHIQ1dqWPwwZCiHZjoyjA
PQmvLLH6Xwgm1HP2c3VOFo2csQ9prLSmRrJ8jvgVYTAxnLC9+3DSwwwKcrK8CTCA
xXS2mJD3rt+qfJg6KNP4gA7hnad2m9LIUVYmioU22iLgC+hAsUum2KnmGpzKgFD5
93afbCtapIYNlNGv8s8NGgVawtqt5+4GvI3iGRy17KH/5ttaIpyZbcmNJ7tfCscH
PFrMuzpo3jsnNNrKef05LH8NlRcLMLOEuqRNQaOj04y+LWzRySoX5tvfG0Pdg/pd
qehXAJqfSf3XfVom3D1hqENBYbUZXzYxIL5VYiTgYVURw3T8PJQ0KN29F1YiQxI/
ggHkA6F1hnWmFvdgAcvQwyfD+NCWLzxwn8KxBE4NMz4CoZHJN17w+k9VEfR3Qvql
rbasKKjgPj5w/eiXwgAeg6kLkRBYMgIS4rd2IevzrV6S5DyJGI3PFNAPGysYJHcR
u7IJWAIf2wLYU47D4B4iYLWlhoxFbDmwOHD/KcaNpcMG0TfUN5fM3S5R0xn4ai43
wg1vT+OZhjx20R/ADzy1FOUqqi9odYc4uODgzcswHFD/SDpT18SuGZx1eH1aCfmB
wdbPXpPy6BC2bWlD3LAhalSsEIUdnsvowDKIz4wot7aQ6Xw8GcXmlye6EAmqtk2w
LCNPIJK4X3pooekDa6o7NjoyufsndNIF3XK9k+s+fZlmCcp7wi4mAKuTZCPltplt
sQxMuMn/EHngq+KXLzfDfkihYrNlyW5wsDjymniqNyNrnmMtnJEr7Yy9GZfdEsJ4
ZrjOLBOn+D6lS4mZNNAJoI60VbSkZgo6P22CwIOaoQq3rggUA+luAUeOEdjSvEh2
Y+4U0ziLrYlOV4CkbpQ7QkyHBf4se0Z+Qp5x3W3ME/22adT0jGJpHldq9rPk9Pkc
ATm+PC4sZo20bQTB8zqjECg+2CaqZ1UYJGkxF8p38hfqfNehswpI2SRQD9YTo9pf
Dq4xzqhqMfBMl6y+8lKw03RDlISoUF7tj67sjEb8eQqH1GNbTjsk2RNmfOcQKTIu
wOaZemPzu1kBrC1cPT7kB6j72ZZAD33n1DmkGvNh5i7Rjro+FJkqtZKKElqgfwku
O4LZt2WPHNGafNMUFgosF/a9sfpb4Ra/f6FrqEWT30f+WwNDtaf7CUiw5Wx4Gmuw
ZfuVIH4min9fhUbRBPGPiXYKCbw+5LQ+ynqb8J0xcrLkiRNkeS0ERHOS+KB1CgLm
rjamkbWE/0TxGoZG92LL1xDMAgiOhRQBqymNew+g1N6fe0GuqB1D35p9D9HXrkFw
7tG2L1gJiGH9pKMaWzO07MuLn/GJehb6gQ+KXEmLDTo0OJGGxANRPh+uQfw70wr1
8J0LOZI4bHAVEoZXoplgBOAkcFH19+mbc4LfQ6DuEd4TAzr5PcI67Vxv96/veUwP
+74d4WQ4hy53+A0RD0UMQ2Q23IqfI99wiAV7IXu+IxCtYAgoxZKm0fWX6uiHbku7
J5ArjMgqw816ZsdyqIa/1xlH0D7KFz3KL3E/hfcDiLCf/U4X+R8Fu8IiyxyBnzWr
Z3o7XkKz7djWrgm7xafdoxHHz0TQ+O4CwnhdYWv0ajb+Sm/JdlxjgvxW+FPzXCIt
1G48foxuCOIgHgazPowelNUuYEsmLdkTGc8ClQGjsfn7Gyi8TwiPZOZ7//2aY+TW
qXwbKTqj5igxZ7ebabthgdZciIAj6hlrqb3xePUn5fgpQUXb6/xJJvlYJi/lgjfz
+y9M1/52bsruSzw3+5/HlYfS4lWsu65DoWNj7lhXiyvVNqGxyLDANZtJgubqBSg+
t9z6miJenOzugm4HSriPdV+XSsfaNCGTGgaaWDl8lvfHUJ/SGrMs1kq4033YykmG
dcE/jP6V9dGnBl7GT/nRhT0IDr4epFyL80rfBml2gIXU8w19q/do+yDtThFWSRAi
zegCchdgPfXpyaQiKJ8C8RkdZwpi0yQUF7oeyX7Vdm4jk55zRFvFLlcEjeqFbDeB
ZQzfdBFIJlytJLzkiv7JYgMVnD4ocAPeeXHKEScDiT7MOBtlkHE7n4vJFbwFXXQt
xhShPHLQh6oNWoXmfqx5JWlgR0wsIbVjOVUEdXa/AqLIri32KQ3y7VILNdiWFat4
/O4Nfw3naSuyQgaOQHIZ3mdAMo5SCvNf3DE/HW5r2qRftucy+kbo4Qkseaej2cUv
shOR+XpKX3YG3g3kMYRSV4Cj9rZ6fPPp0i/Cc10Ofcrr40f6DTGCMff99pqMZhSZ
WMKKxT7SU8Qb2kFGU1SC/SMRR4dJ9+y9ABM8mU2mXw2IeHxvJiztk/R2DLTpslHM
EV8KJjn0CAi7K39WrMWIPWE4hioLO4Ixk/SchOLHEZV4sNy8/JRa7guHxIFuKDVz
za393TaTMRzqEmj6E8YfRN6hC6c4loZe1jsz+71h6e0b/KTNOYHurzJ6amTtfi5s
u6u7Ao5JuWPG9wgybkX+BvYt+cT3xthu9gbHrkjibIJncbboT2Phb2muYbVsGWqT
GTdU0rVAiBwje4H4dUz5w8k3rR4AbELJbqXHtIVrLGftA7+NoluTyaFRpaXaamGQ
2tkhRxqmc52ZL/0m9R5VcePAcdlmC/BOZ39sR3DR7OCPzAsKZ1uRzawdA7Lju27u
/hfuv6JGEFH1RuIGguqSPv+iC1qWeh1ywQEiTU6VC5IFe7XySyqVR8ANM3f3jyWo
al8EiUNKD9AK3CzJynM7jBLm7cSsbu+OP9IJR+1S229//Uj4Bdr4VtYj7XLWAGWe
yNPfZYqdNpgl3mchu4CJDTOffoI+Qgc8Z/TWjU1LicLYmOkegKwgee9kWETZNo5y
EFItAjki10OU0YrWfmeXakhi3q3xLtIl1HMOOG8dd0xtU9uGt93HnorjBYsoR81l
V0OSM4DTOuajY+lWAT5WEq5VzuZcggwEEZl7vcY3nYWTwfftnbuetoLTbrXyqmzK
5mlw06eV8Hl0vBl6IXPpOtlnfYBfK8Wh3aeR1qHcSoe9kF3PRKZryzgG5EfRVgI/
TU5mgZ3+VJhKc9W6keywgYgZHXHiy2a7xJi4EtFZctzz63PVbN05OGzccJvlm+i2
ZnFbiraRnDlE8auo9A/utOcOqCmPeOCCgz0x6Y/Q18s8lXUkKDe14ratBs48LZm1
EWTXHYf8Nc3i2oMTgUsWt1pfBpLOfDXSjdyDUk5mLf7lVnHu6fYCwQlbTNcoPqLN
JkSu4SfSBlbkQD0OPoJftCXM599hldP9m48bZGxvIe9cQD0tNfrK4u63vMlR84Dl
NUz2F8A251G77HM59z/dljNkcIQzjo+cTN2TpQ1MAV5cm2uRh7wlzrkG9i0TywiT
p6cdt+wY3/ceWPb+lftcC/dJp6QVprsCeeE2ZivllnOVa7zYMSa+vnJdfeTzInmU
0PZ7DjPx0abIOBfMLlu/gEk2a/DS4WNN14HJr3OveVDj7V2HKipxjM0DGTboCJGK
eypsOzExwcOz/sqJpI0Tssf1aDShvMWt9llsBMA8LTTPuPslTBGDAQURV8TeZthY
lJQ7BJTf9UvlEcYtEiXIrqQ+1puvz+17akglgwUXcy4iK3rx5irF+1mteCi4IKO4
i3fTnVFtQpPxfJn8ywZbcMQ80AckcA8M6tIJSJ9HMFdAT+Kqt7EoqRWTBh/0PygN
tGkLLKMB4Ltb3laspJs5zhPR9SDhsRzN4e3XlDd7HrzDzITt5yVPkk7EdWUduMd9
xFhG0XyaEoVfs0UDGNRV+OnhcYuCbSa/2PnM85EGMFtSXfEsgpiHRhmaGRcitD2M
s3d3Csvj71uu0+S1252rKVo8G7NC7+HXmtdNpHXchjqBtUjqZI0eih+INRz0h/Ps
z6RveuUkYrYwNQjRdcfwD9IWQDDoqEMRrgAOK+tm853VQqg3kz1nPSz+9BXCWIIn
EriBU3EKg/aBmgYaaEYm4Avhe6YUDBR7FYWTLFynO8M6GApjcGnA74707yPaIvOT
U09BFx95iolgC8RV7Agr0j8InyA/uxgSxybwEIHQpaDFHl521yYbSNkISgxPmkNY
6XxyTujFjR7msbRkzoORgQ/1ax6TwvblS8x6OBXexHJCN3b2LQOfZZDqdPEM/Nbw
lZRUtKHlSzvuz9Q8s+PQ/38ZN5fUWwwyiCVh1/MroFq2RJBNaqAEJA8xDf3J8EZs
NE70+q5V4gAd6ML4iA6YPr0J8pvDL5YqPN0ZhlykPJcMtjm1AKCK97q8i/yfK7i0
j1bHb4KFAQJTIo+z680H5Ka/A/0WV5+lf12PVDVf+TY8VBwIaMY/Jqs4hGFaaATc
gAzKu4EQcYLbmRNqDMb8ZReZoVoG/d0aYYZAFdUoLOrBi3FfuaJHM9tXnIGK/OG9
LNft2MoDgt6kbjxutXlXRGCT12RZKOWcDseWwPXpnUxHs6nWIRX4d8K6dlv+ZnrM
/ib3hunTdX0yaV25aLeDvdJYLp0S6a8u5W7sBDw5vlsrHzxmCZaVfKbdSvDI2QpK
jPR1UB0b2ObKOGQkIN/0ARgyj241px8jCM+DdS/NXoxw7+KpK8P0ZlTvhiKh8Xir
Hm6nFmWBB6/UmohGhWnMmsYQ8KJJ/DPlrYPhZTCS5EiSzw5v16HQ2HbJmLgaETS0
R03XJ7rQNwRr0/H7nufbDV/7boYk9b5apbsnBkG5mTDUeyI0bMwq35Zyp+Jn3C8r
PSiQhjmmXmy6QV1BqacBuXvXMKixZ/2NCuClqBuxRhYyV7EV9BE1knQfCkuc5FD9
PWaMHswINj7IkeVdfI4hT57naissH492GbvtHm+H2oONtFifw2oVr5BD+svK+Q5w
zRmryb5ineEK0yTsgIhlHco7rk/s81vOrCO0g43dx3DzQIG+7R3RyAipXEF4G2f5
Fwmoc50vKsFxudVgjfI6jamqJYKIfqtndYiu53bucXiwfDLyQULciFbt38YLoA+s
+vYG4n5QAw7jhxwpZt4QEYRW1ghpV2G5BYnHfLdNL8+6YnBAzHUDbB7yll1uIqu8
bfofNeegKBbXD7dR7r4p6wnMjCj2QslJs/W+NpsobfKMgEQToNEsoS8EpC4hDwcf
yjixhPj2i0vzpyU4DOS+N9TQ9VxsXugqVPouKJbtKZDDNH7BO7udqECrn07gWlZl
+Nhfcx/Z2JB5beUdQnHDeX6Xmm82zFc0jWDjKcw133NgZZX/jwR4bEG+J21NtG9C
zE8mEM+G40rSPcaJ+YXN+mOTxgEV9K/d15xQZ1p0KWt1iCld7seKSCs7QeGCNQ7P
2gtSrJXXTEev6FtU4l3T0BDu6ZS48ZIrTVrsVrAJypZQ470ZTmIW1a1+NWsRARNp
19dyZ9QM97jx6Y6WwZCKkj72GQh4R/YHuQKbcN7Hs+J+XrBGvBnK0Fxl2q6UVVra
UkrPErCrp+E1IXX8yDwdsjvbIkHXgNsV4oH7ZExVuvxFI54OsRh5z9yNIvlTee1+
sJanCzBtpG0liagAElGQ8zsGej1vvHRefKsygDQZwww8kuGfA0ZeU1Kael9K0YNS
LEMMxH/nyyvlusyR6Jrdk5uki3PJKx3L5A7tGWDxxE4lGdLeuKOIk9sF72O3zcR5
Sqoxl+Whp5k+Xk96phWrDB9VbO+2eADDk1VhXnFeXiX6RxYa24CkBLw8xb93nDGv
sFmboF7bBnFm5V3IxGuwZUIAAnNG8U0Mqz8qaUpy4bgKPUVC6qm+wWA0PZzptEzt
z8/Famh4eUhSxq1mj0fATwKEljkklLSQLz0aD0o98nqmb87tDV+861dXUpENvQQJ
nIuinAJZvHuKIV5f1y/LJJVy7c+gvsb9VqYIfnf+1YiwkQhztd0d6k71NwvkE03d
/+pJjJGEdSgoPFN7dwQFWOfa+eJLIiAMyyW6ps8Vqjhh3cBi1XR4F9yoCyhiXPTT
PJTVbzoKcRWq2eBQoUcVQwJDSHFdUpZ/lyQIABd7rGK7bY5p5IUqyrMlYfbguwHM
Ozr0V3UNkLVl4vmLFQocQrfnICiGXGDX9cmkP6xT3XMcfU+0rwaeWQi/BdNOcaz4
TMwITbKslNZckiWS3znJgdkfkWQLwr9e7GOIsb4keUfx7nb9zUgsRXw1PrLhjlVI
pNhKcdHWLxr0Db8FebgTyvITxKFS4fL7AePp5vmGCqwf+Nq0YdxdJfHxDCzsY79C
zXe5+VBszs1BrxJ8unasyZQmgM8dgOWSp9WBMZjxKNk2cLjkJzINMTBvsghqSxFu
h28PqDiGKkEL0ZPMfJLOnFNDqFRZUS4leK4YBGdDzuxvlMwwZGFeitDY18NZKfHT
GGK9ZgJfQS2oyWqvqsJwoSGAmKkxj27aN48u+mp/PMEHiF71d2Zhy2G6eoK7N3ef
NSZdArQ8jxbkENFAiILy/qiUDCGvljaSZU4+LMKgvLtwAT6KsFTj6YhTjdSWijF7
5BAUCH63AdT7mZMOdXpDnth+oh0IaLLiEQAMCh6mrVQGYyfq2vH5Z4KhGmQa47tA
JCkj1AzIqJ9gj8mIuxN/OGRK2VMm0NOcniYY4REeIjovk3cufqhyDzfiATRupd6R
yiCKYkdXqyY5UhMXAKieWmjkwrbSfvNpCatv6odXvS2WEtCN22BoZOt1MNz+4KDn
3k90sE93QHJSrUO6WokWUil9SU1vpzaXNmlqLhOgyQnEnQ360ne5W2gx6GvCM/Ih
qs/72FytoYNYEMC4bNtSTsIil2Y4jO6A24OgWyE1BKJjeO+h/zH8QOSEtc51e9Oj
KWSy3sus1mQVvxxA2n7Q2W+vrrnDt+BjTW6OsELUSzGgBqjjB9TEfeJGCohxVQ79
yXk6+tRiV2uH+Vt1ltTcjnlG8UpHiqr04XL7lhiHrArJ+li7MtQSxH8k/3RNUMcr
VreQtt+3qaB275jHaGs7pIqPmXxXnrcUDLGpnPsz/ljxx+ndXJ6OuCc/N50E3m8g
zCRTxphjSxRGEPf/gCKJxcRSU6Kee0FdJIOI580BgNo4Jb+/U6gXcC/vs2DtT4K5
Ctd0wmsGaIdpqOwZOlouas4CynlxJlDc9Skkyd5Xyc+UczBzS7IJoMCKe6CIwIfD
by5RJCBwjBZYjJv7OGTodPRBbf8/380VfCvO3oX9H6eYkDy0TqJ+dQMniDtMS4kl
1jVclDNazM7ax8Kr/qSAre7UfUIhsRaxLTflA1mV6k2FOLzLxJjdHbr3KzCASBvA
bOe834pT2p9c9rVhGaWeFHtdLsz9txFNhEyJ9vifqT3VmmPmv5qRKYNK6EeDHSGB
f1zuHxYCNzp9kJgoicv9bU2WOJVQ8FvbAYUheKEg4LFbk7Tob8sk/FAXu5BYIb3r
Rz701Kn8F2g7xBs5mlSLYQVxQ7v6ya+RGo+rtS75XrkYJpbmQmaprZDkFSoZaEuG
a+HlcFufnoOlFqNrokceXhNSoYDTSx+WjI6Tf1O/vzG4Lh1EuC4/IZlW5elYVZuf
U2LCjkUk2XohKcbJNSQdlRznzL7nfa9J2DQOhN4Pxlp1CYQygsHM7nN2cLVYO/lP
bYzHWeDsRFMyy7NCCmhZStUfxMRDxKY25SQALwKxBpYqtv1daMmjgqnZlArvw8nQ
LSwTIyHRNVwEXTcz13ADx0YzsSNAnDpJTB9yVk0VZa8ekjKal9J65s3LUvrnto18
DwaEgXhROEllhR0NTdf81GGHB+9dpoIbimObRThPsMn/JHdJS7v6tuyUIKyxI7yl
TPic6918MArZfDoisxtvpwnS9EXj2uD5MmFrKbNQSAIYX2hy9WtV/l9V6qwhZ7Sz
AZMjUlsZYVxx7ciYZIFt1KKq6i/wLnxibCj6nvYdikAYaslWviEAM++fTShtzWf1
2IIMNIi9j0FuNPOvqGGOtBihWuWxGAu4LzLjJjd6UZDHLg5CAxx8M0nNSb9fDS7K
ExE3GSrVI3jkmYzIo2B0NUKdx38rM8c3czfOxcXljOABsOyu9mmXpq+NUO2p/YJC
/+EhetCZGwNmh8PFwfTYJmetHcSlf2i6gpL1FcoN3jmdmaXSl3LUb8QDW++mSsL5
rLMvNub9XUrND+oarRkuD0A+6JqhyHEcQeg9/IvKUyTjrb82dCpEC3kBUsS6WqcS
zX/mXa7ssT9fhEFQFOvDbEWUabFvzuK5loplAG3bT5mI2B4CL2edeetQMCLF/PoK
G/pc9GRz2vW4Wai6NLjoun93bfh5OiRcbFsu4P2+GgHMJxVu8LQZdnQ2PVRYjWCu
B1455hsWUfRVUDLgCh3IVdNDSmNWzJ1A1QvsYqVzHxG+hnmIgKMdkRLNOEhy8PVw
DE6uH8SxLwvD4YmFD6ee2lFyQnoDmgWpzBhfyhJmqu56mbqUlGU9iRtDMHLUNJ8f
ujMc0BKoBvLlyfRPsG01DR1Ijr2X4vSJ5pyclVQdtG2Q3XD8cpKLuquGAThFO9wW
kUJYYB5euJ+yYkGnxxDzro3EERN7kJuUBk7kt11UnVNL8vn6JBGM+HgLCCh7uiWf
4WyS2X8um4WC9XsauxkEITbOJ5iq+aiW6Q2G1ieVJmNWD/BUDKi4iB9r3/PAnO2v
5z95AqTGPn2qtujemLJzr6k+mU9iP+xKiiQT7mkvVi5wSICsLxQZYuYWEOMKGXvH
uEMvsOh1Qjx1GDTAWyI1IuvJVYkkP6I76n0fvsl4l5HfrmymyANXZw4ryjLQy92h
YFybSKxOxq3LrJfr2iky5XHpzRcTBKxuoNgWUeoZChvrf8wlsvLKk/gAFBWoEUlZ
S4qGflb2B+vy1/v7q/v1PRQgARu82B4E2RGICNcZnE02M3kzSSHUPYL0kzLDGcVh
V2590p/IDragoiBITuXKmIc2LY1mas576lZcdLOydHUfdtMQj7K2esMuTECWoPc1
ffSlZdfuKpAcCfkV7CYl266XrInP4Xdmh/Ldnv4sahT5tVcGezvR6gGtXfHSWTpI
wLw0i7TycreknQq1FRxkjmwo3zevN7SiNiYy9n6cHic7erRLMPM3Hy/oKcQOZpyq
vU9aPNsCTpcRbKY9O7yaKVS3uZYsgFQtYRr1zBk9kF/ZIWJeq120+dusaX8fN6jM
eAPYLZDxD+qllJ+OqKX3w3jIdgclY/NaekdRo7fcy2hkAQ+stJRQEs85wP+h7Evy
QorLnIk/dHHtHehfYmvu5xmAtavpEJC30Nq4eXZuM+4pxhHARqW247F7sqaPesNU
AdUIpS3EwiZAgnd1KBD/5El2OAsY8txmbx7VqHsuClXowuzNn/UDPI27x83LhPyS
rM1OqdwWlxAMmogrYWh813kGbUsLgzWWm3qN0JuKcKcxnrJjS83zb+iPPvBVhn/n
aLO8pzSESMNWSXdxmO9xmpeoODhhFpJV8GeMgnrfdqbvO/AeGvCh1pvILmCdK4BY
pRyh1gKlWZ0Tz8AT9zub0lEoNdiQpeaj8UhOsTPHNJfxuLnyx6d3YXhULtyCY94+
/X/SgfceoY6kXTwPjPeIh+foq6/3lAoQVXi5Fu/lnbjhQC73LY3VmfpGqS4f0UK0
531+ls153fyAtFQiE2ChjPhuvv2Z/TVmVNkc8mIi2Er6ZTZYmDdCLGIY/Ff++6lI
0I6WXrUVVHHNPPnOLbzO22roD/o2R1l7zuZuj/fA9+XMmIcsSL6Xz1RoqJ0tz0E+
W4YrYbSPrDI8PKMGV4e2VHV9fjfKpjJrNI1KurWOPHjtnrDE/yLQNi8rmBByWBIs
BZe1x25EMo1yJdSxfYiEVlLMWxZoBmK2qs6S64jPyES7L7Yjr1XLA496aCzm+KPZ
U1G7qXrm1YPnXNSwRrXWgYrbGpyJQOOQ9iGZntn2U/L6IKOiI7M889r5YWEAhC85
RLcuntCm6vr/3OYKEptHiqmDaZ2VhJTdFy9ADiZlFd8bu2aQMFWtbyKTco/o8i9t
xY5e6cXH0FYWDWoLYLhtdQyaECKQLMrOKaJg/P0gkc0kIat2smPVAfJTd5iwEyNL
9kpcjYOg5H1vJa+RSN/HlJVXhZg19nIqTygWPV1OARvX4aozQpVJA9s7NYwsyv6g
A/6+YWuhbyiwDolBYr3hX4iXIKd99ba2vh3UxYvXoOUdfu2RE4hbY2mnzXD68f6p
39KCOsNAk58dMkSCRsiKMBCMJU2Ou8D689LlhI8xQrvXqfSf2oWYQurhL0eLlF4j
IhoBfplkPucTFOHDEmZTLmS2PHEhil3rMjLhcFyRZVwmRQAPDQNBXLgKUqCthjQy
BIgSfb3xcfASGv7V9ClEqSAWEDeoJVInB0WZa0MjPxFSfZuM/zCZkQB+Q6U35Upa
yBcG3uwUM1oIQNPnGgsS3LPaqOnKza+GD/Pk/5ttrjJzl/6rXt93rl1hqGb4CmBI
Gz/eCYSfcOW7f8Z1AS5HLdyVGNjvlxFUmha35vKnUREI1bpCljjmZ2OeRaGlvNuf
jwiD3G19yjN6c/gRQaZjjigE6rHC9p4Ox/P4FPCZAEjPBojN3a2HwvrI+dRwY/a4
sTQh0W1LrshMAKaY48b+KSFUgZusMSZsB2g/d2zGmEtqu6SXnzhaB/bxRBLR3Bfy
AaL8CyP0kr2/x18Kq8PjevB2lPmGq8/722GSz4yqagRuDmb7eS19mzJ/d5mxLEfH
XIprCEcMfPtOfL45WtPDbX0tOY3P9NIms411QtAgOx+u31F1bD2Hnx+8V1WWfWO1
8KpIDtGX5Oxp1vFUckLlDOQXopID74jrmyG9g0ZbwKSzAL7vkTTMkbL3o9fsVxNU
MoZJ0UaGgIh0PS/diKasaicE0tuYDweJfVFnUpHIVtI89WUxeyLSvtsk2sVBE2za
mdnESqaL8CYgwVLK7oi4SXYct7LTZqliJDlBBVFzNW5doXPuMHtZXMgkvy7dRWQe
nltcbkS8Vmo79DlwXJBW2qmibu8v0kReBGLlUXSaoRGyeCaxYJ9AGdtic8Ghaja0
Ex55NAijlA40ju/JEkFI9n8D17nWX7mbVeZnRse3N7/PkyOFs++Sn3QUCRzsu5RC
+9x/NGksxK+OlaM7X1GJeC3t9woJmIcysoNqqRVASQENWZrBbvXTq0hAl5FPgKbl
NSGdtOpKkpYE6F32YWGTGdl4nCA7v06sRn0rmIzlQpzzZsL69vpdzMk+6Rh9SV7o
Nq7Y1XAY4w5lkoOlTBykPKR3xDv0Rxr0cUYUOxzpR8qUlxFGa/H1eGOpHICYyDc8
tb1QWqTs7N2xgsM+haRwyaCxcshba6UD45KbI6o0/4POPyxTIhPBKQc9sYILhCzA
439TeZIMwkWT3PS+JTB2QNU+dDhxIb1/GWkORXtjFw/+xR18OaAGgI1DL1FwpWXU
MHW8nV42sfnrYn3tJ/BmLMyeaJng6YmfJ8AX5fOgIiGgw8PIToPMQh5bJwPYbare
/7VaoWjUO/GpXauV1lCYskrvr1jMTGjHpMGAPki4jXyMCZD/pLMRV7yc9MHoEIju
wLI0vQb7cHf+VKyLxpPRYLDkZvS+xkvp37Z+cY18NXqmeUtT0QfJn8ZwlMoGKx8y
d2Q7jtSnsxTCGYin1S+f+gOgXJAr4cZbc7SVBomFEifs1hLeKi0zGw6hoEuBgC7N
gqz2sX9CpKAsg8gIKvkNL6BQzNbFVhjruiMhLaW12SoYPagwU6lvCBYteu7q363I
w28SEh4oMZ0+Nnskd2g51jZ9bTUU6YuMXsq2NCsmzestuYyPq/0tESWG7W3ZNHp5
Tm1Rs4vB9xhw/L4N4bJdjml0VIsIDqY/1BZRJ9h1xEULW6dNMl1cjEUwwY7KsqKf
D+yDbWBwKpRzmsRaKtogVx9C8w9gDiB1sApGIqjw1AUCbJ5WbBwx7hE43rEpeM9B
Zpd3sWPd0p6Hp6+yX6n2SbEhngI5A8Hfr4kMWCoYV64e8Xo6BVcR5Hahl/2h21x1
KVtB4wPjIUYZTFejlnUAMIJ3alE0Wsg9zIkklgjK4xBz0soAWCIyBv8Q0XuVAkKz
61vdC125rfrxsO4e59GBU/e2caMPyO0T+68fOH3u4btVV+NSmN3p3tQx4B3n+EVg
deVlSB8Ryop1lxXbtJOdxvMV/n8Ofikrwa8r7yEkKwhPkY9SCTIhsKI+uTqgK+0Z
bORrsczkfCO6HaPnJ9GXgLrz2OAlqiZj3OB4HoSKBDCYFBf5QWXg0DTl+zJBYEtG
GfpsWJo9+zt1/Dym985ZWjG68FAs23KUkZ1G6YC82/kbq1T+NsG1PxnO3CmMirYE
qtvTgNQ8XwFEolt3Tm+e1XgUL+yxZRrKynHnV/NRht18NgQzzdP4zoLHs5XeThKx
YHXG7A9JtTaozTPEpkM9oziKd2/Rr3Q3/lRfrdxN5kWDL8hZsdWDibzYRJOAKvG2
7gk3YKVpIWHq2O1JOBF1FV/qW/nuu6H+O71kCeIPpEfOs0CR+1bURwsuaQNFyTUb
lb663F61Gthkr+Fhi0IBYbRgvfSn037W5ZByCLmqUOzw5csOpPcyP94SmWclRxXF
hUFti2ZsUjI3Y7u2jvW3DEMuHkD7gZNRnzQrJ1mtDKERBCLQfhlK+XEDMSYhXJ4D
k2yzmBIJ/gZBs6n48tPgNC1NlTWPWy7uryCxlKgg1BQs1NpX+Bp4KCYQHypxpUQd
U17EeTmJwIbK3cTXMYlbHRSfn4+pwcBf66MeGdJC1G8UFI9tHzj0RmS1LBkWhCSU
gy/iB15oxF9Rt3A2jq8bexICpxqV57aqlOvfmWIi1j9/d0QGFI7qhq0bYNyjqhSP
cG8N497xqBd3UI/7QA12XgVegbUsOMu9/TRPEFf1osMeviCEHYPJMQOB5fHamS3D
ZbUenCVESM/vAF3TeKhT9c+zJWkBvssXbZ51mmUStc+jvhxVHxXGAyOeDCn9sppg
aGBBSWbtUkheiqstC30SO/oHXOts9QmIb6Urqap4I+LoZMHEsOkPCCAGaQW4xfo3
+F14Xgrh+rifrRvae3gwEiiu/kqa3DYd1Pz1lQo3WFM4NA85VEeU1J+wHvux6tN8
KSnQ9+BxSoiH2KW4y04RhvQ/jFU/LYG8oHkQeOcJ7HwQDUyzcd061bsUqt2bNA8t
EtMN6NuVREw2Wv5w6Y+dzWPtnrP0HwlMuBnzAj/x7VG4kYmSQ9e/wjBg4Rcs5J1J
iwcgSgN9oRGfpwwkq6GSHO6LtzMtHE8MAmyJzF/DOCvqyvpKHKDFs44LnCPxe9np
xDnxJQRvK5o16kPsAPsHf26J//ewFTecbWt8Ya9/Uxv633rcMjXXMu27gmN6tHOq
OXNXF2VTNtU4WbIvpRHPBK5MXKULtrK0thcKK1e/xJbxsZez0/TVEwdvANbbPIqt
Taf7iODRYad33bws2dkJ2oKIlsByk3KYxSZCFvQum2NId9ytH78muZ7RPCLBODEx
V/h2gqFTzSH0eVdupxe5g1RtQwPKwofb/7qao8lGlPO+u8EqjP/3JqGdS5VqzU5J
vRhXv8x9WEbvN93T9YeuVYBSDZYg9IEV012ZYYZSjDeHWXtcSIFPx9GduHMsab4G
03ky5MFD89uuMXnmRXra6CxwN9jZwVFrqjVTjog6aPxe1Wc6BzmuMyGpWrKK3nME
znpj9ypK588wyGEwtXT+yT5LKbjBXZifZWALEeLuT38GjWinyD+eUPEQubk1/vDy
mUcIKdvp0nNuJIRG9EmynPp2YqZZ6yEtlvVxfPBYuUC5sP/N//SH4uLJY04bLX/0
gsavjD+Y7M4N2ldnvRs63QigQ6OMPazV/cTPu/X8Kw7qpIN8td6i5fH64raHif9e
oqNmToCExoblIbN+LQ0MxqxGNfoOtRb2DS0q4rhxQ+Cj3sP8HQGxBUxRW5sAUee7
QQbDf6aDyXUNVHRB+mkM+Gc74EY6griEsnuYBcsLAbzTUQXrktFQPBH/+VWow9A3
WgU5bjFYL3SsXAzvqIrvuuN36tNyERv/6PiGF+zjzEabqQ2VVGa6VO/s4OtTB0rN
VtWvBKVJjNjmMfPb/AsvTgcldYGuFySHfmeSX8EqEnwT/Q0zRw4EkT1RAllNUXH8
hVJPqch38gGsUgwDByfItvHyuPhrvyF81olMX3+2Fv9L/yLVUzY12mIO2pwpRLN9
guOyfHdyGvspqJocqpMrAKsFbMz4kq7rHKPTIi27uOmENfox6KTkr56SqMwLZ04s
/wvTjEnhvW9IvIhEMgwPosRsSbggYEXV+NTdEvIL5CvtEKnknC+nCEQqu9rPEuGQ
Bk/9JcAJzASqRkoVZuoPrji3MUqyct9BPwJI/PnQ85GYT4vEUCM/J72Xx1yj6CrL
s/TeUVkk24Dzkrk6X+J4v3v/C7YHFsIoX2BimntIFnv5qUTyAbyBkYvKeTNr6lDy
J8rURKXGmLxFs4w2b1p+H/hyoZDZFol6ZLYhoYz/h8l6GsWaCL6eFqsHzWJCjbrw
zNTSzJBmR5qUTkTfMr4UgOd7P0s1NpiazAXyyaGRu/OUemjCcGg5VMVijZ6gMSpI
vl+7SjvEgi+1zVy0J/hmEMrTGV38KWpPUvs0thjuL7/v0FYdjUbyY9sxIwGvrgKU
7+SJEmBBojW6Dm/bkdiu5q625JOfbgeK4FNXKlOuteog+HwGDkkoCgQz/SU6NCK+
a+SE0/gCi7KHnNj2VSvvokfq6kJ/Ec8hzxe2iVO9o+Quf5bVD30czLWouFFh8Qd6
0y19XXWFnIDDPw/SoqtN8aDkUA6ojNDyB7bGjGCuQ9513U0XQM94VP8DBvY++wvu
5O08A11tt25b/gSROWeK9aYih5hyaVrAEEPuJxvR58BKf4nezq7WbRQUslpZMcfy
DrG/te6y24UtjRgU41JOgAwPIwo45g2phYT9UASa3hY2vKZo6LrkZ4ts9uMyQqma
8+vgA6BFV01FCRit3QyGkwaPadDbMLFeqBNUxxj2DdePhto7YbvJ49lOKCe0qVMB
WHSR5YLi0MVB+lVG0GOAPEnII67yt+JzVSPMVj8WRoOx0+fUEZJD1XFY6sbziUfj
h2R4nOyKje9s6tM1MgyCQtGNJnpTImT9QrJWwksa9fbcFtGPg6rxpf3rsvZOGYJi
3mw4OHZixMwRaR6XKsQDzOKoxLVAOjAPKdT7ZbmmIRWxjyFlYRVDLeoecbA2RCF5
CFfGnavaeMTCN7FxY4Qn6nXxWN1Mrg23ITG8pMqGlN0gEusCX9bDGYKHv6tpZBMU
uBuLcPG56/0zSrVsKtXW6KjnG2GrcJp1dhaUFeD2URr2F44zI/LouYgXRo1OyxKl
vrHGnDcAbE6PSXgAp4zkRhmlliPYdzbbqY+4dXQgF5PzIxgknys64GJFi+bdwrPd
Jf0rrfPudwjaj3C9r3hPsNYE5sCxEBYPt66Yr1g5zGROJRQt0yKVWchmwsDgGWid
ASANYfF7x4ZRK9uF2/svFTqN77q3niU0sEkIepC1TbHLOLgJwwlKQfu/movGVHS9
ZnJLvEwt6KuWTd0YgsrqgaHld4AU5fxsoMKHE9IryM+vT+obZWjpIhWFE6QfbR24
z6R0FQc36xS5MTOwhQJgFrUPFoOwMMp/k1SXvRcpRv3upYYbag9wXBdO7ZTxKeaT
AtuUO7wkxNDZS8xI4ZvilDGIek0BuA/NCkDJC4yLR8wFiYpHUMLSFLzHkOvDcXDk
f9d+sCjv7lef2OYrjn84xhXB9aEkvKd/3iifr3Q6uFYxhIGpBxQn1+BNRUrcJ0Rs
swLS09ULIMzjdezoM6roLUCyUsIbMtpZVEFn42vP/19IiZK5gGub3wAp9PrLvBlR
dN+mKs82Py0zcoY2SrubbmMrNy/kb2QlB+T6JFDIjK0wdgK4yY8LrMnz+PaY+a0P
2qmgd6+wXvwGo/43K25v8+cuLiyV8raNdb2mrCe90FpOHcek1RRpWtI/oGOMGnnU
ZG96zANneS0zTo7M16hAmf4Wu11afyw+RPpbxsJVTW0FB66AJUBVHKh+e3H+Nhdc
EqKOJrTZ1KSlxS2sAsnne2u0MYVHQOjuk1GTTR3E9nt5ygVkLNrqS0dVYDWmk8u9
Ior9ozqZdfUwkzlewkHB35Dr/A8hIFKZbIbFbtI8SLf2knOKVvQ4VxOUv9mhK+e3
MzS4G1qt9aNDnhmgd1kpuTNUwtoiqV77TgIrous2ak5uC0tgPX4NAmelRteglEoq
fKzlekwNRBNjLJiG3lsCwsW54cX85gxMaSL8k83stciW/EOULqeJ/uB1khlQPKVZ
6DYCT2gfD9GpImNo9TFAILnGTHZM6631vyp7Y6/5wl30EannlGwbK3Zs20l7mkt5
7ZZUqkVZKpEOnX+6L8MsqKC1mnmeXTfYz7GQlNlSQ35uOFIpJpmQztTTkxpJvBXZ
D+fA+9KQAO9oudzVWFII0kNEBHZgq2qRhlR7bcr6GZ4XInQcbxt9YXU8DIrHcDXW
9u2NJEWxRMcIeTnf67TDWIjaTswtWP/p/GxA+o1jF9BYYfSNrWQYfNJlxywxljgT
WBktS7/aYz3uC974SaSUuudr4ap3Hd7TmMPGbymisqBTQ96qYQ0ALamQR6zL7JaF
vgnsHZPmQcsH0ByIloGMQ3z32TH+ZL/5xT5aVQg1drlIuXvyl41lARsAmD+7YhSh
2YfOba5fT2yk+p0bSas6oU3tKc/dlbt0NbhPE4VIvdTdSDJA4ANMzpSK9daFjZQx
W2xiYKzwzG9/9vaL81b6Tz6sRBJXIDdhPChvktFh+PkFgmq9o8FWPsmBOS+EHCd/
AuihdNQFotl6Z4YyJNsBiBn/Pou2YscflARQtjahlbA8hVcyDsI4YbvA1arXADl3
yHrX4mHfEpv6ZxlRWng9yYdQZdvgzcL2BLG2YIRiYTOa2lAwLdXt/5zr9T0HQshL
4GHecm29pmkg9FHv9r8WegiGEQOSKUzFx4kavvmwTZn6FdF3Stg5XZcxK1mZCZK9
XfDLKbsOOIwYPpPln+8PT0t5i3MkcYF/V2T2FWPnO5gRXhzkiDA27iQ69kYDWTi8
+0S5Kj65CLDnaAiXhEnNTSvQxrrWMV53bhY/xVJqASFOiibXU42LOtvaeppi2mNU
d8XHxxS8h2hfSkQMj2kpUpNTJ4lm2LXLWOTYw1kT4RQ/WnzMeLb0+Lg2Hpkmgal1
56THQMptDrxeAvaioT/W86TqwCELyvyRJhOzeavgQpLHeffW/ggxJb9cdrVCb331
jRhc2mVnmdGq/wzdWkDLgCWBYiJt+6ngywQ/mprawUPFP8Z7aRLEsXw2w1+7S+dN
9yBDBJM75NhxkbW5NhTwK8CjaapEku7gUp41yREW1Cn1Aut6mQ3Fnt1CVlH4BUsM
gHCnl+6bdaLJ254gYEhE438BdGWKaDAxXQmrEDWKwFBoTHhg81EiUQH+jEsJvxdI
8scgYBykHPyiQEWyTi8/akiIsLpoMB2uRdazyUeE7m4nLjtTm8H13ZMQYiXSmXFd
lfgSzuya6Gtn0fZEQ5edKMVAgBKP+z93Q2C2x9+aEr3u7PfvVwm4Os+LjscLpBF4
+hQGGcpw6sxVlRhBs2q3Yv9w18bI6GehG+DIh9Oy4VAX5rzHtolwF2CU4D5E0SbP
/oIPE/OOOYBxBtn/Z8PwtxS384/YxK2KLR6WRCAqyhAAuP5fV6KeLKJFCE0slJ1H
mVCrQRimM+e1OF/onJ1f6Ko+KgH8qlQqqgATmVx2/ng0iEe4dyue0/28wArC5sCY
rxtF+nLuVoqyCu0GEQ9L6hH6eOtXbHiwllgfd11UYiVZxi0mFQGTTNZumQPFzNPG
lujTCiUt9vk9lV7sCpneqnopbpRRmIXQ09mWVr1MsPtKP9+r1TtcYbdXliFU19FQ
Cjlr2Q3wAWPUXp78pDIqcP0FzrqVIxnuAegV+6h6YM/fq/gisdIrop80gCulLNos
1GKj42YmZSJVMUdm5fu2YgtpMBDjbxMMvepYPDoF0Fwf4brhHGnzReqNxAvO9wi+
RjycgpC4lmTQvLhhDQGTP0IYTF9qs0CkV2UZZUwjBbrvLDeR2cE6kQDbNiGI+Ilt
zGzr8gWKh/ieVcDHEfA+2YGvkYJ/rp2Q6QBEvUjv2d/6vCrvy4KUeMHmxkRyx6v0
fqX/Tl4OPAigrE8nGXovhp/9JfIZphL+eyGr/bCCc7M038dK0h4awhPAWaRT2kR/
I4DEHTVLReQe8Y7kb9EaiFQ1QGxnQWw2wCkNfQIGLgrnqLwdO2IdTVprGYqArRad
DHnuCYQoxtDatqqo+nUxthYFks8JBIHDUz4zriUCEK3F0CNB7RwtlmhL6K1M7NiL
g+DB4pq7MfZbp2uQJ5tsg9vhqhVMr9lW1AZ/xSYfOjN+nVlpROzRykureryv0k4o
VZvPV11xi2dGNpU2UWMqgWl/SLx+QoKz136qNH9ixQSWyW4q4e7i+LTu1uHGiPf2
UowowDwp3F4GuCOmgIc1Hlv/hVMGPKcnChFUFe+eLu4hqMbu22x4SVuK7eQudOgE
ZNjx+l+FKdA0R9i+o6xhQccT4MqqNvZGDXqICoEQ77lPBuJtmdXd3KcTh+86J49R
kluNRLyQhlk9mL660JuuIVl6Ia7U0Cri48NI9bXuezlwxotwQy8MfbeoQIvxxlSr
b9hpT/WdRfw0E0jy+0NFantHwZpzqTFd/Pekfaf7DkwMgvvBnq1WVynNB2RzODQr
qMVg83VzgSSyeRkU73tWc1rvhBZFzV2uuoKqOKY50JhPtsm+kq2MDhW6WXUynakH
hOaWUO1tVXnJFJHrGnSqcN9tXV9UraJQZJmtZnN32tWzllB4MblslsQxWLvQDAe8
k8fuM88vSndbsZ/wZulir8RfCs0cPV4WrzsN9zs+Ko8QOSanK8kVhrJlueamKwtk
pumGwQjOjG/lzof67f2y4shYS9TBh8n6ifzcx8MRYNTnBAJxr52ULmr1Kohw/2uF
WTetXW1Aua5yh5OgpcwO3CbQY4LpWbCpGlROWPnr2qcx9Fzx4WvTWQ9SWr1YHtwn
KC5xII+DlhskxykDEc8BsUybNeGEdgpXCZk9UbuAHm1kMNYdB/vbiR//zc9e9QfD
kGiTqN/b9yv2CqXgViyTWFgEsf1cwnXpoypUnb4S8s14D2NeG6wdhHDGf8+9jBVq
LfayAalKQEsAoq6cpqpDEd2GcyIAz+fSKiRZXKdho4BHE//lJ0vmCDBTNLg5RVph
tVD1Yc6N1K6MU3V8JzDaV2ScoFvFQUmZIe31JCzAkIicrRz5jkdLrbRE/WDoCILT
ejwyP7z4UawRmIc+wQSNdVBEiHIxXYbCcLum0Tnhv2I4phhDOROggQC1gtJ9ynns
xDgpn8vXvV5qrPx6jrTFy2HQfpm8MScv2vj7NVqKMlcYWHu5LJZsF7Yc/3wq2U2Q
XrAA67ePWesa2plUbPIrFLzkQ4XEHeHh1EmqhOwQeocsad82+7kjV/n9MzWi56I5
HJaFhH3ds+i5ZW6dZSRQEDybeWqf0WAGFbi1F7dL2GzPw0ztLCY6FzDcfNHMzE5w
9muBg3pY+q/7WFP2hNJ6pAewTawyJ7FAMwMfw1hSHYs8/TeefidFenM45rSZkG78
keQy4lpnQxZV//4JiXuE+aQJMe/Rg33/6lojz3L9XWJ6uYqL1+GU4qztGy04JOIl
8b+2dQo2IvZkjsO14wnW7rgFYCukhj5521CRUl8z3+FvJhJaPuC6OBMUGrgep6IU
7D+rODGOU/qWL57Zo1VgKbCoRdqUvU0diz8IlCtvTyqPUHeMTTuvrqYZexqnAAzN
NSehdgCfQUazgaLWqbmixtSKcQd6l7D4/b+ZYshsbTmoewwOr72rSjha4eJDJWE9
7+oPzF0O1d/eUiXEgOjPSpCrVAqqIol+eVVRmCrU0EGQpw7EDt8NSZu9EoZwCDb8
N9KzcxltORLohthHNnyAlbg5IrDKkO6R+cUYooSqELsFzEawD6gZ4mlLg4edibWr
XS9Zkmg2dD7rUW9yYr2acLlAZYrylj0+qfHIBCoSA/a+E9WwKn1vA4vZRpuJGdbH
eyiv8rUpVXVUAc7JX4WH8sKNBmRURTRRdN0UsHDfky7Ebw/vg77XnX+j5HsHHPnk
hHA1KM5T2tNg8fh2aEjZ8MJtrS4jhezl1Ts3X8/X+ECbhmpQzSfpVud0Gh5bS1z7
n7D6DliOAF8XTrQzE/u9e0u4Pd5NvoMEZWhnY2Yga6djZJ8Up1l9AG1G8QgJJxsA
bwKW+sVX766EnMRh4jIyhmMXk6DsbultEIsfH6fhzFnWXdSe4vqG3zseBwS4NVvN
WIG3dxEIr39mbuaiHE2imQ==
//pragma protect end_data_block
//pragma protect digest_block
/Yh6cWXKjC8AukVHAxTyQi5na9k=
//pragma protect end_digest_block
//pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
oh09+7QJYSn3wMOYn0UrKx7VpV7TfT9Ij2ewXTbcJGZilR1y0Jyf5ftzskZOaDdysViA1pJry6OT
ZOYFbOpjZ6B6pnUTm10/uCk0+0P0gUdrDl7ISMLjSKF0kRZv0gMN/9ff/ynze/NZVZu5M6dhmzNh
O/7zpjKcIMrx4m2ZKDL1O7fMQ7MW2g1kyjSxkK2JHYqwDJ/sxU1B/zRz1CzAHvmT/ZmAilOMi2LE
AduDBgxiKaf/TDR1Eq69IKqpyqSLmZ3BBoThazwGW7hu7h0WoFbGz5P4KWT4CPh5xmy3bv0Tm0A8
KU881aXO0vIbDv38QG+MlPcNtyRbbZaQtK+N6g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 2080)
vp0FDs3ljR2U9clWacEArGkO98QkagBIo9AcW8UK3ddE6ISETn9Jok6pJqt7YVfM39f5bUr4V3rT
okBxOOAzzSQlDDTFSKCA3zfmLExqLEsg70pOXwQLMnhqMSw1TJ/t98VtLIDsABoCP1mXhTU14PZB
f2/K+PhMQaz02JHrpsfDIT8sNnRupyY12coqaWI5hSOyeOvL4nnuH0mh8/c/iGMhAJkcOpLG8wxP
Rc24f66beHteu+upb6X7CLKN1vQXjVQEgHn+9FwJzrcIP8vnpGlvG/0KJjLfv8tR/6zidX58W8tG
8s3+QDxeOTGb/seDA++80T/5s231RBUn5sQs7mSvqglv7VxVp+5d0hx4h9p1VcRRWdkpUkU+8pXY
4sXNjgMLhPBM1MGrDDwNog/oRSjYNosElW6sc2oomuGAj2aG5gY20XYGdtNefVVIo9cWm9SeHDjP
IGqET51OA5NoY1Q5kwqDK8o3cEhBWrQ+5dMnCwesjOLJRQ0p4cYf94bY87yRvdpW11MIs06xxi11
vn8jvY3loQiLH8gbioTXrJG0lZEIw6tjMTn+3YhZF9jlMH5XFN0SEze09hV7Zz2BQG7bhOlZhyO/
a8Ga8f64hAKap+2HUwvBloT2Lt7jahHHQPeQtHrQHmNa3dPtyxqWGcInxDnxfDT3fUlvhR9iQvWL
GKAfAXWvMwo7/ofTp+KnWCSGITC9NcJ5sVkylzKa5Nxmbjn6tXclE5ETEG3yfLfZWCdmyZwU78qR
GuB0VGRg+NNDmYh1VEOqzEuVfqajh/9dSGowAxzmnBtjC+iEgKgrkpbbBq0VR+Yz07iW8w+n4BXH
NyaQ1fqKORp7It++bbOVjpaZFByK7X2H6Ub5iUg/IPhBTMPKcMSnX5oBNbrC7V77JtOHs1+98NVa
yUGYUsztnVQc+Lm32lDMICEppOgzMiHuR2+l6nQDMUzb9sDCZ2CpZaERC84rCXJyAZzYktjYHKOc
hHQMBtyaxlsAFk/S4Zt8nEjcw6EmruTcxMlh+ZwNSpJbQpauwh40DAN33PVBYZ7rFtXbvogt0Gjq
nXz/4QBQV/a+ejU0cwXcNf+GB7+WFePJWd8ooPJdlgpwbNpK+xttN5E+5BHsDWUMQOvEAl7+hurc
f3o4MwtIBaGwghYeMvJnJ1v2HCERNKjPWSopnVSgdb835O3PTbl8roAHaZ/sv/FOLLWBw2kdNgKd
C+Q5vsvo+CnNA2FPCFaWb/JQI0g+ie8KEtMnF0wFPoKC5Idio1heMp6BDfW/AJX4wThJNYbtujKc
eRsw9J4qrWu131qCPlWWXTya+X4fD5BI8UBHopHXBOoAk+GiCKeoT8DDKwpbHZ0Q54dRqUiztw8/
kuDD9FxpA2Qhqmfeh0nTMmR6qxVMhUJ/RXZ1vsAX8Fewx0kWBgYn8/qalN+leAoFF9kD4lElwZvH
LEFfXFEbIXuPbRbXJWnTjLdAtc2ropR58v6Opv39syS48U/hwDt4DjFDlc5g3i3JyUfjrjD60V5n
KdUm9k63aZMHT5odceyFYVDTe+lvLcd4bsSfuEeRnZlX+KErMASpbY3fpgSKPO4zMJVXWM4hQMJs
+lwsqwsYhddFHgOcHcxiHH85HzJoMUvPNrltNcjNbbLoA5mrwVoQkvgoF+dgN8xZ9kVJcRRsfh3d
yXYXgliBdwZhvyNzs9xJXJiFPDN6cAXHBMLcQMD31Wktrg3NV20wdRcAA/wCrQuI/4+eppNO5bdY
sypt9qau5EkCZbpzST5U8Q9jDs0UyZfViX8bfWwfXS17QOhcL6hINBoy+8t5oITu/trCFri5ZxXx
e1j5/SP0Y0EAkxcQ/JJ0uZ649MT1+MrOdNrlm0M7tP6g6nhWbD1cIosnynNQihlQzDBMek3qK9yG
eScxCMm7Sp2c7NLNb7+X7oPYSlorZ5otsWwZmNbfmbFMmdxsO71r6Hi3GWseFLcMEjoaKu42uI9w
RU7RO2xIodEzThyybnYHRCXuMxgYeN+T1mxpCOMmiOaQSm2aGEtYeMJggpq6820jEWpGfHUZVoeG
nlUmk+oq6QCjbBwNIR5370GjhUb7OIl1QrvQdRwB4zS/xY41miouiaSkHq7T2e1LtFccoM/dnsRc
7+c/YXCcdFXiJon6mCirjFnHvn0YxVJU+8uNwB2IukULO4gGEZrPDmRxPnwxlIMYqdn5TlJIZhrE
fO+EB8UOHS4gkkAcp8ADnJK+F8BHdsmWFOvpD+bhTGOzkOMRnTGdMXZY5AanskXiqJJv8BtBBEw7
OOW/0jImrbT3tRXVDOl0EBON8QgH1jqYN7yOcWmXq4+N/Sl+Nn71L3JbBSaMihghEMG193PJIR4H
QE4pz3N9bZGLdVrZgxem7K4F84Opy9+l2CDxl1DEj29StZwG7w2XZvufy+kohbIZu8p2/CybWOlw
1LNJdO1CgQ74DiMY8ZOmojfhv7e+9IzDooZs3drY+M53vQa46f91RlyPP+UrkrwKd/oLL6/ObLo4
nVwkSWfGIe/LBbk+7ONuLXjeui3/yU/kLiZWRpJbEDFV9BZ/yrUIw5ZlUSxHh/NhFAXk31/nKZVL
boxuWOmEfc63QR9mV3esJo8uJUTL1rYCZ+Ek48lsxxNRcwAOOeEEtgKVXWW5CXpK00QAZNZnxVlM
srlXS358MR+1YKL1jaThpxTdFKeI23yQnVOYbsUU/gKC7vtPkJH3ZDCykrRDUV5fEubSr5/iSc29
yYD/Da3llcqobVtB8agfyAC1SqF4Ho51SaG+2Q==
`pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
VEcv28BQKHon0lTbMPGVtH1wmnJURaPh8AfXQqKcWx9EKnbg6vwWd3n7nAFMGdvP
3xY6J8beDy9Jzt3NI4m974tHZqA8yqPBcMBJ/7dXOhz0KvQ6NEECWGKKywOksY0B
DgPhuUL03tMTRHkt8cN0XbnwUIoFJWzMSy3vmI2HNn013t2XDWkpySclpLaUMnbd
TaumFKOw120RrXxjtBwUDXK3INE/uWo8OjRa+w4RFu12O69BBK1Kv0L2yO5bK5u9
6j2fNDiBhXYVXi2OOLHzu4nBOqnTXrG1H0AX9kSg//aAwUV8VzP6OmzEp4iOOFZR
bjzbllJbF4AhzaU+jBPgKg==
//pragma protect end_key_block
//pragma protect digest_block
MyHK/c2/hY2Ci+IJfruQdFEDGhQ=
//pragma protect end_digest_block
//pragma protect data_block
3LqySyzn2TL5wKlDZKi60etEFxLB2i7+1EE9mHgxOcXs3A1amFAsjCh6tfJ3yLXE
0B02GkkouveNM9qa4P9HO7hKZ4AtTz9UeSqYqaWL63FRz2OtoHr5c9Z7pY4DXOha
gziKVMoFsriKKLFT1orXpN47W8Mfdb7hSzuBV0RgUkR2yMQCeY//JmsJO9nn2XZC
fGfq107kOahlUszsgVWfn8h8aNldQBYtnXKqjgrFNaA49sWsnZsXd/jQmeaEne63
gSQdnX+digzLj2GfuJiAopRCF0QEITZoo10bedOkLTsVGkv44LnTLRQjap23SLyY
Ov3hMAHmUHNc23++HP7dkJv8Y6MlpyO5UTqnmw1UM66H0E4u0YPps0g6GEMb8aNc
KU2f/y2hZjohuu+iHf0NewoYPcYMRtm5KnrXFWjqxGyCmWwVtF+4J+7GTXIivTvD
92rYFfGsehAUGa7UB8k1Fhq5QgIftHUYVp2NA+T86/5UzGY+jF6bOzl4ulC5Ieff
zJ8FgypVl7sOklaN7Gj0ayvieiDeHuj5//RtPND2v21AFn55Zysas5Bs0xDwHDnl
2tro166mpMU9xAE125gsj6nyC5DR0JqbggX2HE0pabFXt6D+2h6evp2HF67uC5jN
hvkiDE8CUh3A/G2ka+DgS5F3HFGe/rS75EU/Jht41k9LZ4t76yxr8dRoR/y122h1
7QJUJW6ih1jZkPGNKa6Cav/37j/NpnIWDTa7Q4997Ibca8LJ5YzX26fqx3ehTLTs
EwFUGN74wO7/mfE2jupvQZPmUuGJs5yaZTgL46lNrLxxgPt83J2g/am/S5dJsGCF
b9j9EYoszuaIcK8Ssqu54p6H1aEsPFVLsxyAe2+LYhTE1mhvfFUjnLEcDlMBTZ9V
Tyw4QfaEokjP0bzbN6PpbToNQ3r191DLJrudnEukvTvnv3hr/DqKO/55AiGu/qL0
O6v+493HQpkNUAtZ1hnrvT73Aldqz6xOAu4T88j4giiPrIWrDLiF86pdV5KbbXUo
VhB+QYPkEPmUTIXRyiSosXIAQF4jnTnl0kd1E3QhVUyNm9yFAhk/yXmF0NOM2Eef
34hIJKKrfsheBJlfcp8c8RSDxShM+NAFrW1tA2Wd1g10i5Ngfztr+cFzetQKbPSR
RxjMZKx/eX1bzbQONBpVOhOHppPjYJajk8erX3XYyLdcy4WHTtugWewzn3YQlbcK
a3/+Fh24nEsnGNdvq1YnUk2Qoh/KmzxKj6CANVnR7HfabCCnkvDmcna1EuFWWBnj
4pH+qwZn0KDGD+PWDhCGKoUd3iHqEC01FG2+3Yw7XZ9RpOUz8EVvOBBUDth/2Iw4
rpmQGV0MyBcDvDonVBruoWmMMxTyMmMuyRCgo14HJvAdjJAm03UsY2Prd/zKTskT
xoeNXMLW5O+q0k2ekHTblc0FMkeDXGvbX8HpfN3LhQAhZ2Sdep1POS74wt9ioOhX
0rn3v8nrQYRXfMDmFDehs6szp07G97yjKTCrcwHtM6TcDnQZy0YX19Z3kPRRMDyH
LUy07mAaCmX56cGMIYwMsTxOUMH4YWbDxS7PEfqwGpgWYPc2VRE7CxTFlJDSoFL8
USRInsNQNddu12xiU3obfMCpEZkBwQWq096KMiRE11NgcHmo/uaTtcCbQSDw3QKk
ypwzNheUV6p1UlQWHF40J5fOtSQ8w5k7Cutztp2/fR3MZ7fz8f4i2xLJ6Q9fsxBY
oJ7Lt7ySgsdPUMtvdiof+xoupLE9S6pPNEwbnixb3lAKZec5bIOeFpZZM6q2lKYr
7SSsM3/LYXWxUoCqnvRj4vVUvHrE2ZLuC0zIXDErpF63fwzb9HQKQ5LQ5IQBwZFA
yR9TH2kZa2THbgDZyClX6OEOYshznARB7FwQRzvXYmIGTLHmizu9QiG5WrwOckcb
z9h+miP2+dXZtQWCaXu/x1iS1KjftybDvrRyoar/z/OZasMJXuOoAz7xnkIzBM3X
JHfkhkr2C8jGdBnr5sV0GozOMxqflLNOvbskH9j5ACE++xL7CyUQpR7/B+Sb27o9
uFbMRcWVjSfW3qLS0IxsA+LC0dnl9qMHLQuFzt4idwZ4eMtACaaC8E0GbMUgJ4pq
bmYyOMj5FCwHqZHdZ4H9LK1FmdWPCL+YOWQlp5G65Q9d1yvrlp3v8XFKJ0V3ZfRu
USR6ijX/f0pfapDOKU4Zc9hOlPPvm6JTTK4IaaU7Ti6X3kCEAdPt6S8A4V6/hgAZ
ldoZXoZd4qZrmvT0ENX0XhwVPNdoqBPi02goUswKCobGuZfKtztfrnH6GQz8VHZs
M+3HZCSse5PHxC/Im4FZ4yjgEEkVWz/WFA72QnVmsSFdyM6seuXdRiTzYSRtbNvC
VEzl1xdKmzOmOCLsq18kiw8ILhUUw8PUSd9ZG9niiGs1fTZY1MULkPzEXTxSk25T
bq7LnuIb1HQNZJaSy15rXgztxkEECs2XPx7qQg9zUPdhNQOq3ctscyOkkoklFf9G
nMqEBHCaRkYVDdme3OV7AdgRqCfFGlC6tPFaN/0N4lUEqMVs9Ru1l4sGK7ONdtUd
pZcOsqRqyn5QHPqTTGKcc8Tm0aG00z5wLSLiITNaIl1299AMFfThkStRqbpZ7bIN
Y9AMeWg6G92pjre3WUa9imnyWjnh2vevCES+uzLrMYfLQJdagpw9kWQJ2asHl/+E
ntPdXB5e/rk0BMLD/OU6J3iFBlFuN3ahTdaVsFfJiesQEP35ho1k2L2LYF+cCuFp
cY59uYZKjOHhDobWYi22R7LAVkXIXee/29uRtGUmTakcpV6bIMb+FElgWE02BViA
DfrYUY73Xvk76xuwJbpAjiQ3V2G3kKftNckGsHzvvMMwmqMWJ+HM9eJhbGAxmZby
/Xh5FDUHa6kncisnCEO/nsGXE/N27+NnmLqytKzT/56JzZy5fI/e0MyrsBpbP9Aj
E4SEzr8/EbIT4LvPh9X86G1wPY+ENZN7dGZTjiZPqeE/YDVpqWpEkLeY2YcHJrIJ
zrCU5yAe6Cld5KW6vf3o1ps6E/nhBhe+iaKAgjrqEfgcMWaD5haW55Xgk0v2Rj4u
nlapl5Unl6k01kSdRFVROuYzh7w2SKfqSzsPuphjrdcbb33EZbublcCYRvzP5MVx
UhP7x6i0Nu3zA0FgCO6kBQTQmrYghusNP0vPOz00ImXD67Ly18zNukhnY859z9mx
ivI+lKio0GOynoP0+TICh/6WylS1X6oYiJ1Q7a6zBcT22H/RDE8iqPrNc5ChbQUL
u0CcVZN7hCBh1YsxNzKH1VIm26SG1NSNxAfHKsQGmp1Lt2CxEBXcjhoQiIOV49M+
AF5LH/D+dxVONX88f2jUh39TEuuQkRBrfwXWV0SQduooQntfXcUH8/LRI5otoF9m
N7Gut7m7vE1AyqC/YFulNKyR3/+ZrgV2W6Bq6fj16i3hI7xe/wI2CW8eYX4KMPo0
YM067dBW2JZ+3kg4Kh96EG7WmeCu74QCPe81KQcXs5RkBn+um8bDuttM7bYLeSsp
pPK4kq1M4JJ9AxTjPXWLWwQvZMmak+z+fWenZtdJh4nVUXROOjJe3WUvauUfIL6Y
MVKVsH+26qqBu6ciEqwxvEFfkSkH+EC1W4iLlEcvTEqsMgnsfmUR5RTflYPhLDLW
wSHNSkVVdwASS0QjU9Hj1wcAEgQOcFGPZYLgFU54XwH2c6pVCt6iIdvVZ5jgIc5x
83kuZE8hGOUKOu3rtRMy/QNWsV8mir49W0GRmoXKwLSSKU1nfBM7HkJ+rhgOpwEL
B7p6ZNAKsWTpkYZcVXWBFfDZ2h8Ax5U/PIXMAemq1bdjOl5IzX5+VjGAKxiB5DlA
VSxiSBNeGkb1cp2c4fv2UDGoolHS1/X4zqQgdlWJpjIJTV4MzJFpHEXr5vAGRnJ6
Czek2BuCLRoa/uIrDePivH9sI3dE+Ub7NImGowGyGwDBnJhJAfTFccirbXrCRR6/
D8ENzXBYA5jGagwEslelreEDutx4fcHMWoiUWvNEbbXC1rUX72zda+O0CSxO10+E
6KQVwM2oZoxtl+rfaf7++Z7H1lgGd44IWGsxG9CEKmzV8tjd3/WJKz3w6+/gOg10
ApqvOGHX/tQcuW/mzXPz4xa08f1uId8nSeL+z+o0Tadn47FTEFkn7k+F2mZjDxt2
Hyy0wxVO3TsZXs4Nqwy9FJ9rCJsvYKjTiYIIF36DeCIZKQnsN+RqtUXYYIO7yg5B
WjQBwAay6LppiOM8BsgpFmpxFNONHfFjGpoBxC3ltRChxpUeKfSFOzGe0JO2dJY6
15rYIqH3SNfz9MWJ68iCcpBfKmzWTwAMa/Gkz6pMruH8vFGAjOXMs22VH+hR1cwp
kF4w2vQ4pohy7JRy3EKRhR2W+NeFmzqp6E1G+Hcb5PY9X+cnq6ve/E9YBf6PMQwo
If+VIFmL20+nWXisgLu6B2AUBoPQYLrElRKPxc8VHbN469clESIiE3LRshQhvxKi
P4qj6XPtLdD2RbJYK/mQVkUyindRZPnhaxZTnkNQkE0k9XMSn4L/Gao3Ulm1jalr
rIGAGZjSpNYD8FCeem9CyQio/8bewl34XRbb08bppWn4Ju0GZ6Db3WJa3ocPlHhD
bm9rAslTwG3cSySfqYqJ8M14rfMSUdHE4GVtDQhMZwk50vlEgkd5ML8F6apz2hHG
Fz0o/zmugpWtqxj+p48LuKUcPZhEnsIPJwhuAj+0EVtOvyGmy58QTpMs8WiOWW4v
HCeB+FsB/mJXNNbzqPTgYiFYh2dayA2B7RO9oI2rxL6BbI92BUTEblUAOmh4IOV0
BQgHSjbdNWjTFFB+UdVSmYvVigkzmid+2WIlxqkd0AkIxYMzn645OTIUfgCfABqO
HbLWeu1YE1T6NyB0YEAY5ym8WKRQKMiKb2sAeeI4CxQLiXwNCIGPZ4oqhLSvR7oR
IT6q0bnAhCW0mRd4oCj/XsPS+bhkD4/uWKnKy4D0bVvBb7Fs4O7haSaJsd5uSV0v
wAsaYtAJTOAQheBUSZDBSZSCNb1s8LB1m3kvgECM5BVUKx5EAv1YVpPF8l1UbZxe
1Aj7P0fFcjnV/3i8O8MPpsDP504bbD+6PVBRD0AZdeAknAbdZa0hVjeGhvV1gfZZ
fDelndGvEcyYsl1vaiXcg9AaSXoKKflQaBIK7HnOVQ7GOicfZc7ipibIKDGYRImJ
74TxuJsApPT8alFSVaG4S9AlNKiLYdYzU7Er9ML+GhdL2+1aVbrgwfhrUMYp10Sh
FcsbB7YDJkNLANkr3CN04vOMWOGPyCYBoVbfamHXUC2Mm/nKBUnX/iHykBC9ZMTY
/LfALq6gF2nYA0XtLXWVAUv5XXZp+DiGAt4UJKuoMDUyd2LsBe7O5E95fa7EGlWR
l5rxqq2wadbjjhCgM0iO0ov9WlNKDmEub5lG3t7B059qV8QqoX5Tt9wQv1QvI64y
FCpWWOvFZWkV0XOkyP12x2XTWH4Ct418IsyTX53s9QlFO1XyPoHeXP2CxzdZWYM2
5NlZwPk7Z6zdBG7RQEIHRGmVzhxBgSiEEQR/T4X5uLu5eKjvkx6Ifg8m6EHjV9V8
WNXM9e3K2Wy4b2yKxgjpaAij3JjBV3l80KxJP9WztsNDLJECki0rKALPgXMQn+6j
qe1OWvpKIhbqpTh7CXrUREjZuVsd0s+Dks1ZKhYoz36VCgSpBgivKa3ACK7YA/zM
l5Wt7zFEPiO7y86/1daQlC4Yh3no2BqkPfNb3/6aPBSyEZalZt1uh5Hdultj4gdJ
m8D1H1XlM6TZUdFyXvJOY6Y+wyAhcUyLvllq+79qi2wM4W4yxqqXrqs9kdfvoVPX
dMJWG0vqg8Ixvb2lxiPYMsZRlox6bCx1gAaMOPiRjqWkrULbOBzosmxTFuO8eUMZ
fpw/magvoettq0AfcdGGcvx6kD8W50e6xgUwsUEnCuP/M5RY7rVAxmK2yZBzmxaX
s0NK4KWd22Z+I+ozsoxlwo2KAbGuszw/I2aFPwfB/+i9nqEGN/zidcGQ/iWu+Uu1
RxKSh5kyYEhIr6LbIylumxP2nbKB+tBhvHO890qM3NW4VggOhEBXPJmJkaxz40pP
fSlf8VBkch4/P6MTQjNmJYyCnJ3wqIZYVvTIEJZfg1kr1bldgqd7A6eHaBQcNXmP
a7IdD+VKw1739k9vfqvu0CQ1Emr252ImnqI0h1OQ19efWnqfL/GKarQOHCJzRBmN
XITr7AzRzZzpyxdqJvqIo+AbuNTsY2vVevfAzb9qaLtbHNoR84NBSiVhFMPvJDu3
jXgf0WB8w6E6zzk0GuFpIsL6qqSCCuBferagXfqPZahizcN0xjwown0S9d+yvg39
UqBI2eum18tdU4I/7buXb9hjl+qqO3Knfy5dU0l1qUpDKWK5qISITXvJyv8j6r06
pWDQ9vBxsCMqPi1N9/KhI8mH7LJGd+u9iXvB1m98/dbYbNmKLPGctTMrzyFQ6MbU
6Bpk2CkLq/KrUix8rp3am75J5LASb+2E0H9aI4i6wtb0M0RamC2GOkIW/J4f11cU
pSXRWL9eqVnmRjsZf8dQlOP2qqt8+R27TJxCNubM5Ih4pu+tTX1Q7luKqo410Vb4
0elDo8I7xLkAGTJZwWdCp2+9HvTNwGy+iZnlfZfazMpoH34WOoi3KukfZfysvSCR
G+gpDR6WhiBSlavhHRzIvfquwVqOf86A7ESD1kgv0r1XAHz/nla0l82HyN/3d7i2
jGdjU+mHruYfqtM5kqs4VCL6pGp4qiA9au87r4Qt5HViGZXbgTsdV+JbaTg+140C
sTGoH+vDHvpgkgfyyV/HfCXPG6yo8UTsTPHHnx+9s86t/qSanUW+vjt70HIkH5Fv
BTZ1pBGfqO8KnXtAV0NGRNPOVx0W1GaBXcGHmvnHD/8PwC+icS0EKqVlM8TCyPfU
7Tpe2vE4Z3T+c5rE5QzNsRjy/uHbH7G/KyMyweEs10DEQPT6Hwd+gR8t3kREE2OS
JOSn8YJTVhVR8vK10PBlgx5iyRsI7FZ+5URtB54eO12dBoaE9g9N6lxNULaN38gH
UbyYTQCEjX9qm0m7t63vtjRVP/D2GGzObiJbB+5SxkRbzg+vQ/OTd8pzRFIw9uTU
rdoBW/1X5VfrxC6NpSSsyRTTHtroQf5GA7+tk6bIrQatyFmsthF18D01PfQceHSK
hQ4b4r16XQXgHiqYpvrdqC6+XOSm1CEuMEf7pU2SsCZTRU/5bG/Nh2hti5Z/Sv9D
ZKq+Gu4+nhnEGQ1o/0va+8Lv90lj0fxLunY8QYvRQUfKXXGqorzO+dDVOVYzyNSZ
sl3wxg8XjJmCWIlhU8RR01LwkDngFsV9yYrK116/bmJ2VTglJHf/f9fzbCzFcEpR
wRJn3zau+eGkayYnhtZhZLWPZxT8hgDDIc5zSo23oU5ns7AbSihFh1O2EII0iyTm
LHfkEa6m1bYdI2QXCzQe3PxbMigm7Oa4ODrYyaoDGy0tUAdFa/w7aA1aq5bjK63g
sWRcu/3EA/SCI+Tp9h6jQIELF0ybcP1131UN11OnTUSroMFP/mP2zwfPH3lSk5j1
Z5IOdeRlA2+H5JTN7/ZDQdQawIeEd27spq4siUBfocFmLISjduy/LfbXbTQhYfkD
IOIrWpbPBFKMejUFjIzr30vhMLuSokum5vxvMWFRKetnszx20z0m4KYJMOnmYPBE
SLYdUcYVNlIlvNPxIW7QJdtTPG/U4/D7dYExz74AJNwz69SdCK8Bdh0vPuEiF3WZ
4tVj74jxC6NxYF5e5k6hzn62XFsLJQUSTkRt+kCeNkMQEsTJesMR6L3g9bGZRpl+
bWZDCRInEVGCLpGyhx38YqeiPgy4MykxhdMyU/n3sKXMjZX8g6Ds00k+z4StQP69
LCPHOMiwaoofwwoitV+BpXqUVFBdXz0uVWM5z9G4tz1f6JFg1awWUYHosJCZgkDb
kNm7HIXzeP6C1vmozyjyBMcF0Bx3NCPkmd1BpQo/1Px9L5M4IpQdehi4Qx5YVV4V
1ALpjgcBGjI0sRBwiQk4SGC6I4Ki1wXarfbu2Tw8Dy0wuXuYM7UP8iK47RtAeCry
pUH9m/DgFB/iclwWQtQuWPVmFvy4YSyqhVoW1RY9DWqE0lltbRksMaVUN8wo14a3
dBrX+zwA6AnIJX4htyiRq48SJNzuxpQ8iqspm6reAqWGBXf8v/r/hkqlds3iHiNv
MAqXCzuRF6vXcllIMDvU0ng4HZELAALm3FZy2hSoRvrvBPcwJcZykCPsxMQuBj7N
LyjMS88C9TaEkp0MBRtNRUUFi8/AvjhU7fUSq139i69/5oiLE4/4Ili/9mHNCmFO
lvqY3mJnIFEIWdj3n8SqofKQyzL7TwWj51N8gX+agL+mv6KIsI/C+mSRdCbYAROw
9UmkoUa5tdb9xKwMmcOtyV6Vsr1QS7Zal4Usoci8ngyMUHNpAAiVECtyQtf6IXfx
81HoxIGD8r3zLUL9eIHAgUu8+feIPy9dZWUJi8TqdlDRFUIaXy1Gv5AIxRfNYePe
hakMvKhafQbpEKRXzST/kUy+o33znL1i3B4mQtAg04BEXfapr9YJwIc8KAZI+/hV
U/DwjkN42d9QlTCuQ4RmoDQ/zPnASsFIFUGDLdLSH8N9ny2iH2+6A/+/BDkDB7+u
AX8it32QyHM5mmPitrxhyRWCSkSI2hb04L7Mxn7ZTOdFv3gUZdesBimTbza4FVRj
TFoynnx7m0t9SfX/nWep3tY6JAjxjepWZQtX/jB2c4uML04pONk206dUEEdTZNuH
ZB/WLHdw3u9duZ6QVkI0ZyzJd2U4J5pGVOyo6CWUsB1GROaroJ5dteLfKqefT4yb
7npVOQdzeHf0psY5zw+UszFALZB5kYnUnpjRJM9K0TS9T2Gkh4YoaCnMss8gFYIx
/QoyM57fHZINexv/immV+QmKPTMMpL5GmoEVULrnOPAy1e9k90zveid/wnIqrz9s
7k2c8Ejz2hkQj0cBJv/T1s23P9nJa5mqStNsbk9qVGUDp9pul2LyFNXGaLU9kRBo
z9DkgXzODRZa6kEADdNV2fLF9pLHwPFkRGDQdkhxudp5VlEsQkAJcQLwbd6I9sKH
300gWFhpgNq2K8tRvF5vA9rsKvoGQer7mDnhGPqIDIPT5kb9zfqOhpQSMl2gOrlF
1yMxrKul16GmP+p3cXUzzzIxc6MrL8tj86R7b/qgIDgfNUc0kiZWnKeMljvOTGOq
2YrE8LC5K/wwqvdOmnPqFjfpR+9/O7Uhwqtu5H5jzxUD6sBL7J4US4x0ei0fjwrK
cJAKQoamFLpMxOmQxXd2tw+AwffPTc1rJyCsRFjR6wRRs8+BURwXMnZE3T7C13kj
TQIPpkWBFKXj3paVwWk93S+0PkFRlQCB+pEixY8aOsV8qrVdrR4kRE4gOElJt5v9
q8hQVtEs51MSRbzhLyRLIgW51arGeSjrt7O8dzSId/aj2Ot8eW+At7dxF8nIfzc6
YBfCNbD2SpAJpWbIbcQVloMi0lZqWD7xfEsz9sS0gNdZTsK/DcALf4VEv8MgJDCT
+aPOB6Krst2iJ1KdyomPtdfZ/j2hEuHpLb5k583gLpEMWPu22StvopZYL6ZzY+vo
MgbU/S3zjQeWUdsJWvrX1nkdVbBLjw5FG4d8zKUkEJmHm+EsezLWIlCMB+XGv5xV
+qiSmka52pxVDDCApQKuHQJufyYfK6fQSMZrWNI16nIr+75WHSAuD96EkYR/jc64
yladJ4R52HXZAjF/g/qmgPCDyOqs+wusTj8lrE71SsRdTiUCJ5Bn4dvCvtfEFMdb
UaTsyaMJeX+182zgz2vAu8O4LBBPSf61dXo1tClBbNHhkE8OFe1IfekGAYxUHIvs
FE55Hft42Gb9KA6uugaTjpNHCSegZYFa20DHuexWeVa12p/t6sgB53WjiT5tyufk
isn9k390S+ek4cDQPApruEcS8Gdmq2Z6t/1mdwnUlAYURNS5VF5aOC1u3AANSd/k
F/VmMpfb85OS2JfoQI4tzupMZhAfyjXtDWKb95mouq6kJGgMxkFWE5MW+fSICtOU
DQ50Jk5SalFyIibxgCRUpCWdDQQFKwAq7IaRRxDqi3oXZ5OXTZLCF448qQb2TwXP
4IIDGKFjiHreIWVBA+ZrF49m08WkjkdTsco4HzOYyWaySbjv+wxfBBPQWJEKP3wj
tPNbCDzqQdFLtNWtt7dzyaf8JH6Xq0GprBNenZN1EjZO08pi+Q79WAbaqhWUnM9B
XarDS0pRUPa/GiDeUsE1ItBnZVwOnwvXGIkEQuSFul558oF2r+x/0yi6LVyam/Nc
psyEMKGG6H992u7wagZ5aSaWO6tvQdU2TpTe2YZsexB5MIxISpDaG9ZhgDeNVBh+
UXjnoGxcaaN46DI03eJJ8iIvHhH7Q6iaMx3KXhTgEv95yUjjw12k/diSC5lJ3cNL
KPd5YIlGonQCOXAFCI1YmjQ9GAq7JYzcs8x/1ELxWUJAr/+UBbnwkBZCoWQCmtzj
eysVWCOrPgpFGR60xFBgJSBv/ahO/E90l2Gqy6uF3b59yCeOL7MopL1TyCKvDMeb
Ft9KusP+RveFPfWnDOqRZKUnFgL9uWbIlm8enpgrh/9aoO3wCxTWWDJipb7w8m6Y
1TUYUa7pKNrUiciDlfLplXaPPC5pqTQIgx0vsrdu+BPKToJMNhmDMqqZEssOPv/p
BXoauZndKmSbDT6b420YgqP7t44mLt+fDEXB4Z3UQR3QSTBoGAuk5bSrcr06p24S
+SgUSAkNop4NKPv42X/Ax/x5RdlUmkZN2xhDExKHWGbEsMsHog4CbmfjtZsz7zco
pN3gSY4PfyK9QVKEId+tGkwXd3BFS0VaKovVwrAeyxuHU/fWXSRJnjxTtjFimmWK
AXHwrZimS0AQiEVh/0pzvDn1jgqeA9I6v0K6sDvUm8J2vT0dQzc68EDJOgUDUBVX
HS4KdwJgTtbZru4CnTd9nkADxYG9dtocUCC0DFeXr3JHww8qRAvmdtkn4bX/0o8j
hkk7ZhZMXA9lfSSeSqqwNr7+cwzYXrU0aE25Z0ZhJOSS4NBfkUyepSd4LTvBrgku
ahG/e3E4lZLnp2uaV5iimLBeB5pNVVwcplV2vVbiry4S4vAI1zR9woAsW9wUO3O2
FV0h6i6Gzq9E+SVBdnjuQHgoNiEz2BbPN5a+HEEbUJ/LinvaYyhY4gY/j1VjXUuq
mh5gYTyhqS57jd0XBOzC3VpUauZS4dxMpNKiQHdWHUYHoHsQCXmCyg0hXWoFVRKt
W+NPuKwXYJ+ieTmKo7f9haUMCPJ8uglx0KXGeME5CmGVkkW6qN8B0qNdAu7VRioc
ZMtRsNOPiRXl1TOLpkvpqiB50A5NesfggzJqVtxKuBNBsjkjZhTl75SdOWHfxbJj
DuzPr/rGU1om9eY5vo4QA2MQXDpXFlsnsyMOuQ0aHXR9ONn5ZFdBrwYju9mTGOXt
3UZqY51PrIqZHn4dIqedBilT/ROv3bQyubfNJgQ1DucaCGEk6QKZASizEmsft0Ox
NioNYddfVUjkGLx5WgAWB2OH1M2rUlnZkbRyLO97uiojaYUDlEhZEVCi3vs4FZ1X
/6KXb1XEcBQ5ZkMOA11Hx2TZ3eZpi9xT34ThJv5AzOx0C1QHipoBGhH57RRPQjbP
k80ujhIxzt04Re5sGAraL9MfWD8qVUfeybzPf4GZ5eduTLcbQQU6Z1ZFvE8xSrxq
txbTO2+eEXE+lA3ivAcDaXTfqhroiuaPy3ECZD2oaiFjAJqZ8yBh57Y01dwTW2jn
648LcTzPbUyzG2OSTv+RyhW33Db5cHW95jIx9G4SUxNlMPazWDR/AWWz065FKVaJ
mJrGwUTSet8kbwL99HstY0dIVziJov5xCfJSrN3eu3od81uqMn8fvC3HaHXNeWYH
0Z9oxT+HIsKV6O3ZdjXfYXqx7f0zawKqxktkHrj9G6G6tQK2TxI88RMtt5z3kOB2
trUUQRsU1DXycKiFgzCgtWag4dQJJEUnspTE5eJSyr3zugj3oQAUnzW5cjo9z8j5
Ybq61Qob9Zm7M9VGDW5KTlTud7yAhC6xw8IXA3ZJO+EacNh6ym+dizLDx/YEc/ys
XwnT/OqavIiat48Lt42kA7Afsd5dTfQeMLPU9V1v0I4KTYCQIWf04L04SaeL5rAw
3XbngoF3+8ZlJ4ZbhD3TJU8vtp6ETzpOSofKf0zwIiLcguGUryLr4VR3ukJJ57Kz
Km7LSywlI/uPPE3P3YTWFvapAXFlnFR1LuPNvkkoeyfZ523cVHoIrqwcynsm6RLz
t7vhhvLCrnOh8tddk0ubSrxh/1ybp9nMNT3XmbKeTaKLbKi117W/iGX51cCp93t6
cegt8vsgFBgP/nRinxXPK63HgFZIQef0A/T78VOCcKa6r/Ir+42Bm4iMp75In5BR
g4FWmGvOOw5T8QUo5wZxbOCdPmbSupusZ64sWmbNQXKThbG590NYRmQU+P5w3XPs
36/LfiLFI2sO6aQwh2G7JaCmH2yBwewdjkgHA7i4sAm9an8NBqupfvxCw1sD2qzV
EZn+XhPY+L3uBlQ1TYNE56ZaMJAvR/ob1COLqjB01MB+fB+q1Ul+YrJ5H7jNtX/G
p97tQ7TqxBJ45oSfv3qqzQVaFgSgXiFDmYIk1zEnRKmIINCtOJs8tjKeNa3diEyM
u2D7yJNsjPWGK+RLHYtF11nakw6IZj/4fLHM6iXmok7ddAEVwzRI6NqiWWdYUQIJ
co0ivBOK7XG/1UC8M2tznQ/QNsVSfTSSQzyDglcq9Tlim95cvWCC4MTHjPtKFGpl
PM06LmaamCTxJaTM01wASxHnFLLVEdpiipEWkAjSRrLHnwgHpwiaxfNu2CsgmP+J
2HrA3YWwtGbQnO1OPeYOQ+ZnrIAwWLzfM71CHR5T+C91uLYPH/WCS4y+rnUB89x+
iPw+m1CdFDsoNcTXp3UeRPxjM5rngSNRo9cH1iRgiT3bv82+PXDnr/9dh4RwzEJf
RoYlGaf+gFF0C86ZZb4rHNFQqg4iuLWxebKw7rNaYToMp3D7SnVbdmnUyWnH32bD
0U6mosUhPLdXaKH+a+Wn2MUOJOL3jyF1S1EZa1VTwSfSIwhHkJzQJeiVDY029ANg
3lG5zdlwN/eniyhCqqCUqC4NF9YkphZ94DM2LEk7qOMFiN6Vh65zy/W59Y3QzRZg
4vleGR+YBr5itMKqBGgd4Ngbabt0UeALZOyKJNIbGNg2vvPWrbi8rnjxhRq1nWCb
m1HkXkq6xSsZQccXViA4g+NWNHNwLJXare4PKThrEu4RFm62Pcn6W3LlQT+eOhny
W9pyCRtpGMWy8rTZUWorACcSTzRId2jRqFxLh4VTONb9ptPJMabn/26EtNzEWSxw
Uu7ZcC+LFjeBQBHrwlS59u7BEa44Q1lmaAEHF7I9iseWsek4WIUJX4DBBK8q5IMv
7QbR5BXfqqd7gtRxI4xXioULImTqXO4nxZh+3uU+0mq+yLj3NuC4zco4fd/Zni9/
zByMpIWCgwCtazF7r9cUiqvte+8UkRrBeQZLyOXBuk1dy7XrRucvFyLbwUUwe/JP
+55PUJxNZhRt3epbl/cJ9L+Le2kWyLWTupOejlRNNykFHxtsMU1iIydJUoxEz/Gf
0SUEZhXp3Wa/smVWUfLvOcpXgzaYVjLDA1fLXc7IIY9mqbntkR7lLvcR07nRgS0C
FwkXNiVEuhsdI9kD5vQX57rVYej5Nre3K/I4Xz29gp4JckaEopIeWvZfBh3QYFoG
zfXiOlpOBAkovWLKL7+kkBA/Ks4Ktgd+BrJOB+hgSENkndzU6+UlV/IF7J5RKM9e
hBQLtXKKTsOFdFO7FGsLINYSTKwGz7jfQH/GpwsBi61Zxolnw8yVkiz9SxGEycTm
QU+DEFnk0EMrlXciP0u3Fq1mXjh49aA2o99H/iiidc0UvaKIV9KYwgNxgCuWxEjj
WyL55nkYjZzILPdhQ/cD6bBzYVlmPieRm+uA7R8tBZGn3+odkiUHMsdkcqt40P9b
ol+RkgzdskXq+h7BNT6O11NaUZPkfzkUIb7Pe78UwkPqneMTnzRpVug6GSVxlNNq
GHKI6nly1mYoaws83sTjNOKEue1nvhJGIpsR0/To5O6+naZ2/OZohPj0a/u8DZzM
jtdQoGgDwbY8fDbP+Fm6/XcakXThaqEKtn0wXp8zECvS6QYfqFmLyTkXMJbAvRDZ
Ie3E5KhVQOlzxilmKUHtN8vnhoDbMwXYkzAi9rZHfuF4nZ1c9jFwrPn21aRckFgF
4arxu8LGhp5vZR+CTFAFMogjzKTMRfzWo9ch45GaI7yk1Z8copDIIGs3BbtpfLo1
umgfcrCCMgouUfrou7PrM7P9xW0KRbROryg/xsk8xSZEbhTaf6Nfioqb0hKMWagx
nxv3DrlszFXYz8k1uGPaCM3doq0aQQxHTzIFNS9o/JDvB1nLKYq1BSiVXSCGwjUh
PWezcEPDd2L7PaKKrStiTWrZq07E9Ces4P7VAQqE0ghef4pkQqW7O1TkAYSjVRQa
4uA2KCfFH9WUnMLmcB2FxQc7K1Pgx5S7WrwSfA4A89KjaKWcAz6Zt0QfHS96xGBy
ACxyN7Us84aT/R8ia8zeAoWDv2VrUv+FAKj+f17JdP9zbyOosafG9ImNyzIvsU4v
ZUsctxGfHa2MOzLkE9DYkiJsQ73mjF+OPyeWXEug04rU8c3AQ+vDoQ0MyT+XAo0J
cGFLHqSJ+zDVs4mF+fySRD7KpqYDDRwXLyvqqFdfr6xt5AShcnXF316pIvZ/GDo9
d17maX2tISSviKnWhqCLdVufelfdOYni+hyJwd9ulUvUgUqSyEWTDVw9/61xbiOH
o+JIEjr3TNJnY1Q2BVPA/Up7L9/yB35WpZmPcTb5/Cuo0WFbKLOPAPGTnN6BlR14
kH+b3ZnaZKqxHNASvxwmSVMPsqKzvNVI9EeNE3pyFs+yIAgF33yVnq1ALmd2RIEY
JO4+ufmX0KR0qVLCwj1/o6wz/I8nSHgRUwoMlSfnlOiTQT9tQHc+xCJEQmAbMm29
xmo4iPIPjql2Ygtg5y/Uq8BwR7W7VTl0syf/ile7folr+A33QatfxKD0qVN9nWZn
p1o2SFTCIP6+zm+Ku/jfYaFvJIJajPFlHeCdvzOsAwJJ3FjmrUDJqwmITc0I+Csi
9lVqex4R2TBz+BVBZdxwPGm9EVD5M69GfkjtXNcfZMWIYuM6T71cpHZDNAjNVAUL
/Xw0Le0pkfrVB4Qu2g5kr7BukE0NOQ9TkbCbdpjunR47hhZnf7HPa0R/W7nZ3o1s
aMoT8IlqBY1IipICZPM1C9gT+6q4h4HIAxdRibLXjrJIEFPFuWuqFi6Mv/KlC2pk
YqGbo6zyPKwYsG6bXVOOIDPDueV3OPXQdh++ZCbpAs1YJJttoDre0/faoXhr+6Hg
0VzgZokQoqUY+Q8jJnOK0MHzcFJDaub20Y2POVYOTfT+3mDAN2qEgZKub94an2ac
bIh0IXpEo5LyNBuqoHzsWNGJ9BT8ml2MNGcKp6/cKm/C1oRfJTjRpQZ0YLBZJVRy
nw7q4FK6UyEPPvUGS7Ohz6N9jVr3wnnwH63pDphhuU/c2M4PcBrpqhBZjBsUMIa5
lFxF0t43OlGHFXF+Zo2mmwNiTbSzSB5KU6POuc1PNi5kfyuQRLgJUt/2vMBRs+ol
LP7KfymDbkFqbcYnlj0VQb4izDn+5C/wXJJSJlKNg+quz91fcBCAdshVpxgXXUfu
v9LKn3c2NK4pXr+z/pH5TqjN7KyASw88YO47bLUXtoEsGT14B2I4Gtmesw/nyh6f
I+JTqP5sCm45ztYMrtciKelHzFjRN+pj8wGc97IqqEjKxzuyCCaExlVJ91tWMHmf
6nMCMI1EIXKIkxP8uBDsH+cmAxzSdQpbvw++/Cc25ZYVGRXkf2QCdYnhVpIN3dkg
TF+B912s9HlPh3Z3yMgxdKOVyaWiWpnXkpsGgiUWjV1jW8POwKis2qsGNVnHoD1I
M1AAYhkinrw+3BVB/i4a6UJhXW1bRG+t3Eu0v5r6b1s5MrODWfLtWAHOhL5NiQDs
Y7GrzXeaKFZvN1FpuMyCYVPuolErB12GCAs6LCTnNKEq0qVNhxSj6Mp4kNQxyjNp
XXg6fV3H1SUv3d0GaiNEoJY6Kg6Ghzhon9ZREa1Pk4AifVcZe5TT0TdIUdOGANK9
1yknbJLPXAjkZEw/H3vZPFO/njwOFsQ9DCULB7hwdS7aGpGrS2tfVdPAnVzAbNy+
WML4l9vvI6BofJ+1n0csc+6wQEm45wyxxPq0eV7ripb4XQqZR71KOeK9tHTeEa/J
VsReXIGCxHRESOVypfnGsZhVmSDLVFeWnpfUXSRPp4aGk44fAml+o+4rY3c3HXnS
4c1tZl47nAgrYeglTmOCMQ0Uc7CIJL7K2c3Wa4JJVg25bRk13dyDJamae6v/miwj
nXT90p9BxNOrpnfhGKIOQtDKgIFpx0qJFy2IwSGG8QNongjldVjnHY1JShL2m4hN
ZW5atUMIwjKmD0KkLD9p3h9mdSav85diyM4GQXagogvkv4jguqZXyymqeNtfo9wv
h1DGiK75LLgXmmjKrbU1zJ4Hocrp1UD1PnCiIGdFbyc5JrBxhYDUf40JP+pAplzq
rmPYgiL2AQrUnW+BiJ3CPMinxObWjsClKQ8df3LadTiryANcq7xY5Qngs8DoIY/W
Q23Kdjb5qZwmvCGJI4066vA8BkkEh7nhYHoFalkbK9QLNoHDnlL9knrYOxeYSQcy
meYNmxP7fJICKXm988Y3STmMuPNKcHpDCcB2mA3xlTRkP6s8qQdRpKOdb6guwcIs
ZALWmsl3UjmS/OYsNmXbQumcFujv6+t3CSsdkR6YjHwvYTbpGesC18/aEJz1Dl4R
vZ0hRk+cMFCC1mZYzgzOt3197ktjIRFsABUzbw5Q2wzrLLno/stCTQdd/tHzdaww
Nbojr34y6xfTvI4Ap2YsyelpeNkg7BMKs9Jb33TSQSF4DlHDJuHUGoUvRTuH7mVd
hXQO2LGi2BK0B67NYLxQKrhQA0vn6Ny+mGduVVkiScORgB6WwP0O46WzlFmKO4aX
3WQvw3yoAk016+KSFV5bLNhjdjwfsg5qUSY/nDDWucwvwzKb4jQnzFpA54rhvaoo
Us6BNcqtlBFnCEO8ETe2sERVrXcRuC35MZAhxbhwUGaF3c5HhPxQXYmS8G2DG0OG
1Guvh3IiVijo2icmQv3LbUvLO9XmLz7A/B6W9dIRbaOJgVLwUUfqU3sUzSZocmpP
WAuXZdDNQ5eD78nw4f4cnVo4KG9/65tg9BdWXTr4RuHk7USI0aMribtrKF4sfsaN
bRgJRqMuMAKBOEyGeW7OBjDqFU2YxiQjy7OKamRub+iBM2W2PVLDqpRtndugYwiV
t9+NL3LtYviGesDKB6XZOCzkJEgLpYMrKkJ6IwJxyjALwP+u4SyHhUiPmDTH3WJS
NaxdFXEpE1LIz+M/GbuyhvumtT7FktpMDddQLpsYUvyYgnKQMa+IRjU9NAcCFbdJ
yAFIxYBIUuvt5k9gLxBFdf+Jof/r3zUhwo0LiupjpomCvUvg1ANpcW3KCP2YvHj5
hRptbJhy4HQH+w49DhQrNBSOllPdu8KcjazAgQ090kM+HEBwzcnoEbPLWANNDYUe
aKLs+lyqZmQ3JynTZ9mf1XxzdEPifInMCvhANxus3iWvjayi49dlPJdfZaDHYpHS
kQaIwfUx/Bk8fnEgs/Novhdvqmyd81gAgmU/V/No1OjciQ3VJOovDB6SQiSlY+W7
Gr06YDmRMHGZjt7dVsnfjM41GvGuEUNJHCw+yxQH65IgQDx7WGiGejptw9iRrVwl
FuLxRUnmB8LtPdWSFzzcwaarE9ZM4iYh5h/71fptDHlRvESnDh7sw8mqW7wuJ442
rOb7AZNbbIOftN1V9g3d25z4XME/kNvyAD8JONDJfOfqkeXl+E44mBBPSsl9cTxR
X2kwPlkVJtFwfkgkO6yLwewu7ALvSxd4tKfqUz8eD2CP/KVbR0pE9TMuEkjCZi0J
pZ4zxz1UMNUOA2bZmVRTQU+3n3YsUMaGGIDmnQzm6efY5L82qeC7T1Fi1nkMKmOg
6fd7Wmdua7ObGcK2EQ6h/kjf3rT68c5ndXG2Mw3rpN6WTCqpo+BPKSILWgYtUaF5
gK1C5uQdQkZ6ca7aIvFU1DwIkCd9GvAVUObvHOwWbhKTPvhABGxk2rmp7IYaBBhy
fhRyu//mdk+7YrIRXXVCTBosq2PfynIHLKrcbfQbBikUJizodGpVBuqbMJGuMldO
UmxP8EIKsxVe0kPrJh8KsYKrLP0OB7s9z/Heiiv4jOJj1QrBuXSBJz74Wr+vEMZY
uZxZX0fNiiOAY5UaG0usvIc/mDBqyAAZHRDB9NOsWBPJ/kxFnRdizbWo+6odeGuF
IztURFNL9WgwzJ7FwlokNUGxNTjk5fsxkYFfSOydNYhCVPqbe6qSUJF/B4HTGlZL
Q3851rM8mF2hsGWN57vd0XvzN7j0jhaF0oBCIUwnlkDC72uncBsptN+QL7mCf+ys
f23a7rjeOK6wHmd1SnO9xBkjfyojwo2a1dOQrmyq7Ns820Dre/HRI0b6jJWPlqlK
RGbW7Nao2xPCEmLi8T2vebwTqATxap5h4+XPehmbofQNtDb9oQhITAiqdiwgqBAt
VXa9lz20AfKJf8vT7Gcr9t1D907wosIIX8dskA0UlFGe2RPhPwL/e3DjXiG4egp2
tOfbDtephEECb9WtDovZ3tOjvaKV5pTvUSohwI5VgrcnqCg1UJfe3Yy6cOpTe9RC
2zfpbGG49XcmeLQzqTG7HhgmIbkyLEpvXi2Y6hRdNyrtPJvq5t9f8nkK5/mWUK/d
Bv9tQ+ase9KGsnVJNINjo3cE+M1JSdppGNLLNilFXYO+GM70+KpwRxUcTmOeIefC
hsnzIVU/dSvrqpin1mXQHxrJ8FyLfaZiz25GG9NNm8qF6dN4gF99bwx4/qzhK3gv
QVUodrSEihUeDzzh2erdfSPiam6DTdAnk/tlrZmaiCP60GMO+PWu2s6YlzKGjjiN
jbYXVeiXuDaH19COaETJG+3jypN1/SOF9AdGfQ9XNF+mtSVDsP50c7gXcsuiyE/b
hhDpQymiBWSPxLZ9ScsJSGWRhHdZH66ati2W18sApXn49ShKcVwYn71ncAbQGDfj
SydY/TirxAXYe9toFwlCSgerhl0IqaJyC9XCoU/WoBdx2xqTnNG2/FXT6mjaFoW+
Q2hy1GGaCk25KK3pFwwDysaxoV4t9JWKbLZXS+3mseGgTrHCqS4EkZkRoGQ1wB7F
g/gI0LXewEnsvltPLWWYCBlbPhsBOl/E+2+vJi4n0cp8Y1lwiBrzQxCeuzVE061n
NdI19oBVbTXWW1fKE3MogEyADjMULYh41Y1Tv83l4P20wpfe0C1a887bYOtTmWoP
P3pak96QO2w8qkaVor3fej/oUY7/ovRSGKUl9ds9yjdAdkSt+58TJtdvUI8lZTtb
gDKyZDLXoiTAM6J1yfXVZC8ORGa+7OczwIAljNp4vJSxoGXYAa7mASPzSe9Mw+VS
Ht270NyMw9zdpME4J+OqYN8fWwISkK/zi8ZN1j6nEiZFnrXqges/wiSdGjshCuxR
rhWCIaDe34HkFGIbafW/laYNOnYHSkoAmTbnMZDdHlFPQU+setfpSdMbvGPRZvd9
bHxS+M7CXndr9AImzDTcXaWaK3OuKyEjcB8Ks0WlKJlNp1H1YBWhn/J6XkqkejAy
1z6ZK00Q39lRha7V7MmEHk92kp9gABuVb/ctaaVaaPHjnN0kUETy7FTZafW25SYZ
ONpgsvRJX74SE3biXxqbu3lfZXzayzd7m1N1CwZbJLpq41MV+5m80VAR3FUwbL6c
00tIqyoaiWayHXQywUckyK/uQ4cEdRN7tbNHnI2ndqGHu0OeAeAh1+DCVTAvSAFO
MHQfh+cM5OExjD0u5DMsmCOPJMxkvm74+5NpZsN8G0SRpv6SUuhmfnKMi45UyIYg
8wX8xL7JKo3fKKvhG5hU24SrNf1Bw/s6sz53uCobpkKfdOVFLaW2jP9Cmo8qta44
b2edGdrPUuIUSgoa7A5zvmGm68L5zmt3I3YMLuXlxxZwPVMAPw7R1ItQmujxan7a
HfujwcyMqvMAtcC0EASqX/pjU6lLunhJbb/KwSG2KRJGkZtS8SHsGeHTljdhwfpd
tsWCCinTrd8slTAoS3Vi0SSqQvN+x8qlj8pjCpk1/TT50YKqskoYmwDF9FXMYcO5
3NRETR98MEzoupr/cNpZF2RxgKg4O1CdcvqLBrKama0OOdlOHyd2QhBLaFdVA95v
QM6coLhzjlhEK5IJi0rXyV02QzucUhGCfG1Q/+yEkJyPq+cgD+T1VdztDICWd8v9
Asoya5KjzHCA1IidT7D1nznS0vxTszrqnKhrF1IHL52W8JLm1phSt+wxo0xLAyLn
iKT+Oq7qmEaDHJoofqMzjXDy9Hq1CnWdS+YBLI0oODdw2/1Nm85N7QxVr+x23Qaq
5yfsSDNhuDoj01Zt2gyexMrt7ybdS3NHsq5TD8uHfK7RFn/2om0qWJ+GDFpOCUK5
kEF24BG8dPpiKG2lQJ4r98GAEhtjkf1qmHN0zCIr9nT0WaExSXHXXeLUHi88haqa
uAOQH+TGXkD4ZjsApyqXwiXxc7NwVhTZPCLuoR8sPFeptV9F8lakeNzihavgnPht
a8UDpiho/UuEFRoFZRodfrp5Iwfmj5i+mCRP0WBsqKynop6s2ed3tkoDVE9RfLlO
uCcYV9RrTGxxq+2a+HuFg9MFtnnjRAVmrBjxszDhSaZ45Cs+1a3pSSK7UM/rENyN
RPikHc3mNpmNFhlkmFi11oA5J4al1G+e41kP+R4kcecDB0eceiV0hT1W1F6G2t4Y
qTG0CUKH3glbtVrzY7xu6gLoo2aesaNzAsqGgKtRBTZvtwjJJWdSAFbEwxXzey96
h+FsIAVRMjFDlgmbEXzuZlcjgqgg5N9rJ5bLD+/9zEVMITEDR5PBlxE71mvfz/85
tw6gUzDtH4T+Ax3lMHuK9Lijmwr1+xn2nUzfdUR1IWeEKBt6Do6XuZ78xj0bvxz5
z8hLPRIyDu2OX3piN7lDeNVrr+hG55qAtgF5L8cB8cB6vaIr0nvLJ8noFrFB2KZc
9rbV51Up8iYfM6rK2LpdGDy1ehCOb6wEN1dokAJgJvEIR52zbNbyaBS16Hq+WgFO
BGPeBRAsNA3EyCEHw6+LF0dQxOyeebVIsXqywDsBDDgw2FiAJEDnB+oDwy79iZOa
zYFuS2xPEWlVhUTEYoRpEEL2hMCzlR3Zlr281m5VKPcbsHRRnbrZSIHMrQN3kvcV
3e9ZYZj/hSIhdcle7jpPQSzgtsIUaChm5MovOVf5isMsLy2+N++wCm+9WCXnDoH3
Gh0Kh1AwMbfU4PqPQyQksZuB4Jurs9PdGBRWJA1vq60C6rQeyg7PaIMsjl7cegXg
wnoXqPnBg5Y2Jx+NkCr7pqjS3jqZaGaz/v4c7B1Ku0dI+uSkwL8NYbQ75ckiKl7q
yPd2WBQ9yMmO56ekFPJiJgx4HX6I6TEMHeuexQM/WM+iR05iCO19IzBAxqZLAHCE
T3ai5MOU9AKiEmAdO3T/0WG7or7i6SnjVL9CVR+hbyhi+jOaBA8AYerNPJha5mAL
H1yQexqZAR6MOr2FLb46k3vv8Ns0HTUZbvdU+PA6ObOtCqJ0nwbo6zj1vAnYAVF0
ZAlsbTUjBM7ZPaj+8jr24o+OPBUJfDmTdIwi4ESgPsfCvvMGTpS5tyS0RTn2Guy7
tQyTc58GC3sv6fX0AFFGdbBFD+GMnK84HiSSYX1JdgEEbNdtPO0fOBqvgIqCKonf
S9R7ZUme4dKPhsEV1D1s5hGZe0AR2D1dL1Ovmd0KwYFYk/OnUlCsoAM8kv6zQF1t
zQiKj/GzLafj6UKDPnZhYgl+xuq0d+8lV4OcnjOgCacFZkXqmMpeW6Bg7DsWHayx
d1rRyY773KVCpFeVzszJxH/TJvGyHHZW+V7viH/1giTiFSrd1sOR1xDJpzDrKxXs
gWNSG3BxtFY9ZbT1s2iBOJT9AFLWgJl2lDKmUIGMchUk43ZRQv9gqjeLjYGRRCXw
UhHB/U+XaPrY+T6c7SobdRJvODUG8oSjs7SSiZvysocjYu7s9DdqCeDWdg/IVs7f
5ddCWPMYL2wjfFdlXxVWYV8X+HuOPQUBtSy65fhCCDlytrDESRsa6aN2EyAVdILm
aHm5yRWhsXSPpk3EEnJjhfL3b2z7qj5Ghh0/g3l9nQK+lJNJvGIvPQjwNL9eFb/4
rHWoE0JmlSyPPD7DTkPnL4XzlIEmrCiZN5sV9bzHo/401XbCAhCO9MEOQhkk3FYZ
zpjjhaMO9kuPLhCo8STr3xa8atpKUptBV/UMFaHOAdkmjFTI6EvX1n2gtc39XXhU
2zZBtdOlz9OvdpagfTns5luG/QJ6HSEjhx6V6yeh37Y5OWKiBxR1p7l/F6Ot9POW
/qufx0mTki8oqMwCPnbUZChy1oDkn8wAOhxmEx5ehGuW51inxT2frmu+u2pJbojW
1T52ybZoZRxGX51u5/wy+Nmu7AxVZoSDSwO0AG6g7gin7zY/eS+UABDZwdlHa2jZ
jyU0UVKfogRj3Ag1a/4FuZ3lIFdBJay/seBQcaPVonxPYIMTU+S14lGpQCPcHfP5
o8sRobqCRgEhiKyVm7MaFrFrpGP18miWQztZfVECZkfEmH7bpbOgEatVsqk+Z1EJ
mGFpc3sRYPqrRt2gpeoGn8oMH/pI//AQHbVvooaJJDJMxv3KZZdTdWAK1BS4trI8
zhzva/k01O9NlgD+wab1/eO0cPrn1IDnvsbaRHIBojlO7W5ioiO3b06iUX0XUz0J
Nf/K3qbYqQZcXWuXk5z5kwUPAOqqIiNwyoT63tD/xCChCoMcB8X1k1+zgljcba1r
mtUnytJKCn/JA3hEOMczIGT2QdgBFZlOC3AdTjLq6pvr4psi5n9a9AAUuG71lv6F
90YRVx8TZf78pCrcLa9PPT0B/XpD8HULJ0bK27c9ofxDXtY4SeoKqgFyeozzuI1Y
9AgYi62UNSBEfvHuqft/RV5JkzwRP1ifQsyOF8P6wHAwDMcupGFAvxbbUhNJ9xMA
31A4I+dS3Ai5zbVnbie+P4rmtKQGQp6lxJ2IC+6orUc496h1TmXc8c33j8XLVzow
ru2vlCQxPJY4g1lPjYjRnbFEQ4PcJWvLnmSEhh3mzE1MKcn1WDcmMQV1VV8QOwmt
u+CNmYS7Wq6BDEzPFltnoUmSoTkNDc0Bz6wzg23CJgCMqvybfqa7AJ8wWQbjqx+X
+FiHUsZoOLt26v8cOE6toVnBnjwWZEf0Z/F9QdqT9eFv6ppIUT+xPUbaIfQATXJm
W3fND1j0XPscql1RuE0aDg9M+CJknT3nkWAaz5vlJ5MByhI7tq7x2Fwhg+gZbc/f
ZmovIYU53oYe56nLsrEVm/h0uBDuB61emq9YAuiv+Mn1MAfRITMddviqRGMDzJl3
QgF1WYEUSsas/4jRaAUADCbE7hwieUyvm2AylkqymLKyzKvVFTPN/Tjhwx+zq/Xo
F6yDS+pm6wrer1PddxWX9gpufBP7boEb/e6ud3jDDukc2dpcTh9Vgyu/RcS7OKc1
vubEv/mFtM+2H/b4kDglyTw/Qmu+gBYJvSBa8TsrTwUdj5QfR3/b1SSM83PurP5n
RjEPRDWZGtSp5ZGI5P6h/mN+UOdtTQ5Oy1WmCuROybPDr1eTA87GeW7V3qDmP91f
YxHumJTo0y3CoOHmeT9bPUGZE9c35oua2qrxWfWP47b2xE9wW+Ofc/osM5a0BX2U
hRKV5jAn+Y9PWzg94d0/NZh+Czv4q+4lT8DWTwQusWHqFk/DbCa3/EBraAFizFRb
p/U/LypTkf2EFhNNPZ/FjYcaNjzjCnKMmsZI0ajk7g97FyJBxQcI5m4SpZbff0BU
urzV6QIQW522F815OPKBm2AX+SdyElLwLUgpsgjeF7+G1C5za86kQtpNb74sUfLf
EMDFrJ1uYy3qVFAphgRShJbyZmQeNQ588/lVK2bDm5TJB++bSSbXrqW6qgpreR5v
z6OkPVlCl8SFOSpNcFZtPDR92eo8+ngR+4veTQtQ2X+tdfl38rHu5xsyQzUin1hg
DbjJUg1TEd2SfXRutY4Y7s+Oj+nnAkoM5rG2B8BZNg26wDxyroSvgoQMVk/PVui/
eHnhBOD25raAA1oQYXoaLw7WQV0yLOqWnbghRxHDYkhvnmR855SWq4oNeBc4HQWX
qf5dWRJi0Judfw4rYqCKLo5aCKYch/TeOsbC2hRJtUfjzYHSYE+IP7XVrK7i7uEM
WlWLk+QPdaGe5n2eFcBxxIcy/ZUQno+JbwQG9b1RIIBQRpg5H4Rj7yCnwwkeSh35
UtJK4OjvwpGykFn9fORXXoXgsn4IiQoysIIj+v99jfYldQd70+L8jqPUWt0f9yG9
UanBTwThnxYxOTH0cPr9YpZIdm63CyFqoKUkwlsoLgjtuNHgxptmYWxaRwpuV8AW
fAtdYaqWCir0Aov9N/+jEGsNjo8upwINLIgKOJogXaVGUR9qxr1iriNBV3ESNQVp
d9m0iQ5cR/EgOC/DmQEvPDzAyDM3/n9NZH8mLGdp9/7hWTfR5eksE4y+eURVkpxE
9fPMhfgsocn7oTvjO0WF/zoMH5fWRs8xaguphsJysFeksYIQNjcgmK1bJCfESCk+
+7mH8j2pYy5umUK4bCl+xGmd5F23AAIWNGx+zUOnZMiTx3ZqReNKezCJxgeNUGEd
2eBkMjYyU3ulzzlYqOT8qTu6eJWCzK3qM8eDrFaAgsBe+G5t4VvwhZBUxeK12FMA
SyCermtnaiIDIrOlIxFVaNvFbrBc4N8RV1Rj/qnastGpRWgySIxkN3QaTG2l+BGl
6slaWCrJecnSDRzLA8V0KPZtAgYRL47LVSGAdt0pPTgRKT7TU/jkM1genQsE6bKs
UoXMoYdEYjbz5Jc2jIQ+s9LL02Pe43IR3Fhsq4P0CUIR6k2TDZdGjg6Z19kv9rw+
sBFB4abdOICNkfsuibnnAWG1KFe8jf78pbUi+JOHZBWjUAjt1LvP9q1OE2ACYgjT
QIm/WCW4QTCTHb4QmlikJxCw0uMHEIbJ7GObK5Yx/FcaqM+Cu6S4U3r77nB3VJPv
g4xUPEcuO2MMzz/eueSPotlmbgZ6lTkmSFPZ9jRJz4K6L7itW0nFdqqqHUaNU7sX
53T7CiM1OBb/qvwWyb8cB8V7qXsXYwpOTMERpMwh4zgpM3m3nmrMWVWXuszBDCmU
uoHh2MXHQzq7wLqWYGODycVHnqz1TRBbb1+IdyqCiNc+mVTec4/I5Gl3Q3nGMTTl
iv7OpwbPHqh6nI+JDzuDoYy79rfjsN15QUiJWLuCxwonqY4gyhWYHbPoztSmwfrU
L+wjbjsi9rXpktIBmIxtXXFoVD9kugWDjavTBZQr5/Q+WGHsZcxL6/CqNPzIOgHN
QJJXlAFTleS19PRZZPB3uRkI/aI1OeNsS/E5cuFIX0PFQ+0/8+rENlkro+ezUoy9
BnkItDBtayiOFAyuXNdF+U4dv4qIdO0LpwY6h7F4SXy2veeIQVplsZsp+jvC+iJo
GBdHSU6BsGakiutaLTBf9ENZBeCluRyPfqpV3unYnuK6m94ngQN2Esr7SRGh75u0
tBzsM9l2ocXPHFI88E6LsC8DcckZLOb8j1dQEEKxd7gkVMSYbtgyiikXFgSkG8jX
y4yd7NWmZxz5tPNDnYj5Fu7pu02LhyTVZDNmxZ3AateqND7GLVJIJtn86LpdR6b1
te10NmJiYDBFiDDhwbE7t1I8tmRc53GTcx2/hw6Chh2Z3yt5n1MMWRfkkqz1nXoW
GTs8xv5Nn0y2/N3u0dm1kPHB6roMPqeIpLTxISH/FiLemXbS+k92W0aHl1DK80Bk
DZflMet4zcyUrUzKAzB+ftMjnHQ2mPETBP5VpMvgYQivTXbFhYedLE25kMlqBU23
ssa2n4dtGmEPI/1D81H/dieRFSujtvV+RZnSiJENYQopKH2l8KXoAvPQnPZfTS/A
MYGtlJeUeEXHN0eusmZnEAMuAx863pXpuLMhm8MKY972f3kFbOLfmd5uAVRunSkD
/Nr3vVCunFvnHHTGzVOEKIMt1YcOa6/q/rJEB8Ntisr2qtch5JujIr08TciDrWVF
y++JaFx4Xch/RdE0zQ+8QB9/QEmU7yrJweo+DbWRFvCOckrKmp6yXG6rzZ9RjWPz
TMvU4L7eKvtkZrU+Hgw6GALs+21HWui5YWdvPApZlZ5rxDkKJ2a3oRWRWTQbC4kJ
rR/O5XppunoM7pY6+i/7dTkOi+Pdz8/2Aj7ixIbm46z4z1CYx+E1QhLMniXcBtIN
rVEL4L9BTMrXqJ65KwxysAiFskF6e4sVbnRFGsHBzD63iAM27cI+3O0z5bOnLWMV
2p4zUp6Qlv0P5pewwKWUXeedBrsqerDoHQtgu94ESRLSZEiVjViLhSBm4hip4Ye4
BD7USvPR3zR5lWskyHogSF8WjnujpP4FbcwOzNfRYQR7c4HMxQpdp/imN3uMOxz+
y19btv3c3cBtPX7Oknw0KRRYKeO8fSERSUXmencYMHgqP5BOAuP16lax5LaUU3co
WlGYDUeI07NDTfk1TBd3gwWgi18ZxoTQVi+jm+BqXuxmxxANYTA0KdIqBeCeMDe5
lEbZywfMAaCuLfINvv4YhqM2at11v7Ll+cKWoBYEUhH4gbA+zROiPzcpLCjGjhBk
jSwZmRh9bpPVLK9SQUkq4Jki11zOeKNNa/jTKwq+2Bx1Dr3eFs/52fFj617k9x89
2gQTQNwhl5flXnkY8ExUCQ9fRda+ms+GoN3mptmteHt7Hh/lYRrpQ1HvEQzUrpqA
U09m60PdSodIgInwQkUhKbGs5ivyBwU5DTy/eoKp6kHxc4S0FGt7ArLMXJQ0GfQB
bc+fqfrhSoNTqFnm3J41yU/Yde1Rfzw8QrL8DQPw6j8QueaHmf5oiqa23/qBb1Qh
pR9oC1XVmKw2Mi6x3xzaQLQxuvFyNU23A0thiTk38KaNIhY4EG0k2C7lMXVfP5GH
i5m2BqRdt0uXTzvGitTmHK/UFhzR760X4PFdhzqmt0g/HXkjvWReFPxHYqxAxiDX
iSPHIYBMQNh2Lqz4bM2f5FJ30YoRI9WDlVsTHgKvCREMiygNj20R/sCYCnNdUx8T
HYu80fkBhlq9h5yvMlFSS/HTBHFarnclDzNlY7HB4+mG5s5H1GXquXYGqRldw3M/
C+DUCXk0T2hVl2B4j/2LAXPjw/5KUejo40KKYSX6k0JFUtmoQr96e/00cHdeEfPu
w1kdZaIyXiAcGcTtVm/07nKaN6vqw/fDNYHivX1xCmMxiWRG/6hDFGJZBoIhwpbR
1FCu7dPZglSGDJNg1I1yG19xt4AXXcy4E8VjQUinI0eGyLyKJlZARV+it8dKs3cz
Zn3FgIgnhAnBXaLe0XpQsqtxcybBZHYEbatii6+Qs30mFRsGm3ef4e6q5cc9FdPP
reD/B2lbcz6fWDOeMTl6tFIAgyaWn+ouOEs4jFQbPyc2ZRpITyy1lLbDfu8qCrqI
UvqoReAnFjfl0XSzsvryB6yvr8yFgRiB9w7MN/An98fWIzgM3fOhWQ9O3zXYxhhS
5zsLFn9VRP7LskQuDHVRgtujvr5PcTgKfGu+0XhhcgmXAhZW9qhZEW/Hy+a0M3F7
ajXTOIOQ0QmwQQou2VNOjKEN6gAl+uQL/nnVfLicgsQm1JdjVjoJ4pUgwpEapxLf
U63pcNiIjdoNvymgG6qU+CTzexZOgSlrBx8cLg+rfFe+AcAOhROu97FYpVJPzm06
/4/hk8jAiMIu4CExdgJBhuXqKSotw7EybvWcDEOM8zHxdr74i66bKwlTVb765W1E
glXHB+/lKVMxUwWS8dS3nl1gzYgPwl6fVTEi37NeCR9/ukKeYx2ggh43AYM5YWog
4eNbrTlkaAqZ/CLUaxj2aSYfPn88rPPVEIntodBQ3g7tvYc/mwVKbf2rA1PbQyi+
rd8e0Bkg4098Neq63rdgAxD3ad26zpli01LrYehLrf3v3m/ev95tLwnAurKVq9Tv
Lg7rW3mOvNqu0YgRMyVrnwSwq1KqH3kQN12N4eL+U4zKKwEuegQ7Z2PFL+ycFn+L
dY+pOSWs7TaT6IKK3V7TnWIBLoVa0z/VX+XBdP4yVtbsdCM1coE70FeXsbRYwhGn
vOuBZPCqsdtkkzl+TmaIqpagse4ohnmvGKexLKJMuclBujx7k3mR202tRNxZBBJR
+PBeNhajox4AclAqV0PjX5S7bhruKlBXMnUAlCfdViYwdbmCKOwZ3JZ8z3zCL59D
cfRXa3hOgD8CKFYShDo6mR4X+JS++qmRuvXHvfb770FjNX6Mz5XbXP3KokhGfOuX
g3M2JT12AxlOhJHER5aAxr/dSUs+BjqpAkuoD3jXLigpqBfveaOkzkGc7H4PUeAp
oUPNppsLfdQNaZub1uzcShl0Ny8Ao4RDV4ffCVYj6aCoXYgtVBCcja/5HxOBT0mH
x8ETknz2V1O4KkZ4kkyCJtY/76y9AVRhhoI84y1WibjBEk+PC9t/ch6QriJcTt+j
nvaq0tWJA7xrCehq2+3Jl+0pqTsFZm0sEML5kRiFq1uPJgZ6x2bFvHRZIYDuiSc3
y0gBNxL/NIZSJ6J70CW+fwTbBMNFPjmRT7WAGYIvkwFXJ7UQ2s8mkXX13Cjm5Unz
00jLjAaG+ROjwJZvEFRq2S+r+W2J9O8OeWmk82H7oVLzv6pPYZYUGLEAZDEtxztY
qn4ciVVivHvA9+ISbdwE5wvAIw+Vv8dPJsGtXqFideflrlpOEC4zurazsztTgQTQ
t2KIoTp4JhKgShmsU6gZ66V9uvXYtfnEi6GDOhZ4J5HMpQCy8IXkTn6nkj+y02Nk
iojXM0ArQTPg6kJYTcaqEkzW2eCXs2E7SIWJjAEbn/vLkpOZerrUPk5gTTo/D7FB
vXKGQ2q3WiFETz3kwIHlFFK1ZPGlxhNqQY/aLgnvGN1kXQSSp802HL9AllLGrjMH
boZvB7klVr5yoET6aCd0gNnmMAs4J0mldm+62zZJgFtwQUW/jbkNRGwBhVscrQJk
HZ8EWB6KBoMK4VY1WWGjdNOwdSMHEvgIPLIZ6Z6J2HTSB4GTnU//VA48BZHV87KP
Mo/6mP1Dx2JpXdTfAVopMkxWZB87BDQVOL4fN/fhBPdiSwzjXeRAQknggw5Thvx7
YY37CfErgNX1LhlUP8N8dz4TRk0keQSl9n+o9mrj70ga6CzZUyqJ5Rk7LT/v8ofL
O6Hoq3NjSWoPUXeK9AtQlo4rlL4AkUqYEbcNoLqS77URh0oaBC1RnfKpuR24x9pd
E+cH6noLP9CsQ79zrJ9pZGuv21spl6zCu8W7kksDTW2usxyJj6HNS2cK9QhH+yDQ
YiSnzhIUzr+jcgyJFCucH9l2tP+aBc/IXMZiqukkkxFz1CqHE+0i61iuRZIJCzGt
szcwXSJWl6S7rnl/TY4iemLQVtprjsHRGMiQe4aNTSO6Oz+SExJA2KfVL+wKPnzI
ThT4zLe/zBLKJli+q5HYjnsaSyoRcp12bMpzK3ckSgpVyrbb9Muyjt4G4UCmSN8t
iPa2VfJH6/zkgP17CfzIb0nrYmSDszlsBlM/YO2hf6JmvPjvFOPVEpZX8ZKeLKiR
07T1ey/Pz5vbJ4hspakS8g==
//pragma protect end_data_block
//pragma protect digest_block
SD0bL2FCYlo/kV6rzgWdBN1yebE=
//pragma protect end_digest_block
//pragma protect end_protected

// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2019.10.138"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
t9Cogn/g5rFt8vqaSvw8zG5sll1wRUiCR4dmVWlYndlL0VCsID+z4Z+wkTaDMz/8MJ4exGtRw/7Y
7i1LaioljsmXfyA7Cnr3I3vknwpNGob3VhfzYChcrXbJxXSS2afE+RFVW8Pcpxi1T0uDJThWW90H
IiDYWjU41dr9aSUV1SMBR+RVg5PFXc/3KIeAh2Ykd1I4+l1jBVAvCClfrx1WEXDlTojaBoNl5wup
mULV38T2W+L8hVbzy6czNEyyqXgS1OqiZy3HDUen/EiQMl18KQwptIqfX96+WMJmeBKi+F0LQFr0
EhIDIxl4ZW5wztf7A7KXm0EusqKWcVO1WYvDTQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 6400)
0hTb1ZYYW3fm2PHFDJOFdJxIXHb/RG11kWnPBkCRTa7dIICMmG7W5Axph1AAO9FvHZxj2iiNWnyZ
Hxcoe1LokQMoc33IKqMA/g0SqxeETQSKXTyuDZIoVg9xGgIuKuFEx5pLsEBRivMqz9U0JYENx7wt
K/2JeqbLbJUGNcgMetrDhyHjbGEPmoCsVjQiHE2ztIPISmKTYuDMfNDoUiQzdLhi3pfoXG/w4j5f
s96Ul0oryVMTZY6CsUyuOrk/y2VoqBDvnEDhtcEEIgh/WQu/w6rHHtoJAjqjWc4toZtTvEYvRmE8
ivilr1UGGHFQ6V5bruF5Ht63qCF2V0S6DD0iUrUsE7i+E+VzqYoMw5hRp7ys97D+yWC2U+cTVpw9
TKodBcF9VuENwHKdFwvq5/qk1FtIAYqT2cGr3ARJjMbm8Rx71wTK4eq9tg5nfz3wxI7H3b1mED9Q
6jefTMCamC7z+zDPM9PwCqmEsFLp/qPmTEqKAJ/3i9BluQgsskMkmAhs0Yo1tFiEXuQ+ElSBJOLa
FCDHIgbjiVrfVrRut279Evbiz03yCw2tc/mZd0S2GSG09l2xM49K/xG6plyvAs+r6ZfpOQwLvLfz
ss4hcx+BgBJMy2jlJOItb4rTQ1RgGorwy2VyhL7+RGmgSo18X2drakLKKZ/5tQhgqDPerbbR1h31
x+ID6RCBwJ2kzh0CyWXBZzf4PVsD3QLANnKFYi1mype2uTmAu5JcBi8FIk3UjwKTZpymvLIGBwpc
aWQzr6CG0ial4wwMA5z6InOozphv7dGz0nCqFuKk3AByF5xexha1hp0gSptMr98fb2Hy4e4RndWU
v3jGcoNIkAuiaflNS8ruCtzME+vy6tLxDUqEM+CA6S74VwzjI4FlCqH5bz8GoS1J68TUfZiunnt7
U+pULQuRM2ACmhh1N3+zV4d6LoTJhJETJL3EnnKRxObAmQ9bqrY5erwcWQXHByqwa97HpRyouIb2
AQFJVkWSwCKuwfwVYzKZXLP5c6tPQczuFKeJWFI34xdWDJamR7KGuDuqngMPziffzZW1hiKcrsZF
TOYLEnRxvvshnIvlCc56FCdclKO6D4NwTc/vy/SmprwW0PfCA9creSDJihBLkmRpF6FaB074XDrz
RUM4nqcPwu6z3+evwpjrzSoi0YlIBNLkaXqGR6noTuyaKRzzblGXcqyrSqVogttVl2Mrm3I6y2nH
0IHMXfe49BiqlfHBP8kBptBu6NgxlrhP4B8CwlDvLbNttZk1vlf8Vu4WrmLG7V7jQr4TFimgoe3/
ykMFw4eFsJSHh9ZCP1BOIn/gJcUv4DTovrkJS1WnAe6bLHpVjouKGnivXhA9E5HcUS0u4Dcl9X1p
IAeuwwrfn5z0FvV2Ej5Mkn+Id9vm46W7sXylODZHtEVBOycOWqFRdjpJG0lVD8ZViFJ3EQXgsKDH
wH32C9qWmxc/plCMQojii3ae3IO04SuC0qPHPeqhB30Tpk9M/Tvt38tHf/WI0p8PsJqMRBXZodt/
R7m98uHVsKf8Ij/cDaI8fuunWbOLFFHHhP16Qz2S/BXtD8+6WSGzJ+/rklmGmlOk3YglLlLfjL68
oOuCNeBeGFj4QnkmW+hhpzDLg9w3hYU52+ZvQ6teCb1r0HMVKJLqNxL4egXHBqYoPL6kQmPxokSW
EY3n45KqhRkdvjmoE5OElI/pdgAbhMcPaXvKh+iM5d4hHu02eiNvyULNgqJGOjrQS7igJuKfQ6Wh
HYIIDsKo38ErjUsbU1AWh/XrqCLiNrOUL4syr4Zvvr92X9hTT/ZGtnyBj9Z4XWi1zw6nNzaBXaOn
VZWQ4DrDTTEMnwajiwUR67mbAFqNqL9QTCq5IB61NgkB/cFpuhCAsz7NuHf4WRs8g96n8fwK30WS
O69MKrU/kNE0D4BMKLoS/gboa1XnilN0a50vUVFWkwgu/noFgGXWM9cV4uqXC7Aa/VRoGqQbXz0Y
uy0XQPAfr8VxY9hWblRYJyAqWlsdOaja+rzdd8oKV2LtMtD9msqULsLYa6aRK6N5ktgpLnukvnP+
WmJH5Jq8EFeqYLb96k4S2PGwNnLI9f5VZrDqBdF2C2Q6lwAzBmzzq1WwqHDb6ou0c9TAEhDXkq1i
q0D7+jY4Ocwmrozn0C9ypqWPle1qJX3rDjA3dvHJi7K+PoerdKaz8ckJ0L8fsKsTCTB4pGeJ+79q
nzCetF58Uh2KDs1+/kORVc5w5TWdrvPUJ8JOkXpnX7b0npUuSyBKkMW6O9zVa0Syw7trlu7ieRfE
v2aKKfr5p1f7hPdwOHCNZpqDT36ynuLJrDWGV83ZTbn9SZgT3qNYMTtuDtYTGlkOBpTOkfKXmy62
vEGqtIwI/L+i4hxInLX1zpZWveEhe0u7UOi0N7w0BCQxPUQE8iNCE8TLMWJA+sh5xg1NUW6Kz2XH
6boofUhNBS0lRIeZPQcK5gOcxIe1ZkH6knfkcJJjH4DamGMN22MA0wCwxDnjt8jKdVxlZ8dJnx7A
RpqElE/JXMq5ngpUR+NA9rMocJ9xRqthDbwbeqf2qVhokiNdRt/AKoDb+FNvrd5Ytmo3jPAylRI6
AdQPcn6eNzBEok83e34e02Ft1a+J1k46lgFRArz6KcNT5t9fv6uyTg4fLEFRHKtorSTw1tHqrqIQ
dNLwmx5WqnRz55xsbfpUQ0N3Ua6mNpk+m2hqhifZPckkbIymFL7Z5v2bdFL96uepnQ81fYh3N6Rf
n2XNlr33foXKezi6qbDgMnUh0/tzzQVH5tx+roXBBFg6NZIaitskT9LgrO2qdXUTN4rTr8c/nrDK
IlgQn6ISwLz5jfAzVkQVwjQK5J7Z7a3ExbfocRB5cvpMGvyEC3hGr/KTD4hseAKrN7p4pI/qCRZR
jxG2lQ8fb5/iH9zu1yL1DBphLYWDku7L4ZakMJV2viupk7zK3VKe81KXEscv2FkjboDEWUryZbpf
6hE4e8lAfJClBR0MUW5P77MXy3Hq1whrLUTsDL7L9l+BFdp3CjQgHP6hyyVD2DSAlv/1KlmX56i4
EmNK+Yr7y+MOiDK7+IYLsGMvUaQKlTjsy6sSGwlxGo9yPzWJb2beZeSsxjZMa4bdiHy0Vr+VsYZK
+J3dz/2lIeeOXmU8YPPBjVxHCpNEFiARo4oCj0ci4jZxG4cfzkArBAcrow69qCu7WbHppJFa4Wa7
zwzR4EvwbrZk2xVhUo5ETfeYsI4qrjmPBPzNLxsSRXmA3eWbL2JQBhBpYAkrgFOwl6igSn8fnDZl
Pr2mQAF3Hu46brOL2zbQwaEFq4EJdYRlaNh8I9mbg35hrJfSVXMrvFCvnWuQ+biE9EPQDSMIYypE
RpIb5d7/WIWCHTCd5TR9Nfwy1Ez9b2A5f/T2ucN4pXLngqYfM73l7h9pjmgnoXRCLHBBK84xD5sO
VrTyjTUoaKQS7WPTrPQg6ipgiypBGTmV3yq3JEnGV2f6p2jDd6nW28UMHlY4jWDV4l/b5A2C3Yee
guomPgS5vjEw/WjlaFQt8drBeFw6xoDn4fHrjG2Nvz+19BCVrSdgtFuHUi+6eWJcRYBJsW5qjkox
cgeWOlFPMjbtY+yDSKJW+YHm8NHuZ3TIP11K3pPEEs6wrbfFiSSnR3GFYu65ulwk8wpxwf/qx5Em
ANsVpMz0xKVBzagKN509ur90qSBbJQEfeKgmyklCcAnDi9C2GqCPvIWnRlO8Kwm8l53RTbJaAwWX
qVCGwX20/VblGcsaWvbWSQncOIWje9LcdcHXOr7CBXIFBqEJ04o/FaIvfcInOTzkjXMpcQUm+rDu
LTXdoq2zwVuM6fFb4TTsDbireOlp7c4PsNjLe4VNgr0YLV/YZSWmI0/PmK2RL0Tc0H3USVAsHNNI
OM+NtkuUrjTcWINyIgDHawxY/BQjbvZbD5/7YlVsH67ffjaTdr5/AMAFqto4jfWqGse+hFfo9DQC
BmhrE9WX2/puudQl9qdLliELJWC8gd1B3gCQJ10xNoc42RvIQM9/vKfcVvF9rFc+UTqn6fQXSgGq
LAp5gpmNwucO/zXs+No2UbGdzN38peSQGub1FnHFfAMXQt7MeU3rNWAwmIv/QTGiXRO55bVAo+FA
CI8ybCiF77cs+ffa41Ha0PSJYKoEvqffYx0Ji4JtZEkDIfxEFb/xwRTNSzyqrjzhZw5p1lfRgEA0
9pY6MiSfCqdrc9ApJDYmw7GTkytetFyEcFeYH5zZq4YBpRKJzz2DgkNFXVr7gAOxIk8MfK+8oHeQ
Os8933scb84eYW1R8JHQz8KtRagLM9FUD5XAQtaVWpZ/Iv/5lOjQc7Ujn8fZS0EQbHjDGND2fzfh
x2SNTa91ARQ9sdoud4QC57Y8MXbS/Xj5SrLt3a9Nc+n3+XJSglcO+MTMD28WZPSRSXyMOoodTg1k
Wku50505HxmztKp/XK0QbuLNCmbIlYhquDhOB8zcKPoZ03rHgP6BrD7KaR78CwyJdAN6ZCK6RNKI
+RDSYjjdbja26kPFmuVcBs6HeRsTQZpV+zZVJGS3xri52eQ3Ky3Z6ugtVtpO9pa/E8S+YVWah9zz
5QlYG5dHV6/MWRTGKhmSBisYn6tiLoHHTBe2Fs1Ntfg7ipVmIWpd55duq1Fx1th4q9deI3Xrd64X
T9eYOrVGlQ6RrGyPyKM7OZvGUbuYWmEBTA4NaD9EtnAsf76f6nBF/ZguXrtaGU4JZe1+4fHK3XgI
UtpCqzsDjQiTiYeZCn6hZS8AkWSL5p8NGWfL9+U9Kkg7ps9MlmDuFHw3DIcqv/oEsO5fnQ+3JvKR
A/JNOPOA1iweL8tUJVqg9PpUUkjlJh7anb18U24FiOOv2ceAI8EBAmkSupMhXdMK/PsyB4KUYzc2
TUpyY9SNXTiM6I8ihUlR7vz4fI8wCbLF8wFtZBtUIp1eW6GGsqP8eG+CO3Fm9B+Ww4MLqCFBS+l8
8WJs5ILA146oCpL0HnoI0KIvsuUT8RgimwbLe6aiEZ731nliTbaJhaisjC9CXR4fXcwL6qwYGIcd
1hHfBxsZlVyYQOjQiT/c2k/GhCjoP8RbbX6w+D/CNV1ZAgamQSrTZZQ9r7l0XBfJZvccp4YMo0QS
sFyx7afYvEZozMCrxZociJSa0OgFNuoDBrmvoBjUERzJ6cgYkBcoSnUev0zoO4GbVijOBQvphIgf
C2czwCkrckt3MenZnsPvGWl9GYlAtvZ58UIVhn9NoVSxug0vQBtCsa6kkLVlGYq5bx2XmzIl0KnY
Nf4og4m5/zwnreu04iEjm6TEXQd5IguW5ki85Pz03LoGADDvSinfFvjrJXkEqelL1qNsug0u8PiE
TNtGI+K3xEEszEcJWWkFAXQKrjlA6WDnAK/ki74HTOqLhb1T96t30O80Do6iNQjoLtpCceejTgRV
lYiOI6ydcB5UFUPDDZH4b8+wxJEUD/03REsLJ7d43DoDwoDerkebmcn/ck7tGyXNR/Bqz11cwkl8
AD4WR8rqC4v+n1Iwn2J3W1En1/Lv/f2oqzxz/sc/epoadmmwmiPb3yoecoXIQr4V6JSSNpKjM3oL
bW0YHwg6YMxbGtuqQVgTqFXZNEY26dH2I1yYpXokiXZWC37Tw4H8jOAEjoQxqL8p7HydNeVn+VPg
YCKu8jQw1335QF/YHpPUMFF5lodo7FqgLVlb46Q8L1LR1l7yBJBs3OPc+cU2ZCHyOmhoEJVNgFg0
nascnCXuS+twLfUN4T6yeCO0O3M16/YsC5LnrMT4JBim++UlRTE00ixEJxKXMAe3Nhu9fuM+yfPG
KUvMFX6PwvFoZHoqpOOjfdp8FRhHdwIb1X3sM0jHD3GzqNfo+Tp8FnnmQxIQ2J76khcTHmIRzOZD
W1/iuZ/lowAKOUHXzQKaEv1+Lkx5Hr44wM+5MKODKRdJGqc8QehJXtBK2TvrraJRtw7t6rSuzNhg
WHrFeQMpEB6Mh76RnOY7HT5AKhL9/PPkpm5G3zI5U7tFpDR+7r5fkfutv+fGq51GYFqjXOkA3j9U
1atoR0rCI7giyy7+70OAyJ/e8h7OE2jEBccfxR9DBKlp4vM8rSvvA3wXOB/UsxfnLGGfoHhbgJ2j
G9xgBZW2rNdxnu/XUjd54P4GaabNKGl6ThJmwSaMo5HJKPoywGGnamSiIy7KQUcfAtGJ0Q1qR4tm
7YD+zPkDklK16aV8ExrFPlCn6Ftg/WAyuhaWaSq/nnpvH3dryxXoofn+zW3BKxwbZ4wCRw8DOCMv
pvxoAfN8jiSSikAA2TLAzdaf0mkf13BEjFrS+L3iFkQk3xUFoFkP0vr0cfGnShYQGhaVmLoa0fjh
HahEXI1DYt1nZgIV0hUSESzEdBkT12ikCwDjwRlNjig4tTku6Fnf3V5pG0ZkmS4kkffP43vwgyj0
Ys2r/MFZpaQFgyjM+naswj4dmIpiN2qaINObsfZEvkLANtSowpI+9FFPFTPLxEmRpOJzCM4YRtf7
Vfeb/humEXWExxEAi4M/lZ0cXHPsIq83zeADrvRm4jDSaiepp3y+yaJvDvNJDNgo/UH0VnP9/E8C
tPNxwyAG8pT4TyimTNoMex/UDzOvg+y6D60uJ/oaImV9EMyotA5Jjd3l3NSV3nviLcRD8bRJhWtZ
uUOP2iovKrlE8a5FaSKBdfwBzpUnE9gWhmgZC56dqPBMfq4pvTSSXWn3kMz91HQRkgxIeL88tBFp
OkMAaU7grxlPowxbA2lOOIno+Sj81guLIZP5Pl4KzC5KjUQa973CONFFWieG+1APiEBLmEwACPaC
PWdKP2o5sFseskdzdVDdpAPwmHRXMVqTLq5BhdjHf6EQmhNgqR58uCtama0W4Laic86AvIO2odPD
fy+NugsYMdMbwKmHnORicJsXAnHjmwdKz681BWHC3XQr9OCfAtewzQ1yRU58gR8gn5vTPUf8/0/B
p8W74vghxXaqRzwlHc3ojf9Wglr/8HV6q1PXjwik7n1OVp4Tudie8IBDsJbAb/+IePW4shDcO90x
NFfq9Nk/Cn3j6Isf5mf1Mh2l6D9VqfDnp5FQeo7jzW2Tl1COL8SducpHE7Pf8HUmssETeojwK4+0
BVzIc90Cv46afz1uhfi93GJUrczLRAUc35hheAdf2ym8c0Ksrc2J6ijeaF/IzJWpoba8I2MExVqK
YHCaaYE2ELfT+oiFfxfP4WA8U3G0ol55uYK8pHAB+8qgFaC6dTWn6g+6UAnhJbcD0LrILKwz48QZ
xfpSJ522IqpKAbma0AJsctOl04riLwLSe0bWz+UOdZAobihP4O4T5OMbcIlxAZ0ZkO3TDBk1zHEz
1hGdNbm3/RiEh/QKmZaIqvN7yRWZygDOzQk7O6QZPxNMjHEoK+jvWavT+4DxuS02pxv6QKxd+2G4
t+0hwmR8vOfOxIrnGeTibjzVFP5kjMq98pNPY0RcicbdZ9b/HtCkyO2pKZfn/zmYRQZ0qt4Ru16e
/K62f70Wzax2D3XbX7ni9PjJrX8hSdVCxZpmNpc7FV4g5ZTwHiM3puOUZWZ8wmhgEQDS1/rXbl7s
d3n6VvoZmUs7ZK9ZJEp+0rAO+cQ6WXg9nRQ0S2xJ24q/JdW+cmgtw6cmMaSs2VW4CGwSFHhZBKIk
2viPYXQx9oyfgEFmufh3ehHwSlH7gZ3Bm7+wyEHL3lGcHsOYJ+k+yx25F61JoXP8m7G9OLtPIV3t
ZAKvuy9KcTPej54GsMUhe6LkQR9RiMaP1GtpIJkHT4VOZy8zE+St3GcpVFEKUZH5BSl/uda+ntt3
Db8cDkkBWtJnDJGU7gSG3X/mXgjvT5Gt9T5o27GMUetlxZD5+CpUO4BU1cTI6pjMwczIyMo6lQrc
Z9CMCNvyV8uuSpXGS/o053ZJaCktL5VtaDjOnCyU7c9+/BVD7m+v6iJqRA4pb6ESk+WCzeG/YxmS
DvQgXPXMz8ls5ETqWfWzfTKH0cWEWMrIBKwt8n4K42zjXQqe2QCB+zMGhrC7E5F7NNBClncVfHh2
cS/etW1pLgEgJ0B1t6XwUK+RBMKqwou8Gw9TJ+YczppjXoyqo8D4OL24t6frXqyfBkxCqvry/PtG
+yf05EaolBR1nfvejPHr6DlQTZ+Hta36UEnRqSn7xrWmdtBs14f8IzwbVrvF6w/Xxz5B/iGSfCFF
dEidVbf7aQJyWDVfLBOnBpReukDmCJVf5sA4H38LP1L2B0RwYondXj7QvjMl35LKSx1KG6/l5DHC
JSvNY0rkhuQlNKKJ8OSIdMe8TrEOE4Jq+pcnQCG7fsAGNjnbvpUYwFAYHPmKqD4CP1f75drXrJeo
1V0DXZ5bT5KLgpsQauudbLt2fZaP/aVTE10M+awkfVgBnhhtnz/cjG+jPMJJjV2dz+fuJajsQ6Wk
tbfqRre6kQ5Klb4znQYgT/xT9MVrhHWfBhx3kLSVy39kD+VIPUVz5HcDUIRYTKsSAcjwBruhUzbS
4XrjJ/ijEYZhJWZlg2SUbNLZdne2TBXL4akyzxeDBZ41jTJiJljq8vG/zo0LRglyvoWb6SS/Mm7B
9EZ5nX7XY/cU7VeBQ7N6UQ==
`pragma protect end_protected

`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
SmaS+UMhy7s/8g1Wj28d3O01DwUOFW719lzULnPL6DsxKm86G8yy7hJNR+FR+6IT
3h5WCR7/ukOCm81V3QKggLQKNnEl76FJI26FlwHTspk0/y6LGbJuhVyGcZGgzkr5
Yl4Xy3to+SxrJ3rLrK5F7jNK6c+nfqWPnOFWFjaZzH4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 14448)
Rs/pCApnSuaqiiSkDV8ygT+cEbotsProNN1QMWI9+sLKt6C3fzkB4RFuLeRyAWbN
UKnu4nhbjQz9GovQZAS0QFPlaCX+moIsZG/rkqlBiCfMhzGrbdABscQ8tj4kxjWf
NqNYzxAm6eZm8O3P6MPdGeJmQbPB97sl/J3x7dousBHrIO19i0f0mTIxdkEc77PM
rQcjqGKLnsAA+WU85o/dlMZQs0SagOw8Q2k5IWMFNdlvNN1kbdO47jDYcUQMg83C
2A03RTMMQ0BJ3Dx/91GO7nY9yCQOpBoFKmTW7ANd83sxZQPDdgHtsyJy7Xkt+u0W
kaEAzgsUI6n8IZvZncAGHBZhKqgRF/QRZpXJflEUrQiiNUOcGB13dcM2ieNb6IYF
czdhvbmWxKtlH/InH+uP5UJ7t64y7c3nFtW1ZYCiAcRjh5B2PLmoJcNQ1A7M0JZX
G0ZJcN/44ZMG7HETBEAANdvmljyDXCUBCl8k8lHlfzvqdhv5Cwd/KKzO5bzrvHzZ
VpBiVk/GJTASB3Bf/LLYwrwujE4Uhzz6uTB12OiurdBs1mXbo5LKhbXAo6fCTtx+
STHkvdYwmo8lPVnynsvyCzicJjxUsELA4JIsjWvPEvqTtqTNw543aQiOEqZpv+n7
kLv+lSZ9ObdTEHjYnYD5N0CVFnhH8fklIx0oF5qiuiLbw9g2uJHsuFbz6IHvOUTx
xic6Ba6a+4GUu/qv5QdPhLzTbDHYhbbwe1wN4X7IRGU2Okp35jnlk+3VkhmkXCGl
nuMHQq1EvhvIIYhAVzyxH6mPDg0jkdSQOJFLtGntEbTCCTdUgRS1qhS7OosXmlnt
1Ls/8TQSF32Bc0+miqOts4kjJxlkRZuNV6REhYlCuRpy9kMl38GIxH8ZW6lfff1M
eFt7w06JYmVVez08SO56/aaC8NHpX04Tu9bMeSpuwltVdBzbUszRo5D0McbdPiP5
rLj78hw5sKCMwmONlSkfEles/A5xqfv2oB/0d9erb6Xe8F1x/9O7HOqyGUfWYWYr
wVRz0mg61GCnyzJFz0Ao+7SmgHZJhLb79BUZ6FdgzBGK+Gz3MDLmWa8QF+rqOhET
vLlyvoy8nJwu2r26y+PUws2wSb+XYNCWCmAT57lUKY0Q7GO6Xlx0uYfmC5VSC6Yi
uC1nn5yw6Mdj1ZOqYHv5DeIQmILB6aaSx7dLMf7tPjfFK73nfBxnvp2dW71CS9H7
d0UEnH9FeLV/CQ0eO+8vLRJPimVSppXxE5Lwb7l4bSdMzxLXfSLlw/hKOx4uMhWG
9U/ibXxBaiXAWaMu1bamDq4Abf956JUW+xXAOIbVNOdbksRKWmccWZVsj4SULAS8
laOzPn2WgpeLm9Wpe+m1dHwX1ZBRZHY0fI57uTinxzUSN5MD2lqx1FI8vFXmWyqk
YUfIarZyWGK+7h5bfFt43nu5ZHaW2bzW3GsjgXaxEhYE8AcTtQVJfTGhoXnehk0F
HvxtEM0gaQtLJZc1+4UFRuacFYX95S3rBqsumn0SPOkl+hlMdKSk5Kp+xNwKnjS6
+YCU2gmiRYFsGYIaAlGRV0zwasHqqwtN86JhELToOjQ76db4IjcQI1hPDfSoxm5R
CVZSUScbYdsdcj9v82M70eyJkygCs/EenIwvo4wBpwJhSZpX8EbkDugJEx9w6bHD
rQn0ReCTrO2NZP+6FojNWpxjHIballoqc+DaaFmiD//zlUYblG1aVurUKpE2eBxS
89U4OMwubKoVlckOMAeFjkthQR4eiQ5Gz9gSIixaExa2AMQFTfBBMERR8YKSxnum
qYHSr9s4YuFWikC8+CpYrf2xdQBIneSdEW6LM9qqqe+2zWvS77Saa2m/tQN1E1eT
qGkYxX0/eedRz8EqcGA60PrI7N9g4DD64swFQkq6DddgIMvl9K5mWr/P5uyiJFNS
8sO9j70t+fq6rWa5hOaPbS3iY3qkrZA3C/VtQ5RqmSU7BKGkcwVhQ84zvsKfhdq2
7xCxWX4F+1xCQc+9TMYzG5Wx0oJOYwYOLW4JLG0BlCbTE+P2wkq/gI14DEgt22Ws
sNL/5eH+vQo6kQdbHUgy4c/iq9mbJfKI6LwmB0gJILjxaZhDm3TLL+GFvT49Nmg+
Xx89Xsnh0sOlLnKpgvtts3zOW7dkmlC9DFanwTY1v0xtNMB8zMheghgKScz+05x+
L5+tLnGiLn2Cr0D7+hNNBmtV6lN9DHgjLEna7eHw8krXY1OM0wcyI7YCOVjP/WE+
ynZhCamz/XTFfFoDif1KbPgEZTS7+UOPFMQyUbq+DQi55uJcnGuRULPDTDPSg8/L
8SuNh0Oskq882/vF2kYRBFyuOpJhqOlm9lNOYRbvQnBCQDOCP+4h2Id0Pm3OPeFH
8UOlqshPekD1Uvj6yCoAy+1SfVBCjPwBIaeQBf91W3erpDj2OeJ79Rn6W4aoOEgz
cu/q6WYmBaxIxjqrSKMDXqSb1Upx6wGDSfSfuDmjj1DZTEBAy8WgvQmxPiKfpqt1
4E156XMda/3CpLhiXjGKwKL2+0rGLPaExIahqVOO730BjfiFtDPhM2LYz7IUBHDM
lhQJU/pfd+4yZmIyOjgUzhizngr/KNMSLmkrRUfkIZE3Ha96Vvb94TkX3FHip9ER
Zu0hOqWsMTVkuFzmYlh7ZfWWHNb7GHatkpd5+CmOAy1YuvcN9IXZV3JaF4/oXAcz
Kw6bdF0a8Uw2o5wXG1c29XoYwEQ9/7wJKpzPPkIOnFjG4lt3vpVX2wGlgxnz9G0d
8Bg95booS0SpHBvDK3LTCsDZlZmgjZWLy9ZHmhknb2QEnj+iFI19p5lTuFgy5mHH
ifHTovufyU6sMLvAilGe6o/PWZhlcVKw3UZK3LT2ewkTZOHCfS04vegZ9xd1geLr
4vZCkhBdBMiop1qil9X9cFi5rY4NtXlOwvNjm6RO6MTY70pjHP5AIlOzMWrmtgMs
+05h5vqxnCTRdzIIwDSgoSDDUL5syMkoYRVgW1avvpl5J+moI6YhB9Fs1uRGUMMg
GDxbCzCfFXUf5Tj+M69rFl3ULrPg2kuSPCiYS96GDRmVAK7ZmKFFHgEPs+BIW4Gx
U6OQCJvVdxjfCSGplCow9NcN0iRMne4xGg+9oGD847QoYghNf3BvYPWS9fEvAfBp
Tfg9hM4WmcN7mLIKp2I/UFaatWAb9wWkSsYqTlrtCUyLtOUXrMM6adK629Ac/NPo
/wKFHWmIDCRMiWJaLSOfaDzGivn8dSXBoPg0oE5OSYnQbkbv1jYT+fJieWFLfxhc
mAQcxrJhSY3agwUKbqLTC+/lZFZVNELbN2Zv8wlJep4KV0BZYI5d9+2dI2LeE/ct
JU8YSx/MnpqNIhgmAQN5KS1aeOdi9vQ08HSZTQ2jfvAZfZcfhtcGCeudPza/ynhf
W6xMyFZ7W5rvNKQ/ZeRuc2TvFs3vAd5AgnwysMhOZtu3BqxjonozmGylXo9DVlWP
KaRHoplc+n7Sd0zgobQpnhjqbPE6roY+foWq8C0Y6PFLabpXBtPedN3Z0wnEyvlQ
FsFnHLFFAxykeNGp5fiTpVZPMQ9WegdjU5itpc/sYuLpdhmtbfwD0cpNbXOBlpJx
7BuhctK1ei3/5e/wwfvRNyZPYIXvHEsAVU9tAnxViGJXnDagix9eTrQ/yQQb2SXj
JWPkjnAQrZMHhMg7LhBfW7cu2kX58CU1MN0Hn7hGWsddcm2w3Fueb/PGFlXSDIfV
MaujC8v0kBhD4LVd2036hm0oqXJ54uurGLKVNFyrsspi6AcbY97sxc/tak9dnQfO
CYV7Qv/usVORaW7lKkJGXlNixPrDAWNgG70gjI5umSmtF66GqOAQPEiNh5KnxoW8
bgzXc5P0AioXwnmvLMFx+1Zcgz8+G4PYB8VfqJd2avaq2eMeyhXDFhk1x3kS1SoZ
3m9fCqxXHW8Hphk7ItrW+jw3/6e+vhOKYkLH5o+8MvZCpAQfJgQJaSW4syO/24kP
LR5lUYYGZonDFZrL1+sh5KxjX4nPB4mwDp4RGJRqf4YhKr2R+zet9ObV8XM0CZkO
VH+5WY49V4s7w/zg05NN4GtqHa+ZsmeJ6gBdL4/jz3mMhPTSff43n0w23SzH5ue4
Iu5bB+biOwIlCKvNmgLVx0u8Gqki22Vpxxr2yxgjHBCd6Xq2T+gPcfxKX5NhnpU6
CpWSYk/6OJ5SXPNCOny1kJ2U5nN0PYPj1L7jQVUmzdNPJFoK7bPx9WLLx3V9qe5i
VkXCGcBoREMTl08de967L9K01VXvKA5Gg055TkEzhuvsSSsZChq7iB3MNNw/7Gki
Q6mjuEJN2ZLBgJZ7HyL5yTFcl55XKKvLfABpt5YawOb/Zd2LAYZFOjyIlCv1QZeS
uSyI9LSKgHTCDj/gYLIbfuukC4/w9EcY+gv49UnfH28INjZkjdXoXylMYfxgO5VX
kcTnkke4HXkeWpr6TG1u964wK2cqnMczdtcWcfWnEYzct7GKQwLjxy9GYNk3Vlzb
d3DwzcoffmWUzxCqn0xDzFkjXSfaFliVvjEm7z8bqcdFUFS6y+4DVTgq/P4WRabK
dAAJELP2Y7vdzf26aBY+lGG2cAfZ+qn8vLsrpkAI+4bdAVXTtdY5lHDmyTtRBiHv
1Lqv4dh6P3FEg1p+FqyuN8buajaDtJHAGZv7o9S+EvbrkfK9O80XbE6683Y9dET2
PqlVMI4Pu5n2A8rYJwBIgGTJyjNpkXsPycnnvd7A92Y4jjUVTZmc9soEjMG+LR/n
DK1qTEdoRaNY3vxix2O7LJhPad8fodKZ9ZmaUGYobQKG4Xm3tQyNrFXVeCtIdkOm
6qLzZXEl9uCkgiuQKqN+D0VKeKd4S3aAepcYRTveQJa8ORq3zVkS2Dkgz90reJqS
ZxsrbbkNVaIHdUBRi+rEKLbhmLfSw929fWNi/wIVMNVryUEDnJFEhtEnWy7y4u5d
DkAV/yvtE3eoDR/n0c0wNXenzNMojKk4rqS/QCCTKCdDfczaP+yCb1Q1DiYmkq2K
sOJcCD14x9W+T34Wwy/9/TENXfKL3bX7oadpHseAJ6/AggmRPCzrfgkERtBDy46d
CW5kidosJuYZ/2GgHQxkXZ/65XPd0TZr5AmQjWzWJ+bgegfcscsr/WgoPXHBcC8U
1vpctGTYYhlub5v46Gv7EMbqlDugHuYWkFHtZcLKLJ7P8myYGer1nMPwfgohcWEv
m1m2Ln0z32aUlWI8A6qc+P2NBM15Th8QxB+0Noh5lceCvNtUWGrvAGw8ORRHA32o
5U2jZUyY8qRLueHanyHz7J33VUz8kypKMn3UKP7C25ABpMppwk40dPoKvPDz7bIV
AJxR9rjkEosdKQkhdNvrUilBJMskmn+DfcvLvUANkIkWgdrdTyITT2HMTE64GIML
z0CQF23WjSlfvFowU4i4kzcn+EYM9GDy4BCc69a40FsWVSGCTo0Nb0zDghC+Xkba
xN26JaovC9j/bI6TD4/beLAzVHyjGtG5UvhuXXhWZL8rvBUdS+AHf3pyIGJ+9QYc
pMJ9A06qhFLbE7Ge52yg61ulAJN0mRfXwka/8REp0tS9z4qnMaappyQuSrPXoPw3
LB2eOEIiC1lXvDK3vWtBX+iTFDhOFfH2yDXMOW4iBZ54ggkywwWBQNj7hiJIm3h9
sbAWWtiR/Ls2RcVHZ7v5a8rHqSkdIE9fBeivtOCM7EPDN3oeF30nF/oFnB1EKjKb
UWqNF+N2MQL/Y9PuZXl/Ywxunao/5AwpCS1ScGxJwCwqs1zpv6PEggclv5uHghTd
m/5fTAVg/jsxDgElWBMHUV8MH8L4dRqrlM9VPTDLS3oGYzQxvCPOH/xF9S4CXnWv
o1Ux7IhqMe74gf9TvLQVMCqbJJnvtTbNjt6O8ZiTwcbncg0OQBoJw5OotBF1Si8l
1cfYnVheyVtkYkA+gDQLfgSPH6gapB9ubSvQT6RkLKZwz98uDneML0lxbaqc5+qw
4YtKcd2i2EvWUBTaD+xob2QD/lbFqt7a9K/5djZzwIfLnsh+UHQLWGWcEi7ljRiR
/N+L1B8DJzn1ZoTKci/6QhQzXvnJqhZ8g45vgA/0/kFwy/leG7t2OJf0r4QWignC
0bG4BZTzbGWFVJcLCCyHj8sSWuSwXvMAEZTO1YL64nUdzfodxfvryt701fU+a97x
w3Jy+WnMJX7CjGfadK4/rWFyLWOa6omWdOYz8uplMnLbnYT+WRXuFSthSpPC3MPy
mFcr/TXV5s2JOFQLnZTj/8NtHd8m29VBAgpQ01NThbb5VMGBJ7/Wj8acN1tUyaKx
QJJ3l6R4262YiNU7UuCd6VhHfaRXFNUapefwEc8W0to7PSfOl+dbDTu65mkGSPwo
aPzq7U0geSSGevFvwcYmSKNIif38B7tfGEkYRU6ap3oPxNzhrAvX2CLesr+q+i0x
kbsUZjCR8WXXlBoiIXcRe84KG+1AWfQMyBLjuJYmPjWGlswAv8VB6jdAAQiHM74G
/G1gjxH2MrOk9KPvevj6slDX/fwSre0CayVwGZgxsm/3lBKjEFOEf5diCaaKWnhI
pdrP7v1xaGJ6WOLPHwOvWxtTO+gwnprcwsuRQQqHe4IZyCv8hXFo6MQiAkqdW6Me
k9zy64J6svpF8acXTD8kUelvN9Iq0tfSUQGLGaxr6JRs3QiXPzJso17lNu3jjCN8
2adN/sAq98XEQqQTBsghvCCj/xkPWDYoa5l1GpUgQ0bz15qlseRnHP+8T9u6UXfc
uto5c8106XKUbklMAnTOa/XRIcuIIT7mMEkxqbAkpj7OOTBVRyAFNYJoNC4ei3Uo
YiaqOgkm55PoBRGtRCqOxDpX2AseqTJV9tW+nkCOsHfr3avzstuKFV8HqtDr372R
PZHmo84gQs6j9VuY8yQ9vLJzHZQVpT3r17WBBhJQvctC/t3mxozfTIVw+1T4OsyL
iTpT/1+vk3xebw2zsIcb+ebs/JDKkE6IU6sOQpS2IyeSTlYsjHxTK1k6p+mMFvvT
/wkzkUyIPsPy3+PgwYtUmh+0Tkg4hJaGiUgnGjBdHboPY2uiJIEzeju6QskkDVkO
oBpblLaG/iIQWNk002Bq3zOv6SRljZmKPUHqsiYMrO5jYrV/yssjSAjdS9jDBbAg
2+ljjg2ccZZ5abWshDhkydtrlLXO85ZvxfaK3gE7+nLDSzQa5leWmkLdbBmr6lAx
xRgawLdq53/ZJttr1i80rzBk6lV9PW8EKT759oxL3yObPw9Pr11R8GqGSn8hKMS/
9ZTpeV8LUcDhXlwyAPugzvPeaF1qNs0WuNioUeHbeOwI2wwNth9WLs52rIw04FlP
PORpVmuig7qftmB3jbscxSzm5aUs6FphDXPB3/acik7irVwD7a7Ha+ApfB8qRNKt
LtD4guGYnbJ8VyIuGFAiydVtZZicmCVHSxAsdaj+XlyVQ/QRpekt1euMPhpQRI+c
qGMlQC34A80DTN8f9Oil7uJKi5nzNf6WEGG7qV5hCrO7X4L5gzcTCJIKdDPUI68l
y0E2+vSmn3qu7klh2tovqwt6+bXJ5OciTkzbGAgF1sXFbw7ZRXjEDiAkJRyis3PP
tmgSecogjRZ2qUQ0aFRjfmuxfp9ljct8o0H+UzYQG3Ljtjlb2z7XHkg2XvBLzSbm
qElAlAYT9w+kibheYJ9FHzUr7Rwg8qdO/Ht0w354NzA8PMqePm+FszWkH3n2kt0N
yrZfbT4WPBohB2fzszBOMJQ627moq5z7BIPu92Dx1yjhpxKhMNyAvor64YbExc7n
VLU5Z/cdSQbxjTCDPFV3HAQG2FL/LYnKBK7KKQd0tGNBFuBcInak7CZOpGVKXBRb
hV6I8kIBYMETp4lDTZ8nFoFOti/MyxlXIXGKNXzJSFHg88H1wVvLdMGyCzbfs1jv
S98ly6j6nP0wZ3e8/gJdLIewS8EvFozLslK5Vxayytu7rP4aPIz7Zhd4M+hkZRTq
I2Gt8UnmcxPXG4IPSbhoNHv92I8Sz4Ndp6sKMAuaglACGxdyxoXHl1jksXOY9uSG
pTssSO608jCJcXvaTxujQ00duxsP+e5Qoq7IfEDoVlpblfs2O4RPzQ0MACHp34rs
jlYr+X+K0IOdR/ZiIraxlDTYSp02lEPRmWnAyVGbRgdIcFYAtfx0iy8FkWJQFuIY
NDTOLN+YqJwaum0/cYhjFoSmEUXNO8UnbcmhEe30yMpxZGa8kBZZ1Fo2vB+WB59y
k4TinjiGfwTDaHh0o97sLp3ibTNYIPUakM4b1bGYxqvbmuchQ3aNlGZLjsLS2Hho
vWYbEsZ1uDQfktnotjKsGFop35XuBnG3oG5J5mHH0Jm0x097ofdnjxHZvir5vJY4
IJDL3xG9TiUqzag326YiVYhoMrZnqQSFZgdeJHopQcWaVSStnE/dPmmmQSHksMkS
42RVIoHvVTjok65YuOycB9QClVcIwpNzQ5FwGX4hP4qFK/jijbFw35Jd0ySbQsXs
4sZXi0g38RmrhJikWtdZYKgGLI6hbwezjzowAvlra2AJQGGD+kBsRIoSQz7W32PE
zmDmpjZW5tOEGRHpZAxGxsf1vPSUVP6E9iyyHPq6ZFG0/qGlEMU3hzPkILq9ewW7
mv2MkqI6efe24t8PtjWnD2KeTdCFRjj2b3GL3U93dolBp33uAGN8y2bjyYlhMlEM
H5mOPbDZayiuBJNINhU/Rot4MHfMEMymbRIzuL/2A6kUnH4Sk9Mufn1xX0J80sQh
B01vMNRX7e5hcGjgB9g7pN0iSAhojSB7qPQShjDGogphDM194nR45Qt6K37Qtll2
rO3/Ry4I+ZtUvmmimya/L9p23CTAOIvQmR9/v72slzAJa5c6x9BcdanisCS1wmHJ
IKr5iBXFUyndhaFr0r7cDD+M8/tCNvxec0glJVjrD2ryUGjlEE+e121Np8OXqBRz
QlW6vXuXQ1Pnw4l4ik8KJEV2/HaGMgqr9ChlQ8Iqa95Dxnm0Jf40bnvF59XABvga
YtobmgjODge6bX8pmXDEu5+TCHpHumfYY73zDUKj/3qpdS37MEKW0F+uMzIqXjiq
RM+5NPkpdItqr7TFE5J3JUHdBSSI5o1CbWab1FAU1FumhAozxYoRt9mUD071HlDb
mPM9F+XtcoVl8l3UAPPYDmRJbKkkFKtbg8f3QeY14pUOd3yWGM20SlrKEsNboxPF
gujcChiEvFsg9XE6gqMFwYzaVLJZTk/FSIGRKl4kYBLUwspVCU8TnhjNrFnd7hjq
KPBBQB/S1mL6167KP1SqasY5qSZYSctkvg6Ew6IGB+255JbOVb1jwBq8srEBrPq+
+5hxDpC5qLmGc3NgZXSy/eL2VfaxAPHJe1bkokvXfKRhcSKcjNfyB1iJeekCQX+t
ouYf/DeQKEGzIpv/nETZ96EVu9g44eoqRI0i24h619UMwuX/Iq7p9jRGr3hcPuRV
MlUT1sgmLLBr2ORYV2gBEYylRqsiHk3PW+JMtn+HZXA3+9W5pA1wLabjaawaJSt7
UIYoTuxHGDDb6NAGduM8hY2nm1kMrToNI20KqOYlL3Tc2iav5SGdwtGrPneMJn6u
oR9qI1/AkC3gSMz/Wx3er5uHb4s4Oe+IIPRzyec0szp+Oqe2iGctqQ+O0g9a3pje
wPFSB/UtCcaoZEh2ta7ZuaksgY1xtFyiabzxSKfy816tgBJZRnWbL2qrLslzzY5S
HtU5Npd1ADisui4nMuBnZiBN06T/WgxbeqCeDi44HppbFO+DZZnoCAmOuktOXwR3
1PF8E3LBCjuRUqPFT9+VLdjNh2xfLXoAC4sUtPU3mZcKurgGcaYz+VxfZucMbCPf
BQvTun/SsWKZjasYQywZtKi69E/ThyZR44WazUXyQ2RzyCqaOtWzFn2J4Zl9+1IP
B8kMKxI8GlMy9lws8Wlvy+RpUvBfuV73ISX42zyili1SmcMGf06rl+ZjijPtcGr7
FPL1D0sgXmL/pvlyQVxhBxW/JUX73xH3L8d1pJf74e2riHnzYR2urjuMmM7kFPIu
u8B3/BTur9N1s2Z2+ZOoJTUYcdE1rWdRlQUiVsq9yIZdSs8MWv3Vj05J5lGfiygz
rScVnLTJz/zroWPDrwYljY6NqiuMlDXw+OkiuKXE3kAu2wbwh8U53jREhhCUnQci
RJSyC0i5cmjM7PKbJuKyD6ThuLVHf4DvKFKPiz15bXoGaZvzGIz67XQiXuzVK4aF
6G3MMcvGS43HVlHHN1+Z3QlyIql0ptGHfYtiixUNmz3/B7PqgcmriaJmIln/S0WU
+AhpVx+eefPnAqIV+pypjGxLqlGNG1Jx+cm8Sw91b/ebzGnPDsuE2mivGpUmjCwe
32mFvGfZ3Lh3msWbpvjjLIvn44U6zFMghTEFSf0NE8Td0eo+E9yBv9bjii8YX/Ae
zx9vGM2IKPMPiQWaO0JJPZfRHICryFTnGJ4KcpWgUED52oOg4MENr1H4S0bn379Q
zvO6ysbm6UNkYxdREHwHPy4LnsKwwBwSG3b1AfH4aiItmE/RaBIdv5yl4cXIWBEa
wsTkYOL7K/aFVhJT77F4n3p1LCblflkP+3cx8lG3b9Lt+DT050KU4iD9OIIlxVUL
49KTQ48kIX5Mv9khzkxP0N3uRHz+lFSYAbga7VxX4AFr2zTNqUrMTzUbTvd7HMyz
78AOY5k9PH96Um6VwQFd9N/jPTR3/hqjo4cHTXO0ct+LdRe5cZCTFdY/fgWygPoJ
Cs5j+/X7b0wgyzhcQHhVXnURh5L68mtJZn1iK4X/B3PATnasg1jWXFonUrmanV2p
OHUYAqbbpNyx6TGvy/AOTRRVLWSNsp18E3EZwASLEwzaxVKzgQ7rtbQ83V8kzQ1k
g6GHwKTq9s2+gQjhcdLlX2SoKgHKkWp9m5s9XmJije177Kive8olM+KgqeUYqZCU
d+NgtA/0ow54qgQfXixGl7a5mgJt7FG2jW+m9TV5gC+jRhvy/8fQKnvDFwF9M6mV
n29UVwXTHmE9I9hdWxLtU9QADg+1dHGRu0odFAN8SlTxhytLjmffdFwBQBEaxDzP
MN0056Q9K3/V09Qa6A/HtSGd5bSlo9gAAXb+MIEk1Miz4RxLhwPH0wAJkWWODOpY
HisN7nj9xdiwaEEEBtydvIuXpDPxZ+Osn6Tb8dhH292kAJfooFtXU7a9j9/zMeFa
NbmYwSdTiunbB4pOeVK+xg38ovgtpHo1bPJ0Vdt5sNe+B8sw8NCnnBRPBduH4tI9
YIXizeUjQ3Ac2XSmrGFMUajllwPREpl2bQKYtMOaVw9OyMYgQWxr05S9mACiNRUD
2D4caQvS7TMQsqZYxwumOrlsW3O75afMra5CLmG8roJO1ywL6cRNBwzZ0B7+At2Z
h1LvnyoOptIU47/oZhkrNrZcIYkt7m3QsQw3ckg655dhnF7wuaaNmCsf8ElaFVrP
C8teMlOIKE1RCO7vGN8denva+SmfQnnNJXfjQzOlVznMuUosRsHG3/QO2NJxrW+7
c5CxOTQ5wBAw1cSlplLogpDQTYYEMnOFkxK4QAK2HOAGCL44J8SMl8IBnhpwObG4
3ePweAi4Yv1T73nvw9coxkMxrqtRLnhVDTmPYfUqbkfKtPRS2A9/S2Gdq6ER2hhD
4Krtzx31TglbbLwDaaJzdImwuaBeZomR50jTAVKr7KigeFbpuZjTED9noET91uEN
s137aHqscDJdedz3gG6UuAEQOuzUVHKsH2cri0CBqq7c1z64v/7xSSgXPLBJuGHF
iXIFY+KoHVi9FcKFfvfmxip9GrMJUBj5UqQV7L+lnMR9fwPkpm7vDgIDZGVIiAhg
vU4UXnZdsEAqGm57wKMtFjP7ZwXD0sAeOSnomvc5aTaXtmbmmn49v1IEIDqEydC3
Bu1Afpqyc3ooOxFCXYEIN9ZNgVBGXi0ipS8k1o7i2odO88UYNZChTlMAWlJc3uSD
LblPO1t0A8M42YsV7ninq7fwr3qTwQelrPE3b2sXwbaZqhfK/E35w2s6VirT5cHc
wNMUfe9moW8aoYWNBVZR+XMbx9Q6QD99oomlkw3Yskp4XsPesiFXZrSgv6exeOpf
4fzPsGE8HnWmumUZ3gGjLyOPZBzN9Gsr4A2Mc2YjU4Lh+h2FXt2XmnLWnzNTJFn7
w/h4biT0rPhkiJ0O/YPRL45QfC2p+FTOmKAy5Yr+Zi1GKpA0sjeKhENRQgb3Hu14
7B7ehIL0Ei5IUXcwibEFBS7lXiBXu+qSpAlyOBOlr+aR/mh/0iPaXjXQl1H074K7
faHWO5xTFG1+H2TmsQ15deC6uB6CN6jHC2kOV54/yLcpdYmWuFUkwtFw9URA+idi
CeB9vO6/H3t7h8aYu6rUJOgwLSZyts1EnDRRvb7lNKuN0eDHczn9HuJ9tqLbpLSC
/4qa/+whrfKuk+B9FfRIgwYAjLDnPLFi3YSmIHX3cPXuIrg6d4Sf3NvDxPTmUhd4
0s/QgwOul3LEJsP4P9PLM6HuO9BrlTWY2nBFc6oCQUTc9dZ/qWZkm2Pziporkko4
P2j1Nf8nue/XAhwxi3ZiJQrUOmeVWDdxcLhYhUNQmVMUPKmyyjw95AwqtC1UQi4C
Ipckbd4GUYPyI40qHFGl+cAqwkPtsl+Gdvk6VjY/2PqU1bpS8/xfnqB5W6DhPJZr
TnGXhByVqAfglbyAo4R7eMHa9TReMiBuwFrQ7LUvnMgFnZ4kH4sCbaVQxzclYd5K
pVNPPoGu0Wp1ycU/SrDSbwgnNJ16TnGh3BmJPUZUy4ZUN5Z9lQdE+eNkNOwU922g
LOSzbFLePZBwQS9364C9fInQyZEhNfs7VEEA/G2/uJzrqhslnBtI3ZWaihfChLzU
5nuMjIVS5NfbgDsA8lW4VAKacpnam9R4dlKGfej7R4UIffuR3XIPkAJaKBIACIfe
94RmHvVZnakKiwypxDQMUHRzzLAW12ck/JXrwHEFosgNulGwNjKb5OH9bzHZRC4R
RSv4e3Pm7jr37K+9gqPMVDlU8YMkL3ypaGwo6GOJUmxABv3tojsGcRnS7DHNq/Kt
BUwUr4gC+JEElw1VNxTOZzRNnmKBTcmmzvicNLkubazihR17dD9yhG6n8xypL8FD
O0jmhgpn8N7ZbFTmrsJgfnGpKcHyHu1bGpUbdpB1hEMbwZuglZk1MRQ451rl+pL2
KdTIKxtB6vNL6vKn9HSeb4EWq/uMLdC0iUlmR2gnJEsgYJ+EIOcLdNqzkI5c+1cO
uach78kF90uOixFQG0rGGpWxGJCl4sk1FWRi7MmHFD4vbe84BDqP8/7Khh5x9q9V
KfzBrHAGvHHdwGj1sjPGyayGstJ2HFHNrBrwRwdOzYvvzcG4s5rkiWFqnIFXK84Q
fjLu85s9LWod23pgdKdI15t+MbdYnzdPbRu8wQwqyMTsMkXF4xwHDkhYbQ4rOkL3
Fk9UVhxA/88kftb0qhnBQeJYFDrFJvQLEG6Nx+tOW7wYMt/kasBWF7u+xupEDdBp
1mfs0bpTv5XFJTPrTu5MFrswlC6lGqEQJ49R7kNk84X+Qg+b7G4s80aYbZ6a2fsP
nhLp3CxvYCqmRi58Tuxnne38jxWM0ieGyZUqz7ULgf3vV5QJkqKxgxllRw+XSiLe
MpsC5ddKlQqsbFnJWbP/vxhb0rO1gew6+CXfzE5WUrrUacEktICDQBpMQ6HDltBM
4SiBQdf/tNliRu8p/aGVAuYjdgZViDwFfWRfr8X25j4IBBtWau0ZQva6G+hoxI+H
umZNvoyy4VLjr/2G+fVJut4YoqOVfdvH/9RLYg58Ubnd9ICWYbEapRjhDPCQ/0E2
T7yzofTGHrLzf9oJU9zO8uG2efIqFHPqaoG73M1a6KI3jpWTC6TnFeywFpv8HUK6
I3lQiYYaIsvsLmLvoXm8YVNe2Cy8zcZydkrDZxiVl0V7ZnpNBLM4oB0ksNQ1VE9x
UtYrw/2azbjStjPFFZnsVkZfVGFIIWKZK/Vmo4cl45UeAGDWWSoYZlarb6yH7MYq
a8QPKCy0m3qwmZCTHdP0ky9HRtMFXsnRIPfJA3S90eHGA5WvJYWtgCykttaQd8Wd
0u3dKKM49JoR45+bPp/SrLQN/OTtmx5rk6jtGRR0/KfJshyB+vdChRSeY2n8CRjk
Kr2oV3upOrOPDSdanxnutM2e7gdWaxYDjaPiAB4UIS21MMzNgeWpMo7oemZig7MF
s+N81vUBS52o/jSNNCZrjeMGUE/M9P5C0w+LILqDwLF4iO/qpCsivcFhGXv6amd/
9MrDY2d5z7aGjm7NEYCC8EVrkaJ0U0rEDvwMMjWVF8ZPG0Yerh+PvOUEDFToU5RA
6WSCjXZcmeBA78Ef6y2Qb2nuZv+boIPcb1HbV077g0yiU971Xlp3HCINidA+QgSe
cNuLRaoZJp7AxsBaduJ0Mo/S4lt1KGkEGTKBM+zKutWCqo8ZL06uFAOytb6F38Lu
suZZ1r8CtIE8incUa6tqI8RO+iAaZqs1b2yLRK1NEHJbHuHFnX11Q9usaur5rAp7
1vsIyf4I3rXf9AzEVIHEtnVP/V31QyLI4TvwtkAA8Y310n6v/ma7HXegWfig7dPv
E2pduXwgXqRlRtFeB2XgSXmYjp7wxvBl/O+1CWRAnXS4nG64s2t37bh1oor7VBwK
PVzkqpf7epE/dmg3R9hRM9caCyXYjN1QZimIO4IuKeE51WbbF73Yx5CG6DcHNfFa
3wNP+fFlS/gXnaF0kVY4bC3wfLWed0f4h09G7YeBSUlr/27sZwzV/4F7oWReeRNZ
303VegV3UoCytbMwXdDGrE57MSCci3BqnY8YqU6SpXHNU+wEnOHrZ0rudT02xIlV
XdqkB9kdYR91NTQ+DcfkmKngv66BbNEhBRPHytLrfJfGRN1mNnBFUPL6QsiS7v9N
7pVS7XCbKqsYoKnXY3adGDSpOy3WAq+vnfsBoZV1wl06rNswocWBPKHL6/1m64ht
zxA2MFhdF2s+T08ogQ8SutprL5ivE4Lvbi82G/QiSNrdoGIO9jYw4jokvmw0GAj2
eKi3UaZnw0nOhdzLZ9+CV9cqV6oQ1pFpi1KEmK3m9ZSCuvhH5n5ah9HSwjxN/DZj
OsBWU+dtiyRxvCGxy3QbPAQ8VGq/P5dRWlq+Sima5l49D9pXPAf1/3B14BRIvpg1
dRg18rO0v5p/uO1BVT8Mj9yXz0JPstJFJEd85v0frcmuyPClIlr0uN7qo0D0v4Xz
VoyGwuocZbopaKv4AZx0zho2gfaagHy+dfFjEp+dQz4N/udHyboK+GN/V93hJQx2
ZhIDOAR+kX177xg3FE7stoFp+3nqg9SLw3p2j7CAzDFD6vHRTprsEiaK7y9HE0Xt
dySTKK9iV8vgFVr1Vol6kY3cCrtiPc2I8r9XAMp+/O4jlP2mfPrfaz2bNPFwdmXE
OrnYCOj/qGrVl20aj5iUj7TadEvOwS62GhaTtPIhQ5UG5FcHahRo5dhf3egTgQgm
sb200Y2fn+WFpTGL8oJY4UcqiBessbE/jl4fcqzTuRj4OqAD+fmXykpR4kt8234G
yZ5RpF5MgvUooE9YR9iKU90fh+fw1X/lJrGjXb0MBccW+WXhthMhefGkl2QB4ume
/MhFytTTJ/reA+d42MZt2/FnrzhHskb8pDJr/QDv4C2EJMRj2QBfXzVtCqqLGcD+
65SUynuyNNiIAgOA/DRPlAkB7IUVTJWjFU2Pvcx4eKhuKamwBrrkkdVllwPIcbBk
c5+7tbGHOpaM/3aDraXNDqfZ+NG0QmLqDZ7iCztcdIguBsv7jqhYhQdeOWvE7vbF
ZECvx/U/A0g0g03Ttt6A1yGxr33dXBYghcubVik8ejCDnpYhVz000HqeaQkLIpBd
9DWJaKuKHuUisF3SEzWI+gKVqTB4ZOL2Kq9FU1Lrqwfw+TN9JLZ1EcVhWgMJwc1H
yIynnxJjeiT9CJsiIpCbEPtBMuDr3noq71oeO9rKvcsJMVX/ZqwmLQls7Q+AHbOq
PRVDmCcryfdq+/T9KwehgOruJ1+Rs+DtI5qKjO6s8meBnjCPuSK6AZ1nOyYW5rBG
YqQ/y9vplFBVhurasAehz+BBxOrvax3S9/k5vNRBx2q6yRIuGL6xnhU54rLRoyJR
IiJaP9jnc2B1DzMqZskByjrpkYcnP3tBvCPWN4otfXD9tXKIv9pUcruM8c9Lw9bE
Ef4N7URDmCdQCwanz9E/03SSYPMjoauFSjxvkWFCBw/QfWpIQJibjd8aniI7urcr
wNEi0db+MrHNDyuaz6I0Dh8DCZax5PcMZ3XzD8zj30tLVqxG174hXnacah9QNMHE
OGrfwdEXrR/3yo63/nYkfzgPgcaVAKKsgLo9kGMjxrQ/1MAfUUGXc6+w0tCs+EPt
wTcNoZxyraBZxWe8j4yhJuzsxFpsEsJvBDcd65s/cEkSwkS02z3f71w+Cz3wqO7b
FCIjHK9lgM8Garh079Z6102zGgoYWr/y69b5PethvK5WP6SkGufSlT8+vkeQF1nq
gyBhyrFZZBPFcBwjGZB9SrBL9MJ37B1QSO14kT2lAc2Hk6FNRw4BqM9G47AIpurv
0JAzD1+hNIE9SfojWAxWkVYA9iXwt7Jo97WDTP2Yt3K9vhhMXRJraDeoUYaNyOFy
ICvO60GDK21+aCYor0RESKb1oKJE/2Nrt7NzjKztPxbOXwpNYAprZ/dI+bXiTyED
0nQeBO6+j3aYdCCi4M+9aU/qQHMZd/9+gWLXm5S7KUq8RmYDXKIh6oU3QiKmsdD/
NubK2BAuAJiFLqb8KTsUQTSQ8g98a3ajfGaiBldDWSplInwi7/pBVzgJ92/q6hlJ
p7ej3TAwVGQMg7zwxhk1jyQmlDnIbmaPiywG68FRSAwjUJHlgMvYckYcF3EoktMX
PJd6UbcIq8ZVjRBUXB5HjqxyA+IkwNuLUimMT57XZZbsvcqP5z7heLMlqX/FdfLE
EHdZdn2FQQG73d0413VxPhYPX15msBCPaDBQV1lJNqbL7EmPrkM++s9Lb8gOG50U
BP+Vi86FF++xwscTglwNjuTJScS+pnu97Z5VTaTPri9D9CkofL9MM0drUqOlHcrO
h79AiRQxsc8lw7HDEXuDz4CxEaqA6izEuYYnD9jnEu8xAO6jbBLj+O6ZQrQpujk1
vKmGSvANLXVymYkHPWsRz5FMn8N2RFCSoUPFYnCxAUThWj2HNquiD0lrPkZeV/s0
5Y/6oKR/4zfU2PfDD6/T0j3TPGr4H7MAIWc3VD6k+tqauRIfnSV1qCGWrXVlmIz7
uQdbW2CZqvTxoB75shfRF7KgXeH/+/h0zDBKIOCTn/KuG0NYqdIoySzBYf+FapoS
BvZE1oTxwVmfGXbU8oC38/DCxEEWSp4r7yOFLSMftwsGs2GcG99ozmvQ8s4g2rdy
X0NT7zVbvlFpSgX3aDOPhCRjeQyACH1ELyctvn+j0O390wGomUKiTdyIaIwXrE8z
X5vgIrLDGbA7EhF7a/y2WyjZhKl8aIAq8zIGP+2jIQFYdLkeQO8xvzqL36meeFgC
+5JzoeS/QFsfIFQ3up25W6tpAru9VVRlN7ziAxpJFNoyv1NB9rEec1Ib/81+JoEt
LqeAnnii53lj4bTjbUQJul0PDq5+Ykpsc8v3+ZOJVu99pJKfhIfoBQud3X+CoLL7
yO+FAPv06lH+mmlFhtJLWGzdfQH/Sd5Qd8aC6Gd/htEVsB1cyHjOoLfdTF7rAWLN
ewOE8T2KvmiytiG4R8RTLOVqBbSugkQBVUcXRV9YIK/hPX8Kz7tvICXpP8M54qMn
aNEy5E1xFaPCEi8ZjXBFkh/pTsumI+xnTqORIxOk0WkGs4pvHGaWNoc62GwXtrvs
Kzf0+Bn6V8EM2wXSaJTOOnhdDPfRDJKnf7kb27uwHEvwl5aHQ0Pv/KlDmNBQ0/ln
kgPCAUVFCo7/wNGzCcK+BlWKZixW5ekklX381Sd1eq5Fo2rnOSqj5R4r8pGl7/F9
Re9g1IsZv9BfPS2HHuNakgMP/Z785uii2NVHg3GK2hrk2UoL2u9tdMSsLs8TOQWK
g9/y/ki2egXyZFzM14eRA4ZOs7cduXPoXKUGwR49H8IVUWoagqNRXTxijKSKUktf
nnvi5BTRn5lbFPpU+g3POKf50WclUpJoT2hJpFEzEiqz8uiT61ZtgXWg82Q+5kiq
8yp/7uSZCClmZ2qRL4ouP4foKmY98iISQy1KlKkMWrj6Rh2x33PD2PqXy6Amg4Jo
+Sfy5yZW/1+nqFfpRa/820JrgcmUyQ1s/mZ1PtAYy4VXkUVTBLvBGphV5AX7RFf6
VB7ofxdj2u0sMz3uEm6ss2ojSCl0kL2ZP0PduYQha5Odkw8QDukAXFWL2xTK4JgE
hq506RZGi7TBh4T+Y/HnSf5V1hdW1nnnW7mQ/IucL15QgGNofdhMRrpQkgAsuSRO
QELtthYKNfepdOIyO+9GYF5aPPf4SeujoKi1K0esikiOP2J666sUQWklfy1c2HMI
kP+vi1NbPtRdmsx0p+08nvxtBywBeIPaWgsH9hwAVPrppUTb6PiYindXSEO1dLI0
UbELmvWhMRTK4DOTL0GBvyCUZe+L/PXQEjH9r4rZrqiX5AVc5+K1cM5MMndxAzz6
481KTm+KVT7izBgNC+3vXorU1xjZnMefY9DCob1HDlpVNlauvJC+HYZjSvgQ9wtQ
3j0nHVMUUXRWRLi5Az2Ym7miwiKfm2mQ0FCshWf5zN0rkUzmO4kyGbSj7ldWIBR8
7DOQftND8KIhYe4QZxvIcqF1tPpLfy2cts+jfdfW21HwT0I4wzmVfju0hts2PsaZ
5nN8VVprINT5vv06gHa8jlkK1PEIyza6ulwCg9i6D1jhPLz4pe0rHUR70s59x93D
Tev55B3wKQ5dhos93CKTpnJhyqWEJO/6dbjRmHm3d7fBxjkYJjKazHPR4/asWYki
++fRuSVCPXVmw4BfvyprPcyAQQ1u3soo4gqlAKfnK5yMSn1HacnlIfnIJ0K0xzab
qmTVGrWk0LmimOaucHsk6aml3tChkSnQCssDKNr7nDg0mjKgeoWRIsLJRwYZmkRp
kDZwAtpcJYL9/pFNBML+jjvKYjsANClsd/cQw5Xdv/3klPb7ooI+BZMLFwm1DcCq
I628URvOWZPDu8Hef9UUneXSpTvIg3ebXJeEbKpmzvAILF2jR+GXZIdjxnaMMNob
l8mYwuDjLoSZCb1VHjDSk3VzUwGVUm4PT1BwbwtYZ6IeXZWLexzw1s55XkmiAzCc
55axU600YcHsJDRnMX9zSPxrtiuPwDjkVpUQ+shjF+5KknDQEjm4ZF731GzqYQgo
`pragma protect end_protected

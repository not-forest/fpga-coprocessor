// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="N-2017.12-SP2-4_Full64 Build Date Oct 23 2018 20:47:29"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
3FiV4Zl7XgIxhJT05zO3E1cU6//UmTVZxj+6FPksbZJJRRCCXAFIKZMePoKO0bE9
Kb9PwbxfLohuRjTzWwPYckkSylgk6OY+EnGNvGwswH75jjpaXtmRy4AbQyQaVNaQ
YUvka/rEDFn2bjLE9aMsHG/+b2SWt1x5tEvZFuunotg=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 52352 )
`pragma protect data_block
ANykvEg+ap+bW6fkamcjI6KO9WIIjY9MFXDf564v/8rj8lkRdcikehled6ZGPxtL
w1TqFtPQjmCyqfTMr/W/ZcnFuL+Z1EykdmGwfzT0V8EeIuUmLS6vTqMRgKX4FwgJ
TLVVrsRCIdy0zVs2XRFNlYMLoRqjX7JO4+UnN9Xd7q5+ii61rbEO4cWojEptr8Nq
vzALYu1niIBymdPv6KF2YFwKAhhdIgQyP0+0WvLB+rcLsilvef+vp4xmYbEn3oqA
gL5GwsK3haU3myLv9enpmAWb1ybXE6VHo3GUhbC3lP5xqRZKgxuMwB3lwkK/6Q+a
od2u/zDqjoYquDYNl7WI1SlcXgtH63zRs6bO+oaCojb4tL8qKDIgD3x7sWj4S4ob
gfbEPaWWaPLltf2pW71E1gLK+4ytf1NDYRD0v7zfTdEMPvOnuE14pmcu4dpUt0WV
jq+LCFlrkf5NdOZY5UtSC0/KjBZiUpxlEHzTz2MuZWcNRZor2YausOsvFT0DgEEY
oy94EKrZNsFpBQLzosD76c5PWSlojHnfndl5HemEHZhu5qrmoQfXPcv5d9RKcfXK
hzq/Qbt16LM+ZcyKPCA4x0cIpDc5QSPXBIvbMSWhn3YbUvE+5qpxwIl5XDYf70sh
b4sxTYqyLRDynf8q9M6oUsBC08jlM9+nIbYRxcnCfFmSNGNSufDWa9ra0y6zhVF+
bOZSC3W5PDTkQGCRfAtQd1tiohwtKkO2x1cC7U/A7BYh/9Ei4a8309/0u3f6C9ed
wLoGBu/AQCJHbECX4vBwFycicA4WwoxHX7yv13oDggsQBjnEBIJLyui/RQPEF1qH
ruvG1JCxjmgiCkfjomIjBdVWKe5tOpZxS7Oe05tDOwSZMVmkMJdQesdasiG6TCw/
Ba4kSIBEcd7flMyNY3GGKcc6p5mBWt7d/6ov1hD1ynC7LvWJMiIjgEpfZdQ4bDJu
Yb0iOWkrACdtGFaxPgCZRs5bHSyM44ISwmqenRQKLDCgBkckQSQOtsN9Wv/oyaXA
0tD+LtnAr+6K1a7uOr4GaZap/ZYk3voqbM7nF3oAh2/6JNJ6qPn4swka+dihZCer
ad9Ow/VoOHLIbfLjcvugQo+iyWH7aXSEaT0ezygI+BXHMcJgwFhAbBZN9WDOwCbt
STiWKazNULyE+AEIty73/sACKDpWeFrKQmvFVSbwqqZMhE7MGuBLpeRo51U0RnZF
Zc5s60jxkEPoz3r+McvZRPXp/y5CcJesPxiCmvngs35CDPi183UqNvIPS9mFj8nI
iHD62L7AyHfLliLhrhC5Yv4s1YqXWYJJwW7fQx8ROms8gm5GrtX0SMaHvjovTjeJ
oiPUTWuVO+BvCIbsriRZDXEjsEpmQdwILwyxsWR90rIaIP+LkooxZTi0kSxmnMep
/xTjyv4ZURoQsX6g4p/b0AiIm4Sgh7/CyL4jX7wAOeAF+JywlZxmWqO+pn28Jyay
U2xGiLwfGeYYuflnvF8uA0BkwSXLyuP2mG+1lEDPJ6mr++buTDuHYE7POUGdQMuj
bkc2bIdzD21Nq4FZKXkmU9PmwHk+SQrorfYaMCiazkMUeEcTyM9Zgx0s/p+hGGfC
HkrQhQU7HCo7St9/GVRnBlMRKtTS6HEStj4Pq2WR9VJ8GuLjp8PW+b+4/ijcllzC
nwVoIdqYe92SZIk2gPu70hea//wZArKUugSrCyaD7AWrHu30isuw3strAptacpKZ
m0dl0ZM9Bv0ByTL05DvTQlZBt96/D0YUXB0Vi+U5wxMmdpTAP/44xX6WJzO8gCjR
+USkE9uaIalwOanBVLtQ46530kdJFO9UHmp2abyKKYOsCM9bl1bJAKjS39bMG/cG
kjJ5OFgmYklXL2CWEMWo9ldFgbzmPfsPzzyTY3SNYQb7BXN+3TrVpPC2admXyE3J
iocdf9Bgyb7EC+DZkvJvLuLyz7p3SsQ9VfuTKBiaLgqNQoy6CinEMDHPSRigHcZ4
GjbZVj8h3MF/Zm2dHAiRfFfZ+UnxwjHxYlnZ3ni/c9gGxAYJPZGTc7/vPPI93Caa
RwwCUP430kHiP/kDkiQ2cglxh4AlNr37PK0xZ3u2/gLYOR2a3R78hAcpQVIeX1GJ
gxffQn7wD7w7uakmBhNj76wgDGQnVs4UnOkut7917YhysIgf9Q9H5VtCasAZVxLD
YEDKtZvD3Hwsm9BGRPELk1RLh2MM3CjntJHEOD3eOA8blTMjtpFMkNRdqqZJ6doI
Yk/iGUc/omMRYFAc0OgPAIhU3tc4LXP/RQL3A1GuPPQxI43/D33dk8T4KF3j0XHx
6wIAI/HJXBcrgq5+w/BsYZw9lH/iHmFtahr1rNAYFtWfUSLQC2v5fK5AvCVv7dfM
e8H0RGbYHBcylKd4OFrkMD05rqePcig2SeI138zXk0oo+UXM+P5OEfYHkaMv4COG
xIcc5YRcSa4di6RjtgnHMkSzHguD3x0y9UN0qPLuehmyvkkAuSzoaLXBSk6dKDs9
7hrBqnpWI2iNFNKDg+Mp6liNQCkz5gveEnaxFMlgXWvmryBCpWKE7fY+jsuIhAW3
c1mMBrf0paOtSHIA8F5o9exF3jZp8Q0VZDXj0rD5xKqPgZBtmngK1q6ujbapqKUW
E0JfSUG5v2ZKvqNqCLNmKJmZ+z0s/QQOC1fA1iUF4t/45pPwX2bLW+x0HS7Yo90R
ls8CrP5wsFxBVGq4G7xqRK1TbCEGm6J1cTRsVBW9UtBj6m1LvhzRX0o4atlwJ/O/
t3ZcUGu5JvCc48tO9yq7l6vXpyQiTfy/cs8pNHUqaS3UpRa0StTFXRXsosfOpPTk
T1a2jjm+fcHC091DUpegiUgp40gMZe9zDrDp+igcek0moKvlA8HohHadgHqLEP6J
fNvX7M4nOrPNk8w6tr6tyzyJuC8kR5xChs2sqCiomkoxvGNsRVIeBZelWsSeprpX
9EwBD68BqFXc1b5Wzg+mxfKGuHEutrneXYM1T8hgmG68kiAhW5kpshlAEr+c1+M2
whFhRSHpoMNNDlemIlcesFqZay0NPJJLQmXvrhK64kALNRi4W0Dd9XU8meyEPZA0
t8BuzOmtj+oSd8LjNrIaIXpMXTyAYsdrFiHUL/pAj82Y5CDgi8McH6KXHlwnKYM4
vnG9Eh8f1e5S//Mx683grcTGBepEmJrztxvY01yMABIENccJFYdfhA3jJ6sgMUux
UNGBiJH1pYMXdkZEOrCj3yiiQCXyv/WIhqyKFwKG3LgLvO1xMCNx3UFS9sZMz/+c
akI3jgDzPanJj1wwRNpW9Nlpg2BL+AJXQ9p9a601Y3WrahRs3z3lsHESKT7wZfsJ
RMUxiCtZTV29pL9MwyfL9Iy8kuBIGui7j/dbB+9iMA2hrqCeDsIuPEVr9pNR4P39
LNVX7GlJdX444ckHZC/AAVNS3kUysOpHs6FGcO0IfvHgZUvZ/nENovX7qlmy2Kzf
VDQvoYhhkt/UBwdW+8iasmLCYaIKYVtBfJ2d7YZ7pAkiYspG3G145nOBeLFxDwYw
x0d8tW/PGqDwwH5656vK8n2YA8lL2ofqKajyIM0KDvCy7Zc+P76/hEyzwEV/NVsL
p53l2KxSauTC9WgRP6t//iVrUa9ptf6Dxue5S3AOu1nOxCqc+gsHbmH/Iw+bePHE
V51UaXqk4nZRfLhd/DCX8LPi3zOFwroEnkzFOyBRKVlDhf508z8kF+wuhEJo+Vh8
t9Al3wU7RYDNEi8NhOQMCcqd8/NQCeV6XWGp33H20unElrDHYr4SVdMNhWxj1f5a
hmDCAqdAJxkBiX+bpHRlciEYlFYEZz8OUF0+OerzMZCfl0eSlVoGwXVLqGjuHaBe
dDlCjJTC67BsDzbzAofCLW5jb5vDT6Tyl7qrfojnXRu0C8chzirdrL3G1romkwvl
g49g2/+cZGQQXlvLRKEDARJkgLRBJuHqyJDpcDYk1dlGIe/oya2BdswdteEm8vNd
OY561xm4RhrCnehkYzludkcR4ZlqDY/l/eRHEsmXjFwFfRS9lAaN5/KH8zQbITiA
dVklVUNJj50tuiI3sjEPESVGIgz+8jbj3m6/rOGeGhf0PCg/DdrI8twtzvjRVpfj
rAwvCGPPmTyWhqHHLmZ/lpRi6IGcjuo6u73/LsyTM/mqu+imkDiFG2rAKCbmB5ID
lWh0MN5Jo/Dedl0RUc/uP9MBoGxsVVOpODMsOkMtzoChYfbLYoS6ujfPcw697DA0
Kh4EROvCm+FoieHrQdRsECGo1GaCyrsFU94MwcbN8MFu2bAzvHurRgCj5PyZXU/V
W1DSZkct7F2M5nrp/8trLrQiCjNe5ua3q7ZG6+1L8uYN9fZrtjXmjK8eJ6HLMSE4
qdbObUaiF88NAJfUDiQ+YwtpiqhSxsMYAjFMQqjdYmzHMZHxKf95wl5wxTZKeeg1
K3SI5hxkfJppyo5PVt3KZqa9yZX42AnBkJAG4YRWAOROHUjh8CIefRQc0K+fr41W
eeZWDXNZQX1fAhHSiUIgRsXlgfNAsQINe//QjEtrjVPYc0tgcjbgFa8nBzA21MdR
0x7menWc9b9Al25guUfRIwsTDg5zMQkqV5inMsaCCgh3c7RpeFyeNexD88AptYP9
klMy7IEEcCb+pvkfHP+VGloEr+xdr2HIXJ84m+50IdQ/jwF61pCpEct+v/cnY/hI
iMP22fe3D8s8X6VfqrlYsX5DxPPS7sVqdG0CIabB0YvAOOKrUZFtPWIXmD+4+K/p
VyqlF/eRqU3q/qCGAWUxP7lyt+bBmtHg//mYm3NHgOd/RJJZiHe+oUa5hkKwGjgi
fO90gw0RmfC8aNSv4oyjjC5nLPOCsUvylvwPaDqTHwrhQ7N5g23S36zacTrMefP+
zMbeUkfMPTiD+AusXn7veOBcjmUYA4ZTIXTz+2UbZS6NCMupg1yDOujgPmFDj+HS
MBToN6lksYcFvY1sEkXN2gihD2T3+x7KvbR+Kj49TiQ5qQ8QWuLmCxA+nbGQBscO
KbmtadY8TJ/4iK+7UjAJZDOxCzGjw7AoMLhhRzWHhqfo+JBIsEJzTJB+BXrllwER
ZdCE8JHerIfPJgZ2HNmMOYWI0XQzamZYA3K+n1j26xvadeihAwyFNGy18clUwomf
B+3sq1no4cESHtnldgfiwQ+4b04SoGe+cjF4poLN+nxlX9pehYkxGeZCpARwOk38
kmlav7V/G2TvrSa/QxWbi5yhwsQjCMx7W1bKyBShZcJrcBbMj3G/RGAYvzzWBA94
PJwkhGk3tvTlDYFn1LRYdzw7EBjK0KOaqSXhJLJuqCLfAokCk/6MCMXfralf+MxW
R7MTe57dJZpdCuhSRsZL9/utQFZ8bHoqP8YX7ucM9aj5qsAW/POodcpuXFoz/yb8
WEFhdrD5V8LotYmzrkceiqsR45aKgHUPKOiV2dc4sojHKV1/2VPlBZ7i5AdWV2Hz
1UaXZXwho240Cc+rXyGmC8H6EWDhGUMrMh40xAonuiEBAUtc0OO9Ee+ZLoOBZg/Q
rqYYkaWJUaFZSb9RvC9XMPf+V5219vBXF1k3sbIRt/ttPUukyMQXOZggTX8c9etg
JX0F3UGrar+hWdnRYk/muas6r23k7c8QLvGenuKxnGn6M+1+0+l0snRQtiSegLWL
a5rG3tW9bAeQVgjaLLA/eYadQVneR2Afo84AyKMqdNRRauMu7NRkX/qvhXUrCZC5
NpSW2gb2f+3Y/EkLwEkIzQ0wRPPsnVRsu8827AOl4d7XfVnzoMwMUS2hpFFm/AvY
VAp+HUsQLKSb1NjwA4GehhiY7tM8lqJzUMlqFXPfiwwSqyfXWJ+9bzBuQnUWMWbj
ZrvmAuE4cwoniaNzYB3OUIo6hUF9w2QIk2X2Op52OiL/pQz/9CCuaW0ej5uurzH8
uZCC4T/bRAGbkU9fjW7WBs1Z1GVye4vLabk6UuvQ4LVPabk7gVoyeYWxAKACfZzz
MqhWGPEYmxwKMRGWbtbi9xeBQEEX70ycNwW23i98Rn4s9HIk+B3O1jyPr6pNOPnh
kmbd4ouVtwn7ZnGEAa0T25t73koiHbruSffz+h1OkUG7zkVAr0lco4WZvJyk5ueG
U/VAIc2KMYwdUvR1gKWLtT0cHMPkds6ezTgzoyVGDhZehXQV0ahwuuULL1U5Zk5I
UCCWfjf+H8gDv8WreXeHv6o1Z0TsT+AAR81NdOr415QcpkxUrDoRvIDGbXLJ9aGT
iQbu76SxEkq2q3F9fk41/z33gxhjs6vOrHffSXWpd3thwKQ//4W7IWP+uCVSmERW
SnKqG7d7VrH6PyvWc7QJIFp4LMYYuTC/+pq6rdewHRJovEL29RyiK37y3totOgCA
UEsT468eVMrolkhu1Nbbm2pqlCV7U/FVpZT2uHPJm88bX8JgyOv1d4/GYBaHdxaG
azbkULe+7DzrwnIeASQcfDs9V58tnaSJPLP3EgK9EHyn0Pr1l2HPgDiljtK64UBt
w6lft51w5eNFTjXzfuBHcbPQ/NKhNFlzGgwIZCLVwov6O7rbH8nnWSK5bGYX2HVL
fIqwlqNCu82dSJZ0Ezo2R/Im79UvJG40Tls1MNTiLdkF6imSZglsR+6mUTJVDUMb
tZoC+YzSzlVXgi1geVX4znX/mCxnKyCb+QwmHl1dfpv7hyE6w34I9KBc+d5o6CuL
wS8enrBum2O7Iqxe8FUcC8EEBwngDqpD+Mpi8fXjNLg6pv9UY+HDglbJmflPgKyv
HGZfJM5/Np72a0zRdfkEwWq3hNusxH40wXrKuM25dxFlS3tyQgM7sow9kQHoYP2o
kuxCWA8wXh0jRApqqiCEjDmD4mPcUvluUWro6r0+QOId4QPQV7H8xLgBSV04EUni
H8eopucElt4k0Uh2qSgQ1qxBLv41f4BKC3gXqEkW6f46+KAMqcSkdv0ypi02Hm4U
29NeikwGWZueTPX8kR2a8NirnJfJm3UyOR+xWZ6RRPYU0hRoyr93Wuzt1sj0r5r/
OwECB1QMfuXU8OpFiIPSwXAr+/6POVmnOJBnI/mWPfwhMYrTTu5cBc2/z9Hd0drF
n9duMxFVhUNdFaloBbX8J5mtbfVBbnovEqUVvAu37Zr1RojUBzK+zFsqLzEFXAmr
t+FfdJTCG/rgnOenT0BXTf0EE/6qi/kAi5Pa/gkNmw0OIwpR4XzGww1NL/Erdz6m
OPjavHLAAoLTzwUbYbVcFWRhik2spL+cu18zDtX1uoI30oFdyNmeHXIdKIIePM1n
epbyp2YIzWveoGpt9I1MN97avYs4uCKPxFV821UXg8t4hus+z0jSgT+TIxsaBFDa
7nuTB/ibAT14UF3RJF9C4gUzcHPibpewumVsNcyzxx+e6gMGGwVMq0xheLtCcY5+
TTSXkoQrclrVFin2rA0TRVQLL55LoTUOmacu6VEu05s/l/4mH84q7EL6OUVPJTSp
Ssx4Oe4+Qs6RQUDVl7UQ4YdCwRNK8D5qQvv+0GPJUJLU2ctvIHLN0AxaIUkSM4I1
i+FvET98K+XiX2dxFVPnJ94J56v1F3WpZS48wXdM9FmUZHAv5PLR+GPGrVNnFo3w
9sE0VXZ6+DBGorbMqOp73G6xSUq8fWP4MZQfFuOFwgNrUw9C5RW7pE4JnaIJasJW
ZElYXbX2CB4KDuiese7aIesc+RfxS2aWvAbtPYPGr7kCrTwi87/BwyA7qXAMxfBS
xV8UKnJvVYlZz6ALbgndwO+IAX0KbO87ZTDcaGVcYm9zXgmdC83N5tCXXXVsnYll
kY6QifFbmZK7X4SSNnRbYBR/twdaT417BOBNdgYdy0CuNZe6Gb5z+HUPQCzqavPA
lwJfj3Tijt6XA0PY+Sk/VElyb9mZpNPr0C30MmKSTEPNdlDQa6vEh9tboaF2rkzO
WXuY9w517LyS8tRWxaSfsJr0v+s23rYXRKFVYkM/0mXsX1WQc021vd0h7hV3/+Uw
yPA2wHSDA+4DnolscgMG3Oxe5fCYOlb2u5II3bVccguC2wrabHceBqVxYjspx219
ySk6jtvBIdbln7MGDP+Xplflm5rY1y2KJ4Wyu2JJIpCV6Eaps4NxFF5SLGVxviGI
/ZNbCG3IDJZr7I2xyemY6nwaloZQD/0jo5QKl9+4Aq0qsK0lwQ5RuQ3lUH+MJthm
gpfYW1/gemcUi3tNmYwjR/B/0oRQ5QVtQAN/OuLSkrJ81zMWA2wUPjyr3DvU99Hu
t5Sz7NZz2rEUXoLgVDwG9+RwMAa3NX5E3IGHOhLwjfuTW8iZOebE24sxLyuxK8i1
XFewSOubbBog3Bb1/UptkqUrhM5arkVcNgGqWRIQCH302LurEtxk1zDzMkJ3o58c
HBHTOU7h84wylhzFffAxseWtWiJnoA18EztwYP42J3v113uqraPj5ee7MeOQbUUi
gjKOac2nooelH2rcHutBfO728mKyw/L1blCNs8vNngM9i8trZYhiuqY1Plmn3yb8
vGLOP+Nb+VGOEVfMtBqItmQ9/Pke7rK38O63EiWsiORmN9UW8KZxrh7m41XskUO4
UzDmLsTcQ7sCuAAE2Ih51s5OiwN90sJIjfACibUfYun9CR1GWNY6PfVIYZ8lZ2zn
KYVGD0Nc9Zw0+6QCaFjM94AL3+6VpbCk4hc0421mJvuC5Rdm/gUIcYr+yll7TdFm
cLtKoir2DlV+r4bdanOe1uhcQD+Yzol0Id+QqM7FVxA3sq8IYed1BSxFpc5gAXxj
CR8Ccup7q4qnxAknkU2tRD5b5Qocwbt7XbYksLXfUYz3mseNTOvnYyf/bDbgcqSv
x7HSr5wF/T4GSEmPp1AlCzrWNhMBvx2wTql2bL1VV9BIPWtxjIDrN0MrVyiq8R5S
jhVqqmVgwPHtp7xkPb3NZLnqIeb2XhvbpAcgPQCrDMgRAbhOkOQgqDADBO/Yznr7
LoL4ARe7jHZEdWikN4bj7sZxvuZSMXQTj0ssNdLyGqQEdYrDl6dlET93NZa04a21
HbCnK1Z7EylflQ/IpIWQfF6W+VGIVtaCE6jxJ7eCA49KCn8JqByyxPIHNTcZyGwG
s0MwpG2Z7P+ptPe4ODw0Ol2dxBu52HuoKMWgP4tch7dYy+J9hX5PWRXh5pk/kgvD
cy8TJKrrZohinfikY3FY9MCFeXSJKHuTEgwtZavs3PovESPc/jDJsWLpHLnctGoe
mYXlxMnNiNnnN8TglrAwaKlTSan6HESQXa21hspWCFERCOoH74au8G7FE3UePaHg
fYdAlOQJntJfmtc76WzPgpAsO4Z52tnfceolY0IzJhweb8+VDdGJmLqCA1qyIijs
o6rEtcKsz6brzUjed9gbJ1BGy7j3nFYydhNMo8IZSt2CNXLY0cBt+zPkrdmSBH9j
iys5BaWfhwCXmc35i1pqDmMxOs2LxmO8I90s9LEKj+q4za13FCxoRKs65a+MoAA5
eXB2bISbRKi5pT/0I0IRkJpA5O6pCAAWVc5t5+YU46x/yjPKPxv+qnd0VqELssjR
AG+Y9aN+lgfhDDGetS93AhSt5u2F9z8WX3AW+qnkOP+Fm/pWNnVjs7b8BzEMb4S6
a5EzCwe6zvmQa1O1Cl5ZmIrZyma6DlYhgixK8dBBjuhtVmf4+X+TICD/y0gGM9rO
g56cl38gfinmtyTvTA/VEeDPIjYdV0itgvLXi+LJusVbh+uoQTv+YYSosOwqJFD3
4m56PGisRfAIhxmVRyGlzHTSuUOM7WWCBbtfXZs3ILJX6PL4E89hTY6FaTRJgq5y
vJNOlSVdnp3gecNDG+NN0quer+0KliPosM7Bti0pHaifv6QTAdN23U5Fz6wWMHkR
ecBDMbFh469R9+uGMwTJEbVkvpuX3xCA8Ir/EbtXipXf9+tqJ+mK3Y60tfcM7H23
JGmrYV3AHIspMXx62emJNdTPY0bJt9kiRNf1Jd828/B3Yyi6wVaLwCOeGtOvvPx5
ZO9I6gur1ZGcHBafGCD6HTCaCFTbXABOuZhVQ7ItRx5kv+D97xX288LmA5qUhGoD
IRteaSgjgIlynfMZn61bvRiSMxfQUJ2x2l3yAhyEJHArpZTEanztmF67LcZIO1ZW
dRCJ4GT4/qowEPb8WJ4VR3WlcK2+zrInrTE/mpI6TMQgl08RLZ/fI8kstnwszHH+
ujg/NFaBobI/TCuriMp52bNHzh6Sli6DzksiLphAwLdBu+7J4TgAUJKxTidLSEH2
W7fYosIfbT45iQptS2vWCokIVqJYENEXBBlLED9Qoy5s/oMp3C3lRsXdQyHQdizd
cRhFxSswGQ3ULnmn/3fyIaf3Xw2DzmMCZ2792wH9Bl2xEx5KegiJT7mYFtpM2sGk
ZJkhCpsncEvbep8vb85QJ5S+fvuTckMOSXLsH0dd9AiOiEuSDryDBsNBuLLln4Mb
9If6qRO1cK2coyIEP5jjho+jCg+Kf+MdJ6pwIc9qLk5Zm2p+/SDc/Jq6T4anA3FM
BzhcfkN1mO2bv/EUfmjqTcA5yP1GDeNARG07gOIkVnyRVD1Rak5zgqwayc1Fl3BQ
oyfscPF7k8YT+gZ9I5Ub91Bh3aq1UlonL/bfZIT8YiAhPl5LQbm9VVpYt8cXiCsD
w63xjzB2zepdzMDetMeaQozArlAOdokBGUR+KYJdTkP1GiiBkKgT1OeLa13ltkEh
3DfHyRlNGXR+fBXYJBplPuZ5WPZCeIXao4LAdqC2O1vzlnWdRYp6DNpfHUd1xE9C
cfJcPGpCvG30E6jxMF7mle2WvAfe7qZ/nyQyXkCVjf2cPHrWAbccePdSoUag4LTp
EA1+bvVsKjhKeUfprNGw1/Bsfqrmlnz8bTPVsP7bsMwrYTlbWWqkgeVQZzoOj8d5
00UvIuWOuEpQF7+vlYL0lzDJTsabOpIPWOI86ZDwdvdPXPIM1ZJRHEjpRhw0Ldby
CNg5FF2dY2Qsf1zGjW2B8OcJK4bPQIVXfEpiPFyc3LyW0F3TTwKvtWDjVmaY41yd
lh050PLjig9tZR94VejfN8xD3g/PhQJSeaVIri7UoF6MEVKQa3NGevF2us+bQ7+k
tZZlRKGYH00RwiN4y+KANcd62s4xlNiDBsM1nFW4uItHWCE+zC5cSO+MwYbgpqIV
tyNOE7ibeCAxt5TBnc6QCzmFHp4UlOPQQpz3+xHXuDpjmWutSH4FWfHcrdj+4x6P
1Y1ZHMLBDAAP370G6OWIFimFarRJ8ONMXmrHktoh6brfaUQHAHlVBerSE7WBICz3
kxCmZyief742GvF4wzloNYgmNQZfedbeUM6QmNxJMtAumQYUL08h2TW3gzc5UYR+
aqCRUOVVQxSvKIGgnmUpjyZFIqX0O2xc2/GyOuhsb+4eGrprsrGgOcSfQs04Cij5
iJooIT+PySrAc5Ovw91W7HGWKy4eZbe3cqoJsK9UpGPEzUR2Zwhi4EzGfMVMOJEB
KmpBdjTR+vDtaGldKCXIglJ3MQhGsUwTQsfTJyTyrQVLLuzdBS0BCrC44z9dAv7p
90wfoI9K2Ou7ySo0lvBCxUxF48DYHdj+3v++ctm1NEIJs+y5xSY6pfDnI2vl+xHC
nLyPbWfu7wZd3fuRlbHoUAplzr3xM1hUfpA9RcIP5xUfsS/5wU2OgzyOZ3JX/s8e
7uT7asfTeFk2Lnx3cur4hrr9WqXE+oaXOco8JauVpWUJbGXcJvnT0gMg9oEmrh0S
N3NjZ1+tI+6JM2Gd9gOaazcZloWe6qSUHHFB2sMLxLFfTHddKUo1HnYL2+0wtFZD
BT3BaeLFkHXVLeuRxmiNUUu1Pa3fLirHp9z789c2JwxXNgLShdPMqWYeEIdsTg8m
EAA9o+Tpe8Oqmwwm45DBq9o82k3dtuDZU1hpYtgL/NC12Kn5cPa4OJxI/p5pBKx8
6RXdAKB+0HQX87a4gSm/9tXlPOx6pk+3EBm4gWEAa1sdaP7Mrh9iXmKd4iVcRzbN
Z/p4tI+TgJifLeVRK2hJzt65ujhAhFoBIE7F9kGvPHuPQRIHHLKd1XEi8qst6V89
eVdwMxyRfOeEabTVYX+q3QYmmZMmp6ZBOhI1LoxxrOmoKgV6X9cvcgZMqxWOKghF
8CYDPwEHAFT4LhjXncWvFS/K8U7ZXwVQe2astzs03+zXHpboydQP9cZAfkLl2toq
0eYQlERVrZKCTk6EkX4MtYcgYzKSzCRv4CYCjRGAOY8MhA2EFc0lZkS92HWzA4tk
aHZ4YkIb+rniMWjtjxgMPjVHvu81JkaC0wJEqHWnlDrM2Nzyj4hPsv3Itwy7al6e
alkABX/WlPzmqjVP1c95v44IzlxZ+SibMJdlLi7oGFFKUFXIpddcWDWiQKcgU+jZ
DtICMX7BojnPyv0hxJQUN/ow+TgUutg8T3vOaK4ebY+Vf89120odomNqVjJIca/h
SS2A9/mBd1pSTel5czg5fnPK2mOD2qShIgamjjplKTlznFrb2rJ4lgMPAJRibtw5
xDwMQ7FGWejyJLzMfYB+MPepOJq+ChAHcF15rodHk2qTULq+e3+H0eIeByjQVnLJ
/lND6nufozeAAwlmf2tl1+9t7K54El/Z60mb95dbZpbhpGZ1gY0xMqfSUUnr0saG
iCCDMJkZPtW3UwNJBJ1GuT5trmyIMDGrBDUZoY+ppmAyJRHiN7cd8+Bfcc5biOe/
1L6wl6UGnxOhsdUmhhnEXvqXLvLgOmNR6AVphKfAlTydEXwQ6K62Xb+TA4aK5r4x
dWcnADHZjoOv0FfcGOSi9lbchdeiPgoeUnJRRtaFIu4Xu/b+pTXFjBymFRbLG/WB
XVbz7QlZrwMmNuJ1IDdtFx+qL/nx1Eubotg64HBFYc+FEq3S9VZYW9KP/mK1dE3A
igME3w2TTQLyholy923nFWxW/W5yLHuggWXFAzdaaYrT6qYjDFH9L0kNZqLuhOV9
77wnqj3B5ryqjpikqqYwtdM+D0ftIS/qIw45PsZ2Oq+dnTqCB/ifzrH2Nw4X4gGx
o8n2rpzqLc1justbnWqyNR65q44hArhzgdPfNlcGVxO1GRU5NLzeQm8lks45YNx8
5gqwmhjyV0wgm+AurVlVSKFYUsTsU4AJZdYxLnxIt+vQmElV0MH/yCgPxjxwi1mU
iuglNkDmboR1NNVNdUQZ5YfXHcR26O5qR0zSl1ZNTNTTb3+pk6ubTMxJiyyuRnGU
ZWYNmk2UYAP8zwbNxKNx8EqTlfp5BbqzDAUUvPw+vdFtme4lyOgm4jkPx3jZPi0q
73IiUqJiW2d71/dNpenZEH+aVF88yHS9smIr5Af37Qc7E+W5QXPJLeFL6j/kb7F2
MQNMBM6wx1OViEJCp93Iuve9Lb9TG26RHQQ1WTkKhPtxOnQEQfcZEba+bGCkOuGZ
9MAWqgHs74OwRT3y0Avle64cnJbCm0rXWVY29qXObuugpnUVb6oHcO2rxmeOoUWJ
nTPG3nSoMm5J43WiGZ4mDjnuv0Tst9R6mUekpIqiHYdalecB1oS5D64IzfbM7+1M
E0+8HjN7xA69coO9k/6aFx9eoqF/6MD4k2tCF7bFRlzqBE2Y+1gHztf3hExWR5kl
Xtr/3u8qrJBq1kDSdGxtpcXT43D4RWRaMxDeKshgXjZDJYmlAH+js6DpkouOMa5q
bfgpZ403kzuSwLyESbJ2+FlRvSJcAA9PoRVAb1HGjaLGnXU+z7/DBb2vHKDcpOxS
yPIPJHpFNzhG9lvfE3X6lvSGRYk7aO/rW+OHyzfM1mrTG7WGUsD0YZbbXNNyXKum
GEUGEL7JVZCXzkPO6apZDW+CiqjTXV2KTfSvssEnRC5j83dWB8yYwZyHThnPSD2p
GXz+qYVxCddmjVReRhqNfUnrQLCKR+e2Sw77diqqIgzhrDm+E21xKHwH7vIHTeIi
QZf1NO0bMdZql9qkvDNu5KJP5/RRmHnOx3YwFqg6V/tR3OyYelff2bzCwlA+mpXZ
V0NCY19AovEpcuHfVuswl0MZQne5q3G3IZ9WIdGk+j56P+eNbwRl1ibE3LYb8cLw
zymgnfbDuckwn/CSS17AXud2kreQjKT2g/LI9TgBqEZHxfDIFYXyRVYiCJGEr0AX
FDsMq69BDOlnPObf3CXA3gPZzFUqH8qzl4AQVhVc3NtuL32OKqk6bhca/tCQnX7T
Y8yMtgZh/Y04ap15veoue0dm1eNtRmC+pb10D7Qkt2vpzgf5weiWdg6dWQtiBk2B
jH/rtSpbPMIh+79tPpbb/TFQdYWiby9R2FNXcpCw56lqxlQrzo8fM/T/XqwYOZfA
W4phGjwUY9qLVv7HLdM5sBSa9hGude/JItfW+LeMnYQo8F9AHiUpDnlj6mkVLG2K
cY7p0uyv7772GBEOsi05avqzeW8R3iU8ADHJLNxf1MwbfxM5HJJ1sWIScRpF5j3R
zGKscxpiKUvDyuZPkwCeDmsB6EO8B80Kc+Pv4bdZNhnecJUyQ8IDzaM7cvm3ScGD
ahanBDXP+hqTz6QBLk6uYFntf2N659KZc2vI8JZcpZcP60VyedkQT/WF8eZU3yT4
qB8ctgeIn6KTw3R2JLqapxRZs5XtVhmUZH5P79u7JQFRCektVg2JFqYbZ80EyP2q
NIeWKI09MRl3IgmuylwV1qmlCgdMkr0J5RvsjyVTXjnwpj4s94sMmfEzxnEYtWi4
fSM5TXj7MzQlqa3SADoyOh6C9jbUeH0mPc8r8hcHtwuH6QV0cZTaDfoCJzfyWnq7
kTPVhEgZjW/MEdabQZZJ1FZTMoa6QjjfChAbXTzF6bhSWcHFwkqyTwVV+tPBWeH+
PPMCMVYpFLKZUq1I2A1poEkETHy6TRTZ3vnu+DbijcXhRVxGqMI/EGixhdweG1PK
TXmtYQOHaxJH/zjPG1ETWNckWhFqigyG+8Bw3ctVzrjZEx2hNfXw2teMFuPL/gXC
fMyWAcl6Kvl0uALZ0eLxnpInynKgQCddBV159FxRtoEPm4agrGv8pXr4DUeKObFq
1dW8mH07HmKfXI6T5ZMxLy3pxF9XPaZmpGlKxKF1pfp3WaxaE/dAdSHDnModm43M
8WMTssydSqwqFAOnuKU6v1moTajhPlAhU+jntYtjeqGrAstcdi1zlWFnuKSZxPCu
RiE1C3R9vMkIYpw23QKUvxhxkxb5lSCP9QfbUdi2MByMs/ILQcElsMk1mNs/Vf8z
1pgdLctaC03GnVldbL1mC+YIx/Ibyu4TsuFRcUi0iLtbIQ8bFz/YWFwRefPnHpSw
0dertnAuqgO1xv9EftI72z6e9bVRNAGAgt/K1ebvCRkPFUNt8YwKcNlt6YZqLAEv
GqsHzpAwGW+T4e/Y9APa72rXEcDMn361fNbrk1ordahqbRLLMQBAavgFjgYec11o
PEnAN+fjrRYNGpASrsa/elvEiQ00WqBCXNqR8wSGSyxD3w3nRJM2fYsMezhNDg77
N8Mtk7hsgUqftqKuz9kExm2GzIsiH4pm+zckL0XwTTsu8AzgZ5b0k4Iy1LKdYrTx
n/XUWSXlJosV0UPFTgP+GvSTg3cV2qBoFbzCXUKVKwKG1RXy+DI8Xe0mi61UPZZH
qn7xd3G3Q7D7GN6rnExdbC3cWy4nV/GhSLPQQllIrpvL38WK/YECnwcgeoru8xFC
7SpKuCr/YcWKnDMjl2MMSl225xyueKSQwlDYCnUgwwyG1FDlW+udGOqeg0wgbYBY
vIfJ67P69NvOtx66NXeDo8nnpuZsRncNQ0vPy95F8NqxqfMYtCla8zoeV2X0U1mt
QKtJKXbzkPq4/LgN8U3JbXegUk63ApM4j8jJBiC0AdQWgAE9ce5uwHdlI47avNzc
iNl5unHMIVCwvxCJcvz+b4DaOXFLu6nKiXrw+mHzlvMVuFho6DPiqI9A7De2SQ/C
VLQdWpqJPg9WIRWF6xiZmtKQ+/dorpm8Y2CAi5nInfox9i22FFZucOGyJUwrB/x9
2U8yGcFHmXVX5YOvQQTal7uayGvYkujbXHilMjvHBYYCAQOyuwQIZxBV5dP3ZZaV
xoZeGBDEuORT3s8EYnhhigHoiBfd5PfdBmosX9rJuH5jnwglT2wi88tJn0/dGoMe
8Cr0rmty7DJI4MyCfaTRm64lq1kWX19SdG0NegLcAhJflyPVHlPrL2eIk1eYvPH0
ZTNHjMb3/4FvZqHTlFb46/NkkOzHLl3dkieeU+PnlEjM042n/sLxPXqWEs0tDsYz
EffCgUy77PnyeP27/PJJyfe1Zj/Ineaz+RnY/W75zNMEz/VSQ9mbQvmbGF4H44IM
B0NGm48V+I8h6N0XjQDKN2xHDWCgY1UA82KjLC73627IofFb321x9mtmiZVXdWBg
o5d9THRW/WPe2lTjevqBBdAdm/94TGgQ8PKY6wGyWNRrfoviSDNCLNsx8jid3eu6
/ERoVSyzEibO6A36+vBguqeZQSSWMBQhijHcY88uYtxr+bAlIC3CZhAsmFW4c2Ri
tyVirfw0h0oqvSQ5vruxTJ+U6CA4xD69YG4aeyeNMeBOmG10ax3Agfp9b8gBICcP
iy7Bx1dzyShXgCLOmRCgqwI87eaFzLz+L8Z0CBc4JPDmUMiqZ44HQ0ui9YASUP3q
C2zXllHlW3G2O3tScFByfphEPhpl6xeLqnukPYnOxSyUSbR/IB8katStdtKLwj1R
4/Be4uI148O9aH7Rs5gM3k+SE84S/xNkRU+874zqqVf+tJB3bU9gpE2yldMUhC8c
UqfX9Az3gysohF598ntCwERW5F73K4tNF42Nup/uakj84RI4SJPG0hYkODzZ0G7o
uDBVT8kSzun3B6WUXD9DD82MZ2+h1169M+SBoBurizkswuhRAHMUhOztPPj1DsHz
jak06J2OA+VGs5xMXQoU2WP8tLP80SvL11HtM62grLQqp42nW/zZ7dJWaCYNwuZl
WlDF2bp/9obQWlCpC0QdyLfJV4b6Jx9fQtGm+f74QwjHUMw8fIGj3m6ODD2lJwYt
xlLKxEiZbWS8zDaP5d0pXRJhMZyznwpUlmnuoMomLIUYEYiFo3/aFiBhADZdDFKZ
APklf1nN7UKOx/R0BZ1uphnbl97BYjFTXaG0P9zkF97g+FCeVkze/PbnObsGHb+Z
TAsZyECq6IXYqhw7yielbRSFYSe2uAKdJ4k3OLXdYxwi10+BXZ5oRAXTNOunrRGY
p1Oinjc+Z8u1B+2JIaLHNkvpNfuTF8daiE1fvQ0UbBNJcp2ccO+0ugR0BSbxRYOa
utFsaS1BByoQUSYU5AiR1dmcRl2ORK/2PV8mvBU3IjsOC4W63++duH2bxTsYNBj9
ZVs80wdlpuXPMG2IlbzLfyFRYY5ODP0WkeaGXS/GT0PLZ2BpVGJWWmqDwpnc84ZX
u1qj6MnhUjl51+mP61HPmPnIrJ51sUEioDbVP1OZO0N8pwWW/MD55cyL3LnfPFFf
YxKko5Y27NwqaR9ABuqMYoJ3Lkvz06RZNyt40HOQ3s7dc1QXQaz2ZU+Yh7bKMGos
WaCVGkIHyFwFe4HuzFroSIB8kK1wQs8EwdQQhevnudNbVVPhg90KgoglwjJQZ96B
exmtx1qvn+A3a1f5mXQU7MejZGvRsMt147LBlcXWPI6nh3PZRCN8F11tjnMcsYus
WYraF8vgyAp/aEOS8I8yJDPRJrZNgemhb655KapWo4PgMwjebgt5fPAtr9g6zLmc
dnaf2gB5ZgGKM2QZY9cov0YQI/kjQ3ZJTKNHHZyAqSuLsk3fCsdHx+oM0FK4zH+E
A626zrpqX32EFZkqFAla3ThhWSCJki5jW8cKk8xjSGnS0ZUk2eg1dJadfo6n2UrP
z/1zUAm6mn2klxbr06+eT90mvaDZCqpuNkUFlIXZ9gMev6eeHuRAg4ncMTDkcYfg
MaK8S/RsX2AqPG7bRz6lMIj2w5CvDH5wfVzuZHQxtZBPekMx3gGhe6YHNN7GiD1J
mN1C9GBjyU/2+V7mPPgp6L/8FLclrvMl+VfQdY/60lvyaXjPiHul0otnFPrGq0K2
r6hlVgrhTtjXDOMbqPEr/ood+0823LGYsYez3VRGvrgrdG6F5cfEpy6zww9Mgpk3
GnOCuKM9dzZiV8SQwmCE5QvO0+/StsBMx5Wp0JNS9xNbqjUEKsUQVs+mQAa4ZrPd
gULeNDh6kz1jFmf+54wUcjBwfRPHHccyO7wcmZs7/I+dphrkO9MhhmbwBdxUrOvJ
XPkBuxBuv5xg155qe7m75yV+HAHq3QqLyJ7c46UWnCKJxew0pBCcTqaHCASMgBrv
yWk4FGbOcBfNIfcvY1ipKzARPY3igc3OlrSTBfrq93uZ7n4aCmMmtYJ9G9Viv1dK
czCV3MiFt6jfM3hB6XRzoMq6iPp4ZggvhQ27yJSAzkK7yMXZNHcESZPv5Tg7L+aC
YTnrXf2Fl3yOsSp4ixRaZcoF4wWh1OG+OZQohHGBzXSQ3ls0o2LCMG6k7wL2gysT
lBVhi3hnS3sk71SgxDZUbzey3LZLX+/nwRYvUjDLeNU3EkZ64m1E3ERc7XpExOVC
BEs1ohni8fZzb2XHo1xsUld/kZXrfV4Yfxaddh8GbPR9DnYWAySK/84FnqYAtrDF
Febqt9w7bYifYW1O3u8f65iyxPR5SAVM7NnvmmJN9b8xyWpD/xs4u9o3MqsBISz2
tYsCE3HHtb5bWeAFVRiDSyImI1SlyyQ5puCkTkJ0995W00WwbbvzjODpHVb0aOvx
C39gVMNu3v1NZ3/VFMFedKpWZNitZPoCgYhD1tYSlTw1Qy8i1/MjeBxjdwp1V/hZ
vtnSROGggOLcB3LQaENZzA2WbgxxkxXq/dELlbjPPAIsLqQHylOXMg1ylLlCgBGt
PY0lXXFerB/9I+AIgQzwJKNgtcdy66wXnctPEaqmACMW5Fqft6ZyQ2Gu3Li7frJw
HgPz2lfE6c12RVXz99FAtWToqhLlinS/KXqy8DUB6+lLRju1ytEsA9ZQ7HUYiXlX
pKQH2LB4BWyXToTUrRq4S8OdxkCbYHTaWAjtCGibXMtAE8xhHCw2e9609jYQuvMz
IC+Z+T/0+Ra9QX4VQKZTpIGcoyl9R5ph5x+TGhXxZgR+j5Q9mhxf60NHgupP8jGE
V/Nb64wN92cCUW84qdvPb6KXqlbfYZu8UcemgkTZGNfLLeYl6Yz+egv9nGct1rpA
AwkQHW1DY01xukaldLzgYXhB0td1xs5g0xr/zkoeEmfm0SYTaDCc1qb9n83ignKH
GtmmZLTx3cp9gjwp1ps48skWe7JH1Tu+KinJw9/uUH5z7ToVZ+kUKe14ZUBn+lDO
+11N38hnF2AjNINf4HOzhezgm58Y7Kjxqd0i4Hpe37S8IvyDpnm1qGn2ZOb71cy0
zK5D0BAM/Bf8yTSpqtOYTW6XawvnKhJxlaieqfUV318O7XU6xRI957boiPJesrTy
aCyff/pS+vExKUuT1alaaA3PmZHCnItWY2tKbe0bu+seckiARPphzQTZfgPyvkX7
zF5P7gJuEBaYrFuvIGeNYGprNwd0FZBYG+3lEcFYtvGaTEfT4H42Mz1NiQDfAzbg
dMyYcyWoShHqhchSULqcw5/bgCEO5HLEQOfW/qnLcB8XmZ4soxMew2NYEKmsyyGk
Cl8IRbftNdIZTNromxCkARYzjayxjFMIG/z1Of6J9k6OktTKr1IbN1xCVXCSdppy
1TLr3laxfi2pknp03Sw29Z1+SYpN5BoEaQt8XDBLVx575fN7ATk381lS6c5vZE3P
v9hGCfw07IIwpPe4LktPwQQqv+R06jYNw/COwF4L5BoBLCF6r7dk/sXBeHZwg+dC
/MFHkLm+pYPbvlYBmIkAwDt8TWUv2ztkZD/k0ykE637vM7+QaJqZy9lPonvZ95To
Y7dgCxWfDMF8S3RLLcgABQDoiJ8JsGM/ih9Qfw8Zjn8oRYO8Qz1ndOz3fnDdy2Zi
xcob5NQxusYg2mw/Wb7pbZq0AvwHTsWuLgU+992kwxlaimiIM3S8NAGR+8rfgiKK
APG2OgW4hcyS74akMfnH38HmqkbJydH1v1IPqDFGbfOWhLRGM+aVaeL7VcM3hozm
YNzF4JIIZAt7K7EfTfrcJo0v2inn+jvWtvheaSIM6fYWBbhHV+xMzdcCObA7elwC
oa6K+oIm1ucB+f4cWYJuJveIdvvS5wJ0Ju2zLOdVlC+KuJTJvfSdG8PEGW+Ic5UQ
xXnsaDVfJO43MQKO7EhLagqAbcSc9S2UbYU2xTe7ddApOWVgHZ+J1GSsErUuwgAk
OmoaULI+jH5nQcAz2v9kPPcfD4hbS6+jQ0EPxvirhcgtMDMQULKjXKzl6e/BA3oo
65ePErXG6fd1b61E9CAktekDUz4z03dfe4wt3YQE6vsCdYfR67v2rNh9MD5W42aQ
TTwV+LdpGhlQ1uDyf/mldOGZWNXiptghY4u6uQquIAqXhYdzByb+MPwdThMiw4gd
Wgdp6auxNR06r43AqK949PRuNZOwPw2uWu0l4t9Oe2pu3GbEDCEFNGBV80C5TMaq
OD17gEDw0RV/OPPzFgalmgUkzuY6aexH/RZyUVGXXYZ9vYN85IsgNWOji+70eNIN
05vxMUOs+AktVNiPIAk2SvjxOEd+/F7b2BdRoSCcIdO337ZvHLkquWLbgua58Esl
vZtF3n0Z7QqhJ8UptJa6aidJaPGgzEiqboTpPCHrp1ndxuxKm5kJPY2GDoaYlRjx
iyCBK5FX3phjyjuAkOkNntx5zOaKgAF86SOfr50bfCzAFZuUErFiV64rXSPtXRhV
Z/R/ZKRDHXU9+uDCVwY2LjjhR48hM7YO60CPNQoo/fIMKnsbntIQF0QII7MnJNF7
/U87jQaS8sJpCcPyEBFwoNEZHI3bnnM/9ZOPi+56oeQrYWByJ3/w8zKutg241yYj
/nspQw9kJgssmnnlNgxyAz47YNFnlyKs0rKnPsC4eFHGG/1+MZsnVgW8DxPXUHtN
MaZZGnk58yOLsOEb0cijTq87f1NbLGNJ4AfqAr+s6t3eJGVyANma8KF8txK99zyp
GqGR5kD9jo2Gbr7FXLUfTvXXgCSOuJ+jq+BQniHE6T3s1oJvPwUCkKs5Dhd9MsA0
J0Tryohzq/S2JEK3EPrzS6yxsl82cuTACs+x+hTdIVdUdL0D6aErcwlqT5QOwczk
T3kkuWx32Li2nkY+UOAJaf7s27z+pFklXMx9oo+1x1GcRyXxxkTMc67S+6AUS+m/
CND4vQt+eUuE+n2hINKZD7SE4nxLdlSoB6BHvPjnAf03uaX1hv3D3WbhWr08X8TH
hnVCa+O11j9sQn9f3gnQGWgYcTjvPWFHZV0HUJFJRdN3kfR9pFw0S9r5cZtwF4fd
XhvqwifSVcYSfgeMFNJ2oxtoJ+OZZhmUWQ2Tk9zuPYVqq6lTZylU3iFElSZHOfXd
Vf7c+nLvLBN8XexEfFGUnTB7Q7rY0Fn9+spu4NMKS8q/2qynT3mCTopfPAV4UNsA
tMIOpEDkGsJ9zIhxSCn7YaMZyXNE6Cs6Pp3M966vgbiGZHxp8563jS18SdKxr3Ew
ZT0ki+w1Ml+8CAD1XY4zXQcGkWETsg+eStqUvb6DW9JwVs7aoFDbx7yDsTjwYWO6
wZiyTwcr38OANXGcG6ffAEVs2rc5u0LmmeATjPoz5ZOW4IPtaSCT2Lt5dTw0wGLW
SV1ZFyyY1E7loxwUIYVCRF9+xoNpjGLx+hYZf7FL5mQbjivWJprbYMVZ40fCMEBH
U9RNOaWS+sNIZBu3yi8mafmoN8z+0Num30B+ZOB6eToIhBMrwEcPwpeUjNw3hY5/
pP1h3Y0R1oS93Le3n8ojRkvtaFheDTRQBLZDxq4pYFp/RYUqe7hZFvfLd+oDwFwX
bEyxxLZXuoqKSDl4IlheFn7iotyauCCsyvf7xyTtSw7wcHR633oIu5yqPUTxfU42
lAPsbBJvjy8mHYwXM/mcSWuLXepyclNy5qP1zazL40Ztnjv9hdSt6z/meVytNJZm
ZFmRehAWjW15J2s+Z4YVQm3xaHQ8CtvZwYCwqAKss8naYDKvbxcsXSbEtyDqJ7cO
xso7TydufFgRF0bR5HMg2XzCu4RDon1oRaONjgJ8LNjgQztsc4hmQiyONuLQDVmG
Eqz6EMElFj2s7Zvs0RbTBlEsnMBSfsCgKeGDm6eeBZHOrVsX49VQ7qvgdO/4J2ef
c8MqpKsZ5mEPb+yKDGkfdf+Gm3OrpgdnVSptzw7gxGVp2gXS/5lcUC5m9GANK6LM
pm1mXSyKILG3bSlz4pgGC/GMmDgDH+CkbuHLj8Z5/cnVBELCX6JsC8YGnr9Nh/FP
klePgAjcHsLHYMASmAVvKwg4pAUzE5Yx8Wos6vF2di8opkBno9Tpa2mVmG373LHh
KTOPbefvbEL0IFgLU3bo6okexKyXGHT12/nAKoAz8ivzFfCRW6WKy5xqK9G06vG3
YTyjhj4XtsxYdrspp7EpXQtIE2+pgKR4RlWUaNFWozenJuR9CQqxyOCVo805Nntz
9FC1DUufdo7axFehNco64/L0r3cTMDaT6rrcQ/rJn/Y5NfGcGw/+V1SVNSt5ARyq
rmwV84Q0fVuXfZO69+5Sz+n77iVNK9Oc8wuS5SXl6O6Edh2F4dT4sgAcitDU/iTg
fXR5WGIrsuBrlZ9Q6HhOjBd2ChH9haBjiMM2/d67czXey01n9RSMkBlS14cfwe9r
CFQIymL1Rt5iqd66RyVDs+b7zQstyQ0zaC5lh4SE9v93FqwnUNTyStLEnlQpsXRh
8NoMtQo09gGTRIfA/JXmgcL1eaig+lJB59N3O2J9DW42hf7foEyRCEJHW+4VywJ7
tQt72IGAg6F/oZTc34+NpfToPdqO+qOjvujpx6FcqqDKnb6XZkleA56pJM5l4+Mq
/kwTBSNM8T9qFei4ieik7gGkFcG9KQwifAnioeHqJlE08+Q5tLTTJt/LSkyaQ2P1
7NSiNV+AJKjG1wRd7XBHOhAEUrDyegayVrGglIm4S+IeU1mxO4Gl5DBI/TrA4L2y
WHF+8ZcvTIr749W45qewR2PUd8Ltear7lWM7Z8pjqrKsmGbMgN0wBTKc8yMlx+Og
H+hBFNgiiq05Yhhxn+wI2GyKiMXR6jf7dmd8OaCHF5bPP6zcKUJ+41frdH6YUGmC
zlsTBp7Zn+u1aYEsGemfhFyemHR/JFNZ7nVJvkun85tuaoKdCO3zUpxIc9Tr84kq
FCMLmeP5xhFJXVSUJyVYNNKT83ancmwIVfPhkZpZyLW9c4IvxA/kpALtVztjB1AG
3eg7whSXjpJgxhHkwwc8eEZQScf0t3nfzXKxNsIne4gj51PMHrlUjNyHsoXYGs4O
8oEuPkt9Kn7xkuwGJGvKAixac+N6GlGfWiX3pRbhQ0tnUTxA7KDzhCCDTw3JxAdB
Z7hOyQQ6PvLcW01l6hb7Jdv5+l9jmT3iLcJzh+m4HCHwlbNxX9R0+dSz3C0bgCkY
K6Ou3mV0Lg9Z3zeUbdHoSTLUEVvM9uVoLf9IKaqGn9+hqTbbtHvmZZ088nA/pk6z
Ed9xQeZtsCWWuzSb3HiV1Fop7ujG48r/L32pbVeILNKSDV0D0r24G0ylWAEcXmrz
4uYYJw86se2dg+uVklmba26VqHUZaY4amwEpa0q7rweqZXWoNgyr79CEQ4Lf0Yea
sUNxuBlfOzBwhc7v+g+IhjbUZYOF/PB0xEr7dGjGdhed/61dXT+l/d1s8eALZzKP
u4x0pj2TkG9BiFeZ0A/oSIoOlbDrOXRsexyPVfTfpqQazjpEqLqN0tO46NfejPW2
Y3OCdtvoPJ6UlP9IcIs3dRJjsz+d2W40/GvFvBl1mEbyeV0DCZz6tbfd5xdqEGa0
v3nLoHspJStu9NPkaQ7npzRHZLYrSFKet9tLZoNlSErSmNvR1WaXJYws3Dom6zCg
aRKuArErG86q+XWt/Ic/lb1u8n3dtxb53IUn3IpSGNYE5oV8u5/ZccNPEaItoGM8
utiTFIqHCM0VenQb1HyZL05mPMQo5K4CEd92JGq8OGktqkPW1ZoPEM58uxKl6dKl
ZCjErX6SJU/wqHu3LK/qYOm+Sm2XDd2RQbA4vtsXCJ1w8v3VrOb/Ar4inIAutSxc
pRhPtqrAM0cs7zbTsZNfrAgWKWp8+5hmjE3b1h/G+C/RmSBlIGiWBl+/U58rSYHq
IofM3CPSDhl1hZDBEcxdUkpRFhGscJ4eXWscrnOyqp3K0TbgrPiZ0iPBotllOhrL
peOvCGdheCf6/3AqC2DSHm2TMgRv7uRzLTXcXNuZPJMxoEOTI+ECXJukHyZrgIXb
FC54/LMUXrLVO/yPHOs1S0uRB71L1DLdML0P40Sl5z648mqtO6YL6g/D2AXfrzg1
TzxGFQSMSIyjRFmPrBvyWkYeyhx3ksWtztxJ1RIjrRAcuE67bjnKJT8WwJ+wrJ5Z
QPXb2tE9PvI9bPvAvxHnbrvEvLgXkDuVvQ/P9I/URrhfch/draKqFmUZxQosMD0s
JJBXtXshr+2s1dUJW6PZHbKneyvPNzHRRqiQ0voVMbXt2ItwVhULNBWjAmLOYUdI
jieN5Q6LDq6X1GBh1XnV7y+CZ6DTpVKcbHUoRZp3ByeAXp4blNWHjPMpEqrpX9QH
W1kqj5LdpyHKSO+m1Vj2RLT7FovnEfyjrSER1J0pOu1dZFPXcN80HcV1eVWZsvp7
nXhgRShmwUvxdilKcVd7qgXaEqGnd1oLIT3z4Q8S+OxCoihhtJn2vepT4GH+AjeG
MSK2czAxU+iddcbehwAsxjf2JybjXVbAX7tspSg3cA2g/jfEql35IAn5DgsoWtOI
J08sx8cJ5TWEENSwyplUNQ6Wkv822SzQg6nMEeMDobdJnUp5JHc3gFL+hWjb7OhZ
PAlawk6wY7LhdDn0EbSBwLxySKD+8Vb5DuarINo9kOYC3S7lIASP0ws67hf47H/N
YXnknUz2eeNCCj0f/CwT2cYJ5bDMHiIadx1B6tLex3+bfqGenHu40PYe1GvJ/Cik
/4XatAt83z/aEWHjk6qBZOYdot84ckmG0m8xdaN4odYqRdCrrnsBJEazY6HXUXc8
qeshzO6p7K162a2CU14+jRr7nagMFpU5KjG1L+1XDbkWl3n1VWc7x0HMCl+Owt6t
7HfTzm9knKgFudZfvSPqONH8MXGWeFHe0tr6hwgRrvIXssdd2dSzyQaAzAzEjQvG
kwYT5vqA+Aq9i9fG2SOqjccw+orFwtz5ji6GOhy3DMdeB3waESCqyB/oyed42L4u
m9gbWEMpZvrVoyRvohkBmH76G+H8+oStX9wrbkvhH1mZlDX81CpyqoY+qNuMPKuo
a6GQdGlwh2pt5LKnpBXAIi+DT8VPp4puOgCU08sIc5wAxCBT6SYJBffxy+JEA9Sn
+FssnkKcZGZUMQ1rU28c1GxoLLNsUnGbAJM7JtkK/huoRjGGFSnjBEwkmJiZV21y
k84CkCIN+w/OGpPRUMwlz0WaRERiWAOhWlw5nlMEQ63fcYHl8cz340NG4g9c5I1F
YI/1kOIfnLoxQq1MzrhBJnbZqYa4XRbHcfh2jgGjMA6KerjfHfQsp7WrmlQD7B6p
ENXTmvedsaSBfWCvHYBYWZ2LUC84tpGbTvdRXaqzuHDFC7VyfRJVBd7mHwf5pAlF
2n/e2tDjoM1t5OiZMNMx/BJBPCgzMJWHOkx1COzn5ccvotq2Alzyw0LEK1ZDVpnA
26UX1AH6I0aoTr2aojClKAXOcnrF+02gepDp/h6vo9rHr1h4M7mh53nxYCdcUO9D
n+jk0WLCH8rEHa+7Yz6y10Tm5yc/tE3utncEA6zF+p5MlAQehCb409OMu3XJINXu
qvJaYhvWWpMxUOgd7QpVtgHnQy2QEr6kiQZHGYNWvt52pPZmkHmbjnEUwPIdasrr
asgF0122ZEE5HzU2MJDaEZCY+e3NdAJAN2HzNJBMfMg6ben2g7lO6LNQeoRD3XK0
cCaVIsSNKpqs7fmPrz4prZo8+q0wV0KaNr+Sf7D6+a2SOmKjPOoNUHjC0ccpkx+7
nuxNDC2qxLCgONL+Bf02UT5R7Zp7Osj4rhSVSv2cu9iNTV+4jtyOxUPq4tFfs7Ai
emxVKg4rt0IexeUBNxzYHYazNul+NMM/zOOc9ja5sKpcKT0Aan/VH+d/WRw3KId5
aKXrhmtMCGhG3I8t4gUZ5TmtHmNyip5S8kWgWO1VRns6vEMpCapBdjgfd8FWxrom
KYwTyEdaaJ480FGwj3+ybCR0S2oLHzlSzWEaA8112dnO8tp/M7ejV2CYp+e0BuRf
plUZvmPwy39RM6fddXJic4B1g9hyAHyqmiT1viLTfP4FjlFV+LZworvOB2OPEp3v
OMTI7ibhZqScmpG5fTR3o6JsLE4R+G2SgfosJ94YSk9+15iQhftYoirFxzlNqR0G
yBmw019PA+QyG6A3mKnkhJ7FF0zaQ8Kjcf11bCG7rOcEH93eYzdtZJ1JxJcdNVOz
om+2ioma+MpPJYuAgojK0tQL4II1IODQN+zheKsCaHwIaOQftwH1xnaU+/RPrq9E
D92cz8tRd7pgsqchmADXxGy1yl5SXgPsWTWHD4F9023arsIm2QD15Csm7VFvReAy
BIubtWaOuAIbdm7HYhyyB8K2ZfF3LgWD5nKtZzRHkHLD734DuNkd2CyGEg6TIN+4
7NMXZLXL9eNCyuFIDUTGxUHl0H2rzdknRWyXUBXZCw5hfTHQaw5C1wIm/LiRhUjY
l3AVuz7rC1Zvrc5I1abJ2vRWWwKg3NLbPWmJaM+BjoB0ssKBE96lHDug1zxRrHRf
HTO4bZHPYfapnbfMsEMgTQoAmFuXYzD1onHb/HGIRKpBq90zSW2iFjbz+yolkhtk
o4mLbuGk2qa+VMw7yAKWf9oUg9bwVl/qvuFLi+Qi3eVcwynAr7vu6xlRb1rHUZlz
HiEa+GP29hG2bVsjEX1ulgMMYo7TXLPxdVL+GL8O9w6iEpIU3eHHxcBk5i5ZaN1I
FxuTI+DO+bBI0KX6UtEf2XLStVoQQg7TFRTI4pCMVNHI2JkbwTrZwouZy0IWmkSL
58iLjCTsW+OpfDD7ojoaNjH/qFNtxJqIzMJ6Fvm/V48BX6Y+0g9vc27a9cp/SOlm
/OyTP133hIShq2LwVRv5dcUAg6PiCps1SMKH2X1kakD598fM3FgtJKhCv0xLXj+N
J0lGH+elmdULY7UglsyYxvOElo4Ihw3bO/T9ZWL/Izdy0JF2jlH+rpPdiSvfM2Bd
gep3xk8y/KfBVW6omO9LZRxLihQHGpeoP/u9OlSa0ANlq/f7vhOO+C4m428U3SWo
2TfjF5klLIXQyTYYsXkslVxHmfHYR/3VRUJ7TrDnHcZ1XRuzzYIi0gOQz5l0LE29
EdCLuLWvd6qmdUr2gtfBmvF7Rn0m0pyNc1A9xnNldrXdTwGdeyx3p9bq4EEFPjuv
F5VMA8ncI7WLr2aZHaJBFs4FD20l0NdaX6Y1NgXO4OZWT+z4rtEiAhm3+9vNDm9D
VnTgTVZjnaLc6OCO3UnR+oBHXnAs95LTN/8v1radN4j0Pg7+Lyh9iEdVvrKW/W92
XA4LOHIvPj1l7oDhwo3qx59NRmc/vxsgYspg1mjgME3cXtz69i6kPASTNpXxezhe
cSAkEnS9gjGICEvDfquLQp3Ubd81bOlYko1mh0t36rwoz7WXmzxaz7T5WYbpCYki
kWvOK4yAEaZZu09R92QBWgZtGddTyb4R8Fw6yIlxC8rxvuxDCj5LxJMpcV41npSr
5HBD04I/vyVatUl8JQWossuInD5FNtPU5KbmS4PaF4aw6vyztDu/RtpkdkkiovhK
C9qaWnRdOb7WAIy/FvOoi9NJr0fjsJeqLUH0XyEE61wGVthpvNtdUXB8z70/Bwby
NTkC5ecwNUPYtcWQRt12KCtAje1TpTRLF3l/91YM/ZjIQx65nJNNAIrJ1fOIpeCJ
0aA+pQ+R1kBLyPUg/JVcPdsZIigEk9imkJSlXGoGKEOzuph+t0oUUX78mhV6MtFL
vF10BXbAk60rXz/2xL4+XHZ0sHuxSdWdT3OxnsJcDB6KkejvSuNhB86DbyMFPmYQ
orcrOo4xCPEVwLBFcO3dOyB+LGOhFm42ZKAdYMBIoaPtWV0XvE0HKdfTREA+vGze
vMngGG2ZlGmtLL8YBZuEwQNyRy2ry8Bp0OtFpxrFKVb5RIrFpa3F29fsR8ZPYmDr
MSQ7VoCgNsdCKOyi+pptUm8d5SPFCE4MibfcDP+pyaVGoGdnYUEl99U06yY9LXqb
O9oI8FCpZBm7qO1sNWb5wsmEKwx0do0GeR+s5rEbhGoDJ3wbTh9u/SezmnE46abz
fWM4gx2w2WaCJ5FukkS8FmPEWcqlm+YsHurXLuslVHur9ZbEQcONJj8VRLFq694d
O0xFHxEA/fkeYYgiFCSpFqu+3KqxcVlqorrWkvbEq1hXbjSOO1t5PHJeamJFIAvm
YPEM+ezn5EhvmfWfmPjhEbz3n9edTWK8nJ9X1IyIjpr2XY+k4EJvXn0VxBdrHZ+J
0Yy9yVJ9dOPpRjFCDeK7HnjpHMryiwo2jyXrvE9+wCTQQ/H8hNWnV5G1dzCcXwv6
BTyLVF9TaN0/YdhBT1JQS7sm4l5z0uLopzvW8koFTrrHqEc22HHHKRSftBwMEIKZ
OjrLFrfRhvsLpRYBZ/yf2rkMl1ty7dTL//XcXB7JYLfk7mw6V+7cHDOh831dLbbE
qATCcRuQqikCPDXC51UH7iImHOaLbRUw92UdIToVAlNjP0YTYxi9rD7v5aJ+kIYJ
64o1d5wjGdqUz+6iS96f4eYEr3lUfZi2gLqBGZ8kJPaWT285KH61O7a/bf7LvYSR
iJlxMv3qprnFJ5ncO40AkXRMg01qY/d9sCUGDeQ78DagzIrp78mcIvn0QfUTB2T8
pgJhJot5d7Bu29nidApHsrtgtf5W1JGCdAEnJYhpbEdAbKOdbI3SE9qUPzlMjBba
CTukYKp5tbxg4GhfFb5FLXRhAIhbRkakE21Cglg39Q3gnLJ/oUTeGWcnzy/kNvJ/
30ZvWT6woO+dXiVLXqVk86eYF1hyEAPfTVfwiI1uTAY0bTroV9COQT48KDjmsAaW
pEG6ztvHoI5hL5JUIFwMnfK3T3NP/Uw82EvUwLiH+M+dmaOxg2aRJO7Xw+JPF2gC
MpsolvRPe7LfE1/onZVUrZD8sqEoUfj9Vg/+GQCQNjAyie1G+q+lQoeoQntdfQot
hwIyqVpVtOPBjKjGAbCX6Br+qMRrYjNnpc/vm5JPMpzycOkdEtglO6X6Lhcta0qJ
AkUQ4DvvITnzSwAyDEfK7CNZzy2HOm0M/tF9uFQqQ2sFwtjjMvmjM5w/6HqVCe8L
sn5oxPXsd+nmRVk2dkqAi46GFKTCp9SpcepxuzT7ICBNxk8nalyW0aNRXBjQaZeL
dSXK7mVM76SchvvcpuHaZSt83Wls6GVwIMXokQsVFMGCrG7BjI2/LLFMoAf10D1s
nby72Rq7ytOVA9ZO6Osv5F6iLP/Yr2VaCIXtqbx58DZL3YqqZrFrAawZr2uDT9+y
eLafllB408YNUtzbZBmx5TQYkrdTKks/2L5bRR0QGmpHPMNFlbIXWaykgidT1mE2
ZsXP0qa6ju2dc+MEn0mfuYHbGyH5TWhWPEH0wBoUJOtIeV4fBMfxZznxInN2wCqQ
yhA9j1PeiQu6ghwpD2J5bmf7f7s9tXt0pvVgCrFZRSy9zwqOliFL3zyRAKj6gnG2
ikYMiyvXrjyLunXxoB1gDzExjzEds9/Gv3eP1axB2+zhopmpqU9eyZZgPqTL8GMA
vkpEtLJZDhiVOuPhPMNyyO+k5luWuvaAmDPm0woRJOi/ISqkF1BlxyOw5+SV8rJX
ih7Z5zxpp7ZkSd7ealS79pcS99cv8+4L3zELy+gO/oJdFajo9BmVUwOTowqyB1aM
FLAawB6o89ietyrItsWiw2sMyriVmdMbqEbFWgsx2nZJeU8Nk9N1c/KclNKGU0YL
OLb4T8jkkC2GDYgetttcK2DaDYNpNWiY+JlnXQDzmWxCWXAQjvPNZmuPngZBGeTm
eNsZXZxvM76IWoRscaruna3RNVEkXMS0fhkYxG5Ezux/kQ17GP98EdK0yeogzZzu
Ojdwz0bbAdEq3IT3x6SHkaGN4yhz1djLwfUeoZdTXCSzmh1Qfs0K/ZTESpQXa0sp
IjPS45+nO+WpY5hcAU09LyvUX/tI2gwlks0wSucEKB9kEFnNELI+aZ0buFYczXjU
iTQxqPHG+sRDYfxUGtzBFTSRBsUUXKcqSYDwGP6eUZkchXOrDrI7nWeW5voth+qk
h76yQqNn7xVMC8+1ZM/44DIR2KBU7wTcLB63FdVqrM7y/n8iTSGrecL9Rc2/mcgu
AAliIKDiM/YD7na5E6gqfkZ/bymVqs8Anyhm7vMqjiVAR0Ew82aUyKIGmRVqb8iX
D3/yuJb2pb9lSNQiHOAY2pKAl4Pmy8OtWtH9gY30B9S6CnFTuaDlGTDM5/Ue13zk
RZG9vS4sMO/nUdduf0Y8tf8CYO1YZDosATDWnXyFC94b+dsNmKXLnkgAT6TqDmFa
EgPOHc+tZhogeVQN9UmIxH1/zejDLnPUTkDJaJkBBDR2EW7G34EMf2+rElBPNpss
CpuInUzOhttVaXg3W5AS6iFBMMDLzyKsBBPl80LPEUVdoaHHcJ1JSq29HsV8+3Ja
7ZmcnN0lxruVM4KImMW808oPRaN30poH43mfG1cZZU3zkGAZ+M1JIcs/q2pSYCI+
vDVyG8f2Ckmbg7db5qT7BRHkVDVWWhKHyNuu1ndwEcexDr9qUdBwcmVHecS6LTJb
ebfEx603Rz1lfMn8R1kRQp0SL1Zd0f0oJex68xdDAp1POsnsiNO7zwsZs3fT8HJF
3KnBuGSFtU+nXkXFNniDOia4iDIYc4m/dhBp7TmpOEMCfL+GfgnWLsmqxuHnvT8V
hukFH4HGSTVV0XFVWNMIUhdcdAQMsqW/oPTrllFr3dp0eTG5bIN+/UzwHzpwgXMB
ReH9LjcUK4k8HKErL+uePEp5ToAjmuYikQ1tKDoA1T4JOV6MykpD1ASNEZ8BSrdA
H0VbBGoHr9Ps/Q+vgQlbChXnntM4SIsCp+UmEHo8uuTSaN2AtcHV/2iujdgP6uzl
+zIbT5ebOYJy8DSmOJRBngg6sA3ptoNE/VjNIxIYZCqzpGDr9WjSsYoYqx96J69k
J2A9sINEXrF6clxB16NOODUXREyW48jhHeq7m81KFuluKQFe3Oy7syJKIjK7QIWi
9o3kEPwf3SyHdTuatSiY3VouAjAddHsUctX7xyTYlIvJDDStWHPidnZDvERga0Gz
xp45B+WKSpAkCjsCPm+WEivtQtj9Kqe/FqkRJLfFtBt+0awCrgvpB6HUNTLlYAzE
zgMmvi0Nu8Lzvov1zzMBU6i/rT75ArYLCqVOQGZL1Zv79GBcz5LUkAiQ1ALLm1IK
5QwifTXHkITsBTkqJ91rGXsGYX99KGaEWcoCbK0TjHArTk7JBeF37L1sNzCoe7ep
+SuJIuz2z89mqpn61Y0th+hbXXLf8PM2i3YnfSEFtYdqVRYPe4bKAh/CuxOCyyLk
NkdukZeoSUG7CX4uQFPxNT+OLtFMQvV4dfTOdF0geQSrloD5MPOCKCwqhtOFcPDx
1iGSsPCkGEdM3iE6/M7HnUt6/PaLkkkzJQuVJLcx/ZC77hH3p/EgKXirUW1psbPe
4z392HuJNiCrE5O7ib0TV+4ZudUTRog4RZi4Zj3YzjSRPCl6cxZBsgM3z2qSwGAW
sUwNFnhPSglcAaw7Zhj+FwgpBfWwDDEKNEPUBiIbq5hVvh/Y5ggihFM37DKcMUIP
rHybvWfPLsOlFg4THinHf/2eJQRnSD1hZHG/kx5mkih7AEL7TzdqVuRwajXdWcDF
Y1wMWhr067YX7JMh54pFrxeZv6gex2ACs0tch5+fqUBd7LspWuwwQYfSjK1Lc3dx
jx4sGolTMACkAAt2quI2nxfphwkTryW4Ci3NP6cRwOkbeGAZMSyt03EP6KZjObNp
Q5VCYmJe56IFKi0X6LTR/tgr/6Oox05tztlZ2dye/Riu2pa1mXUi4z3LegU/cVAy
5mzai1xBNpqIJativ1dSV6t4iezHjbdOPPTSezgRLQpXKe3ESzWtWBB4DIRETwPG
99+t9gtDy+9eqsC+Ud8Yew45AJh4nrSk48ivB0RuCyUINma7+ULbgkmivfI1skmp
6rec/vhLe8gy48bicRl+g+/f/+0VR2cOfCsDnVuzSRboiB0mqIhlwF21+0+J/EH3
M6FwBmq1gWvjDGIfohS8Ie15q6VsnE4ImyPvQydNcNrSFpdW+G/GReZW3TN/imy4
8yfFe82Nk0B16Z+V/SOIi3CNiyTDV8FVYM7yxIDc8c/TxRrLZ4C35tPjBRcszGAS
04KdB9AwWW2UmWFB7j64L5oGObacztXLhFdWbWDGA49h99zyKl/zci0ErVn+nVpg
cqtjPrQ7dFqxuf/z3rb3t0Ug+nsKB++RwhmtQZk28GEBYCY+FULVYunvbgFTmcY6
L5+GD8FkuT60ktfvN/1rApwURwaiTbQTXr/2iKQlRsO3S25ZL4oHzw80UDD1A5Xf
039rhxPGOn6GpSjnA9JqQTFGbAZecMsmdrvjqPB7FMbX2HPET5/THJBvmnSO095n
EW/9PbUNVW0F3mq7qEQQmoAWzhWzRKdYm5es/BgUlrjD27dXK9kR6skbK60H+9+P
jm1wIQNoj0wC/0wtZo8YAfRDo6kHTb3Pz88NPntpDKG44evdhFMA9ZxfbaPFx866
hkcQ6xT7vQ5RCf9K3dApsoEGM3REtFtE6sWzP4HiTkPnTxoEZwMcY5/ZK/POMi78
BwdctHMA/emqej8S0wAe9nTpUz4Uz7/f3/qR5xztGMhLG28X4xzW3dk30/PnsZzd
jG6kiar7ZYvhbcEA6SyKJ516qUcWQypQBos2/EmqryF3uiBOXkqEKUmKURCZy2mc
+sN9Ja/f46eaU2tCf17gWND4U4Dv/7SE7sRduHwAalYsxSf8LgiPFiUxxfqcyzvf
sYn0eL5ocEAR8bPSEt4S5KWHnpX8aN7yofxPH4C1bsbGGVFGckevkKeQlt1TESTT
ZoqL0m3bZ3ZkHdkV8q/aXTQlIuHV9DWJiiqTZlkfLs1CXabybexGUiQTNMOmfIVx
XDv/cd5wKrgxMr3S92yVzbUFBi3vAM98+BorXL/MesRx9FZxWBnk6YlHw4F2FvIo
6aAdQ52r/DRkPofYAOlBVwtG8QgAAbbfFVnTVKIrANYb8pIfvCi+TgtGBGLfW6rK
GSg5uzzMBfjtw9Kbo1L+m9eMMqyWDVYDRsTAXYox7bVZcDmn2xoupzORoK2ZH8j8
D5g5k6gio68ZWrBTrlOHBKEjq4o8+ilO/pVFB5x1GzqYWZ93Htkaj/EJYbmPJus3
SYlP8sDTsVvRhHJjM2mlkQwnIyZxkhQG1a+yGYXWveQUDl03DxUIXE4jO5cBIxtY
V1DY0BFiFlbg+jyv/qGpStre4BUb/UkUkv4g6XppxM7a2pRrzwkzXNnAupx35JsR
7QmJpmtLSj32ruqua3VT8BCIrCwPZw3dd3/v7ViR72W3aN0yclrToaB2sjw2Uhkj
nIpMqZ5QIqmkH24YR9nZxrzIeHWzo9EkSdTCaohuXpZjAGYfBwXbxUkRFN36/0GG
mRYokyLAkBW5xX+soONICcuunEjq7BnEKNbxFgteGMjo9gyX8UKVv3WdY4geo2Wx
kGSgiNcLTcA6Gvy+JkU7+SpXTO5QPmklxcMj2dAyzDHRvhTHYFObzxoVd3dLdXZF
c53ZmDo57KL/tVY5YBPbqoYjCaDQx34W63bz9ozoOwZoKGoqf4ZBpWEJvThW65GZ
kSuRhCy5XcVCqWObSKHMRnnrlQ5QoLx2xfOEMi0XLdUKtSY1PKg7bl+yXV27bBoS
4Yi08cxq4dp9INZQ/7pzbzO+VGPMqLyMsWqN13OClqZmp6nJOgiehUIk2seK1Etj
BadvTXH5cf824Bam5JlrAZWD2U9cc4jLloSuTEIycz7Lgyn5JZrcSFoVlMGTQUSE
6otvCkUJt7IUEm9RRS5CqvX9g+PMKwZG+wMzuBeXcWw8LhAMfuP0HliXXSO5+dmP
x0Cf1PCsRpxIj89oVpKRji4stZm17ZT3SwsHRzvUdDbf8kouYOVYShHEZ+EsFJj2
QM+S3bL6w79kfkVTW0n6CoV48KhdhZZAmCN5O27Swx0LqohomQw+wA5osVaL3z8n
B7zUlqmtgtpwd8bjujgShaRmD4o2hISqTNKRG9uC7coutpPHdDf6/L5MoY5G21xP
841a/RmXH7nKdWtPdIIwIkS4i+VgKO9KwN/EqRIsdRKCAyVKWQpSJ2uSLFZwNtrg
R6yQVzzcy7ZNVBs1LkX6FgO3r2CrV5FECN96nnx1LiAoskdHQlEsB4ikIKt2OlvV
pzC0cC2CB9B4zzjz4IKQA0QA9rWKmlWCJBLdaUVNRTjKWB6hs2xk+XiP99T6TfP+
wx0QudnjJaYbqy12WtXLrQKyRuB+iZID1CYgx+5v7T8Isc+dnX3rEPpqKgcKxqnS
ABUEEnXdZK6g/NjvJsUkGELC3AeGiOFjBWos+jhGvm7HAPhQMZPRazXOmQxUanui
8qvsGfqRYMu1YvZViDPB0fgLqOYdsdEH5PyGtO+OSRkPJuv4C3EFQzTIhqOrztqR
94qDDe8JWk+zFmP8+H2wQJhQu7Hvud2+83EyDrJ5Ypg2GBqsPfLxPuqKu9zXq0Bv
pbN0FW8s3N9XapAyp9qYrpSmCcrED19mGOCPZu4HzOD/0f2qyLjvyb1KK4EPHabE
WaN1/+lUsYPEQO0m1LSqU+wL1qQOJYfCg45e2SjvJwaruv+fIqQToGwQN1OoD5ZF
C/b4ZfLNPjGDiMQjoDv6H8QkaP46aSl72jtvgoZjohBtdG2L2sJY7kcNe8L9DYWy
qQM6aZWCnutZADHCZLoO4dZkQsnGtO/4vTN8qD0PXhHPF8NsMCCV5Po9hSEidOGG
oDlUb3m2vaoKIuHjT9GAvlNB3RtBJEHndcFRTZm2uigjNJFPPr1fG1OHn7MHQm6J
cDaDriLlD37lwiZJVLURtTkkV0rYnoJu7iK6a8a1d16gmTjWdKnRGcq2HqZp9ryT
/lwfFjWfFpl/rgBzrLxhei5Rf/0GKC4BKh+/1I5dz5req1G6GEVbCqsmCjP9f9+c
s44aRjZuK4wkYOVDDBwkzXC1LMRYxncjgFOJo75e2pFTGb5OmQyYqs3OYo1eAhfz
01A0IKJj5ZAn3IzXe+W9xF5TqJ4f52brwrf9/vZn7Wy0Iq9qmN9WnpgR/Nuv4UB4
kws+lyg0+l4UdY0W0lq0xwRCl6WDH976H/BYIVPSdgnJmcbmUWCKgjqg2ytKzFKm
+AET1A7m8hu/EV7xwcDAgINMSACDmDe6ZnFZNEU8CGfWcJ9mHJ5YSh0dPHdDa22d
X7koCu/5KUULxDGpBxX3td5bMtJWYYv8Pv97tPOrcjgOnTAdtZiDR6X3/wwcitlY
UzxGyAxI+l2hYIirF8duy4C7taYOZGYh56KfZVdnbWFHlEUoHnD3uSvPr7d7Iklq
qkRADzS+VuZce001Fam+3sA6P9L9sb6ZGizhDmlSpT6mGmfpt6qtJ9DTEO5uPiKa
IGtONDkcpTPRiKAnlOXyzbyk6IfXOqWcE/awuIGiOErkbcuDEDxz72XLuYdvrLd2
ECx6uSB2olSIBTMirnz2v2qOQnPAHojWuIgL79PTGB6sA2X1yOlHBsTE8+SCFGzo
7EgM3+CLa4ReZUgH7U7DoGkovhY7SqhqlABaIQT/cY0tF6bXcIS+QDCHuwij3ee2
j6HiJ8c4GaDI5b51LhWr5NugcJAq7RgMoS+iDVOkK5lyrVnlRowlhEsZgirWKPY8
wY0M5sOlz9tJjuK6tC2lOyvt0/dj1iAr7Uo/Nn4mo8S5xJNez4Ri/7/MBr7yRBll
5OnUNQd9dbnHz7iRlvG/mHo2NEU3giljJ/98OhB0K4sfq9PlThqBAss0CN7gYXHV
80hU64zcs1nLX2qJC4VCUnhNEVyFa2vX++GF04InqQP8fI22bTHihrcKWeMIHdtE
e4iw3fM7xpHJzEyndB7Qm2jp59SM6OQU0lKhlaXqt9IGLN1/QhHER0sGk98MMlby
7q6YUFbAGAmXCDKc0OzYfyAAI/whPupVM8zM8ust3g6TrNCc6MoxcV37JBukVYrF
AaMJCIDL49edI+WMFk00Ttoeeb/xdvN+DH1RAFwVdmfSSEFCXRCxBwrn5zwND3c0
6KuXIQX0BPj/x7p/5bIwSbziKdF4oQQjlt6GNtgjIacXOFRn0U2jaPi6ZE56BwyP
OfKzb0LXshLgDLyKgpb15d0ipt20yr+kxhhwIyLh1HxyY/ZlK3y+DtklefjGjGLu
5ZGRnxyVzC9hebluseHfp7Xdky9gq0m4kGOJEmiKueoFXdYxn1oc4eOVNlDgvN5F
GITPmj05AzGFiV3Us4SVDjBW7ixXjAZBeDxt/7lyrpZuGrD/nbOr7vdh5583z53l
K7TMbTajA31jeUJO8sk+WS1NpW+g+NW0jI9FXAdR2H0YQyEFGPF1uvX7UVSZpL4O
dNg5vatsV1LKESGmuwpRCi2jGIU+onnaBpYyXXA9EC5SUAKK6wg1psEZ0g3N2mc5
t1wuHfAqW6UjYwB2XzafipMbCJZd247tNtEkf/A97XKrQPwydiztu2AEkvPK4JGC
nXP8Hyeszi0rWkN/KnDOejjKK7h3wJxtS9dhZmMB4ubl2oGLF0glywaCfsTHPKkI
s32qn1Pjj+0evaiuuVwbXjXRwJ22hyhhhCTJ3fgEeLWD3a0ULSot55TS8md6G9Rn
Z7z/E3Yqg1OrXlYCL+zi8j269/W+XKBpVPnze5i9BseQRXrjHCJ2Y6MEgs4gIZNS
soSnmI52tYvNyh3kmjud8W3iUGokFSYYynVxN5wI4jpLCWw5WTcb7uF1QNXWmb9d
JopcDjqSWl6pqaw/g27/E9LjuGWDAD+DfU3j/C9YLB8iW3cn51PaAbC3E4w1u3Vm
SssuSXTTR/lCFfjGdizvddo+wCq42bbSHKQKYji9VNwajp5O8NMMUGo2y0cejM1D
ZcFwmkbahD/7dqxS9IardnPKCH08LzEiMoxmn5Krl+gCXY6M4Qhz3ue8/wRdSQWf
7ZGlF5q1tvSD6gxGXJfCu4Hq71mNFo0q5FSAYfMjPqQ1a5wkQeTzb+eGZF+LE5gw
+bi9Zwgyz94oAffll+4jVh87DYgSs4O5j2d91Y7DrNrcfotrj1Hn2IB6K/HC1Yn/
FcGCMqswal4fjdcscou8NQ26Jc0EczkbLMVkVmXFbkaS9cY/WJ5mRZ9e3zy9sNJw
nFm/gJs9tFoY6TIHQSdr3F7IntT6yM2pGY2HIxxtuyjZK3HKF6xHPy3IUzp2SVpK
THyRED8mxE4SDoGWSpJ08Tt6gM0QpxSHTkoZZ9o7YqF1O5uXj9ukpQyU+KENu2Gu
fgDq/ZBOXZTTiQu8+97ppgIbbbLWEU7++ohO1GaQoi+TdorVuMPnjXTWPHzFtlrE
ssUB4LeRsPgMc/ov5C1Tvu0XS5dvcdAg/sYVa1SOhwgK4+oL/Lyxy2jiumu0yx4K
CI4iGHN7uBsJGSZYWJotABAOIKAm+dACQan5detbut9iJXYPu6Hs6hbC2Oba31KB
27NMFgWwR4hKDPhE5lEGmVU7Tg+Bci/FOMd/6999vj8KKio2lUDNR416NaDwxbvR
vD2g79nFSNEsHJwvdBorChDICWJbg3GfqEvVtNXRazN3lWhGaWJ4Frgzj0X20Fz1
Ymi/s6y3FhnIh8pdCRCnDr5PIOdvkXRCYJWZ0/QVogWpX78mvwmKIEGgctsdd2Ve
i8RyEJRfQlVvfRWT5EJ1Rovl8rcaZ3zqwL1P9Wiy3aMd1rabAAfxuqVBDDz8aN6+
pdltbxdh4mktitmBo7i4U9WLf8gSI8OeD1Rk6v3pyD5u17SSrBmSgqGSOcPF/J4A
BvFmJrBIu4aY/9QHhPj+xxifSjR49JmpC5+FELOqNtPBeAYsSjieplMtKB0S156L
o25HeCq/3Z5qNq+Cq8Tp4QTJxJe6g226iNTD0+YGeEmMvDUKzEwGB1ij8OVO7YpS
/FqNmw4KEucKhAChBCXRFVsYl34NyXuW2X9skxV5XLY8lCPr4g700N2aPfPz8MoP
jKwm3TdSkJL9vwAf9c5GHwuyl7RFXbKVjY8j5MPSsvU2wGNUBJA675Faej9UZPG8
W7KA3UbNSqOiPZwMbNBScHh/myGWKr/7kIEPEeoipVWsbG05w1qY/iZ6B1QF7Y7c
SZPyCuCR9v7BKhFmoOba3cma4LDMiiboW4S2deBC88FNCLtXbHvTGXrQnuJrTnsX
Os+lM/JSVpNa5E3cffOYXpYqo95n1KibqpClwYsLZoD5yan1277yMQgJXJZda+Nq
n2ZhXxDpq10tcip5WZPdoNwr0vqhvQ5INVI5OGu8S+1uO0TRgVKGeU9645EMQOB+
HEIbN381WO+pRkgnHPv09KTCy9FDQ4Mm46E/+HqdK/tptPzM42KKLWYGx8LGalxc
R02F6qn+tZAFRCmb9kZwEkA6Fns4bgNlZzT/HPKUUBhefRxnBQNZ+JjUn1WSVHVC
b5X3HpQgIf1Fu5dC7qTVt150yQ8A8AjqidZeK4CWfFzz1BGyey5tVF3Usk/hf4E+
rIgC+X4Cb0eruGoBkRlR5TeKEHVmMOwq3/jINDvJ3mwlH9HDgCNCNttH5hVB5wiH
/tTb8IvprU3YWB/OA7QfjXZlKDFPdiYYKrRKi0vH53WBvdXbD7C9obNfi65ImZS8
OKAlxcyfdUjH69LLueWQ/fYHK5zC2letjyqODOU8YNGE5qH+JAzflxo6jR5XzO+L
7a1B8jnwe3KYGyy9QmKtpPBcB24p7tceenUx8uYtwuvC/uZ162MKO3es0+2t0jil
VyoFME8S3dtr14E4WWHVg033T7SuCptGs3Dno1xTv2K15hvzI0WLxT+dkAmE6gKE
31psbRYKVi3VTwgF5hqhI+JzDJCMbv4zvuh+OZ3wY35MPTByeDzmblEpQ6gxlQb5
A7s7WO5b80fnyh+BihJCuyXR2OmbR3fWvrEoIFKWI7Uf6Rou80CAf3epgwJxHPle
M7NwJZTjdwr7swQDBlmu6tn3a2l+OVeKHkZt2LtG6EK+xic2GpfBpCZE2wOqf7qn
HZGOuJbFppK0KJkmU3cGG1Lzd+7KH5ZoT+pGT5DDbrFy8NvHr/TviNE5URR/XO3g
AfiLXGtYfFDstTgizcxC3I00ClV9/uARKIE9yypia6YhrBkspC7BybAf64V1nkWd
Fwf1E2fr8C3NEFPWcjcmnGEQisR8ebsKfIrwwDMbV8wL/jGgwyEuB+vnXs2yeji0
T6pAMgxGJpoFtAduq2rCpkvns97lbICaVv7vwwxJgOxDIV7MS2FfC7YUlsob8Ywg
OcJF2uB+aTGnJmLNkreYvDyTvgq5IiLpKunRjNdMsvatbxgL0JW/xQt+6T3qoxPl
bGMAK7cdYyRfogJzr7a1+FuKOnoJYGnTxlxmRIT57sdPW5Sp6REefx5hcOEN/4rO
UXqXkUoFKQr7EwFzI2UQN4j8R+YnjNwYhzHYh4sy/dmUFQpakOa6vF3S8gE+qVMd
xCHRjXhVTRFWEXnv6VCasOqIrExI/wvSbJZcqq5kjVx1IWcH8wlpRF0WOn12SKO3
xL6neq8VoBO9SgoWjqFKS6EPVRB/84u99pJwdK38XTn/X5ktMOAKbxDbsaKOC7jd
7UdgJVhK7vQuswoGzZrUqAFZPz4a1bjWM2uiJgUj/2pR8if/HMU5PBSP86Uv6cUi
xM6VvMWNR59K06AM58c/GMc7mFCY9RNuC2KnQ4IhnxGOhENHjBPNtgMA1PBh/rNN
3d8AhBTDOfGp0AidgMW8L69upFDVaBKO7iaqS/FwmMQ65O1+iPazjqF032cxcSma
VSbZRl1ZUJS+hFMTOVdyaWF7blIjtWSt0bTWDLfOJeNkpiTVwAN2J850w8PGVIqL
t3D4JEEJ/BSq8vjLPpjO4RHSONn3Xpuh5xy2m2Ufal6hYsei94p5SXZyGHyKJwkR
Ie25Kk3A4C6JK6iG6VYFVg5fwprW1CR2hfl9JUsQgjvFY+/rFTM4+3RB4dAJPaZJ
m17OuusCFbU48bGd6ZheXubsQlqFgLc0B2JkUOUuWBr+01ZN/r2hULG+JZCPFIXM
Brb/eV8f0IWId/ApNXe0DfCJGOpVlo88fYrtJTPvQgdhSxpkc5lS77paFCw5AoUd
pirHyesSMcjxelJ0QxX91gLI3XGM2uoFdT4SDgXzTlBIU/ct+zr9m7xjN0XCgy1g
uLKhpZQ2UpY8hcwHJ3KuQ8r/Tx1TPDGyK6N38hpK7o39nPB91JNBLiBTywlEafmu
O0H4eCm2sFRrkTtxlL4A00+/lZQG6Tv2q8FimnOf8Xww0NNQGDoJj+HhZINBa7iR
WftRVQrUUNxlFvbBRQftWjW2srpKt83jys3C0tpiuRdIyQ/nAItIGU1jt2TssOm2
/IP5lwvHrRGC9ykHinXjQFIVve6b951IRRTgyzNJ20MSG3iYhZypmRcUfpapCQcS
XyaLtBnuSFEfyLIlvCT5FL4ykUQqGi3AdvOHmkPpWI02sb6a2Yt4D4SnyczAiXcy
CWmu0yc9n9+YXxZGpsIa9AwBYnLh+wolnmU6iV1OVyWNHTKo/8Zsb2ufPyZqKFf6
0SlykhOIQNWZuQda/FSArGc7Fhurzhs/gFLwEAd7iZ6t6mOpZ0cafQ7KuBrm1xEf
LI8KfqlDFPmy9k7iFtblpnZDXrmIW0U8/YgVjOqboaDiBpyx5iQKZsDlHheTKHo4
14kyZqF9gFAO/uEVFK2ZJUnXMWT239T7FKH0XQTMMkZZrTNdEN2sMAPxDyhiUH2b
PioVGNzHMVhbJsAdQWVK7yC70DgcUwb+KDpHobOxhBPwJBYro3GIf2Mno4Wj4WbE
xPdaQKkNCqrNxIampsB/DJlJKBt26IGO/qrnV9bQrL9NB2esKNRZVJyIJkYvq90x
fG5FC6rkcbqyyn2BpuIZhoux/mE45kmHPiCobl6m20avskpNE4M1WA53UDOEtIy7
u5wEw7ntopuFYALRe+0RffJ7JpG+clNhji0CEBq9AS+rfqkRucIC3bV+ggSLWT0O
YSxxmFGF1Qe0+Jk9tXy47hOf3irLwsfm0JYh9ga9K3iBgMMJgKlMXXPSizA9iLAS
x+xvAsgO0fPlMspXrSA0JriQaTQJlURdaOpLoLRFoQ+scJSVr6PVrP4i59eenfBP
1eiatI+w/mrsdhCbZ+OGdAWccEh7Os1vF7DpLrEryXuVJ6ziRMJrCf4cdOOHoYdi
A59EHbYR+K7XVJoJis8s3OKu1xxfwHL98sO1g+wDqT7rO0rndukA83VybMufCmEc
5WPrFgH9m/Jag8ym1F2mCqeXkbZsqQTGNUiTEH4KwPHFEH9hsegUNYMdZb2gFGU+
F1XPth1IOt143KouW3PSv6JQBZzA1HBH3t7BtDv8tSW5W21TrYj+smCRp4rWMEno
/D7ntq9Ajp533sxrQl5gZ37sVRZFuuEP/8vwAJFfDNEEuvRlBPahId5t8FgodBvk
HSIMxQpq0Y1+04N3hOxMLApucHYnFS3kzCQ6MDjQ7rVECkwMxIzHI5sAmXmuLSHi
CHbo9bvqogQUnJq5eJIem4yvDaT6JM5vd11TyZOOFqR4ORgmmWXJXNlGvWWR4s2Q
EPIxgJgOecXdqaO53loQN6oKDuZ/rGrZVgDPoNKwHdy0Ms9ft9R74pUNfjceTlYv
zhrdcm4N1d5J8QoeipYYBW0CBXMlD71TJCAJIdNrf6yWYSm4IWnfyitBjoGeQadD
lkBRh4KKV0bTUdJ6/atZLY7d/gekceqIpf0Pq8p34zKgP2G6r8+4VnxlhuuEhg7d
TKdzSwGCTguxdT6iLFwnGAiIjg1fSTP/kEEqjgI5zVWKnb8+KlQKLiZF2Tc3e+Q8
n2pM2DiX55QeIcvrs44RHLaUot5naJPmSero+0KP4yvpf+wnu3PpYi+1tSdG6Ink
rkfq9koVJfwhirm9BHua2te2bdE69AH6r2yIUhljv9M3NwZriJ99i3No6QUfgKhp
dHSsvObddOESo0iHSWdOUHu+ltOT9QTTfYi+R4PhOEVXNUm36fSlI6pqLBqNyUIa
ylbIH4DURStII3OLl/GbK3BTP8Zn26J178YZzc7JHJEqCDR+SezUBREZdRgPvEfc
ZGyZEPHLRX0uVUZVSZ8jnkB73Y6YJCN/QvBJAhuTeNyvWsktBaYDC9j+4xILGy74
Tze2JsGuTKsehw8iuvfDz5tMKxXfU90S4qiJa37v+XTl4/sw/UlkwrLO0R65eYlD
Xt7mV0iYIuG+skxvh01QOIJFJbfZNrtzQqfExqjbinPWiS+M0JrpdcrcQzHNcyHp
QBFjj2DsKtR08+Ckcp/PPSdrERAbg5W/W7mM5Rsic6x4lHowhw8urYxzeZ17JRH1
qV8zeYO6/ycrw3JtyaGFcSJmwRw2CS9KtjB/cvDT+Rn4KtqnG+53vJJP4/XksaQY
ryKcBNjTtGd1X8av/iO13r/kO4mrw7DVIVLWnUMTvTpkEjXsXszIW/nJk6Oqdlrv
dzq3AD1AH4G5gLp+uIcPQBt0a/p+ZYEjWfpXzaN9mHLPWGi4ZoJcnLVJ1lgMxprU
plkNG3MI7Y2EGrtgbGkwbkmhIsgV5yZ8LQLrt0u2WDNIQXsezpcazQ+LhOlZm8N2
jdBJD/QqG+AKTNyuArenYBDRv2VUruaa94wiOvQWKT0KJudXf8dFgqeMDFwhAxSY
RLCyIxlq/rskv1BTkMUXIUuzDs59j2bk3aZJzq7iLQsit4A6z4+tI9TRVGz5Or9r
4182sys8SY8yPg4oobxg79E+yqDhmu7mzWM+QVlg06k1LudzuIFDWDlgRcltd3K+
WeNGW5Od1EdBKBhh7CCtVnTTDktd7z87D3U6sN/u5rpwoUwR58q8iLacqNIyjATY
Hi9TAFSeOCHuR91Z+E0y/pQCeOVZcfjG8ELDvb5yEbHg0UvCNubCaI5D6FQOJSqo
kAgvkSToYwAf+VSLBOzrUif4L9FGyOl5I4hRQ4ELg1IuKPBei5XpDAcUS47wKIvQ
s19s17cKcCFcSC7GuwN9rd6yoMzd35gnoS67CpRjgUXmlRd7HOwUYXDTxRS0SIW4
Zirn/bUb8jxOWwIJXkFfuOFVDh5tjRzwDckRUPCvI4en0zFsyD+b9mlmh6seK45H
GAvxtdRzKow60H6t1ZIg3gxc/a+M39GKpXeHArE80AusXuTe03lL3Gje46HoXH8q
wtEij01PIS1LaUH3cBwpOt+FgMeWgsKyvz83GK/jv6UGZvDwqiLadpOZLnGD/g5n
TZl8pRJBpYZH/93nt1l7OizSHOvm2SrMXM4Q1h1X9KmFZJ7uoPu8eNuHtWuD4Mfl
5TAWke3VFCRX/dthSooyiI9aUI2C+V0tYs024fLOPDTG0sduwoxutanUydDqby9m
Hx57qKLMYwjyGhfUNAIc1kdyWfvsNDblxbY4RVvM+ePtWSNwEaBKqfLsfoDJ3yQ1
yU94qlbveBc1IfEcXPJHDa3hNf0A//qly3XcQVqVq6KXe1xBppbNV+W7f4N/vmcj
TNpD73Dqoud+SYk6kU7DrY3TWpW1buZbPktK8UcK4nvIRklcnkoZBYQ0ta+fs+sl
mxR35/WPNVa314+VJxMIVwFMOgU1lD+lZKrt5t8zMKCaVIaFSEJ3Rgrfm+MBybZE
CVtMJrMdmG1WoMTqFD/hUPX6yomq0GP/WtFtGsGiLsEQlI0zxBQ15rbIew7bPlFD
65W0L4tIsMy9GE0GPXyCwkzAAZe8FJWbiu/b2XyHvfAt6lYAsEQvEEF2JO9ZwgN/
iA388FRhfKIeoLN5dX9IIN3B8WEozDfwyY9Di6f+UGCc367+wz49q79NPDhEoAp5
ouKtTDDWEZ/JukHREQVOOijW6uF/tVHWGY1HWPbp31cek3pYSYYTbhiL51hJDins
ZFbShA0prhJNSjbvZPENBqpgUOnmVYZew7/Bulnz6oWlegvHQG/xjsIz8ZTYb+9e
DR+0WnlyzRmli6zrawH1SkprwQGfSTjqhwbY70SPIMhW3CgiY5a4w/r+2tucD+6P
v4MK6IhgqA0aKB4UNlmZaoIB4pnwwLe3FT4nz5A/JgDsvc/GFKmMjgtEvq53vVvh
7vjuTT6e1biTdPGXjNgNNk9oRFc8zXXdd4j19IWRhdkb62wbEMBn4b+KVoPIF6+8
GHfAbI7SN4Zmd3EvmIbapgPGhx2rfOXhvgorOVf0LIdYASQX4QIhzm+oIHPAkglg
h+xIYxT0eo5XjNgbhIyKJjjOehvQYha9IhzDaCkdR8VpuMQm0CGWxBA90Bb2O9eb
EwevpiPqUyvO4nrg+lEFI+25XY0DKl/vPMAluzezltM2HuaWgQp3GXonF/d93es+
73sA8NJyfWrDlghXI890iUFfRM36XWrVKViyWOOLbOYRIjNW7uDJjXiHNHyK299C
mK+oJ8CxDiV7+0m2wZKqggRdxw8WXxLSnEPlAOJJLvosFn0p+P9GstydpdzFcH1s
mo1LgKDlKcKpeIuBpgNehZLWA9SKKfPPCM57L8/CtxlKvt9xx31qUj/cQ3c6BPy3
fyJitZy5wM9FGfmSxaVRKckT772FF2nZ+Euq0PSeJ9VqXeNEzJzoBEeD4xw3WtVc
hxLKu1L081wCFtGyMRGsaZ7IfGRQbF1OOkNwbfL6lB8bFlce+Xe3fAp2Nio8NXfr
ePtWSkq4H/A0i+DJ9864zqdMqVjZ8EcokYmGAvQwHY4AEwzKxVfM3h68EaYnyxn/
ugDQ00F+tBt4VvfZMMG4BLmQsWnY50Tkx9/sMT8yKjgR2Wg8IhgelXt1dYbLDlIp
wQNvjYxj0OwJLTen6uU3FqOFu0xXYgj8G1j11oZ5gtJRBl+L5MHc8owxdzLEqzze
P4kYF2xZ2a5aNGPQh/1kk75Ha6rNdy11Njh+yt6PpRM70nnt3Ui+yZKi9dwy3FFi
wtF5mvfal1QF/7A/gAAY9lyk4mneYy9pr9sP/rotPXpnpQ0cgIqf921flJ8tz4qb
UiuUqEOsDCmTibTTgtFIEotjSYf2Xxpf8ZxswKTuATHkjXcqqiSU2BQ0awAS1ZK8
zI9Nq0TXji74nxcDjuao7U3RFnhg+ehN+hGcX1D5yjFwefzWf9/YxG6ivgVEufYC
XVEH5hl7pm79gynELQ7VNdgKzHKi/B8j1w37k/vM/m7bRbl1NZ67/rFos0uW1936
gN6I9mzpfORSHLOhKG8tckGyWqqR4tM8QBAPHkCBYyoYVoBtfXyg3rsYj+C+Hzni
BmnDxZQYtUpr2kM1Bo8+pi4wMnnNvIG26aLmr+z1HlbgHr5l72AZ/zGoCGURep1G
IfHlVSsYdd/wjYYIbL//pwjVGqs2ivtJIR2UK6Aq/M90+/QOWa4HCFQYQCwPdpUo
2uvhMnoKvVt9Hi7z3ibBkUbTLULPVVZxt+8Gpyz3oSIryVpLmRtNPNWVZ+TxjNlV
YkspQQ4szU4ccgof1dkK3M9X8LhIfO9ZzSh+9juaI8KPPjf/18BI3/vxGCJ16UAC
Ep59KEk/rlDa4dXyluWqiLGRK5cU9gnPNoEOcaZ85BtC2q66QPrT6cPdWPFJs/tP
RHMV0vnuuA3aAkLQHyX5sK3VSsYDr/aeHy4AiWTeEZvoQ9u3TuO9vUkK7YaF0JyS
haGLeH9e4bIUzLD1lTuZQJpLI+0pV/eDzNyrBdOT2Wj4ZsqxZsRdO+J82W+nUhTi
AdVkGeBiD//m4PZwOxqxF1pY2ip8ZGiYKy+vfvmVyzsN63ra/RCguAttJQMpMros
GnWuc6bET8KToaDIDLJi5FtN0MT2CvXvJ86PGpgCw7rmmAufhK3u1cz+L3U0Dzie
kEVhn7hgBINoXYbwA8b3iBWqN0RId1pM/zHlyBtV/stL5p9kUTXX0bLdrcKawhES
lonLCbej/KuiXRvid3TRI/ojO34HwucNZhsR6x6UllS2wO1sBoMfaGajjqBCjjHW
PHJA1SopNK9k65hM5cH7leZfQYh+z2cZeKaNCrDE5Hor8jarz8GIWAeit6jZH/f4
WG5IixZ9NMnKcQ+LvkRzpoaXWSoPEU+L/+Q2ioZkCUl28Il7shdu/8XS7/UHlYQ1
VUo8gsOgpARDrRsctF+0QzFtMr+DiEhGl8tWMcK2pOofqI+brvsxv52Rr2s4wpuB
5YdHzSaHdcojkSeYxxI0R6/TlfC2PKHfn9C9TFa3/oX8ZbpW/ml3P2dqtm8koQN/
BMqc/LSwBwfu5NCVFgqXcNC3L1lbllK7aSjJo0DyUY72RXXhF47oKfbdxcoNRQx6
v9cRjgJwlSY0XtBcYMYWGSWfo4MV7luCK07RqmKnGBe2ZvNdOivdXPQ1pPp/x53s
OzwAGgP1uI8oUXuNGhDJyn+6uZXoHpAmdFJCFydZpOtWA1jsr0PINUANHK9anWii
GezHBAYc0AJHOxTJrNqu5DUMSiJnsOZ3XYs4irhpajip9zXlzX25Q2EnIAx+FBlZ
1RccrONFXtrf9gElKxeFqYFwHDS/YJWTev/FuRVJ3LsVaSxNgl7xt1aO8TTPPkiV
O0Us1kW7uxVnCZpQs/JZeKL+Fl2QvVQ4f35RbpBx8NC4izbbGx71G8lHZBu59WwM
+hp7wGl5+fBiYxXMVP6+tSjXnriJqcI9wUkumMDEpSyuaJ33XPYaLhbvT1aAXXM+
auaxgnqrgPsx9UBtF58oievfsSxz9+K7+N93AE4CS8z/EbD0ejFA63H9zxX+ep5Z
fIbBJbY8mWH6dUwQe7InVEl6D7X6u1UNWAYsdXaRw82XsKdXZfAjeol7TbSWOCZz
AT9U/vdo090KB7NjRmkyaPZ2aKUie7bwShengJArFKFN3QZS89fnRo0KF8tf/PIl
DyBzcha22jWtwII4CXjAZwDn+Vsqk6421u9cYvpqT+zSAr2hwWQXToHfDS5qWguQ
Sr3JCATCw0Itj/hApdduooct6M9iyVTcmNV1lxSGFZWWha60S+YxrBD6YED0LahQ
2H/mQxpNQjobVyLNWxDEjmj3Aq3nD8vNluk63sKwXwTaGxhFqXBb0/Hy3ElktQAA
y7BLhrPeV2sTMz+OR34Pmd2dYBj7XbobyMPQn73L+6EaacA3ZSvlnOd6hHrF0h9x
3zyzMR2NurezqKPexSUJuLgrLCX8tyxtWtE89qco030Fu9Pn64kbR5XhwwZYG7t2
294xJjZsJa54ZmvFzoo5GEIW9W0+hAID8rHGDf6jTdS+2E7M29h8mD9B+sinkPmd
iCQETGikFccTG/IhMSGILs1bOywmPLN6gt2q61ysCYnOpgpjig8/Bj02hnvMhnk2
zEWJpsMwkrR8itEAEgnlfJC3bis5dztaiM/e1TuQndB3qBROuOURhNquz4jtCw4c
+EWyHEqjhWnFY8ws/Fd8337ZEfiBQOtbIPwbc0QSB9TW0bFzJVj1i73j8aelQbVk
EVmXETEDb7Inn0eqVTT77BdACNhMn5xgwgB0JJfEJdx9v8n3zqhDZJ6TZk9zjP5W
M4iHSK0xCws04zdpl4C0nLNs3E6HoOTyhwBu+RgNjueuwu3D1PhjRZp+BNIZFryu
OgZYjsIktt0Q4XGDlsgIAuPslrvZiuCCexD2cXfA2ZVvL+P+Gw7nvGxjq8z0c/qw
Q1xBN+7KfLNaVWgtO+kSX8vWLILJPNP4LQYaNZeQmafm7EYFYMI66yNee4hJmiL9
04cs58mI+wFko9+u/eofu6bDld3ugreogPRafHU7YW6yR0KUu4C1+arwAWtuXkbY
sTL6Yy2IOvm5cHU4kxf6koPMtReEs4tRLh1W3Ls/9jcB7TtQtD5pFzJJ9GCkhyWz
VTMQR2FOnKTnNMlJNRfUlmCiCeS+2UZlp44+mT57jXxO6VG6K8XNVtC4ATBVOZYK
9oix2gVedtDjC1T7hqUUtpUAdUdOL+qxv5vCHJOAGHnN5SiONxaf30VV5jt9J/uX
a85btpMj+kgsu5kyS8CPo8JVG70hH2M/N7LqynLGS1ul/INOxc4+b4/B9Vuto/PV
4xaZ8+D62qFJZLcqUpKfJRoXqNHX15u4MDw8F2ZGZtLKq6KBi+al5HzNDv/EiDXA
l4jMVHC9idse5lMLC4wM79n/bPm7BCxe8Oz8wSzF0wEfNYYhe7oQ0lU1ElJoaYFK
W06+dqXCT2J47wMmhLLe4oM2M6zUoH8piIcz5RBqmU4wSUh0gEnwhlz0S5P12MZc
w2ZRO9G5Inf/EtdV17j+X4omFRV8vieto1KHVDBkE4vd4vh1H9D19bZOTkIqV5Ev
xmA5gT8tfGqCXAYtTqzlNuWSrrYAo3ncSrwA6ppX40Lpqrnx7pIq0nMSwdqoO1qX
LVr0f4PxvnYHemkFqZuROLOgAoxuS6x8CjTumlhV7h2PC92V6biXqXV73Lp20PMb
My3GUxGPSX6DSTc+97jMAhSpRTn4ITCysNLYknJN6S3yX6dSmXCo73yJDIZUyxYB
6qm0JhveCsoduX0bDSmvx0YxN3io0YmbtWJh4ifS0djqScdrBjao61IgZKutKMO7
7TsmIQ8zLnOBNfg6c8ZWQJjyCzxGGrnJn1n2hGgXs0HVriWLRn9cXGyEQ6gW5Yp9
7ptsiIlQ1TYYUrVtaNTc4/uHQdFP737APSV6mQDJVeCMMsJxyAHRRhydnVdubXEr
WnwSDwThyW6IPY3jrnf/u6dWoo6PaL/ACKKWdVKPAURB1UnnE2QNp3Q/frEhecR8
7Bs8FPgIoahv9wls6Cpx75JBRAtDHHCAiJUxTtXPIggFkZASjHO8TQoq/5hz9LaE
8ARFXPjru4eG3z1Pfa/jf3EcGRvAq/FQsiMJp1z4GrAAIBN/h+eXTJKIjZYvO7Zf
WdDbeo9iVKhVO42gFerxecwRKbmX+cBZQG6NVxJvZgknJJniSjg1ENwJv8rAxvhj
HSOmtz1QF/tpF8B0lSSxUIEHuDqVJKmSbCcJjxruVtZIUvuBGlYzqzKNslaUoGYs
cUC2KK82PNFh/6QX2Pt9HVn7zXQB2zOvv0TECIpM7GWh7RX1SFGDh0yN54iMtHii
97KijkoJHvgArUO5JshCbAgCJS+rr7VrmRNlhLAYH0waCjTT+GZ954Zllo6kz0y7
xElj3xOMlOdG//aEJNxYTBqJzawqn011vwEhFHgJ18MInGyEMTW2di0fA1EKUK0W
In4ViLJ2Lfvg3ZL9fQsbwt1/5xcGfSV6ksxy8yrRl70Pwx9iuhk9jzm5C4BGSqIe
a8Nb8rU9jeLsIj7PrPCKL/1JzsiGizL6dRU7F9zgVk88LQrfsAIn6qIGjF4MAziy
a4qzc4hYV1ztErh1H4rVANeym5WfuiIY6NqeRAkd8Z2rgQsP5/BEJwc9VyO69ZKc
LpKdbIUj0M+XtifETuqJMuUujl0cl5vpet88coScYL6fsA94LJTb9dVYwW8TDa2r
NartZcubuE5sgX76lKkOxzNyaAh3L+cntU/qMiVgFIYH+iyU8PTv898jQIJlZ/Dc
2kcXuy0Ha94E0rX5yb16VLS1c2o3+h0/33pm9puKSCaB9pqtUPVPjI31rErcxXMD
rWlO95adMppIjwuF8JwEOdpwaQZwd1i/onS5xnOPNESru/qfnMHLMr5hCbVve81A
BPE5h+c+oXjYvMRZ0N0WGO9BeNtWsZXrca+YntsXwMI3DArstnJ4WMrr1HGhTDIy
TElru/MRiBeK0OE3H7lN/z42UOf9ePxNPIyoJ//IX7LL/P21r3JOj4SRwoYjC1x4
5t1bPutA7ApdVANnz7tIwj4tA9L4w/IVG/Dp32sdLR/4eVR1kdHehEsl1uS+u6rb
q+CrQAwmIWpVDzMuqUXKwjSoMU0FpLjARe386jjiLE0r7JhOiLWS7943nndHsvOb
Gej1zFWxp50OR9QS/+4gKs9FwB0RzB6bbsx4e8F2MjBtR6v7xU4av0d/lvAbIelQ
Pe3SkVFMSGhBr2mOqTmed0vWmAuYkYD8Pi+y5xtdQdlaRB3O3IW8eLH+pd8gGtfU
YfjyhFJmBRGtW47/cxPrmosNJ3FmohmPk4i5gQGQn25WiA4RggVc0oeanF5yr0uO
jkxIUyae4VQyxtI3+Hz8Drkj/ybAh8FCw+FaijhJSUOSDMfioqYgPm2lLSEVgf8O
NCaCLrPCwohNKCZ+ynDtyIer5pBNRA92Fuhq9mhct93YMlL7UR19y64gubJAt2em
CK+odV2rl/oFdyC9/RB7y7g1019Z9W8vybaYryeLp/VcFPoesdEZcrOmdxOTevPY
SAndi2MW1599H5uMp9eqe7ntQ1tYo9s3ora2JdYeV6U1kkWmtCA739H2Nx2iTPXl
9IEvb6IypQ80+FD0bJvxrmh4s1QpjgCt2S6SBecx1+45EHrQXtzbfzDMKn+fLqMZ
deV+CWBS/6duY0eV2RuIutAC2QjFmzNqcreO0n1QvynfG6RYPHiFmcJcdN4kGuxp
5O9PHielyUjDNwyGXZsWL4YvL0azJqj8R7syYmF29CdsYpD9D0S0HLerifiG1jSy
28QJoVuE+Ey9EPI2Bdyu5xryuRNRW5ntEc4DHQIyxekuWZIpd7dTxCfkQ107piI9
Q7F8KF1cZRLqyT4J9QPqXL1M/1AMpiyK3Lzuwcbe1w3iHV76UB33nwCoX8qiV+MR
0aO1pZEa6ahqXlvigh5w52XHvMkvMFaeQ7isd+bC65hnu+ryikl7OMc0rVvuxQC6
sN5pPqXv42N4QnH33TKk3PKeZrPA0GwBvnFD18fKV+RQI6t3cKb9gOtvSIW5A0Tp
0pu7U2p1eosntGfNSJwCegv0TlimP3jAtGtR/eMu6sd3YMB6Bnvg/jk3I5+v/ikv
bTOl4CmYEFJ2jxFThVICAfdhyOJxmWBknYI9d+1cJQ5Zbl9G1ZMPgF3FR8hfjjAd
SJ5v43E1Ksj1RDezxyEPfYJfaaEROrB28xi/RUylBW7jODZsnPT89JuruZD/Ucac
fYo1QQ2AutBzQjOb/WZ7UizxXbM4ak1EVVRouvxcDbjw38HnaScxgcNr3rZEB+HU
C2pVd7ro8YTC9Jx6qea0A8V02ADfsEQnOnuVZmZr0y34mSl85TxWQJr1sLFxHM44
QF3lEFo+MWNEvBP7jmgA+4+KjPteaCgWv1aTK5FNzPMRD6IkJErAi84peT3p5Q5J
W/PC+J2SXPvq35a4Ri6qn8wnxL96pbaZSKTxUkt5FwmvazDC/MdFz9+X4bvQZSnr
4JzEp58uIKlfN9eiPldsVbbgDhBA3BUrG7WAtAA98z//7RF1gfzOAwp0Hs9ViQi4
OlqM0+WaSGCNRCIWCOBUsu7j5MNhQaT+dqmcunSBUxKx5hBRXhvv6IKgy0V3D/jy
Y8zx0vR+ImOILInMlDvdAKth6odhfjx7m1Fg7SS5w6/yTXYPRhaUXaNnvqrh5yaj
VVrJna2aXqkewY58v47rO4WIuuoOF5QAi/Tf92qKsF1kMUGU5nghRu9HS1Y2N3Dz
RRXlgvGi91o5o9ocFUJCVgZgjlNn29USjzm4rwkyLmh8+C+cHkOxiM9vYOKZngLe
1tW+Gx1LBAllV9LXsjtVogTuyS/OFyFb0XLtCc8VBggJnv6HVn9kDxQJpwNMThxV
kR6DeTrRGFrXYDjl6gZijPUa/Dpih0qTg8DoNfgLDPhH5BPKfeJgNXxE5twGG9nq
Ai+Kj9xGSUlR64Jnmg8KwGU+5xd2Aq8HUdocYj/2w+mnYwGP5p+s5J0UzZnkD1rx
Ceu9cxyeDUsFOlZajUiPQDrQP+NFgL6r2EmhcavmyOC3mzOBBBBSuo7V2nCFDcOs
j85pow+7emmMgG7HhMPapFAxUuhBW+SIR/Q0ztSGuh8DolGz4sQ5DBeupcp/Kjro
bat4uSJnYK5nS7oYdRXiKPENzL5DEA10LdY7zRoLYL7/KPTaqh6ymJjEPkhoVycS
cSW+e+uPoArQ7iFIUTtO23z03ri464YZkT9CqR6u9BJcF1wS5H7EwXX7c7ZVxBP3
Rv85Kvfg2lzljEsNDJ2rwSCLDi9ecWfHymUxRkJfwn2BrantIG6EZYDdhfE5/JlF
yGnsemN+mdwcUW4bTjRbv5RdaYtTkeFciMk5NM2oZujTdJ9p2t6ItpPqiWjW2uG+
a1Rbu1rGPUvmehvo95608Lm3YZMblAO2JZ03oqC0tT8MlUG2py7z0uy3IvIHZleg
+rZ4gSXsRiKJ5OBnB5aes2ptt9QQ4Ffk2zAyipHeOcxSY7C0PN0vSp99UfBdV9pm
2kh6O1JRRM1wiC7mqE1rk2hOLQn93xm4Np4nTX00D9B0B3On61s/ZV44gMOnLrW9
dG3r8OLtcK8dJUFlvjjf9XAzTghgeaga3cMxLhHbuf0PMgM1v9VT/4uVKXYtxLzL
MW/OZ8pns3MBb89LnHA7RKL1QwX1RoUlG6RTIYE1HkbAHzCwjXbSNsBvYIJjVZFS
YINAki6DMpYZ9qJWbl8zxuGFaI7/gmYVDSYrJFQGrnxe3IF8zicD9rsBwvwk/YiX
j3bSlJWXCJECvV3RpRCI2uIyVIijrPNiWBgX3vAy4qeuDoCJQ+DgHF0z/LD8DUcQ
acZp7UaaWG4Z00NnZ0qWmldSptCmyHOLmRzNo0DDaxmROct9PMu6HhtrgkcLMkQc
NrsUxSIxBIPv5k8TSgwHYXPP8vP5BnKv5b1CTZPA6rr70o3VoSI963vBoFclXh/+
yfwYTzEcF+aZuD9q/iSJIIrSF322jxB5HLLPJ4TnWsYu0uUzzDb8iifjLMjvXq3h
kdjDWAW/8gDFAyvoH7gJmVUHgv+rN3dhSYJpMLHkkty/OutDVyfcVomvVeHIbzKD
xlwNvI9AVa+XVf4QAJgxLNielmYeaeqpMk7CFVsyxRvtGhusyYtr3hwEUkIhUrCh
yKcAxAsmd33FxLpY6lL037oifFE7prCyqb4BjU8Xnc7W4fWrjEjG0cdDn/vH0bQf
2x6QpBY1GOZ8ZN8g3zbrTZO3+HYsvI68pqZBVwqSQzfC4LExLBMX1SdyTZbM9mla
AoR3x4fNUf4vIdE97Ww3LmR9YOR9IFVrri1B5HLfiOOC51M2l0+EROY6WbUuI64d
2i48N9cJGfnjL0Dsi6UM9tndRtOvqRomOYrVsa4BSD8MKmAFKyl0OJowkz/VY9Xd
szmpHpapUOF0b+HZr6hWv5tQoM7dpUU5cyONH5G/BLom5zdO29ZvgoMLXL4XbkJ6
3cBE0dsw8lnAe3c0wjeoi2GaabRA3Pjc5yi5LImx3HbdA0Pf9CLNaTtRa1DtqUK3
WPMzbYDPdVswFJIRolChcAZnVpLuTOchYs4CTMN3IgQSKvk/cCh8uP7461fCKVoI
UQU5n1a6ttpNoKeCthvO/Ktcjh+hDI3S1YOgk/VG39jf2AOnWoHpSbZ01q/Lr/ea
x0A9jYCUi5PobTx6tpJirjHOaBgiYPbteJVZfXZkBhCRfnaJBIsnund9WSdTLIUl
U+HkfWW6sVRrXhgXVNWPN66g3XpZYG19oWAe3JPPjMTGfGCR5bikfhyy7RMY4z8Y
MmmatWev/SezV5QObcdeGoqedHEFVc3Zcrexw2EpVn4XFph4u/HZxcjbiJiVu8Xo
T3+CLSEcoGk5l3546171PH+zUX54/CmiwHb5KGAR5XhuBFkZ+WLhSdpDFyk7qEBS
zQeWYUYXsAUpOkYD3I6FU8MWF1rtBKfqL9UuI04b+Vhj/crIl/zoVkreReSjEqfo
3lyNznLcTMVwTwPYDk4no283omQ5F7e4w0Xemso3E/KFSeQRL64G9UeIM8RkE9+t
OCtBnQfWK3ZYK0m54k+/hQ3qntawr1UEHlFaZosBlUbzyjbegDh0k3OLpdw1rkOZ
fkDluEY/9DJXyJWUYiatZxeCGbYqJfxjbM5I1Kg4jA+LsM0jdBxv7bJ4uH3Nc9p2
+36MTxw5XZU0C4aSd69o9syqF/r+T+eNsO4rlbW51+/cTLaN7TINBchxdy16iTVI
RDES2K7+ifY4IDHHI7lzGR2e1KdBuw2EdoyVlW7yKGUR0YYXzwqpEhX5Fqsobjs9
//cJHqxLNbzwQPGDH4yJ8xnBhhBDveUL0rvd0v3Qd+IwsuK+NO5oUwunojdcYlim
rnslp2D7dqlE2rzRARDTAM9TQ0yY2NZN4+xPRBV3BU7Itn1tnc+onNuHVbqpNJKA
jsqgTzMNjx4z7LufHP3fYjTlwPrD60cZyRA5XXykf+OiF6fd+UcQOXpXAriqNVWy
wMWloj2ztsFLfPf3Cln/MFTRugRp74jpYbA6G5nFmJwUzP4dcCLO0Uc460+vspKC
osCgqqq/id2Pxl5lNWXyFPju9yfH2dnq4ZVNstkxlXCbu5/jlGgKycNVF9haVTAy
sfgeLLuq5Ksk2ytsknTP0s/gAkIkcqr5yZ07bjwXQ0yZan7I+Tk6WaASY3j3vLfY
/q72X4+D0/PUANSnzLODC0e+mv2eMekM+vDOWHaKs7frIoO2UTrDGodcmRsDbx7w
cWLHpXL3VJ0mkXyIlOXNb4Ju09Gk6wJcDgVA1u+rk8fFclVK4ZO+MBn8W0bpElXo
0rO22AHdT8KCwm2eo+8nkudN7ZWNJhpLFr453qFb31+r2jskvcQf4H5z9Z4gaems
lNoywpkS8BjcqTJ32tIA35qBfPopYqfiKCJJbh3TbdZ/lPKHwRQ6xOHPx1NBgQDv
XgJF9ws8055CNS8WwoXd8Za/Gq1F7Uc8+or0T2S34wmrotgEqS1uK9IWz64Zp6nb
RKhMnx+nhQuxebzRCUuu1PylJDc+hmarkjjMTNil9nzOYQL1K8x1/S9R+Jrkzzmx
s6EywE/lhck1qMJaKK/AO76XOM29rq7s3VkN+Z0+emejUs2wxD/FgGaQlJKrSqJr
CjaI+BckrxqlEbCnFwLcrSGo4P9xH3mBFEGnpAdx4QTjKT/6wRZNgnpqGml46PM2
+6QrrAZkdm5cA/yEEDIf7OT6XsFbjnUoojgkuWr4Zb02YS9MzYoYBNiDPct907JY
6JPQBsKNaqKrLoIhqlA3oQhNleN3n7Ka+h9w6nfYMabNRNk6r0IR8UdhfqJIsHYI
XcErWfeLNb5JE6JUaBeZMmEq0pb5q8c2YewwHOcJ2YP5D2nWwc7XwlLRyAF+epsr
8yb+kWk/DLUmK2S9W7ycJhE8zrrUlbShUi7yrmvbHiRZiorKM0qMxR3BZcKFKtee
k7+sDEZdGSivPkwoObHaizQWt8hi750d1huj7uMSXiDhgCNA1eEQ7DLlRKRcOioR
qgyWmxKCwHGL6ndn1fUZ+b1Z2eSZT6sqEecl7ZDcqvm2N5Tuys//DBkHhYE733oC
Nz9Py7wkzhZIjGLEdz322VzgdQ1EQlbYE+f5WiuzFZ58+Sod6se+2oeInjD4E5kv
1i591KDw1xcw396RssxalI/+DlvUE8epVdwayipHegaHU5RahlnKYQJKY49EfJ7U
KRNlOR5tfWJ3pm/1elg0hPEst58U95mxgE988O2C/3Az2zwyGuyGCZAxMqh/E4L+
7N3wp/uiNXltyeSHOSUp/X0gD8ivPf+V4FqBgmTnyGNyKJjbcXTdnpbQGTEOmzEf
gKZdGDc7tlIjJlKmYdZiIgRjXLERrkLNuiUNJMNAIna6GD3ThDkOvcNPfARTqV2H
1YmVy1Kbl6QYlP1t0ffDpQkJf6v1wNZh+IHqBl8oa0xBm9TzdDpsZAUkhmJ158NX
oPfua+HD5mC9zCb+wn7hMfy2nUp/XCHQBMOGeo10dVUYyU2sg6ZiS6DwZbvTFJtQ
tZ8iM4f51C4zEIVnYf/ZpUA27oYqGjuO7jjhtnUhsCRY03ouy0szxNHk7qx0BGya
GQ1yzc0G+4LvDnuPcmQewtzQwl9/buH10dHQX8QKyi4ogc9N1OsPHWBHv4nUJjul
vutmYXp3+0YsXIFntVrlf2htywE8rKPoxRR4B9T5zfK5aG0bT7ThLHASY3Aq6jQ+
aqqro/9kmPzS9QQ2xhxWxo+c+Q8gy9lkdNrNqeCd2EpN16CuIbABEqr4Std7q8o6
6xx2wXu4HhdWYO7MCXmHKKxeokbCD+ooseLiwmIzPQPrFB6nP8EHMcf68Wf4K3jx
fFiRcPqirqxIcCTAqrNNTHAxI5lmSVYjfmxeT+j4uYln4NSs9maxe1K8Sd4Zz74T
GjY0uu4begSLdjttVKF/H63F01OOZu0SVhZJyPLrSUp1WJ+fNcg4joEiNTqiBv4u
VhvirLHmcaA5amBybwsmzEEsHq3rbbrOuM/NOqvIF2i54dvYw3HzeuDgstHvcwX0
w1/btAvp1L5S7Qlx0QTXRAUcJBYGUfH5tZeG2ux1S9/B0x60zTF1R29qBiILjXWK
RECSm9Q4Hkvqri43f3D/09vfXUopmXeU3PTIIy4vRxbGNzJmSS1cBR5aIxbJEFyG
YzLXx0eiuOaH/54CTP6THJ13pYxOCtLRjGXPGw5ZAgQIEx7XAJSOgcIT5725aFHZ
su7oMF/dyS0JYbrFZzDnuo5UXv3kcuDOLFOqYG7rOp4cJ2yn6uTgTph6quqnqCBN
0djKJFKpzHAWbWcIv6DSh2kpnJBN5gekcv0mF3twyuryYqU0zTiCMSbS8+qnAdI1
zAEx1ANc6dXisQFxqVenEeQPQTJlV/6eUV79EJ9ftn6vXmJLx109rMLBokCXiNT0
wvUWMffbWBWLHTU9sEaQ2LWaS9hZKF2i9Rfz7ADn+a5ilmRyuCFd0FAZA2FtPtCc
usX9/1i3B3tNERpm8baWseqwYkm/dN/7GL5MvV3cnWu3ny2MKZoYyEeun6gtJ6MN
+8ACpiz9rDJBJdOMbG2u51WpS8uD5Uhp9adLcsXFcdFWJmlOXMVozIihshiWIJeJ
bEbL31B268Jt7WMJMEswvX44SJeJV6bMVmMiz7sMIBgr+ZLqFw0QAkqnJDf/3mld
12stGveTRSJIG35qMfba0RPx+WRhEST3bLWrSlHuniyJtZlzqnCxZa6Wreb/7mDc
EyjJf9y9+wtW1d/vYRkcGTO1Ud++EZWqy4S4UIKmf1tEGE0kEf22vv2T8fMI3AEw
ASiE92bI1tQ+jzgXVMQg9MJduxw5QOgWOEu1YcwhmSCfJCeR4yNza7pBMg5jpwQR
n50KmdWNhB05lWLLe1SToFVlq6BOgk9Aprs05lsCOMY1z1EM5f/mYzO6c/GpUw2s
OJ0Ev+5tfwtTu4n21qVg/hR/iE4z4bXZDbCYHoW+KyhH27eE6H5TnhpXqRKANEVQ
kc6XT1va/kbgTQwzaEzfm5dmA3VcspRDLvmUt7mEJj+mVN1NPFgbUb9Qj7oF1z4C
tiBx3QJJy9I401Hy89jllEUAlRLLNxcJk2+MZ52Zl0+zXf9SWPdo7f7a+xdRZpJh
jSUe8hR70oCI9eVtLI4wGE1ZH63kAbxZywNDgZ2IKPvwa6iAAy/OfbexF/eKc58L
p6QPExakEmqtBvfhWlhKKaLEa29Si1hlkclY8amBxvrpqXmxRE8DXxXtPqdXz3yN
R6Nc8cpstZrULvA16qFhR1c0QsUjZoxQ2VyNUnSy3d+ArNmpNjW1Ml6KKky8501e
XR8dKzRTwixljcc6iqxAZFyNLD/mnsJCFsL7owolu8ptZc2as40Q3f22I83aNM8o
HCz80mFHCCEaXg4WeAba+2Z9OrGMfiyvOOrwr70UACN55/isYwPCO4yCBWb/hHle
9jcBsmjtG+64RW/I+xm3DV1R838waXNnBWTilDVbU8g0STx3jDZ77ESxUTudf8qL
NZugJyMljI6VosFWb49LqjQ63N/bTe20lfifNAMx93QmG6oBcJaZUmamBSUWposq
VuipCYuiS6K/lpKRjZcSOlOIdlnIausVISnw45taTer6XIatOD/xKYWlwYIo1YBl
swLcC3x9XgybgGbL1nlHBUJH5jScSgz3RDpyLSUtPnuT3tVPiLoG0Y2Xa4yZ+gbC
EO9AVdFWiolc5PYt7isjxtYCuELq/0XbDIeeNnkZX1jFDmhVb5jFDwa+0aclrCnY
e4vuVd+CLQB7Yn8p7wXM5iOND5YMnxmxoK3WeWkTaROusUCQFV9D4rBiio07Hiwx
8q44TgnkEee4NPGHz2Tb7bBw5Jnt9aWPE135G8bBf5tXy0v3SzsP4WIScTXHcfP1
3kQWvk7eaLhdiAL3mLl0YljYY4+hnOSnYWjY79rAQtsvQoMCLivKr2WD6nuORdFy
8VzqZQ/OsdG7pS5pwxZfaUnLjW90XeySKw6BZ1fFDg+NnFBHFrJ+U+UHdPU61de3
BV1Brbyt8xQUThwgWw7y93zKLdihh5bNuHX6FIiWm+NpUKn6A0WOoNZZiJbFlx5N
VeBmTRG9Xuns2QXWZUccUd5NL2v5FPg2jzxpDcOMs1t6ShN4Qe5xzosbrsgVS9Au
8x89Lm46GqVqSmipA2HYCS1MPDoYQM6DM354CDqQ8xZ/zRb5K6Q2lNONy7QngI6x
AIcjqsJTE3GwUTg5yO4TlNqsyYGd5xpRO+BG1oUqglSfcT5YKMn61VNqn6Mk3Ov5
845MHVe4RU+nG91UCf/U2PzgSPT14k7WJhXz9Q5tLGKWW/F2qjEzJOaOGfCvj1ci
k7alti6J+8oFQjF6YJbiZZARrXcYeuL2fpgXmWzwvoyGixC18NHU0ygw9LT/cCWA
UNxODS8MOQTr7Z+xC8rzdqBaIXVUkVf1mEcKTC/gR4yrslNq7gtN8E2aq9MxQenX
NtvBeBwhM0EbB41dXkHT6751IgMKq3gdkYNn+Fd40qYVBOLkfweAi2XkteSRxDBC
+VcIuGYdC6FCmv+MM6V8KtCfwzyXfzu9orXoqGc9B9Mc8S58JGDjSibG5eTUSaE6
z9CqPWx3i6cysVVk0/127eJaN1PMu4mhSaZ/gXrpiuMLLvD3tLmQG0XoOF59rJYu
DjsVJd1ZdC9IlwlUEtjYOK69RQ9JjA7YuViMB3u2cZfHrX5am7N2KJw1bccHNuGf
twrz5Yu9/Y6CV/LwqzAMUy6sGZC+M+E1uQL2sLK2t11pJwGoNFCDHsTe+WjV1yQR
d77GoLXEFmZxNKFh3K6066Y1Bu4oTJZzLtsPZfes60dHT4KtCZxc7DUqQ12y98iB
1LilLKJ3Gy/2Dj6ug3nFaGHf0JW1W38qqxB5mf823Oo4M4/sjebYIGFHdvdf55A/
RP1+Hr6Z+k1Pp+mdwnttnRtbbOY/ojVUTggNaciFINm2lsqHwc/KbdeRdjawt/t7
cW/bEdohqt7A6FBarKmxC6rWI57DpZTqGereI7/+602yjG/4z+HmkY09rwJwOW/z
9SFLGdrCreHgV62EzMGwSB9BupiGx24W8+xeQjJ84vSsvP/HKZg0S5KJuM4LO+Xc
58Dl9R74nnHPPQoTqG+XwMSH11tNkpgMltAUXTmrox+TimCU+2ddcuhPbL7/6Z8x
8wThMhaBVFBdDtyCScB13u0U+C/Q44ksjm/TnIlY2pJTwzgkzZIgWlr+NZUMpd5Y
aHPEZLfObcTvg+ZjTGsrWXJSgb/GAkRrsaER4YX3XPtwdjnLn/AVz5TzRSxGNSyE
EzCuk/mpH79OMkpVzbt8DpwfB2YbJlVlPwhXRVPPV+PYZ0eOJl1b+Ef8qbUIMjpr
X8xkXi+CuAFauOMo2ntJ5J6B1e7URX6fUep39S+z1Fk/aYUYCdaBP73LMEPUc95F
823HV+nvrzE4Xb0lSHFqfz3LbxEz1pYgipC6PIoZoIXwalMgu/JYcznhPzLlm5yz
bLD/R93GW6L0wutXalI9Ftz06mqbLtbPiRwZMxsaolNevLty0+LQLUZxf5i+abpl
zrgFE0duvzbK+VcvznNDDIQRH6nMiPphDrDtQcoSwMH6WFoNCiUL7AkwdMBQLRuh
LMqwqtUvnJ0e93ej8i6fQDRNBBFmBzyX2sHfb6i3vwNYLP5rIdvyxsbZZRphnUCT
JAktve5kROjhPl+0qckoV+JJj+cFe2DL9UsTSOYyHyXncNOvaU71SbfHJUL9wm9J
awQAnhxjfjWWcLBwbRfNTY0nHIPf4MlCZyFxnyKPfz6tBxGLqkHEZ51+DyG6qe6k
Q1xhCRCP5YKOq/12C1cdGQXc21FhBukKDgq2rwjUl/eANiWeH7x++05R7OcW2Xk1
WTX+5deMfPjrhlbdTO8lahLGnqLWgGCDj9eqyORzNy06o3W/TEnGaPjvwVUcD3vJ
SdSsZ15NxtMIRaV6Gv5MbC8oCvRAMjS9LjfaUg0u9Os+G3QOM89uU9bQ3RI7+rjW
wnkV8NO2bzze4PePz1CUaDMUVGbqLqnOP+VjXBBTlxEypkeEoBlnp7Gu9GnyziJL
QzFhJulA6NdnWChcarP4eRbpd+9x7sV+RqnwUU7y5JxJVJsYWKgRXI8KCRsjLb2n
2Ss0ROtJYKLDCHQ4zEL4GzOMKA1Ai3MqJfh7vy0crWG3CTTa8UT414x5Gp+CKER1
C8NxafKVxRDpMZJ+lh8RMFnvGpJC4tMMxMZ0DvtuL+aC828r7nJiJkWGGHw2gOds
i1BUY4Z9bOsR/w+ckO3+Zt0++zfDdMkc+V2/tlerBAiJizicfu+z7OVv0hscU3v4
ce2wafdE9hzu87BekBMg00gn01MJfn5sZRhDfgu9R4NEjMPd44g9vCNQJX1t14W1
vRqmzFq2dFFyOzDCkUVQc9DueivjJpIJbhlRgNYKV4o2r6q7UiPeR8Qw/5+p6ohd
TYvvOCxuGUEwCRVZtAEspPElw6Ejo4SJQW0ti3Vt5AJZxPNsFHmyKYh9MV/YknLJ
ZL1t8bXmOuLqfWuMz0IDjcqkVlPNsABAku8dJQd5bs1ikCA2GvHKnLEn7wRGsu8b
DyDspWKNo4WzL1kEN7FqbqjdiEcP8SEU4/Uyk/jKqdDFix+iHBH5ZkqO6iyhv58r
Axv4kJ64BdxD8GNoZ7cjCRVGrHV3QJJr6RhNYf8YnnzXKUWBnfa9WWOnwNNM1nBi
AMddZ513KqFkrBlB9kRMcxrQgX/Ixgxywu6oS9TzZ1dvDLNxI5uRvRAR51kLWYgE
174ggQZTQ7NFB6gSrzL6z/jNzJedF9buW4ncJpAjLeB4objt4mYFdTAUA7kJhoOW
+VxvdMiVSOVJZPRj7xr5wY2Eoeeb26nh39MqvS1xGxGz+2mOda3/5q8jJklpeFaG
+3g8+9J3hSyEgi9jyKOweJ+jziWobQCDC/csGzghMqH9/70r9fzQwU1ToARTbSXp
+XeJJu9jOBd5yOAb25UTUXtLBuDnTFAgWghiCRtRLKETay/DfjE0NWvhF0buuWIx
jkF8b/FdPanX9YZKSRuHQYt02gPNp4hos8AixQ1EpeMhwL2H0nUiqYh3Y5lqlu1X
vQMHC1kahPbkz2Eqea2eTbhJoV7+V3okxkw5tpDsNSr3z9vC8/vmc7nElD73EiY2
Wtdu5OnV/9J1vMByCDBe1q37/FouX2Ou8CqHdKAUVeL50sJZK1MUdPz+rnKDAWxQ
ZrjlUfsrbd9HOnOlIx/4MEZcGlP7RIV1g9i7OyoIPhuWLmxN0zpophWSVmIk4vq+
qhpXHFDiqoQ8Sx9ivj8sux7POkeh9im3vOqgbu0gkRvOspm5oYL4gOEznWBeTopy
yFxY8EOZ3w9Q7mmrUrB5bxg8nV35wE2MTnbN1tlo1QyTkwzLg4p4yW/Yc7v2vie9
/CksMQta5qPUZyjrOwmprbARlqguyPI4Nx2tL3i0lexThJZvUc47BH2ufxVchix3
pUpK0k+MpGjeautaFIVA60KR9OTLBDlKnaLFYz5bvLrBKi0Y3lT4myOEuwcsRq3y
4kp0dmMDtfmqAA0PVvEAQ/v6VZiq8bv31bi6oITltmRuc7iLB8lDSnbd542FJMZV
XdbTerGPwbcdPidI2yDoQXsw0evNJ2tlglTuuqg/J2ibIkojow1hseTPoPOCJnH+
3YXxfZzQovrGErmCkXqA/h+Sh67GZEh+r6/3TbUGRQ0BOjHwEE0RoWJ7HC9i30LA
Gw7ENSVq0eDi1hXJPsXAVntHq7n230hVx9UN/i+WDdKt8MLsah0hjtoXMvFJTPOc
Jq/lBlX6ZGrD9+/BFI8qoeDb21XMUjGNn3PQXS8SL0VKOApc0RdrAM6MRLPeXmZQ
S/9NbW4FXKsN24efhgiU0OwMB71SE2WLsI38oYotjWGlxe0y4S/PkOUcst0AfoiS
ptgIbjgU82/sYuDV6URv5Tz1JbQZhkbe+STpZrh0RIilIvSBv5Fha5b0G9Mh/e4q
Dys+FxPztn5z44N6nk13c+d00yRxJtE7/Jr7HK2pmSJh8ZtrhXCEHir8Q1mtsdCZ
4PvejbV8mNjrbuSiDlkwhVcknTRe8BmFvLXZc2kphGIiqTYX2BGsINrotfl4Zup3
TwAfU61YLTINcJQmq6rjA0/qNkaALagM/VMgxsx1j11G9XdlBB/YZy4R4kZRNjfW
v60+3y6yLbXzULlyUL2BZnfCSjoXSY6ef4rYwAeSyrnnBxf4bKPF1eQps8H8ybru
f2OTuQJgOfJWm6ZGhtNaVNd9g+oyL6O6Cc+jrwTF0Pr2CkA1OBpaKovywYKDwSwQ
gxJ8HII14ZEF7AIAS8m/cpUUj4Z61hAAry4bpwulutzfqZoH7XYP2ykZKbI4xd3a
EaRQSuCZeEAQgph1CtMu/FXJv4ab+eLDwe+uR/ISiuDuAGU5AScFccd9lKbPi4xk
Q+LIsulVJO946gtTWQHxqFyBqocO+jCQkGSeNZppWEhrf+czHks5DptStqxk9max
I9b1OSVu326K0cZferDKBt67j0/cBBbmF8ZIJMSJ598/DJd7rF7woUcpU+588Y72
FJDFdvZbokXCdHsxy4KPKA3/hS12R4YUPOrBEwRP0rMRE29MRbqcsTicimDnqrqr
gBKBbCjPKdgWIOFWWyc5jkjkX2xiuTnAapwTFvJim/hsu3b48tprw8anX1HDpHht
vBRymnVds9hNUolMiAs2aUkofN1qqo0pBYNHhXsIPSBtcdKr41IiJXcDqy135X2J
73VB28iURSOnSmgda2q8sTAWZLfSlpdaMfoN8mPM58H9LZ3mjUyi/ieEDLJFBa6s
nftJVHlwCAuxIP7pVAAtmPbWyufdd0bA9o8mf0y+gcXyYv23lCFexWBbYrApGB/w
5zhO9aUaWxchAaHXLOkCt8DJJgSyPZjBEcoE49to3c7vsGuxRJvk7B6WsNjs3ueo
h8LockJDmKP+BdykYazeOLGx/f+JdU3YQsIbEDiuYheN3nNBmEp+to7L3A7/4NF+
o2VqxRlPqSLVWEP+AWlBv2yCUYLnmq8oLRlJtw1Rl76zWwZMUhAYzr3dJgQpjqTs
8EC6VR1Zjgmd1fw3t+G5sMaxZH0q+FfKxuky1NVUdXjahZE1cTgAmUUT9MXZCBIw
GbbOXAoGQGVu67dUGjhjKdDQmvh2h3wU8nBlxoXGYJwQDfAAF8pdaXVk2SOyrukO
5otMEaGMkVqpRYp0jiYoIt+36u86gPfG2hQG8yU6qx1byEu2hHl6eZVcmhQQm5pp
D2lcoQN1GyRIytmXUVPs3U/IYYl96ecIRPxHxDdGGDVqzvDCjxjfAmFu/zJ6IBuZ
Tb5BcOK5KDbaz4Yg7kL/FApBcZZlZRjGPFZMPUWZMitarIzWmioMT5uU46d0oaIP
EOe8RaVvmacNuCdkNpQQ2qlMLFQuvdqCE69DCzc4o97XfrW4wvcmNAtytqSy2Rdu
4l2SfhX15CY2pNaOQiMNZdsq3YdwmLn3919D312hN1leNCjT7YLN54zkDYhJbM3+
32umnvpUGlq7/Yly7ytp3grfaIpL5R4np7fHwoTnsd2mHCjcZF8sbKNAgrlLV9H/
B/58RRL/AKwh0EGL/PkkTIMGc2dNr2XxCT/SCCP1KSiYqVOWbJNmq0Vgn0X34t8h
K+QGqmR4Xb39MqjmAVckj3EERPgJDYMva86Xi6hAbisxFYLofGaQMGeAzw4BrzgT
hRxEE6Hkjunz3HL7vVdPceQuhmaEXNDB0li7ySG+ZDKvhDoE1oeTNq3VhgSCpVQw
2b0LZqRTwH2fie8+oRPs7YPEGthaFYBJFX4R0Mt7tSLRH8wtx+fEdeR91xy+pNIH
fTzf88jvYoCms2ZADVIW8C1o1QPdtDE859IL4bwRqYSw9Y2Pqt0DpoEehpm2sNAO
YA5pwI9JiW5nNA3U/Qo8t5ROC0dSyQGuv0txuMBZ942B5nFQOeRIyt1XSTyLK/qO
TQAf4k6TTeqOXBVbzbDXs8XaBVuWJ8nNdn/QW/zOOVObKthXZequ/R/DKBnQc1dQ
z0GLuRRiBhVPfuetr7m6WGHUyTSep/IV/DW36MNXraDZ5PjZqG/3zkJNnhV9j91i
dFJEuYsHcPGmp8mai2BpyvYKzZorQDNsd5PiYYuxeBaaYjpA6kpsHT09LjDEBL7m
TRWnQvVbxuDHvj9GRN1ueSnQt9qo6cAfkgmYsj2PYI15Xhch4CpeeYHW4RJNIZXC
KKIIbeo3aFPKe+z+5jUti7MyD4gVQpn5vv3hiZuCf9SvnNzTHQ6gcMyD+y34zM50
ziNBHt41zW+o8JXSwl858HScstGNCX6xTcgHzCNESeUeWptFj38CnvJEt5GQb/PI
u/QxfcxLr6dlQVsLjjtjVprcrLQv4TRUaLQpiYhthvFlDfAj+7MRdYZz6OBniOmm
A8iBxjH0kWDxkq0Nqc2QYImFjq+UsVJUXbnB2BgCs6cDM6IOZENSf7mhJvC8+A9k
xxsvDVHm82NQNThzFURudo+0ky4urU0xwwR5WjIGn57bBEX6j4ti7QTR4Rh0XF3T
gzqMtFzQmxJFd/vLGtmUk68a/X9tCiKhLvtDS32X0Fw+ivHSuuqJ89iSItkAayEf
WE8B0AKvUf0qC/db2GqpIA3hUeq/jBdvZ9Ek6bjAR12pmTC8K+/YRym3ORYrBO2V
oqBck67efPQDTvWo7lvpO3W4hUP5ppszXh2lZim/ylv7Znsp4toZtm4pm9+ltJN9
uX5KnyO2tS0kMlEwZ49NOiZEtlB6yR7KMXybrIA6Fq/7eEghxpeCBLKqwHpeIAYM
0IVuDiawi6Ia+rcf1tLE+uTGA0btjHREyU1RHsnQ/6VgjgEwYiBeGgL9/uopBgQO
EskqrDMiHjGrPueWZydqdcl9lDN3SfI21KEK8sTLSojFYMEOvC70XS3y9YqKTzpa
zE5zuBDIwQ9/HRUHORWF/Gjq3Xv5m3xrh4gaqQRPD83fmH3Ff+0tEFheSLNsPtUm
7UPUosmlsd6iNCrB0Z6jQ5WzwvYk4IuXgDg/KuLT2DfCQg+5xcraB18xMdp8Cye1
JQn9xOA2nwChPv2+ScnnlM6CTXXMVi5XasRnOmzjG4b5i/ryjYvDX57hL4NQqXo8
oJccysRyHeN3BIReoakVmibYuAaNqbKFuBlGWN2BoTK+3Sgzo/W9Wxif9pn6VHYJ
U6cYLeTzquk6EDXWuVt4izPNm5cWtYY5A789ubgnzT41HzijXwTHmbeucxJYrelG
LFBHHTNoKsDOJd/EuED0zJJ9qALu8j24agDx4N8KFfyDC0IzgW2aob3ysdgC2j4T
YE7jZvpW0deOGXQrTEIjM2x++v2t63K7yVP8SoB2Y8pH9PswpF6Vk4Fm0XzFcikW
z9z50SBu0rDNxLNBY45BNx9Z81wegxzN8/w76ccwGyzJDQJuSlr5N1m5R1iW/Yx+
SVhVD0UK2wzYxUM/whkjAUPsNfwu5FYYPQLfPjMC/JffXg9spdsiHeffgh1blhbF
/yshT4DEVOLRVAR9OZUWATQHyE0G/ERX+zYUWdhC4bzx6azZycgVPZncHnjmHiMF
TLXcE2OzojYpDh76VPDldyy86fHZRdc0F22TJNyD/bQci8V6OrOM4x3S5uOmYQde
2844ZJYKRQASjJBNUmcoWTSbM+S3ak9Q/DYUa2dvO7dtM/OEvGzqq1+DgZITIXPY
TMFdSaLhcZrUsM76QMN2pB7/BbB4TX85qkmoLkq8jGmnP1Bq91yGOMPhKtZWY4P4
Ih6s0dxQcvza+GGFWEk/aMgol7flJBvTYMannFFxCmh4tf1Q84AhUskeXF58W094
eHFaXMjYkCYnLPUebqO9l7H8cx18K+RHbYAZBG0iDEtgBO74ivEANLvbPQ2/JNkc
oLYQp58atNl+d/NRUKe/ufbe7ZBf9srqyjJsO2HX1xRHDk5/V37Uv9o4RyQTt5ve
DxMKxAJcF70yY+Wfr5cd1GGUZlkHsmvWVRp5BAQMNLdRTkjUMvsMfZnMhtHRUEUY
SY3iQ6FqyL+Fr1/fbSHawJz3cK268UpFTIRxIrHF50lENZ74mSgOHBUx0rgd3QXr
U0AiemXale0e92Sw9oU0IcmffX+Y76F++M/JwWdUiaDuy8Lh/ktteHPZuLYdmUdW
VnWSCsLpG0lHi3nvh83lUJh8sVsXGC8rUYkQL5hz3mhGFk9B4NCuelo+BLanibx5
oTgC4ezJfMkB62NgyPEsy43OUpyBA3gd37No2/pA2niOg5ORZgVRy+kM9ApeK9Tn
EiLymXC7a2jYp7i+3VOhKLHaYU67FSaMZb4I+a0BjJPZOvyT9CIW/0KN4wzG0Cc6
3fYwQfCBgP+165ohcn9L8XBcLYk6hwG9LyRdgaaopqHxmtt9sdgplPNQavw0bMbe
8TVigVVYNeZTVNG4qXN2v9QfToJ6Uc0CtaRJbA2RDWg+MyAqmTqyCAMqRwGXGrJ4
jQRlmgZfBhaMOsJ+SaVdC4fXEZWsFMqe0k+Xw1uInuQKpE3K59z7wRzDDSobzdDp
EOWeoS2N6ILNQX1i7S7PYfALOuFrqiyDa46RRqt0w49XFOs1cfUKE+lfEsm5t5nN
czxbA/lSzL7FZthWVf1vdHzAMSVUHWnerBibPqWSsFAbMh0wdMwj5TiaKZw2uO7R
xad33bk6HRz9IyvnOOxoculWwUJ51o1g7wylLpoyZNl9EZvH5+SpILfRf31n6F0F
tDAMBX15LCEsNRspsik9czW7P7EkwAaS/NB9WJQlZLhh65lp+IyPF/PyNSLBHnqM
Yy+18J5UDNNcYd1O04XmSu8x3krJuD7jv+Z2XuH/3U5Xxgwf/W/e43M6y1uTDaw2
Fn7AKqZWtS72Pk+SBddVzU34vWVBDjIj5bdHqwho2/CBgsUdqa9PmvqFGp2OPjTX
W1MpjGSb83eIxDlKeaza1WY3704i1UPnYpPLSL3iqBqQCTE3I3PYiVGhYELrUdMA
kIfOOWwyLKlmCMRoOgq5w6mloP8gzI7pulVzuAtBrvrXgZ15/Jkala2UETONx4+H
zd2iD3HV74Usv9Hf6kargROIjqlatAhvZT9mbMflUo4ub9q5p4zrU4aly0CZSg9Z
+e6yl1sMP8ZooyH4qBZ1HV/8dd+gP10KjO4YadgQzWCQMp+c7Or8GGlgXntmLm/C
R74pLVGzKkEIMm0NMwLLe2Ikg9MG+x8UiF6cbYibSeyolkkjlxea8YTr2giv/BfC
RNHBaIX38ecSQ8ksWScNM3zBFm1XMk5UcyLhTrFQy0PaiLR8n5tyPy0BCif+YYXY
y4j7z34ElSN5ZnOcobAYCR7tXg42SCBEbR8CKPNtgOVZe3jW/ucWCi5jouNz8h+I
Qpk+NnLK9/iNdJCBylhsKtL4fwsKlA0OCnntbSe4y60v/+MejNJFM61HUOK8OyZY
+7nypBqpTWpC6ZeTATZ1T4U78OuubuLWiEEtwpVuYRoeFHhGovwa8rXh7x0qxLvs
GY31GUIDhpOgHCPxasHelARA81Qc0diQCktTRp5LF+b5Bxi/+56cTnV26nOnUHR4
HdatU56QkboVom/uAN5c3Y5w0AZTq4XlIaz4Le4C2W0QTi50hG0RhOUJmwGVeUPo
TUKm+htjKT7/yMObR2tnDeiD8QpmxJOy2xAZImxKoa1gyiW3BQxlWiiw5y9ycT+Z
nEWzv6nP4PLx2NhlRM0MrAdAu1DcEftGn0vlVa25A1F5fVnoG28HgF7oGsQCcApk
L+DzUxDujamAc33sa02PgY0JCIKQsXnggOvHRwy4sTp1BGLV97lTOShD9FSTTZ3i
tf8gHSZtoVSgiatCeVItLVeImq2j/JoXQR5NXjYmBtXu6suzmXSMjKQHHHve/Ywy
+pc/xHwWqTt8kQTNeEesBgwQ+7ok4SPBn95OxUF1bZdeIGq+lTNtDa83fRCdYT10
+9ui/jf/LTgWudlbSR59pZmX/4LzirEzk0UQc/RYLGVco+b1PO/VZJ/NPgn6RSVG
eOQMgBJp6tQDzHPxQIYTCoVGdP66+cA3SNED6xrYK29YpIHwVT4543nYh5oZCShA
RmBbntbEITC0/P4EqPtAIrrTRjweHxpoMJ+7NiDBl/4KlYnz1mLatWt7aeyUkHiJ
OkxjxBuYJ3R0XdHiRFR+aXZ8sjXxarOXP1//keNP7ygByUkqGTyZsXUsPpbO96Qq
GiKhnTy6A/JVTGIuOLIRoWxd+7NKbvAOursVp2x+5wQrPMpkGarCiiA6EBPfUONk
u1Rv27kxlwNPzFLfP7K3YVx7er58Sz98k21Fl/05wxQABWXHyTHpP+Xy9RxQUmol
7cFhGvKtXVINnApGCJl/+vGVpjcgfe2TekYrUlQm1hwVkmg5gSqDP1iTDDYur6Vp
UDRyhAkMitgiSnAec7N0/gohGroN6I6rPuDiDIf7i36hdi2jCmmwSfsj0QO6Wud8
1qbFu/COJ6PLALMJ46DmDTrvAQ+olK7Xp4Q0wiv55c/QY1RWC5OdISbpo4909oIU
Ir5V7vLxbdAca3aWRq4UPLIxnayZexlWY5Nb2TCLcGZCF5djzK8uq3gzwyfMeOiW
WGf0PeLoh1s5S1nJADRhCn74u+tp3+bOtK+F8uGOMdmrhw0HZmD4VKdNPLR5bO+S
bAGMbfiP5iYwm+W+mpf9wDsemPgcK4X0NuppUSv9GJaC3oiOwy0a42SGsXu/UaGi
0ZJaJGLrTmxoDLxcW4Ew10eghE7DgMuhT9jM/WqxOCvL1Lgib2P+rdN+v8GJaPNn
olGddNyltdGS3aYERNSp8zCoN4Xh0OtVwsXsd03auX9plAbR9pflH3Jw/HRlVoNe
Fxa70VpqnLMo78FRpBoPplmOfi8zLCz+9P2lkt1HcLlvX3NJ7ds31wC2Ry+0JX7d
pms+n1dymPnTTNlJQYNPPvRXnXr/Vi8R9wI8HgHF4mbffMFC8wSZ4Eh2PDJlSA8K
frVbIgLS4fbNDm3WipwGUJ0Ff0hs78F5bqqoSPrUZKjZy8WTKmctDHfIhwFzp1FO
S84ipOtPF8S2Ly/oL54vKegRFcyBka9l+7zbbJBLDqdYhL9lw8qpMnXQykqfw55w
4Q3lSLNiUarWfVx2b/VJzD7JEn7pbe93mXXstd4KXMdi0HIK96Ll16eVl3yjq073
09WSM8w+B1EeIbSJKpdkgZ/joVNVSqJyxYecO2nYWTJP+4UfCo17gfPSSxH2+rjk
PDr2hnMpPKleDVBw6na6T7TLGgp6oIomJ6xmTkHgSre3ZESwlEFVaCzPm8TxXsc+
XUv2luct9ML94qZbnOX/V4marrJEDVMQRks/O900s8bH4KfIu/8TG2XrVe19QJ9W
A4kH/lhFF7iln6uB46BZ8moo1k0S+jbjei3rMhYVEdneefU6CdpQXAZPobz6RtoW
1FS2ie0U3n3BMhPV2bx/9PZbR9vYNnxMa65GZMXekq0=

`pragma protect end_protected

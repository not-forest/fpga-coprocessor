// (C) 2001-2025 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 24.1
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
Rgd0zl+gw/A9HPS/y8m7oIdhulAjodTZ9uVepzSuZkEl32cNfMawnSDohJ8DchCD
4/Cizwm26DS+WE6fu+q7PODY9Glp7plCDQ4ILj20s+xFuCAe1eTpw7DLfFmdo6zh
1bbx+QQeyrbkfOE8q5RZd+Pu52+wjNFqzIdDNvEwWNrqEDz/eMLa0YuLv5zFbYPs
jk8P2BPdqK8B8ITHqlM4k+IEIFMxcb7CKYLlMIBU+kqGP2Ds5hJo8NtOcyQt2A9n
8tcY1e6vPxwDbAD2SuM2diJP+6hwWhR8fEqW3MyymV1SxYW0kzrf5ADDlKqABlbo
wN1UmdgweMcQnbas7kRb9g==
//pragma protect end_key_block
//pragma protect digest_block
l5WHAqe24jul49MKL6DuJ9FxcxI=
//pragma protect end_digest_block
//pragma protect data_block
MCKNky0nvxMIOXmjaUCLSaUzJ/VX4lgsaLqdCOLcGHGWzeRbIOBbocBsKzKuIDsa
w6OeDo7Wbj+LgigeoYpY6KP0SYoAzyUmciRUnbBuFGHo/PwE/1pQZcS0XQOUQ706
6td2PZ3WMCyJ+M1n/884NFygE9XV3iI7x9G4bR/ttgyM0AlPFR8UIvRj2fjID7JJ
kfA3LII1q9PbbJL5NdxSKsFYaQcnbzO28TPUHx2KYvF32EnvsHa52+8uopawQ0Lx
Fw9/N66UOk1DIRokiRf4oOPOvaNrLzcKOixRPlw61hfIj6xkBC2FszIwQW24XDMn
3wZjbFmoxgHXi+OtQpGpvVnO5MTz8vPcCt3IYYesS9cdXYM9tmRlLiBWlwKcVeh1
uNbUmN1t9JikXz2zeUpt/75EMhNHRw4v9iojukmJcD67hAI54oS68LfGfxym+mPk
nmoI2jcFkeOnCqskVd+Hxc6fPMHhZysxmlwLCjgBO6Ge21KpSp3hN5g/YpPM5EZd
GpM75whiDlRKY7emIcQL6XPmqi7soMnLwg7XUyqyAWrEHxCcxlW64x4+NGLylUDA
bamO6KN3q+NqHTVSozxjTG0CFU30+/jEmcsBThy+CQMJu01L9SQc4gygE4JCJtrf
7c7qH/HcaxqlnA6RpAQS7Ou4gz64tV3jc10t8UxZqpmB7jt9ZvQLan63sQZKJZjJ
ycHipUGG2EJDCc9R9ijjueo987/zf5C79csqAg9qKDcp3D3Iry3t+ZHXMqoXvhXS
VXFkvP2Bv8D4XnTeLGthf0JI+arPzO3fiZcyvS+2wje6Fsny8qizeWe0JBupp233
aIiH8U6aM529XnnGQukBovk2GylSqx9haX105H/esYqDcTl3BGEg2HH6QW6cg9mg
X76OhtgvNi+cA6wzZLKamiul7sHjJaqRxtfNY3EoDHoNWtlLasyjdOQk64O6LYBh
QcVnPxuKNiKempjkZtd6ZJFGRqHOAGliF4ex7FgztMhqVJF328A93NgUJpNGAoCt
OX0aQnUISmcWD+QjFUDR4S26VsMxPjEvADfLlI0Qd/XD+SOjn8ygfiT3+TCutIsX
8Ef6y/1qbdCXXhzMNpfOcJ+C4J5eYcUNzb+E2wh5wErlPHE25O/5wVInNlRGtyPG
I7QwqUcwcC+4zrQXp3rHE9lKVSjLq/y652FaMScvj3zzGXbeh32lVktRwtzJGLdf
V6ZgGJ2F4FHrTqVMB5Ti1Gq+LpzbPcSY1mSDG5tXMrxvujNXk57Amik1ITp5xdW/
L2uFeEtFFYoEv3hGP6TYwsretCBvqy0yrFs93w7peaTbviylh5uqB3pjt5pRAisp
Sr31GHhbetYywUNdACOtWar/CEdruSIOTxv5MZSxnVNEVlhFGmM1ZoPC3+opp9wb
wxb8VKAzsH04qvTC8W2GAaHbdtAevapBcOK2duJGaVtLTzZa+KAfBnz34p96QCu1
EE1BSRChzoRKiRN6QfjXbGbwmdgNn6XmjB1r0RyL6b3Ngyf/N1r9Q+bNUN46clOo
W/VDRKuaGfaTOvfPNlIXwWDVwWzsHdybJgiJaaQDk13jUamIwtCa2HzcHMBPg0FD
RzsOMo045INDLJQD9rGqCqqKC19XmhJagmJI6PBPII8HDqYpkFgUj09lWAXV2pqj
Jqe8nXnfSPihZ6xWXmNGyCMfMaljLEgg1RTmTU6gBxa2EvKKbkYDJoJLzCJ1h+s+
YHV/n5hq0Hs9MTdhrCTURTO0Ni24kTlBj6IunJ2n6zDG5lITrkhHe0XEyrQYuQND
1oCOQ9oPqdaCiqhabVsb2C6RaPsxeI/4i87AQAYlBxUcxBknj4R/xinmOY4v2Dvg
MK9s6OLZlGNlaSZdw6Bl3db4DmxyClYaZcVeewBgE7V82NUBNTgbsYwkj6Wrnwyi
lN1z+NkAK1XPQMm2+nQqMjvgiSGRjKhoiVPkiSY4aTVP2bHZoDXyVGui9HEIBDQ3
OJlirLiBao7ywcXFZayOoIEUtsiYAZ1mj+B16Vn8M874p+sbngFwQmka+ThNZSye
TaJOEb8qMlM7s/9AiHpb/SIbQDgKvtvIYB+AUFC3AN34KvoorpKMaGKoF6vQNZZt
gT7OY6ROIstSfd+oJXtLFSkBofFMBwwexd+K+a3Uzu9ICipo5HWUSgp2u6Z3JU4a
sFHwl7t+/puvQyIfrse2Z43YwMQfQ7dlexLndMAxEXs2MKtgOhWdY1+4OHIMagtB
isA4dXE9wvPqO0bHBHZkBdgEj2C8cclkjBJkmMs5IFsRLHZP/BBXvA+tzm0p3ia9
V+RmpoOoYjt1pyK1aMUUCpudrgSs/d6+INb9JDMdt1EUVoJjrI0oqtWOFtRlcHnw
7uaOytI5C7kWZIpS2OYnhVpbsm3WBuzCObxDTQ/lbDSTc0+a2Pmj7lILOuQAwvTW
hIAl3r9P+ErkXXGoNKjIm9LEo3BAIqgUwLNdqsjsR+qN+4T90Hea0dZfcilD163Y
dvJTpzLmFREH0IRocdPJ1E3Arv4vd56nnX+x/X4GxthQqe5JY55AxZQ7DIy+dF+v
+OvA7q+T88Wm9ReYtk+EgvmPoS3Q0W0mzzrWjR2sDvN1fVg8F8KBzeEIU0jbRNfF
sOfGynAbkNEt/qBel/sBUnQXiX0IG4u80UWncCN7KLRW1lNhXC/rApn727+1mm3n
HkvgDAaAbdMVci2bBfAL3eJEYlQLG7D1POkueDQspAwanhMAx+ZwbOaQ8vwbpO71
ngFUOt/U2J8AEp6xbFZeiqB6r/rkWnFwpF5wK6H3Ikuuw/UrnFLYwWKFg6KbH1G3
OxBUhREs8AwZcfJ+QOdr+qqTfQ32SGxcET8Wu/TlviwJXHOJ9vA3+k9iboz5Z7Ge
6vGN4v0HV9hGZ+d26RHb02q/vqAaM1hKWs5/ISfP9kUWST5deOzClNICEaTNnJId
s36C2FsECkbxZ6Q9gcLeG5WB+COwOYMB2EwPQVWDGPSpW0kk/cQcaaKpQy6j9cd+
7DgrmRw0oIeWHKpDIbnXX2JL1U1BRKCljKI62Qj5fcclHNFfvTFuvk97vRu4cswh
BIbJ8tzSCwoYq7VabNMdFVArHOYRQWN5xAELhzlnSprRNb2XtEkfzTH4OFiKn+Ys
QZ1pyIvCwPWf9WuJIJ9MOQJw/jJ6F94sQtw7ajtRm/DcM4FHa0eb4EK13AHHfTcJ
R7riGUTol6cyPsM4hgZOEIIS8JNrg6/icNLRxsChTZRywCcMN/mA/+rDvLRdBrJc
s4Lh/J2o/5ayopdeGratl8qTmN/Az8woUfgzdG5eHBk2UBeKj4vrVJURTOk/2O5q
0oCAfd/AL4CdIL6JMPE89NhWt4aHRtpz3jzkv7UshXTQdkbdkH2HJzsaj7C2VzWW
QWaLzcaAT48hCZVIPzC15X9GclQPlE71jD5fcT/qZhuYuC2jLfumV52TTtJuweCP
Fp9EkfzsthxjUdHPThDZDV9wkhIYxjtiIciAUauaPACxwVO4gKnF71DLAGrsa/93
z7WOZEPihfVOlRG4Z0LB04HuuhmNx8E7kkXyW79kat8bTxsbfmS0Rupf3eom8iB/
fBL8EAZKLjYYlq2iIe+J3ObBQKblCujQ50MNXFrTZi1umdes3Rqx1FLzzdd7rMJ3
PB2UTzbdsuNKfze7HvRJX8OyJvb9/x+FdDOIBtxtZ41jVFpQZJV1Okv4xWCIZPwZ
9dH4XYDYUS8ETfN4DIKXdCNN/DnXJ0JX5nPn4VgsTr3kxY5lLLywUaB/cOOQMOhM
+lTIu+NsqaUKQl1AdCE/P3Swr/9KHsze8xYkwzFaDcK21IislSb8gTfaD1FU22VU
xKMmxjJo5Y850x2f0yjJVt+ruBx5t5vTvQH83QVm/T5WSpoWc38Qt2NaRimSadMG
01rmaSz0U5qWPm1rfGYv+a83WXKXFCrkc1n4abyrH/o2rurVkIj/h9Xz4e3+l3m+
WaGU3Ycedeh7LTOtavHVBTzYg9uMQOmYVUsXFSzgPifmkQRh0CPCg2f2fBWbju1E
KKil2r1y8WQWkQgqmzgtN/wk8siRI7c3IUTfHxvP08CRH8u+Qz8OnqrNUkitUx4m
a2rXCwyOuFxEV+t400iNAjSsP9nDbZR2+Ac4kYUN6R7UT0Ry/Arc0d/To0eUczi+
g8e3zjOyy/PnD+tZ0OiYJDZXyRPD42yyKOdXpnsy49Q3Jfg+byOLaY5eXa9+r55r
OlELt6tBBDb30vHbM0LyqHW09R1uxVu6NoHu+jMglXGCnvGS9ZDGqjIUVWkk035o
fCX9AABcTwnZc+EOIvWWQJGC+btFm20XSRuMxlhFeYEkNvGomW/iBbBvhjNql6Uw
VOvu3xgZ6WLovBVAEVEDGpGydrHN5+d9jRSEoTHHQcw0f9A7sCSkl8jGm2q20je8
uJ1SY5jYdUkc55pVArmj1mvPKtDJow3k1UUlTJQpaPlAriqHoUoNNjSLi1bVe97Y
yFz7QgnxjbLzZ9sohmQpCCZ/yK+c96vvYHONekh41tsQebzNFNOTNN607sPOPBCV
krvhygESBO2xM4D6qvySI79aSdQuFcpT2aKoFh0Xro4LJe4tAWMsvIqwKxpTfpAe
TPYRLfG6wl7nsqJVNG+Ej5TPx8Az5FJZOoy31TQJWrMP4Oz+/aPYTj/P92TJIsQU
3Fr7KoPY5w8lAGymUqEgNV1mjKLWH78zv4lnrv3yErfeGWaqq37scOHzCmj8HXEl
9+cx+30kmeUAJ4oXF9VjPxaxttTauHPsB0orWox1Ogzk2TM0jIQzw77w7GJX1Fxx
iByAEy/hCRi7KiFpZa0JyFL4kcPxohT6GtmEk+eK+jCxZO1AeFqv7NMAEPDlPD5D
Ce+witieqRXf2lLDY2X7SxIq9CPHxOt7jOCRYlxL62jjE2N85DKjjxie2pWKIjK/
Msmb6gIRNlkRcOCftUYaTxNJsDfUZJxu1VFPo9BnsG0W7TGAGUrL4OU45fI1qV8n
oW0dFVXQxn64awDgou5eFBzxCYO0CS8B2/ldGwTz2igDY3IaBsCHf1MBI2BJ5gJB
Phosf6GRgQ9xl6foNnfaO+9YEWDfou8ZvaVOyCsVinJcYZSvISbiJgCyiG/TCBo1
Xhovx8/wefzbjht0jB7Vn7Z9htCxs12zkpM2qSgsMMfAMwg7M1EoJvDTf5oge2EX
7fQGllKUE/ed2JVAU/sJD3rNJEWqp9Tl/cI+p7aw4aiAFirKutKdlbtu9dia1RX3
VAWuPLMb9OamKv5cI4/PNJy3wvQkqawUdS69E/CW9A6Z/AdYhO3pmx1Tl7WPDEvH
B5uNqSWg7+DK+4WB1+ijnxJc34NitleeWrObGsTvVgDTCIYPKDv0KYSZ3tTbwgYW
8QLfP4vc2uB6ppJD3bmvOp7ip/wbQr7D3bdEOcUuREjwpXsx+K+x0xR3pJLr6ORQ
ekRvgrVvQuqr/5/rLv7WGNW1LvtkARPAyGh45eXjZxtBoCvTkxQq4rEB8GOiGbJy
zQFUqY60MW/8/7l3em4GCUESvrFzD2d6j95s8d6HR7arK0VX3Cr34WzUlqtFdSdF
UQRP1/TZc1TcGnXeSo6EHJi+CjqeGUuwzkOtuh8kK4a9Ksh7Hs/CsxUBuaiM99tX
9F3OaYHFhbuAaa7Gf35crUwdkypmtynJGnVTbXy/B8zB2ZXQTvFajobY8eqkx8fT
4FCx+BhsE2MUC9/eZ/V+WiePSNN9yR4QkX3e4edHW1Nv0y/oohx8N51hNCYUcz0Y
WbfJsR2Oh519sJg+cObtDy+BOfEXHLnxh+RLBRga9/6yykD9djUro8Hdhj5l7f7e
9c9kK9YcX0ySvbwQNZeX3YtucUWlINX73trMiG6nbpTKy9L9xfYw7uO+t4xnqD/8
2rSd6q2u6n7JnRnRcptnqkmx3oqIr5h/VbtSaODEU8iyJPugst1OQAmsOO84r4EA
jVB4T6rNQefeOBBDOYkMDdb8HkbJyPdh9B0XqZe75LJTyA2eBkNjo4Z300dRW+fv
FxgO/7nGTU5FLw76AEuPIFYeRmornfnSgYZTLglnl4a/RmdoJ3kRY+aVlqvALljk
gihA4WPR4HeR+sgM6Bwws+1WnFCEPknHUkbTG4BgrWXS9mdwFNnV1IJ/jK0mhJg9
XNiB6NXC/jMcOVBni4Y8676II0dDH0ADEpwQAKP1JCz+qhZfWGNHqvqPuCt2EQuZ
e8VMJSxAHT3XEuLuj5DwFSGuGsNHZ3/hn/yvhF10O8a0ogAc3cBEK3P+eP05OFxa
+jf+e83Stl+xpQLZ3X3Sqdr9kjwOMSkcV2TBArXeJzz9pP4vmgaS+hrhY02GtshF
Se609HDMeIvzAKZCOiTlwRJhB4O41ZLY37QBrAI7E5Fsts+hHFruF6kXjYSVn1ds
QoDbTpQOFdfO9Zko9v2jgPxJEXokbpKQ2p8zwDfG18bnE5ZCqYD/acz6eMmiAI6m
NLSIAqgvRz5bDKddhy4Qc6xRlcNZAsKIUwvv2+7dCSKJlUY0R3YKnazKeH/h4Tkk
huz21GZ9fkzD67RhS0FDWCD9fWByvXB4aXwDJunPRasVGsstwhdF7qzYIwzxgGun
nVtClRESg+S8UNuSQOw+eN/Rt+DCblLtwryhglhrQDqJP6AXrS6wrlMv4pJ6qKVO
js8sBh+ZVMrLBbXhPnhK/3jWaXbYE/eZl3o77mVN5BYn4sLzXb4U6nPIGx8JuiDJ
ocj1wtHpGSlfMdZAHcVSctulBhSUPsc4lMlH0bhdSh5VZgujEug55KrJzDN/USoP
7gIh6qn0LJdkwtWsRsE+9tWIrkFox9bNIs3MdrRx4BtGb/Hoz1auHVd/MNli4wKO
6isH3S4BRHBa1macPTH6SCjD7/NlifJLmX2Z3wKp3G0hPmMC44eM10mqW9D0oPkL
s3NSYukJAvK3aqN4JSv9Ub8tmN7lmicvunMhw7VDewbK+R1jXQhKGuG/kIb2fYfu
1d/rBXLrp/ZXmEkSl12ZkqALDk9HIUslTWgb3SrAZhuHoHY5WosmAz5nR6DH4LOk
sar+o33paThB/bx1zyFFbDZ3/MHid5oZls52w2L7dU/5bClV/kFQUzv2wfASUdcw
ZE9TnWAvfCVRYFScQZGTof7nRZutWZEXR5fpsViOglkqWZWLktTLerUTNK11SLAl
tkNfUhb7daRfjYkpTf63C4aKG28hd2+fpnS+cmJcTQCYMEzhHsRc4+wE6H0VX0s4
woY9weHJFwQw+b4/RJC4V0xSFzzTZyZRkpvnXy2KstukqOEvacqKZSTaVpKx2rD9
vUvpOJ+VgtuVUR4aFAuzYUhpeax0o4Veli3ohW5ThOM3/n4oN7k/EeSC1VvosYX2
d3W+jf0l0X6TB+ltXGp6LEb/VzQyiYK585sCGskueXdRYJaVwZmeO4RxD4wf03n2
lQiMbYW2dMG7QYwf1JcJ47m9QBb8rwvBjdQxEb71FehKAd1cpdtg3kZNhQxcVgpk
gpcRb+8Ob6+lKbscdIFUe/LyDCMbRlwwIHbu0RMwRDQ4GxY2Ia2GmKtyhXPcmekZ
UPsCKnM1DxIQ7pHXCdlfArbuLkrBriBD/7t4TuW3j7YCd5vzXAOX2RZc+WpB+cmd
QfrZHwR8qhrzskwL0yDr5JJ2jPcEAXxZjh39+wm3xZADezZigsLgdHIkyBPyfYC2
mknag1orBAsxkOyC3J8t59vFhDPU2ylJmmXSQsIxo0/lGdmdaNl6jfPg7vDSn+YZ
w90DYJ8RMEzIdlJIcNkjuAogtGzHIhWOoKtMMmYM0rIbOGplxOiRxt+WV0eYsrEU
BtFhB3iQuw51UPxD1p0/c20tT/1xidXKHcQdvrPIMQiqaA3CcC7AsDnKmW3kLJ4e
vxY/WOw5F0pBDPUdVzVdRH17xCyI0mu5Q6RNGAjFGUFz0UqdPth+7UUb3WtNUMKB
35GHegQp8fUDbPETHQpjNsovI8Q7TTK23JhVriZyzdD3dsJnb+34hykRNWJ8Nd7P
OAoDxAwZYZTjJx1kerXRrsHHTYCe/u5b0Hm4m2xQiCl0yBfLnJwYHw0pmbIJh1bj
HtHKPpn7pZINdq+l9j18f7Lm/MFZ4AASO7o9j9Fz5LjlnrZ9BLprUvpm7ahiP7UR
D3fHs7Wns3Uhrjuje0ig1BJmjmoF3P1f1Thac6HsmESTW79FcVq4e4PUG03DvA5G
ytxNBlZUhognnRcfy7BNKB4CFi4y2IROaJfAM/1IlB+3g+PSdPC+wx3x4TvI22EL
SnD9xEV7dDXoyUBvcQOoqm6euYKuRPx7s799hSdZY2QeX1HE1lUqTaa+/ez7UuW3
XSxKdeJ9AGJsPDhv+o+tqmn1zrW0GNioG11aZjrhK3GGvsbwb+HlMY0evd+i/TO5
MxDx8ry4viaosc+Gb+s9yAfOuMElbdWoF4FnkGTBa5WHKDXSGHR0WuDNoYN4u22c
0wR0j8anbCboqo7PZq5zO9jzttAwbQ56t9YioURqdQmhjCw7p3YB1f0ruMzF3X1F
ZY5yxTKOk0ZRBMFNHLqHiTiuEaCehO1blFDpA/AkRQEUh0w2Rcd/hl7Yt3hdkUuG
xboVjEXZMCEGTYsxvbVVRiLujV4htbFWcAcMMg3ERtLUpsdNgfI0RpmaziQrfO6L
WKgx3OLh/w1GEHj4QAfUj4ukD2u2wMAkpUaZkgVWmYHqSpVMzxpbj4cfJ+twvd0Z
dmlrFkyEsrLJGiSogMLpCmAJju+oOM2lpL70vNIrXQPQjmCMwwD4PfLYZkWpmeBn
mrj0stieCSuOI0v8jzcpj5cuPpzR/5ckn5F9xo9tDJafAaD5RWKljC0orGNMc3Ej
+RRLK/gIX5KqeqJRqnX8IaM44fQAxE3tmQdnyfvfhBQZsWSF1Dbj3zBTgxwkJzpg
cpcgcz6wWlGjDrzgdPVcZJw5TKp0nbyps7DBjdbwUdmZrRhePaIeQxbqoAbrYO+V
PRc9CXEz2d59Bvwpnk5Dlq9JwPBLbFlKY8O5KQFhpbpBT1ljah2bQAC2z40sqVd+
DVoHt63C5hu3Hgqzv8ZFmjT/1zh6g6PbUPsDwSU+ftc=
//pragma protect end_data_block
//pragma protect digest_block
NqQk0XsOyi5l1vMQTo0ip+BI+mM=
//pragma protect end_digest_block
//pragma protect end_protected
